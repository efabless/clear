* NGSPICE file created from top_right_tile.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__sdfrtp_1 abstract view
.subckt sky130_fd_sc_hd__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__sdfrtp_2 abstract view
.subckt sky130_fd_sc_hd__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

.subckt top_right_tile VGND VPWR bottom_width_0_height_0_subtile_0__pin_cout_0_ bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ bottom_width_0_height_0_subtile_0__pin_reg_out_0_ bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ bottom_width_0_height_0_subtile_2__pin_inpad_0_ bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ ccff_head_0_0 ccff_head_1 ccff_tail ccff_tail_0 chanx_left_in[0] chanx_left_in[10]
+ chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15]
+ chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1]
+ chanx_left_in[20] chanx_left_in[21] chanx_left_in[22] chanx_left_in[23] chanx_left_in[24]
+ chanx_left_in[25] chanx_left_in[26] chanx_left_in[27] chanx_left_in[28] chanx_left_in[29]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10]
+ chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15]
+ chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1]
+ chanx_left_out[20] chanx_left_out[21] chanx_left_out[22] chanx_left_out[23] chanx_left_out[24]
+ chanx_left_out[25] chanx_left_out[26] chanx_left_out[27] chanx_left_out[28] chanx_left_out[29]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chany_bottom_in[0] chany_bottom_in[10]
+ chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14]
+ chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18]
+ chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[20] chany_bottom_in[21] chany_bottom_in[22]
+ chany_bottom_in[23] chany_bottom_in[24] chany_bottom_in[25] chany_bottom_in[26]
+ chany_bottom_in[27] chany_bottom_in[28] chany_bottom_in[29] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[20] chany_bottom_out[21] chany_bottom_out[22]
+ chany_bottom_out[23] chany_bottom_out[24] chany_bottom_out[25] chany_bottom_out[26]
+ chany_bottom_out[27] chany_bottom_out[28] chany_bottom_out[29] chany_bottom_out[2]
+ chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6]
+ chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9] clk0 gfpga_pad_io_soc_dir[0]
+ gfpga_pad_io_soc_dir[1] gfpga_pad_io_soc_dir[2] gfpga_pad_io_soc_dir[3] gfpga_pad_io_soc_dir_0[0]
+ gfpga_pad_io_soc_dir_0[1] gfpga_pad_io_soc_dir_0[2] gfpga_pad_io_soc_dir_0[3] gfpga_pad_io_soc_in[0]
+ gfpga_pad_io_soc_in[1] gfpga_pad_io_soc_in[2] gfpga_pad_io_soc_in[3] gfpga_pad_io_soc_in_0[0]
+ gfpga_pad_io_soc_in_0[1] gfpga_pad_io_soc_in_0[2] gfpga_pad_io_soc_in_0[3] gfpga_pad_io_soc_out[0]
+ gfpga_pad_io_soc_out[1] gfpga_pad_io_soc_out[2] gfpga_pad_io_soc_out[3] gfpga_pad_io_soc_out_0[0]
+ gfpga_pad_io_soc_out_0[1] gfpga_pad_io_soc_out_0[2] gfpga_pad_io_soc_out_0[3] isol_n
+ left_width_0_height_0_subtile_0__pin_inpad_0_ left_width_0_height_0_subtile_1__pin_inpad_0_
+ left_width_0_height_0_subtile_2__pin_inpad_0_ left_width_0_height_0_subtile_3__pin_inpad_0_
+ prog_clk prog_reset reset right_width_0_height_0_subtile_0__pin_O_10_ right_width_0_height_0_subtile_0__pin_O_11_
+ right_width_0_height_0_subtile_0__pin_O_12_ right_width_0_height_0_subtile_0__pin_O_13_
+ right_width_0_height_0_subtile_0__pin_O_14_ right_width_0_height_0_subtile_0__pin_O_15_
+ right_width_0_height_0_subtile_0__pin_O_8_ right_width_0_height_0_subtile_0__pin_O_9_
+ sc_in sc_out test_enable top_width_0_height_0_subtile_0__pin_O_0_ top_width_0_height_0_subtile_0__pin_O_1_
+ top_width_0_height_0_subtile_0__pin_O_2_ top_width_0_height_0_subtile_0__pin_O_3_
+ top_width_0_height_0_subtile_0__pin_O_4_ top_width_0_height_0_subtile_0__pin_O_5_
+ top_width_0_height_0_subtile_0__pin_O_6_ top_width_0_height_0_subtile_0__pin_O_7_
+ top_width_0_height_0_subtile_0__pin_cin_0_ top_width_0_height_0_subtile_0__pin_reg_in_0_
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_40_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_82_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l1_in_3__A1 net37 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_2_ net26 cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_43_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_53_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_53_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_363_ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_10.ccff_head
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_left_track_55.mux_l1_in_0__A0 net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_294_ sb_8__8_.mux_left_track_47.out VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mem_left_track_27.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_bottom_track_33.mux_l1_in_1_ net272 net6 sb_8__8_.mem_bottom_track_33.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_32_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net247 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_37.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_37.out sky130_fd_sc_hd__clkbuf_2
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_6_prog_clk sb_8__8_.mem_left_track_47.mem_out\[0\]
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_47.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l2_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_2_X cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_52_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_61_.in
+ sky130_fd_sc_hd__mux2_1
X_346_ sb_8__8_.mux_bottom_track_3.out VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_23_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_4__A1 net31 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_47.mux_l1_in_0__A1 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_3_ sb_8__8_.mux_left_track_29.out net9
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__228
+ VGND VGND VPWR VPWR net228 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__228/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_24_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__250
+ VGND VGND VPWR VPWR net250 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__250/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_55_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net218 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_29_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__8_.mux_left_track_13.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input55_A chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_329_ net4 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_2
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_3_X cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_0__A0 sb_8__8_.mux_left_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l1_in_2_ sb_8__8_.mux_bottom_track_21.out
+ net43 cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_13.out sky130_fd_sc_hd__buf_4
XFILLER_20_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_left_track_43.mux_l1_in_0_ net170 net62 sb_8__8_.mem_left_track_43.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_43.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_75_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_8_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_8_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_4__A1 net5 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_3_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output161_A net161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_55.mux_l2_in_0_ net310 sb_8__8_.mux_left_track_55.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_55.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_55.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_0__A0 sb_8__8_.mux_left_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_bottom_track_55.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_58_prog_clk
+ sb_8__8_.mem_bottom_track_55.mem_out\[0\] net175 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_55.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mem_bottom_track_25.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_2_ net14 sb_8__8_.mux_left_track_39.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_left_track_3.mux_l3_in_0_ sb_8__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X sb_8__8_.mem_left_track_3.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA__312__A sb_8__8_.mux_left_track_11.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input18_A chanx_left_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_30_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_0_ sb_8__8_.mux_left_track_5.out
+ net22 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_1_ net6 cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_5 cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__8_.mux_bottom_track_47.mux_l1_in_1__A1 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_1__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_ VGND
+ VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_22_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__307__A sb_8__8_.mux_left_track_21.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mux_bottom_track_1.mux_l1_in_0_ left_width_0_height_0_subtile_3__pin_inpad_0_
+ left_width_0_height_0_subtile_0__pin_inpad_0_ sb_8__8_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net233 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net237 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__mux2_4
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput97 net97 VGND VGND VPWR VPWR chanx_left_out[23] sky130_fd_sc_hd__buf_12
Xoutput86 net86 VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_28_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_0__A0 sb_8__8_.mux_left_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_left_track_3.mux_l2_in_1_ net296 net173 sb_8__8_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_16_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_2__S cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__240
+ VGND VGND VPWR VPWR net240 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__240/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__8_.mux_bottom_track_47.mux_l1_in_1__275 VGND VGND VPWR VPWR net275 sb_8__8_.mux_bottom_track_47.mux_l1_in_1__275/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_82_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_2_X cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l2_in_2__A0 net33 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_7_prog_clk sb_8__8_.mem_left_track_15.mem_out\[0\]
+ net176 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_15.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_22_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_85_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_2_ sb_8__8_.mux_left_track_17.out net16
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
X_362_ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_293_ sb_8__8_.mux_left_track_49.out VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_13_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_47.mux_l1_in_1__305 VGND VGND VPWR VPWR net305 sb_8__8_.mux_left_track_47.mux_l1_in_1__305/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_23_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_bottom_track_33.mux_l1_in_0_ net162 left_width_0_height_0_subtile_2__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_33.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_52_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_32_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_82_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_21.mux_l1_in_0__A0 net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_45.mux_l2_in_0_ sb_8__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_45.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_4_prog_clk sb_8__8_.mem_left_track_45.ccff_tail
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_47.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net73 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net75 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_32_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_58_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_70_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_79_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_345_ sb_8__8_.mux_bottom_track_5.out VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_2_ sb_8__8_.mux_left_track_17.out net16
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l2_in_2__A0 net58 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__315__A sb_8__8_.mux_left_track_5.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_3_X cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_82_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_33_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mux_bottom_track_1.mux_l1_in_1__A0 net161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_59.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_59.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_59.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_8__8_.mux_left_track_13.mux_l1_in_0__A1 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_1__A0 net8 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_input48_A chany_bottom_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
X_328_ net32 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_2
Xsb_8__8_.mem_bottom_track_23.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_7_prog_clk sb_8__8_.mem_bottom_track_23.mem_out\[0\]
+ net176 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_23.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_6_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l2_in_3_ net204 sb_8__8_.mux_bottom_track_45.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_45.mux_l1_in_1_ net274 net29 sb_8__8_.mem_bottom_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_56_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l1_in_1_ sb_8__8_.mux_bottom_track_9.out
+ net50 cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_3__184 VGND VGND VPWR VPWR net184 cbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_3__184/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l1_in_1__A1 net50 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_0__A1 net22 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__8_.mem_bottom_track_55.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_0_prog_clk sb_8__8_.mem_bottom_track_53.ccff_tail
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_55.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_ VGND VGND VPWR
+ VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__243
+ VGND VGND VPWR VPWR net243 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__243/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_1_ net4 cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net72
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_34_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_4__A0 net4 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_2__A1 net16 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_47_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_47_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_8__8_.mux_bottom_track_35.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_35.out sky130_fd_sc_hd__clkbuf_2
XFILLER_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_29_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_46_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__8_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_60_prog_clk
+ cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[2\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_2__A1 net18 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_1__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_bottom_track_9.mux_l2_in_1__284 VGND VGND VPWR VPWR net284 sb_8__8_.mux_bottom_track_9.mux_l2_in_1__284/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_89_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_bottom_track_1.mux_l2_in_1__259 VGND VGND VPWR VPWR net259 sb_8__8_.mux_bottom_track_1.mux_l2_in_1__259/LO
+ sky130_fd_sc_hd__conb_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_11.mux_l2_in_1__A1 net174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_55.mux_l1_in_0_ net168 net56 sb_8__8_.mem_left_track_55.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_55.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_25_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_4__A1 net5 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_38_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xoutput98 net98 VGND VGND VPWR VPWR chanx_left_out[24] sky130_fd_sc_hd__buf_12
Xoutput87 net87 VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_28_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input30_A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_2_ sb_8__8_.mux_left_track_27.out net10
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_0__A1 net22 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_3.mux_l2_in_0_ sb_8__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_56_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_42_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_29.out sky130_fd_sc_hd__clkbuf_2
XFILLER_54_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l2_in_2__A1 net31 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_38_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_3__A1 net41 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_22_prog_clk sb_8__8_.mem_left_track_13.ccff_tail
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_15.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_89_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_1_ sb_8__8_.mux_left_track_11.out net19
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
X_361_ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_292_ sb_8__8_.mux_left_track_51.out VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_9_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_50_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l2_in_3_ net209 sb_8__8_.mux_bottom_track_49.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_42_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_21_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_2__A1 net18 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_32_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_94_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__8_.mux_left_track_21.mux_l1_in_0__A1 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_left_track_3.mux_l1_in_1_ net170 net167 sb_8__8_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_88_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_88_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_0__A0 sb_8__8_.mux_left_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_344_ sb_8__8_.mux_bottom_track_7.out VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_1_ sb_8__8_.mux_left_track_11.out net19
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_2__A1 net48 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_34_prog_clk cby_8__8_.cby_8__8_.ccff_tail net177 VGND VGND VPWR VPWR
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net236 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mux_bottom_track_1.mux_l1_in_1__A1 net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_4_ net4 net35 cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_327_ net31 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mem_bottom_track_23.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_6_prog_clk sb_8__8_.mem_bottom_track_21.ccff_tail
+ net176 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_23.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l2_in_2_ net60 sb_8__8_.mux_bottom_track_27.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_45.mux_l1_in_0_ net164 left_width_0_height_0_subtile_0__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_45.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l1_in_0_ sb_8__8_.mux_bottom_track_3.out
+ net53 cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__326__A net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l1_in_4__A1 net60 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_9_X cby_8__8_.cby_8__8_.mem_right_ipin_8.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_57_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[2\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_bottom_track_57.mux_l2_in_0_ net281 sb_8__8_.mux_bottom_track_57.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_bottom_track_57.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_57.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net222 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input60_A chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l2_in_3__199 VGND VGND VPWR VPWR net199
+ cby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l2_in_3__199/LO sky130_fd_sc_hd__conb_1
XFILLER_34_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net178
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_4__A1 net35 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_41_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_16_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_16_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_29_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_32_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_bottom_track_51.mux_l1_in_1__278 VGND VGND VPWR VPWR net278 sb_8__8_.mux_bottom_track_51.mux_l1_in_1__278/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_46_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_ VGND VGND VPWR VPWR
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_60_prog_clk
+ cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[1\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_1.mux_l1_in_1__A0 net169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_3__319 VGND VGND VPWR VPWR net319 cbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_3__319/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_52_prog_clk
+ sb_8__8_.mem_bottom_track_29.mem_out\[0\] net176 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_29.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_40_prog_clk net2 net179 VGND VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_38_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput99 net99 VGND VGND VPWR VPWR chanx_left_out[25] sky130_fd_sc_hd__buf_12
XFILLER_76_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput88 net88 VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_28_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input23_A chanx_left_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_1_ sb_8__8_.mux_left_track_9.out net20
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_57.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_57.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_57.out sky130_fd_sc_hd__clkbuf_2
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mux_left_track_49.mux_l1_in_1__A1 net173 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net219 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__mux2_8
XFILLER_86_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_38_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__8_.mux_bottom_track_59.mux_l1_in_0__A0 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_0_ sb_8__8_.mux_left_track_5.out net22
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_360_ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_2
XFILLER_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_291_ sb_8__8_.mux_left_track_53.out VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_31_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_31_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l2_in_2_ net58 cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_42_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mux_bottom_track_15.mux_l2_in_0__262 VGND VGND VPWR VPWR net262 sb_8__8_.mux_bottom_track_15.mux_l2_in_0__262/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net178
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_13.mux_l2_in_0_ sb_8__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_13.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_59_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__329__A net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_3.mux_l1_in_0_ bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ net54 sb_8__8_.mem_left_track_3.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_0__A1 net22 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_73_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_51_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[2\] net175 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_3.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_343_ sb_8__8_.mux_bottom_track_9.out VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_0_ sb_8__8_.mux_left_track_5.out net22
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l2_in_3__204 VGND VGND VPWR VPWR net204
+ cby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l2_in_3__204/LO sky130_fd_sc_hd__conb_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net178
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_bottom_track_17.mux_l1_in_0__A0 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_3_ sb_8__8_.mux_bottom_track_25.out
+ net41 cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_13.mux_l1_in_1_ net287 net171 sb_8__8_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
X_326_ net30 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l2_in_1__A0 net38 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l2_in_1_ net40 cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_3.mux_l2_in_1__296 VGND VGND VPWR VPWR net296 sb_8__8_.mux_left_track_3.mux_l2_in_1__296/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__342__A sb_8__8_.mux_bottom_track_11.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_57_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[1\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_83_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_22_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_5.out sky130_fd_sc_hd__buf_4
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_1__A0 sb_8__8_.mux_left_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input53_A chany_bottom_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_61_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_21.mux_l2_in_0__291 VGND VGND VPWR VPWR net291 sb_8__8_.mux_left_track_21.mux_l2_in_0__291/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_2__A0 net14 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_309_ sb_8__8_.mux_left_track_17.out VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_61_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_37_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__232
+ VGND VGND VPWR VPWR net232 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__232/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_37_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_4__A0 net31 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_6_prog_clk sb_8__8_.mem_left_track_33.mem_out\[0\]
+ net176 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_33.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_56_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_56_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_29_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_2__A0 net26 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.out sky130_fd_sc_hd__clkbuf_1
XFILLER_8_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l1_in_2_ sb_8__8_.mux_bottom_track_15.out
+ net47 cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_36_prog_clk sb_8__8_.mem_bottom_track_5.mem_out\[1\]
+ net177 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_ VGND VGND VPWR VPWR
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ net81 net71 VGND VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__8_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_60_prog_clk
+ cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[0\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_3_ net318 sb_8__8_.mux_left_track_55.out
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_left_track_1.mux_l1_in_1__A1 bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net175
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_57.mux_l1_in_0_ net3 net162 sb_8__8_.mem_bottom_track_57.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_57.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_bottom_track_5.mux_l1_in_0__A0 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_59.mux_l1_in_1__312 VGND VGND VPWR VPWR net312 sb_8__8_.mux_left_track_59.mux_l1_in_1__312/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk
+ sb_8__8_.mem_bottom_track_27.ccff_tail net176 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_29.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput89 net89 VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_12
Xoutput78 net78 VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_0__pin_cout_0_
+ sky130_fd_sc_hd__buf_12
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_28_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_0_ sb_8__8_.mux_left_track_3.out net23
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input16_A chanx_left_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_27_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_48_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[2\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_6.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_1_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_1_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_54_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l1_in_0__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_59.mux_l1_in_0__A1 net163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input8_A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mux_bottom_track_11.mux_l2_in_1__260 VGND VGND VPWR VPWR net260 sb_8__8_.mux_bottom_track_11.mux_l2_in_1__260/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__8_.mux_left_track_15.mux_l1_in_1__A1 net172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_290_ sb_8__8_.mux_left_track_55.out VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_2__A0 net29 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_4_ sb_8__8_.mux_left_track_43.out
+ net31 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l2_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_2_X cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_42_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mux_bottom_track_25.mux_l1_in_0__A0 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_42_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net179 VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dfrtp_1
XFILLER_67_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__345__A sb_8__8_.mux_bottom_track_5.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l1_in_2__A1 net45 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_19_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_9_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_51_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[1\] net175 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_342_ sb_8__8_.mux_bottom_track_11.out VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_2
XFILLER_53_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_bottom_track_31.mux_l1_in_1__271 VGND VGND VPWR VPWR net271 sb_8__8_.mux_bottom_track_31.mux_l1_in_1__271/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_78_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_8__8_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mux_bottom_track_17.mux_l1_in_0__A1 left_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_3__A1 net7 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_67_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_12_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net254 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_2_ sb_8__8_.mux_bottom_track_13.out
+ net48 cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_51_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_13.mux_l1_in_0_ bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ net49 sb_8__8_.mem_left_track_13.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_325_ sb_8__8_.mux_bottom_track_45.out VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_3__A1 net9 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_25.mux_l2_in_0_ net293 sb_8__8_.mux_left_track_25.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_25.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_25.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__8_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_54_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[0\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_18_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_1__A1 net20 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input46_A chany_bottom_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_308_ sb_8__8_.mux_left_track_19.out VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_56_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[2\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_10.ccff_head
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net73 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net75 VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__sdfrtp_2
XFILLER_6_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_6_prog_clk sb_8__8_.mem_left_track_31.ccff_tail
+ net176 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_33.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_20_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_25_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_25_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_83_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_32_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l1_in_1_ sb_8__8_.mux_bottom_track_9.out
+ net50 cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_36_prog_clk sb_8__8_.mem_bottom_track_5.mem_out\[0\]
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_54_prog_clk
+ cby_8__8_.cby_8__8_.mem_left_ipin_1.ccff_tail net175 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_2_ net25 cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net258 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ net80 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_bottom_track_5.mux_l1_in_0__A1 left_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_left_track_9.mux_l2_in_1__314 VGND VGND VPWR VPWR net314 sb_8__8_.mux_left_track_9.mux_l2_in_1__314/LO
+ sky130_fd_sc_hd__conb_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_1__A0 sb_8__8_.mux_left_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_28_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput79 net79 VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_0__pin_reg_out_0_
+ sky130_fd_sc_hd__buf_12
XFILLER_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net73 grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_41_.in net75 VGND
+ VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_56_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_27_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mux_bottom_track_33.mux_l1_in_0__A0 net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__225
+ VGND VGND VPWR VPWR net225 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__225/LO
+ sky130_fd_sc_hd__conb_1
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_47_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[1\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_24_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.ccff_tail net71 VGND
+ VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_14_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[2\] net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_11.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_3_ sb_8__8_.mux_left_track_31.out
+ net8 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_40_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_40_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_left_track_39.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_61_prog_clk sb_8__8_.mem_left_track_39.mem_out\[0\]
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_39.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_76_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_42_prog_clk net324 net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_bottom_track_15.mux_l2_in_0_ net262 sb_8__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_bottom_track_15.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_bottom_track_25.mux_l1_in_0__A1 net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l2_in_3_ net191 sb_8__8_.mux_bottom_track_49.out
+ cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_41_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_51.mux_l2_in_0__308 VGND VGND VPWR VPWR net308 sb_8__8_.mux_left_track_51.mux_l2_in_0__308/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_18_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_19_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_50_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[0\] net175 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_341_ sb_8__8_.mux_bottom_track_13.out VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mux_left_track_5.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input76_A top_width_0_height_0_subtile_0__pin_cin_0_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_5_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_3.mux_l2_in_1__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_1__A0 sb_8__8_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_2__A0 net3 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_1_ sb_8__8_.mux_bottom_track_7.out
+ net51 cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_4_ net4 net35 cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_324_ sb_8__8_.mux_bottom_track_47.out VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_11.out sky130_fd_sc_hd__buf_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_1.out sky130_fd_sc_hd__buf_4
XANTENNA_sb_8__8_.mux_left_track_19.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk
+ sb_8__8_.mem_bottom_track_47.mem_out\[0\] net176 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_47.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_54_prog_clk
+ cby_8__8_.cby_8__8_.mem_left_ipin_3.ccff_tail net175 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_18_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l2_in_3_ net200 sb_8__8_.mux_bottom_track_47.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cby_8__8_.cby_8__8_.mem_left_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input39_A chany_bottom_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_307_ sb_8__8_.mux_left_track_21.out VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__8_.mux_left_track_31.mux_l1_in_1__A1 net172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_56_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[1\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_88_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_3_ net319 sb_8__8_.mux_left_track_57.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__215
+ VGND VGND VPWR VPWR net215 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__215/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_33_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_16_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[2\] net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_14.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l1_in_0_ sb_8__8_.mux_bottom_track_3.out
+ net53 cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_36_prog_clk sb_8__8_.mem_bottom_track_3.ccff_tail
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_25.mux_l1_in_0_ net169 net42 sb_8__8_.mem_left_track_25.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_25.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_86_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_1_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_2_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_23_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_load_slew179_A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__258
+ VGND VGND VPWR VPWR net258 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__258/LO
+ sky130_fd_sc_hd__conb_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__8_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_47_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[2\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_11.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_left_track_37.mux_l2_in_0_ net300 sb_8__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_37.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_18_prog_clk cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.ccff_tail
+ net177 VGND VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_28_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_33.mux_l1_in_0__A1 left_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_47_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[0\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_31_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_13.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l2_in_2__A0 net61 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_4_ sb_8__8_.mux_left_track_45.out net30
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_31_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_14_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\] net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__8_.mem_left_track_57.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net72 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net256 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__mux2_4
XFILLER_42_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_2_ sb_8__8_.mux_left_track_19.out
+ net15 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_59.mux_l2_in_0__282 VGND VGND VPWR VPWR net282 sb_8__8_.mux_bottom_track_59.mux_l2_in_0__282/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_49_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_22_prog_clk sb_8__8_.mem_left_track_3.mem_out\[1\]
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_left_track_39.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_1_prog_clk sb_8__8_.mem_left_track_37.ccff_tail
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_39.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_40_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input21_A chanx_left_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_3_ net181 sb_8__8_.mux_left_track_49.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l2_in_2_ net58 cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cbx_8__8_.cbx_1__8_.mem_top_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_18_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_bottom_track_7.mux_l3_in_0_ sb_8__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X sb_8__8_.mem_bottom_track_7.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_19_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_50_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_2.ccff_tail net176 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_340_ sb_8__8_.mux_bottom_track_15.out VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_8__8_.mux_left_track_5.mux_l1_in_0__A1 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input69_A gfpga_pad_io_soc_in_0[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_6__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__8_.mux_left_track_27.mux_l1_in_0__A0 net170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_1__A1 net19 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_3_ net186 sb_8__8_.mux_left_track_49.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_34_prog_clk
+ sb_8__8_.mem_bottom_track_15.mem_out\[0\] net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_15.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk sb_8__8_.mem_left_track_51.mem_out\[0\]
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_51.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_0_ sb_8__8_.mux_bottom_track_1.out
+ net54 cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_4_ sb_8__8_.mux_left_track_37.out net5
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_15.mux_l1_in_0_ net16 left_width_0_height_0_subtile_1__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_15.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_19_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_19_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_58_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_3_ sb_8__8_.mux_bottom_track_25.out
+ net41 cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
X_323_ sb_8__8_.mux_bottom_track_49.out VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_2
XFILLER_80_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__8_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net72
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_bottom_track_27.mux_l2_in_0_ net268 sb_8__8_.mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_bottom_track_27.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_17_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[2\] net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__8_.mux_bottom_track_7.mux_l1_in_1__A0 net161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_bottom_track_7.mux_l2_in_1_ net283 net20 sb_8__8_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l1_in_1__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_52_prog_clk
+ sb_8__8_.mem_bottom_track_45.ccff_tail net175 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_47.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_9_X cbx_8__8_.cbx_1__8_.mem_top_ipin_14.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net177 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l2_in_2_ net59 sb_8__8_.mux_bottom_track_35.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mem_bottom_track_55.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_47_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[2\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_14.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_8_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[2\] net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_306_ sb_8__8_.mux_left_track_23.out VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_55_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[0\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l1_in_1__A1 net50 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_33.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_33.out sky130_fd_sc_hd__clkbuf_2
XFILLER_18_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_2_ net14 cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_33_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_3.mux_l2_in_1__A1 net173 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_16_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[1\] net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net177 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_34_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_34_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_5.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input51_A chany_bottom_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net65 cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_1__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net178
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_47_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[1\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_38_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net73 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net75 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_41_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_60_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_46_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_5.ccff_tail net175 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mux_left_track_27.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_27.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_27.out sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__230
+ VGND VGND VPWR VPWR net230 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__230/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__214
+ VGND VGND VPWR VPWR net214 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__214/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_3__189 VGND VGND VPWR VPWR net189 cbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_3__189/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_35_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mux_bottom_track_45.mux_l1_in_1__274 VGND VGND VPWR VPWR net274 sb_8__8_.mux_bottom_track_45.mux_l1_in_1__274/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_3_ sb_8__8_.mux_left_track_33.out net7
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_4__A1 net5 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_7_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net178
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_12_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[0\] net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__222
+ VGND VGND VPWR VPWR net222 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__222/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_1_ sb_8__8_.mux_left_track_7.out
+ net21 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_35.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_22_prog_clk sb_8__8_.mem_left_track_3.mem_out\[0\]
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_76_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_40_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_2_ net28 cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input14_A chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_45.mux_l1_in_1__304 VGND VGND VPWR VPWR net304 sb_8__8_.mux_left_track_45.mux_l1_in_1__304/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_83_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mux_left_track_37.mux_l1_in_0_ net167 net36 sb_8__8_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l2_in_1_ cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_41_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_left_track_49.mux_l2_in_0_ sb_8__8_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_49.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mem_left_track_55.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net72 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net239 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_18_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input6_A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net69 cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR left_width_0_height_0_subtile_1__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_53_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_3_X cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_left_track_27.mux_l1_in_0__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_51.mux_l2_in_0_ net308 sb_8__8_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_51.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_20_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[2\] net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_3.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_3__320 VGND VGND VPWR VPWR net320 cbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_3__320/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_2_ net28 sb_8__8_.mux_left_track_31.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_34_prog_clk
+ sb_8__8_.mem_bottom_track_13.ccff_tail net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_15.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ net79 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_0__A0 sb_8__8_.mux_left_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_4_prog_clk sb_8__8_.mem_left_track_49.ccff_tail
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_51.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_3_ sb_8__8_.mux_left_track_25.out net11
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_59_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_59_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_2_ sb_8__8_.mux_bottom_track_13.out
+ net48 cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
X_322_ sb_8__8_.mux_bottom_track_51.out VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
XFILLER_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output168_A net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l2_in_3__195 VGND VGND VPWR VPWR net195
+ cby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l2_in_3__195/LO sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__8_.mem_left_track_41.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net72 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_0__A0 sb_8__8_.mux_left_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_20_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[1\] net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_23_prog_clk sb_8__8_.mem_left_track_9.mem_out\[1\]
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_33_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_bottom_track_29.mux_l1_in_1__269 VGND VGND VPWR VPWR net269 sb_8__8_.mux_bottom_track_29.mux_l1_in_1__269/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__8_.mux_left_track_49.mux_l1_in_1_ net306 net173 sb_8__8_.mem_left_track_49.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_bottom_track_7.mux_l1_in_1__A1 net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_bottom_track_7.mux_l2_in_0_ sb_8__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_68_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_47_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[1\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l2_in_1_ net36 cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_8_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[1\] net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net175
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_305_ sb_8__8_.mux_left_track_25.out VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_46_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_8.ccff_tail net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l2_in_3__197 VGND VGND VPWR VPWR net197
+ cby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l2_in_3__197/LO sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_11_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__8_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_4_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_4_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_50_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_13_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\] net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__242
+ VGND VGND VPWR VPWR net242 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__242/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_24_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mux_bottom_track_27.mux_l1_in_0_ net9 net159 sb_8__8_.mem_bottom_track_27.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_24_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input44_A chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_0__A0 sb_8__8_.mux_left_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_left_track_57.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_61_prog_clk sb_8__8_.mem_left_track_57.mem_out\[0\]
+ net72 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_57.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mux_bottom_track_7.mux_l1_in_1_ net161 net158 sb_8__8_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_19_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_1__A0 net8 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l1_in_2_ sb_8__8_.mux_bottom_track_17.out
+ net46 cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_47_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[0\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xsb_8__8_.mux_bottom_track_7.mux_l2_in_1__283 VGND VGND VPWR VPWR net283 sb_8__8_.mux_bottom_track_7.mux_l2_in_1__283/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l2_in_2__A0 net58 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.out sky130_fd_sc_hd__clkbuf_1
XFILLER_21_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mux_left_track_43.mux_l1_in_0__A0 net170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__8_.mux_left_track_55.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_55.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_55.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__8_.mem_bottom_track_59.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_7.mux_l1_in_1__A0 net169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_2__A0 sb_8__8_.mux_left_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_2_ sb_8__8_.mux_left_track_21.out net13
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_9_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[2\] net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_6.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_12_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_10.ccff_tail net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_3_X cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_0_ sb_8__8_.mux_left_track_1.out
+ net24 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_left_track_35.mux_l1_in_0__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_7_prog_clk sb_8__8_.mem_left_track_1.ccff_tail
+ net176 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_8__8_.cby_8__8_.mux_left_ipin_2.out cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_40_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_2_X cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_0__S cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_49.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_49.out sky130_fd_sc_hd__buf_4
XFILLER_79_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l2_in_2__A0 net57 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net238 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__mux2_4
XFILLER_50_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_41_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_19_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_bottom_track_31.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_31.out sky130_fd_sc_hd__clkbuf_2
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_1_0__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_15_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_20_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[1\] net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_1_ net8 cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_0__A1 net22 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_95_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_2_ sb_8__8_.mux_left_track_13.out net18
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_1__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_28_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_28_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_73_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_1_ sb_8__8_.mux_bottom_track_7.out
+ net51 cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_321_ sb_8__8_.mux_bottom_track_53.out VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input74_A sc_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l2_in_1__A0 net34 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_0__A1 net24 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_17_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\] net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xsb_8__8_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_22_prog_clk sb_8__8_.mem_left_track_9.mem_out\[0\]
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_9.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_left_track_49.mux_l1_in_0_ bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ net59 sb_8__8_.mem_left_track_49.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_40_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_25.out sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_59_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_ VGND VGND VPWR
+ VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__254
+ VGND VGND VPWR VPWR net254 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__254/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_16_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_47_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[0\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_2__A1 net15 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_24_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_left_track_51.mux_l1_in_0_ bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ net58 sb_8__8_.mem_left_track_51.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mux_bottom_track_35.mux_l1_in_1__A1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_3__A1 net41 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_9.mux_l3_in_0_ sb_8__8_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__8_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_2_X sb_8__8_.mem_left_track_11.ccff_head
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_left_track_25.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_61_prog_clk sb_8__8_.mem_left_track_25.mem_out\[0\]
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_25.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_46_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_8_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\] net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_304_ sb_8__8_.mux_left_track_27.out VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_2_ sb_8__8_.mux_left_track_19.out net15
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net178
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_7_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_2__A1 net17 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_51.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_16_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[2\] net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_10.ccff_head
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_9_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_13.ccff_tail net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xsb_8__8_.mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_19.out sky130_fd_sc_hd__clkbuf_2
XFILLER_10_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_0__A1 net24 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_left_track_57.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_61_prog_clk sb_8__8_.mem_left_track_55.ccff_tail
+ net72 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_57.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_input37_A chany_bottom_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_43_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_43_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_8__8_.mux_bottom_track_7.mux_l1_in_0_ left_width_0_height_0_subtile_3__pin_inpad_0_
+ left_width_0_height_0_subtile_0__pin_inpad_0_ sb_8__8_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_3__S cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l2_in_3__209 VGND VGND VPWR VPWR net209
+ cby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l2_in_3__209/LO sky130_fd_sc_hd__conb_1
XFILLER_42_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l2_in_3_ net205 sb_8__8_.mux_bottom_track_53.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net217 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l1_in_1_ sb_8__8_.mux_bottom_track_11.out
+ net49 cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_56_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_10.ccff_tail net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_3__A1 net40 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_9.mux_l2_in_1_ net314 net173 sb_8__8_.mem_left_track_9.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_48_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_7.mux_l1_in_1__A1 bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net228 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_35.mux_l1_in_1__299 VGND VGND VPWR VPWR net299 sb_8__8_.mux_left_track_35.mux_l1_in_1__299/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_35_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_2__A1 net13 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_1_ sb_8__8_.mux_left_track_9.out net20
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_load_slew177_A net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_9_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[1\] net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_52_prog_clk
+ sb_8__8_.mem_bottom_track_33.mem_out\[0\] net175 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_33.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_3__A1 sb_8__8_.mux_left_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_0__A0 sb_8__8_.mux_left_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_4_ net31 net62 cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_39_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_25_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_bottom_track_13.mux_l2_in_0__261 VGND VGND VPWR VPWR net261 sb_8__8_.mux_bottom_track_13.mux_l2_in_0__261/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_94_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_4__A1 net32 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_19_prog_clk net325 net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_9_X cby_8__8_.cby_8__8_.mem_right_ipin_4.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_53.mux_l2_in_0_ net279 sb_8__8_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_bottom_track_53.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_2__A0 sb_8__8_.mux_left_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_15_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_20_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[0\] net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_8__8_.cby_8__8_.mux_left_ipin_0.out cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_67_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_1_ sb_8__8_.mux_left_track_7.out net21
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_0_ sb_8__8_.mux_bottom_track_1.out
+ net54 cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_54_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_53.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_53.out sky130_fd_sc_hd__clkbuf_2
X_320_ sb_8__8_.mux_bottom_track_55.out VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_2
XFILLER_54_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l2_in_3_ net210 sb_8__8_.mux_bottom_track_57.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input67_A gfpga_pad_io_soc_in_0[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_68_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_16_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.ccff_tail net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xsb_8__8_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_21_prog_clk sb_8__8_.mem_left_track_7.ccff_tail
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_9.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_15_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_48_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_13.ccff_tail net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_55_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_3__322 VGND VGND VPWR VPWR net322 cbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_3__322/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_left_track_25.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_61_prog_clk sb_8__8_.mem_left_track_23.ccff_tail
+ net72 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_25.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_46_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_11_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.ccff_tail net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_1_ sb_8__8_.mux_left_track_7.out net21
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
X_303_ sb_8__8_.mux_left_track_29.out VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output173_A net173 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_ VGND VGND
+ VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_37_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_51.mux_l1_in_0__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.ccff_tail
+ net177 VGND VGND VPWR VPWR cby_8__8_.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_bottom_track_47.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_47.out sky130_fd_sc_hd__clkbuf_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_17_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[1\] net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net178
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_12_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_12_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l2_in_2_ net56 cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l1_in_0_ sb_8__8_.mux_bottom_track_5.out
+ net52 cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_26_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_10.ccff_head
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mux_left_track_9.mux_l2_in_0_ sb_8__8_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_9.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net72
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_2__A0 sb_8__8_.mux_bottom_track_17.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_29.mux_l1_in_1__A1 net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_0_ sb_8__8_.mux_left_track_3.out net23
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__8_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__D cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_1__A0 sb_8__8_.mux_left_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_13_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\] net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_7_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk
+ sb_8__8_.mem_bottom_track_31.ccff_tail net176 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_33.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.out cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
Xsb_8__8_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_1.out sky130_fd_sc_hd__buf_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_88_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_3_ sb_8__8_.mux_bottom_track_29.out
+ net39 cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_39_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_20_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_9.mux_l1_in_1_ net170 net167 sb_8__8_.mem_left_track_9.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_51.mux_l1_in_1__A1 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_3__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_25_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_4__A0 net31 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input12_A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_2__A1 net13 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net220 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__mux2_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_15_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_17_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_2.ccff_tail net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_0_ sb_8__8_.mux_left_track_1.out net24
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input4_A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__8_.mux_bottom_track_9.mux_l2_in_1__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l2_in_2_ net44 net32 cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_37_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_37_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_77_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_ VGND VGND VPWR VPWR
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_49_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_41_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_2__A0 net26 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_72_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_1.mux_l2_in_1__285 VGND VGND VPWR VPWR net285 sb_8__8_.mux_left_track_1.mux_l2_in_1__285/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_15_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_11.mux_l3_in_0_ sb_8__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X sb_8__8_.mem_bottom_track_11.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_53.mux_l1_in_0_ net25 net160 sb_8__8_.mem_bottom_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_83_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_4__A0 net30 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net73 grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_50_.in net75 VGND
+ VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_2__A0 net25 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_0_ sb_8__8_.mux_left_track_1.out net24
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
X_302_ sb_8__8_.mux_left_track_31.out VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_ VGND VGND
+ VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_77_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_16_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[0\] net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_sb_8__8_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l2_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_2_X cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_52_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_52_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_8__8_.mux_bottom_track_11.mux_l2_in_1_ net260 net18 sb_8__8_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net235 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_A
+ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.ccff_tail VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_bottom_track_47.mux_l1_in_0__A0 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_26_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_left_track_7.mux_l2_in_1__313 VGND VGND VPWR VPWR net313 sb_8__8_.mux_left_track_7.mux_l2_in_1__313/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_left_track_27.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_10_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_2__A0 net28 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_input42_A chany_bottom_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_16_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_5.ccff_tail net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_2_ sb_8__8_.mux_bottom_track_17.out
+ net46 cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_39_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_22_prog_clk sb_8__8_.mem_left_track_11.mem_out\[1\]
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__8_.mux_left_track_19.mux_l2_in_0_ net290 sb_8__8_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_19.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_3_X cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__8_.mux_left_track_9.mux_l1_in_0_ bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ net51 sb_8__8_.mem_left_track_9.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_21.mux_l2_in_0_ net291 sb_8__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_21.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__245
+ VGND VGND VPWR VPWR net245 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__245/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__212
+ VGND VGND VPWR VPWR net212 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__212/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__8_.mem_left_track_43.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_2_prog_clk sb_8__8_.mem_left_track_43.mem_out\[0\]
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_43.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_15_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.out cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_9_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_3__A1 net8 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_7_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_7_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_86_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__8_.mem_bottom_track_25.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l2_in_1_ net34 cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net249 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__mux2_4
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_ VGND VGND VPWR VPWR
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_77_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_41_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__D
+ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.ccff_tail VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_17.mux_l1_in_1__289 VGND VGND VPWR VPWR net289 sb_8__8_.mux_left_track_17.mux_l1_in_1__289/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_54_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_3__190 VGND VGND VPWR VPWR net190 cbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_3__190/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_15_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__8_.mux_left_track_45.mux_l1_in_1__A1 net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_4__A1 net61 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_41_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_3__317 VGND VGND VPWR VPWR net317
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_3__317/LO sky130_fd_sc_hd__conb_1
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_301_ sb_8__8_.mux_left_track_33.out VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input72_A prog_reset VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_55.mux_l1_in_0__A0 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_3__A1 net11 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output159_A net159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_11.mux_l1_in_1__A0 net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_53_prog_clk
+ sb_8__8_.mem_bottom_track_51.mem_out\[0\] net175 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_51.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_14_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_8.ccff_tail net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_68_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l1_in_2_ sb_8__8_.mux_bottom_track_27.out
+ net40 cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_1__A0 sb_8__8_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_11.mux_l2_in_0_ sb_8__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_51_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_21_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__8_.mux_bottom_track_47.mux_l1_in_0__A1 left_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mux_left_track_9.mux_l2_in_1__A1 net173 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l2_in_3__193 VGND VGND VPWR VPWR net193 cby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l2_in_3__193/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_6_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_13.mux_l1_in_0__A0 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input35_A chany_bottom_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_3__187 VGND VGND VPWR VPWR net187 cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_3__187/LO
+ sky130_fd_sc_hd__conb_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__224
+ VGND VGND VPWR VPWR net224 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__224/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mem_left_track_25.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_1_ sb_8__8_.mux_bottom_track_11.out
+ net49 cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_11.mux_l1_in_1_ net163 net160 sb_8__8_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_57.mux_l2_in_0__281 VGND VGND VPWR VPWR net281 sb_8__8_.mux_bottom_track_57.mux_l2_in_0__281/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__8_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_22_prog_clk sb_8__8_.mem_left_track_11.mem_out\[0\]
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_27_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_28_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_load_slew175_A net176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_left_track_57.mux_l2_in_0__311 VGND VGND VPWR VPWR net311 sb_8__8_.mux_left_track_57.mux_l2_in_0__311/LO
+ sky130_fd_sc_hd__conb_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_2__A0 net28 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_66_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mem_left_track_43.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_61_prog_clk sb_8__8_.mem_left_track_41.ccff_tail
+ net72 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_43.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_45_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_15_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_41_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_left_track_19.mux_l1_in_0_ bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ net46 sb_8__8_.mem_left_track_19.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net72
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_bottom_track_1.mux_l1_in_0__A0 left_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_46_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_46_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l2_in_3_ net192 sb_8__8_.mux_bottom_track_51.out
+ cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_left_track_21.mux_l1_in_0_ net167 net45 sb_8__8_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_33_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net73 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net75 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_50_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_9_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_0__S cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_15_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_33.mux_l2_in_0_ sb_8__8_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_33.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__252
+ VGND VGND VPWR VPWR net252 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__252/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__8_.mem_bottom_track_23.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_300_ sb_8__8_.mux_left_track_35.out VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_2
XFILLER_50_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_55.mux_l1_in_0__A1 net161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input65_A gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mux_left_track_11.mux_l1_in_1__A1 net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_39_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk sb_8__8_.mem_left_track_49.mem_out\[0\]
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_49.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_41_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk
+ sb_8__8_.mem_bottom_track_49.ccff_tail net176 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_51.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l1_in_1_ sb_8__8_.mux_bottom_track_9.out
+ net50 cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xinput1 ccff_head_0_0 VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_bottom_track_21.mux_l1_in_0__A0 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_1__A1 net19 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xclkbuf_0_prog_clk prog_clk VGND VGND VPWR VPWR clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_4_ net32 net34 cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net178
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_3_ net321 sb_8__8_.mux_left_track_53.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_output171_A net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_61_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_61_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_8__8_.mux_left_track_33.mux_l1_in_1_ net298 net173 sb_8__8_.mem_left_track_33.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_27_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net253 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__236
+ VGND VGND VPWR VPWR net236 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__236/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_65_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l2_in_2__A0 net44 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_1__A1 net21 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_0__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l2_in_3_ net201 sb_8__8_.mux_bottom_track_49.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__313__A sb_8__8_.mux_left_track_9.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_24_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_9_X cby_8__8_.cby_8__8_.mem_left_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__8_.mux_bottom_track_3.mux_l3_in_0_ sb_8__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X sb_8__8_.mem_bottom_track_3.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_13.mux_l1_in_0__A1 left_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_3__A1 net11 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_79_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input28_A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l2_in_2__A0 net58 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_left_track_49.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l2_in_3__201 VGND VGND VPWR VPWR net201
+ cby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l2_in_3__201/LO sky130_fd_sc_hd__conb_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net224 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_3_ net320 sb_8__8_.mux_left_track_59.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput70 gfpga_pad_io_soc_in_0[3] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.ccff_tail net71 VGND
+ VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_2__A1 net48 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_0_ sb_8__8_.mux_bottom_track_5.out
+ net52 cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_11.mux_l1_in_0_ net165 left_width_0_height_0_subtile_2__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_11.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_4_ sb_8__8_.mux_left_track_41.out net32
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mem_bottom_track_57.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_58_prog_clk
+ sb_8__8_.mem_bottom_track_57.mem_out\[0\] net175 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_57.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_23_prog_clk sb_8__8_.mem_left_track_11.ccff_head
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_44_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_26_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_79_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_26_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_94_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_bottom_track_23.mux_l2_in_0_ net266 sb_8__8_.mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_bottom_track_23.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_4_ net4 net35 cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_1__A1 net21 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_3__S cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_bottom_track_3.mux_l2_in_1_ net270 net22 sb_8__8_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_left_track_29.mux_l1_in_1__295 VGND VGND VPWR VPWR net295 sb_8__8_.mux_left_track_29.mux_l1_in_1__295/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_9_X cbx_8__8_.cbx_1__8_.mem_top_ipin_10.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_3__181 VGND VGND VPWR VPWR net181 cbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_3__181/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_15_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_9_X cby_8__8_.cby_8__8_.mem_right_ipin_14.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l2_in_3__210 VGND VGND VPWR VPWR net210
+ cby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l2_in_3__210/LO sky130_fd_sc_hd__conb_1
XFILLER_4_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_bottom_track_11.mux_l2_in_1__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mux_bottom_track_1.mux_l1_in_0__A1 left_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net178
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_3_ net182 sb_8__8_.mux_left_track_51.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mux_left_track_23.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_23.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_23.out sky130_fd_sc_hd__clkbuf_2
XFILLER_89_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l2_in_2_ net57 cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input10_A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_15_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_15_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_9_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_6_prog_clk sb_8__8_.mem_left_track_17.mem_out\[0\]
+ net176 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_17.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_15_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__316__A sb_8__8_.mux_left_track_3.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net231 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__mux2_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l1_in_3__A1 net37 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_53_prog_clk
+ cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[2\] net175 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net245 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input2_A ccff_head_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__248
+ VGND VGND VPWR VPWR net248 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__248/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input58_A chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_39_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_3_ net187 sb_8__8_.mux_left_track_57.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_4_prog_clk sb_8__8_.mem_left_track_47.ccff_tail
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_49.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_36_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
X_359_ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_8__8_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_3__A1 net41 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l1_in_0_ sb_8__8_.mux_bottom_track_3.out
+ net53 cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xinput2 ccff_head_1 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mux_left_track_17.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_17.out sky130_fd_sc_hd__clkbuf_2
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mux_bottom_track_21.mux_l1_in_0__A1 net164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_7.out sky130_fd_sc_hd__buf_4
XFILLER_32_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_3_ sb_8__8_.mux_bottom_track_27.out
+ net40 cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__8_.mux_left_track_57.mux_l1_in_0__A0 net169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_2_ net26 cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l2_in_3__207 VGND VGND VPWR VPWR net207
+ cby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l2_in_3__207/LO sky130_fd_sc_hd__conb_1
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output164_A net164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_left_track_33.mux_l1_in_0_ bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ net38 sb_8__8_.mem_left_track_33.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_29_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_38_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_30_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_30_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_8__8_.mux_left_track_1.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l2_in_2_ net58 cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_20_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mux_left_track_45.mux_l2_in_0_ sb_8__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_45.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_56_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mem_bottom_track_25.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_35_prog_clk
+ sb_8__8_.mem_bottom_track_25.mem_out\[0\] net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_25.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_4_ sb_8__8_.mux_left_track_45.out net30
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mux_left_track_49.mux_l1_in_0__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_2_ net3 sb_8__8_.mux_left_track_41.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput71 isol_n VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_4
Xinput60 chany_bottom_in[7] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_2
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_3_ sb_8__8_.mux_left_track_29.out net9
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mem_bottom_track_57.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_57_prog_clk
+ sb_8__8_.mem_bottom_track_55.ccff_tail net175 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_57.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__8_.mux_left_track_15.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_9_X cbx_8__8_.cbx_1__8_.mem_top_ipin_6.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_0__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_3__A1 sb_8__8_.mux_left_track_57.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input40_A chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_3_ sb_8__8_.mux_bottom_track_25.out
+ net41 cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_left_track_45.mux_l1_in_1_ net304 net171 sb_8__8_.mem_left_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_7_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_0__A0 sb_8__8_.mux_left_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_bottom_track_3.mux_l2_in_0_ sb_8__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_59_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_18_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_23_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_43_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.ccff_tail net71 VGND
+ VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_51.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_51.out sky130_fd_sc_hd__clkbuf_2
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_2__A0 sb_8__8_.mux_left_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_2_ net27 sb_8__8_.mux_left_track_39.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_23.mux_l1_in_0_ net11 net165 sb_8__8_.mem_bottom_track_23.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_89_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_41_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l2_in_1_ cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_2_X cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_3.mux_l1_in_1_ net162 net159 sb_8__8_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_9_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_55_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_55_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_sb_8__8_.mux_bottom_track_49.mux_l1_in_1__A1 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_7_prog_clk sb_8__8_.mem_left_track_15.ccff_tail
+ net176 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_17.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_bottom_track_35.mux_l2_in_0_ sb_8__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_35.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_15_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_24_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_53_prog_clk
+ cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[1\] net175 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net175
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_0__A0 sb_8__8_.mux_left_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_45.out sky130_fd_sc_hd__buf_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_39_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_33_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_2_ net14 cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
X_358_ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_1
X_289_ sb_8__8_.mux_left_track_57.out VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput3 chanx_left_in[0] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__dlymetal6s2s_1
Xsb_8__8_.mux_left_track_39.mux_l2_in_0__301 VGND VGND VPWR VPWR net301 sb_8__8_.mux_left_track_39.mux_l2_in_0__301/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l2_in_2__A0 net60 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_3__A0 sb_8__8_.mux_bottom_track_29.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__327__A net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_2_ sb_8__8_.mux_bottom_track_15.out
+ net47 cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_0_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_35.mux_l1_in_1_ net273 net5 sb_8__8_.mem_bottom_track_35.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_2_X cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input70_A gfpga_pad_io_soc_in_0[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_29_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_34_prog_clk sb_8__8_.mem_bottom_track_1.mem_out\[1\]
+ net177 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_76_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_1.mux_l1_in_0__A1 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_68_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l2_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_2_X cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_left_track_23.mux_l1_in_0__A0 net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mem_bottom_track_25.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_52_prog_clk
+ sb_8__8_.mem_bottom_track_23.ccff_tail net176 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_25.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_left_track_39.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_39.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_39.out sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
Xoutput170 net170 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_3_ sky130_fd_sc_hd__buf_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_3_ sb_8__8_.mux_left_track_33.out net7
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_21.out sky130_fd_sc_hd__clkbuf_2
Xsb_8__8_.mux_left_track_33.mux_l1_in_1__298 VGND VGND VPWR VPWR net298 sb_8__8_.mux_left_track_33.mux_l1_in_1__298/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_62_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_37_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[2\] net176 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_49_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_1_ net32 cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net242 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput50 chany_bottom_in[25] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_4
Xinput61 chany_bottom_in[8] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_2
Xinput72 prog_reset VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_12
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_2_ sb_8__8_.mux_left_track_17.out net16
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__255
+ VGND VGND VPWR VPWR net255 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__255/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__8_.mux_bottom_track_3.mux_l1_in_1__A0 net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__8_.mux_left_track_15.mux_l1_in_0__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_37_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_1__A0 net6 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_3_X cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input33_A chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_2_ sb_8__8_.mux_bottom_track_13.out
+ net48 cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_45.mux_l1_in_0_ bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ net61 sb_8__8_.mem_left_track_45.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_5_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_4__A0 net4 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_57.mux_l2_in_0_ net311 sb_8__8_.mux_left_track_57.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_57.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_57.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_15.out sky130_fd_sc_hd__clkbuf_2
XFILLER_1_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_18_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_23_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_5.mux_l3_in_0_ sb_8__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X sb_8__8_.mem_left_track_5.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_9_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_2_ sb_8__8_.mux_left_track_23.out net12
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net234 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_ VGND
+ VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_2__A1 net13 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_1_ net4 cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_46_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_left_track_43.mux_l2_in_0__303 VGND VGND VPWR VPWR net303 sb_8__8_.mux_left_track_43.mux_l2_in_0__303/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__8_.mux_bottom_track_3.mux_l1_in_0_ net164 left_width_0_height_0_subtile_1__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_3.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_24_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_24_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l2_in_3_ net195 sb_8__8_.mux_bottom_track_57.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_2__A1 net16 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_54_prog_clk
+ cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[0\] net175 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_59_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_5.mux_l2_in_1_ net307 net174 sb_8__8_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_18_prog_clk cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.ccff_tail
+ net177 VGND VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_4__A1 net32 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_10_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_0__A1 net23 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_38_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_2_X cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_81_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_357_ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net213 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__mux2_8
XANTENNA_sb_8__8_.mux_left_track_31.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_288_ sb_8__8_.mux_left_track_59.out VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_2_ sb_8__8_.mux_left_track_21.out net13
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_46_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[2\] net176 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_5.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xinput4 chanx_left_in[10] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_4
XFILLER_49_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_4__A1 net5 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_3__A1 net39 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__343__A sb_8__8_.mux_bottom_track_9.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_1_ sb_8__8_.mux_bottom_track_9.out
+ net50 cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_bottom_track_35.mux_l1_in_0_ net163 left_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_35.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_4_ sb_8__8_.mux_bottom_track_45.out
+ net60 cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input63_A gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_29_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_39_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_34_prog_clk sb_8__8_.mem_bottom_track_1.mem_out\[0\]
+ net177 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_93_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_2__A1 net16 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_bottom_track_47.mux_l2_in_0_ sb_8__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_47.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_27.mux_l2_in_0__268 VGND VGND VPWR VPWR net268 sb_8__8_.mux_bottom_track_27.mux_l2_in_0__268/LO
+ sky130_fd_sc_hd__conb_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cby_8__8_.cby_8__8_.mem_right_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_0__A0 sb_8__8_.mux_left_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput160 net160 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_12_
+ sky130_fd_sc_hd__buf_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_2_ sb_8__8_.mux_left_track_21.out net13
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xoutput171 net171 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_4_ sky130_fd_sc_hd__buf_12
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_50_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[1\] net176 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput40 chany_bottom_in[16] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_2
Xinput73 reset VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_8
Xinput62 chany_bottom_in[9] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_2
Xinput51 chany_bottom_in[26] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_4
XFILLER_88_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_1_ sb_8__8_.mux_left_track_11.out net19
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__8_.mux_bottom_track_3.mux_l1_in_1__A1 net159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_25_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_37_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l2_in_3_ net206 sb_8__8_.mux_bottom_track_49.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_47.mux_l1_in_1_ net275 net28 sb_8__8_.mem_bottom_track_47.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_48_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_1_ sb_8__8_.mux_bottom_track_7.out
+ net51 cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input26_A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_49_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_49_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_73_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_4_prog_clk sb_8__8_.mem_left_track_35.mem_out\[0\]
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_35.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net73 grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_59_.in net75 VGND
+ VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_ VGND VGND VPWR
+ VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_4__A1 net35 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_36_prog_clk sb_8__8_.mem_bottom_track_7.mem_out\[1\]
+ net177 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_7.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__8_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_18_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_1_ sb_8__8_.mux_left_track_11.out net19
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_70_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_0__A0 sb_8__8_.mux_left_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_46_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[2\] net176 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_8.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__346__A sb_8__8_.mux_bottom_track_3.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_1__A0 net32 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_34_prog_clk
+ sb_8__8_.mem_bottom_track_11.mem_out\[1\] net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_11.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l2_in_2_ net44 cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_left_track_3.mux_l1_in_1__A0 net170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_ VGND VGND
+ VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mux_left_track_57.mux_l1_in_0_ net169 net55 sb_8__8_.mem_left_track_57.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_57.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_63_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_5.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_50_prog_clk
+ cby_8__8_.cby_8__8_.mem_left_ipin_0.ccff_tail net176 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_59_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_left_track_5.mux_l2_in_0_ sb_8__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_86_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_3__315 VGND VGND VPWR VPWR net315
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_3__315/LO sky130_fd_sc_hd__conb_1
XFILLER_39_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_0_prog_clk_A prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_39_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_356_ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_8__8_.mux_left_track_31.mux_l1_in_0__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_1_ sb_8__8_.mux_left_track_9.out net20
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_46_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[1\] net175 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput5 chanx_left_in[11] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_2
XFILLER_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_0_ sb_8__8_.mux_bottom_track_3.out
+ net53 cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ net76 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_34_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_3_ sb_8__8_.mux_bottom_track_33.out
+ net37 cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_12_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[2\] net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_10.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_29_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input56_A chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_23_prog_clk cby_8__8_.ccff_tail
+ net177 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_339_ sb_8__8_.mux_bottom_track_17.out VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
Xsb_8__8_.mux_left_track_5.mux_l1_in_1_ net171 net168 sb_8__8_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l2_in_3__191 VGND VGND VPWR VPWR net191 cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l2_in_3__191/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_
+ sky130_fd_sc_hd__clkbuf_1
Xoutput150 net150 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[0] sky130_fd_sc_hd__buf_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_1_ sb_8__8_.mux_left_track_9.out net20
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xoutput161 net161 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_13_
+ sky130_fd_sc_hd__buf_12
Xoutput172 net172 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_5_ sky130_fd_sc_hd__buf_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_1__A1 net50 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output162_A net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_49_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[0\] net175 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_3__185 VGND VGND VPWR VPWR net185 cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_3__185/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l2_in_1__A0 net38 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_bottom_track_19.mux_l1_in_0__A0 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput30 chanx_left_in[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_4
Xinput63 gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_1
Xinput41 chany_bottom_in[17] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_2
Xinput52 chany_bottom_in[27] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_2
Xinput74 sc_in VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_0_ sb_8__8_.mux_left_track_5.out net22
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__244
+ VGND VGND VPWR VPWR net244 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__244/LO
+ sky130_fd_sc_hd__conb_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l2_in_2_ net58 sb_8__8_.mux_bottom_track_31.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_47.mux_l1_in_0_ net165 left_width_0_height_0_subtile_1__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_47.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_31_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__218
+ VGND VGND VPWR VPWR net218 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__218/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_2__A1 net12 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_48_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_0_ sb_8__8_.mux_bottom_track_1.out
+ net54 cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input19_A chanx_left_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_18_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_18_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_85_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_6_prog_clk sb_8__8_.mem_left_track_33.ccff_tail
+ net176 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_35.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_31.mux_l1_in_1__A1 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_bottom_track_59.mux_l2_in_0_ net282 sb_8__8_.mux_bottom_track_59.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_bottom_track_59.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_59.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net72
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_36_prog_clk sb_8__8_.mem_bottom_track_7.mem_out\[0\]
+ net177 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_34_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_19_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__227
+ VGND VGND VPWR VPWR net227 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__227/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_0_ sb_8__8_.mux_left_track_5.out net22
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_24_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_2__A0 net28 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_63_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_ VGND VGND VPWR VPWR
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_0__A1 net22 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_46_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[1\] net176 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_36_prog_clk
+ sb_8__8_.mem_bottom_track_11.mem_out\[0\] net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_11.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_59.mux_l1_in_1__A1 net174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_58_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_left_track_15.mux_l1_in_1__288 VGND VGND VPWR VPWR net288 sb_8__8_.mux_left_track_15.mux_l1_in_1__288/LO
+ sky130_fd_sc_hd__conb_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l2_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_8__8_.mux_left_track_3.mux_l1_in_1__A1 net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_10_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[2\] net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_13.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_ VGND VGND
+ VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_48_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_33_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_33_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_32_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__8_.mux_bottom_track_7.mux_l1_in_0__A0 left_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l1_in_0__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net178
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__8_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_59_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[2\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_10.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_39_prog_clk net326 net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_355_ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__8_.mux_bottom_track_59.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_59.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_59.out sky130_fd_sc_hd__clkbuf_1
XFILLER_5_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_0_ sb_8__8_.mux_left_track_3.out net23
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_48_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[0\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_64_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput6 chanx_left_in[12] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net215 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mux_left_track_17.mux_l1_in_1__A1 net173 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_43_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_52_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l1_in_2__A1 net48 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_2__A0 net27 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_2_ sb_8__8_.mux_bottom_track_21.out
+ net43 cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net178
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_15.mux_l2_in_0_ sb_8__8_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_15.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_51_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_11_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[1\] net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_29_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input49_A chany_bottom_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_3_ net315 sb_8__8_.mux_left_track_49.out
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_3_X cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_bottom_track_27.mux_l1_in_0__A0 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_338_ sb_8__8_.mux_bottom_track_19.out VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
Xsb_8__8_.mux_left_track_5.mux_l1_in_0_ bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ net53 sb_8__8_.mem_left_track_5.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput151 net151 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[1] sky130_fd_sc_hd__buf_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_0_ sb_8__8_.mux_left_track_3.out net23
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xoutput140 net140 VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_12
Xoutput173 net173 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_6_ sky130_fd_sc_hd__buf_12
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net63 cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_3__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
Xoutput162 net162 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_14_
+ sky130_fd_sc_hd__buf_12
XFILLER_87_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__8_.mem_left_track_55.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net72 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk
+ sb_8__8_.mem_bottom_track_49.mem_out\[0\] net176 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_49.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_54_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_1.ccff_tail net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_30_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_bottom_track_19.mux_l1_in_0__A1 left_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput31 chanx_left_in[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_2
Xinput20 chanx_left_in[25] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_4
Xinput64 gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_3__A1 net11 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xinput42 chany_bottom_in[18] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput53 chany_bottom_in[28] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_4
Xinput75 test_enable VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_8
XFILLER_57_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mux_left_track_15.mux_l1_in_1_ net288 net172 sb_8__8_.mem_left_track_15.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_52_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_55.mux_l2_in_0__280 VGND VGND VPWR VPWR net280 sb_8__8_.mux_bottom_track_55.mux_l2_in_0__280/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_4_ sb_8__8_.mux_left_track_37.out
+ net5 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net73 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net75 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_59_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l2_in_1_ net38 cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_31_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_58_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_58_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_55.mux_l2_in_0__310 VGND VGND VPWR VPWR net310 sb_8__8_.mux_left_track_55.mux_l2_in_0__310/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_36_prog_clk sb_8__8_.mem_bottom_track_5.ccff_tail
+ net177 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_14_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[2\] net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__241
+ VGND VGND VPWR VPWR net241 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__241/LO
+ sky130_fd_sc_hd__conb_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_48_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__8_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_56_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[2\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_13.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_7.out sky130_fd_sc_hd__buf_4
XFILLER_95_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input31_A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_ VGND VGND VPWR VPWR
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_48_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net67 cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR left_width_0_height_0_subtile_3__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_8_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__8_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net175
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__237
+ VGND VGND VPWR VPWR net237 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__237/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__8_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_46_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[0\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xsb_8__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_37_prog_clk
+ sb_8__8_.mem_bottom_track_11.ccff_head net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_11.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l1_in_2_ sb_8__8_.mux_bottom_track_19.out
+ net45 cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_3_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_3_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.out sky130_fd_sc_hd__clkbuf_1
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_4_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_bottom_track_59.mux_l1_in_0_ net24 net163 sb_8__8_.mem_bottom_track_59.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_59.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.out sky130_fd_sc_hd__clkbuf_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_3_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[1\] net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_bottom_track_7.mux_l1_in_0__A1 left_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_21_prog_clk sb_8__8_.mem_left_track_5.mem_out\[1\]
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_86_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_26_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_82_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_60_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[1\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__8_.mux_bottom_track_35.mux_l1_in_0__A0 net163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_31_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__234
+ VGND VGND VPWR VPWR net234 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__234/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_354_ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_8__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mem_bottom_track_59.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_57_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_4.ccff_tail net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xinput7 chanx_left_in[13] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
XFILLER_91_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_1__A0 sb_8__8_.mux_left_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_24_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_61_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_70_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net175
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net250 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__mux2_4
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_1_ sb_8__8_.mux_bottom_track_9.out
+ net50 cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_10_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\] net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_52_prog_clk
+ sb_8__8_.mem_bottom_track_17.mem_out\[0\] net176 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_17.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_29_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_2_ net28 cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l2_in_3__205 VGND VGND VPWR VPWR net205
+ cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l2_in_3__205/LO sky130_fd_sc_hd__conb_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_27.mux_l1_in_0__A1 net159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_25_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_61_prog_clk sb_8__8_.mem_left_track_53.mem_out\[0\]
+ net72 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_53.ccff_tail sky130_fd_sc_hd__dfrtp_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_337_ sb_8__8_.mux_bottom_track_21.out VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput152 net152 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[2] sky130_fd_sc_hd__buf_12
Xoutput141 net141 VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_12
Xoutput130 net130 VGND VGND VPWR VPWR chany_bottom_out[26] sky130_fd_sc_hd__buf_12
Xoutput174 net174 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_7_ sky130_fd_sc_hd__buf_12
Xoutput163 net163 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_15_
+ sky130_fd_sc_hd__buf_12
XFILLER_87_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_11_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[2\] net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net175
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_7.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk
+ sb_8__8_.mem_bottom_track_47.ccff_tail net176 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_49.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ net77 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input61_A chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__8_.mux_bottom_track_5.mux_l2_in_1__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_1__A0 sb_8__8_.mux_left_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput10 chanx_left_in[16] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_2
Xinput21 chanx_left_in[26] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__253
+ VGND VGND VPWR VPWR net253 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__253/LO
+ sky130_fd_sc_hd__conb_1
Xinput32 chanx_left_in[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_4
Xinput54 chany_bottom_in[29] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_4
Xinput43 chany_bottom_in[19] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_2
Xinput76 top_width_0_height_0_subtile_0__pin_cin_0_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_1
Xinput65 gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_2__A0 net30 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_57_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_16_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[2\] net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_69_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_15.mux_l1_in_0_ bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ net48 sb_8__8_.mem_left_track_15.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_92_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_38_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_3_ sb_8__8_.mux_left_track_25.out
+ net11 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_30_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net72 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mux_left_track_27.mux_l2_in_0_ net294 sb_8__8_.mux_left_track_27.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_27.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_27.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_20_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_27_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_27_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_14_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[1\] net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net66 cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_0__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_56_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[1\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input24_A chanx_left_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_33.mux_l1_in_1__A1 net173 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mem_left_track_59.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_56_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_7.ccff_tail net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net178
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l1_in_1_ sb_8__8_.mux_bottom_track_7.out
+ net51 cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.ccff_tail
+ net177 VGND VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_0__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_32_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_38_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_4_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[0\] net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_2__A0 net26 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_34_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__8_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_22_prog_clk sb_8__8_.mem_left_track_5.mem_out\[0\]
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_42_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_42_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l2_in_3_ net197 sb_8__8_.mux_bottom_track_53.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_26_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_82_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_5__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_60_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[0\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_40_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_35.mux_l1_in_0__A1 left_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_31_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_2__A1 net48 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_353_ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net70 cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR left_width_0_height_0_subtile_0__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
Xsb_8__8_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_0_prog_clk sb_8__8_.mem_left_track_21.mem_out\[0\]
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_21.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l2_in_2__A0 net59 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput8 chanx_left_in[14] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_2
XFILLER_64_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_1__A1 net20 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_79_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_88_.in
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_19_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mux_bottom_track_17.mux_l2_in_0_ net263 sb_8__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_bottom_track_17.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_14_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[2\] net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_5.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_0_ sb_8__8_.mux_bottom_track_3.out
+ net53 cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l2_in_3_ net193 sb_8__8_.mux_bottom_track_53.out
+ cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_13_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_10.ccff_head net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xsb_8__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_35_prog_clk
+ sb_8__8_.mem_bottom_track_15.ccff_tail net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_17.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_1_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l2_in_2__A0 net44 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_bottom_track_57.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_26_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_0_prog_clk sb_8__8_.mem_left_track_51.ccff_tail
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_53.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_bottom_track_5.mux_l2_in_1__277 VGND VGND VPWR VPWR net277 sb_8__8_.mux_bottom_track_5.mux_l2_in_1__277/LO
+ sky130_fd_sc_hd__conb_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_4_ net31 net62 cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
X_336_ sb_8__8_.mux_bottom_track_23.out VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_4__A1 net60 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_bottom_track_3.mux_l2_in_1__270 VGND VGND VPWR VPWR net270 sb_8__8_.mux_bottom_track_3.mux_l2_in_1__270/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_41_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_2__A1 net47 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xoutput142 net142 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[0] sky130_fd_sc_hd__buf_12
Xoutput120 net120 VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_12
Xoutput131 net131 VGND VGND VPWR VPWR chany_bottom_out[27] sky130_fd_sc_hd__buf_12
Xoutput153 net153 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[3] sky130_fd_sc_hd__buf_12
Xoutput164 net164 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_8_ sky130_fd_sc_hd__buf_12
XFILLER_87_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_3_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[1\] net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net251 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mux_left_track_7.mux_l1_in_0__A1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_left_track_29.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_9_X cby_8__8_.cby_8__8_.mem_right_ipin_10.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input54_A chany_bottom_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__289__A sb_8__8_.mux_left_track_57.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_1__A1 net20 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_319_ sb_8__8_.mux_bottom_track_57.out VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_1
Xinput11 chanx_left_in[17] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_2
Xinput22 chanx_left_in[27] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_2
Xinput33 chany_bottom_in[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput44 chany_bottom_in[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_2
Xinput55 chany_bottom_in[2] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_86_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xinput77 top_width_0_height_0_subtile_0__pin_reg_in_0_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_1
Xinput66 gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_1
XFILLER_69_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_16_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[1\] net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_4_ net31 net62 cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_92_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_2_ sb_8__8_.mux_left_track_13.out
+ net18 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_31_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_3_ net322 sb_8__8_.mux_left_track_43.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_19_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output160_A net160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__8_.mux_bottom_track_9.mux_l1_in_1__A0 net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l2_in_3_ net202 sb_8__8_.mux_bottom_track_51.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_13.out sky130_fd_sc_hd__clkbuf_2
XFILLER_34_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l1_in_1__A1 net50 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cby_8__8_.cby_8__8_.mem_left_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_bottom_track_51.mux_l1_in_0__A0 net159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_3__A1 net9 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_3.out sky130_fd_sc_hd__buf_4
Xsb_8__8_.mem_left_track_59.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_2_prog_clk sb_8__8_.mem_left_track_59.mem_out\[0\]
+ net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.ccff_head sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_14_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\] net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_38_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_56_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[0\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_68_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input17_A chanx_left_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_1__A0 sb_8__8_.mux_left_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_1__S cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_3_ net183 sb_8__8_.mux_left_track_49.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l1_in_0_ sb_8__8_.mux_bottom_track_1.out
+ net54 cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__226
+ VGND VGND VPWR VPWR net226 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__226/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_89_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__8_.mux_left_track_5.mux_l2_in_1__A1 net174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_27.mux_l1_in_0_ net170 net41 sb_8__8_.mem_left_track_27.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_27.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input9_A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_33_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_14_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[2\] net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_8.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__8_.mux_left_track_39.mux_l2_in_0_ net301 sb_8__8_.mux_left_track_39.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_39.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_39.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_8_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_12.ccff_tail net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_23_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_22_prog_clk sb_8__8_.mem_left_track_3.ccff_tail
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_11.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net178
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l2_in_2_ net56 cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_11_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_11_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_left_track_41.mux_l2_in_0_ net302 sb_8__8_.mux_left_track_41.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_41.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_41.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__8_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_57_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_10.ccff_head net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_31_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_4_ sb_8__8_.mux_left_track_37.out net5
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
X_352_ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_2
XFILLER_60_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_0_prog_clk sb_8__8_.mem_left_track_19.ccff_tail
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_21.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput9 chanx_left_in[15] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_18_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_37.mux_l2_in_0__300 VGND VGND VPWR VPWR net300 sb_8__8_.mux_left_track_37.mux_l2_in_0__300/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_32_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_57_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mem_left_track_43.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mux_left_track_11.mux_l2_in_1__286 VGND VGND VPWR VPWR net286 sb_8__8_.mux_left_track_11.mux_l2_in_1__286/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_14_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[1\] net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mux_left_track_37.mux_l1_in_0__A0 net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cbx_8__8_.cbx_1__8_.mem_top_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l2_in_2_ net56 cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l2_in_2__A1 net32 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_26_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_3_ sb_8__8_.mux_bottom_track_29.out
+ net39 cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
X_335_ sb_8__8_.mux_bottom_track_25.out VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mux_bottom_track_9.mux_l3_in_0_ sb_8__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_2_X sb_8__8_.mem_bottom_track_11.ccff_head
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net232 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__mux2_8
XFILLER_49_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput110 net110 VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_12
Xoutput143 net143 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[1] sky130_fd_sc_hd__buf_12
Xoutput132 net132 VGND VGND VPWR VPWR chany_bottom_out[28] sky130_fd_sc_hd__buf_12
Xoutput121 net121 VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_12
Xoutput154 net154 VGND VGND VPWR VPWR gfpga_pad_io_soc_out_0[0] sky130_fd_sc_hd__buf_12
Xoutput165 net165 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_9_ sky130_fd_sc_hd__buf_12
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_3_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\] net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_sb_8__8_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_29.mux_l1_in_0__A1 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_3_ net188 sb_8__8_.mux_left_track_53.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_left_track_31.mux_l1_in_1__297 VGND VGND VPWR VPWR net297 sb_8__8_.mux_left_track_31.mux_l1_in_1__297/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_87_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net177 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input47_A chany_bottom_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_4__S cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_318_ sb_8__8_.mux_bottom_track_59.out VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_1
Xinput12 chanx_left_in[18] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dlymetal6s2s_1
Xsb_8__8_.mux_bottom_track_17.mux_l1_in_0_ net15 left_width_0_height_0_subtile_2__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_17.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_0__A0 sb_8__8_.mux_left_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput45 chany_bottom_in[20] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput34 chany_bottom_in[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
Xinput23 chanx_left_in[28] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_4
Xinput67 gfpga_pad_io_soc_in_0[0] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_1
Xinput56 chany_bottom_in[3] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_44_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__8_.mem_left_track_27.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk sb_8__8_.mem_left_track_27.mem_out\[0\]
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_27.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_84_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_14_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\] net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_3_ sb_8__8_.mux_bottom_track_29.out
+ net39 cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_1_ sb_8__8_.mux_left_track_7.out
+ net21 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_29.mux_l2_in_0_ sb_8__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_29.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_2_ net31 sb_8__8_.mux_left_track_31.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_30_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_41.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_41.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_41.out sky130_fd_sc_hd__clkbuf_2
XFILLER_43_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_bottom_track_9.mux_l2_in_1_ net284 net19 sb_8__8_.mem_bottom_track_9.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__8_.mux_bottom_track_9.mux_l1_in_1__A1 net159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l2_in_2_ net57 net32 cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_31.mux_l2_in_0_ sb_8__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_31.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net177 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_36_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_36_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_sb_8__8_.mux_bottom_track_51.mux_l1_in_0__A1 left_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_77_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net178
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_left_track_59.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_2_prog_clk sb_8__8_.mem_left_track_57.ccff_tail
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_59.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_89_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_3_prog_clk
+ cbx_8__8_.cbx_1__8_.ccff_head net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_37_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_3__A0 sb_8__8_.mux_bottom_track_29.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_56_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_12.ccff_tail net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_16_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_2_ net28 cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_39_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mux_bottom_track_29.mux_l1_in_1_ net269 net8 sb_8__8_.mem_bottom_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_35.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_35.out sky130_fd_sc_hd__clkbuf_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_7.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_41_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_14_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[1\] net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_41.mux_l2_in_0__302 VGND VGND VPWR VPWR net302 sb_8__8_.mux_left_track_41.mux_l2_in_0__302/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__8_.mux_bottom_track_31.mux_l1_in_1_ net271 net7 sb_8__8_.mem_bottom_track_31.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_53_prog_clk
+ sb_8__8_.mem_bottom_track_35.mem_out\[0\] net175 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_35.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net223 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_bottom_track_29.mux_l1_in_1__A1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_1__A0 net6 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l2_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_2_X cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_47_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_51_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_51_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__8_.mux_left_track_45.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_left_track_27.mux_l2_in_0__294 VGND VGND VPWR VPWR net294 sb_8__8_.mux_left_track_27.mux_l2_in_0__294/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__8_.mux_left_track_9.mux_l1_in_1__A0 net170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_31_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_3_ sb_8__8_.mux_left_track_25.out net11
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_351_ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input77_A top_width_0_height_0_subtile_0__pin_reg_in_0_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_39_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_29.out sky130_fd_sc_hd__clkbuf_2
XFILLER_49_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__219
+ VGND VGND VPWR VPWR net219 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__219/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_91_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net240 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_3_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_11.out sky130_fd_sc_hd__buf_4
XFILLER_67_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_14_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[0\] net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_70_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__211
+ VGND VGND VPWR VPWR net211 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__211/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_23_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_left_track_39.mux_l1_in_0_ net168 net35 sb_8__8_.mem_left_track_39.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_39.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l2_in_1_ cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net73 grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_68_.in net75 VGND
+ VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_76_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_3_X cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_26_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_2_ sb_8__8_.mux_bottom_track_17.out
+ net46 cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
X_334_ sb_8__8_.mux_bottom_track_27.out VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_2
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_bottom_track_25.mux_l2_in_0__267 VGND VGND VPWR VPWR net267 sb_8__8_.mux_bottom_track_25.mux_l2_in_0__267/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mux_left_track_41.mux_l1_in_0_ net169 net34 sb_8__8_.mem_left_track_41.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_41.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_4__A0 sb_8__8_.mux_left_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_3_X cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput100 net100 VGND VGND VPWR VPWR chanx_left_out[26] sky130_fd_sc_hd__buf_12
Xoutput111 net111 VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_12
Xoutput133 net133 VGND VGND VPWR VPWR chany_bottom_out[29] sky130_fd_sc_hd__buf_12
Xoutput122 net122 VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_12
Xoutput155 net155 VGND VGND VPWR VPWR gfpga_pad_io_soc_out_0[1] sky130_fd_sc_hd__buf_12
Xoutput144 net144 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[2] sky130_fd_sc_hd__buf_12
Xoutput166 net166 VGND VGND VPWR VPWR sc_out sky130_fd_sc_hd__buf_12
Xsb_8__8_.mux_left_track_53.mux_l2_in_0_ net309 sb_8__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_53.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_11_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.ccff_tail net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_95_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_1__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_2_ net26 sb_8__8_.mux_left_track_35.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_left_track_1.mux_l3_in_0_ sb_8__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X sb_8__8_.mem_left_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_3__183 VGND VGND VPWR VPWR net183 cbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_3__183/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_317_ sb_8__8_.mux_left_track_1.out VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_1
XFILLER_42_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput13 chanx_left_in[19] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xinput46 chany_bottom_in[21] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_2
Xinput35 chany_bottom_in[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_2
Xinput24 chanx_left_in[29] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_4
Xinput68 gfpga_pad_io_soc_in_0[1] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput57 chany_bottom_in[4] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_45_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net176 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_27.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_0_prog_clk sb_8__8_.mem_left_track_25.ccff_tail
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_27.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_10_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_1.ccff_tail net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_2_ sb_8__8_.mux_bottom_track_17.out
+ net46 cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_0_ sb_8__8_.mux_left_track_1.out
+ net24 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l1_in_1__A1 net50 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_1_ net8 cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_31_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_6_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_6_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mux_bottom_track_9.mux_l2_in_0_ sb_8__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_9.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_11_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_59_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l2_in_1_ net34 cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_66_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_2__A1 net12 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_ VGND
+ VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_1.mux_l2_in_1_ net285 net172 sb_8__8_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_21_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_3__A1 net39 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__8_.mux_left_track_53.mux_l1_in_0__A0 net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_37_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_2__A1 net15 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__8_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mux_bottom_track_29.mux_l1_in_0_ net160 left_width_0_height_0_subtile_0__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_29.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_2_ sb_8__8_.mux_left_track_13.out net18
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.ccff_tail net71 VGND
+ VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_39_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_bottom_track_9.mux_l1_in_1_ net162 net159 sb_8__8_.mem_bottom_track_9.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_14_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\] net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_70_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l1_in_2_ sb_8__8_.mux_bottom_track_21.out
+ net43 cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__8_.mux_bottom_track_31.mux_l1_in_0_ net161 left_width_0_height_0_subtile_1__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_31.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_52_prog_clk
+ sb_8__8_.mem_bottom_track_33.ccff_tail net175 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_35.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_23_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input22_A chanx_left_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__223
+ VGND VGND VPWR VPWR net223 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__223/LO
+ sky130_fd_sc_hd__conb_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_8__8_.mem_left_track_39.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_4__A1 net4 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_45.mux_l1_in_0__A1 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_3__A1 net38 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_20_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_20_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_35_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_9.mux_l1_in_1__A1 net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_57.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_57.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_57.out sky130_fd_sc_hd__buf_4
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_2_ sb_8__8_.mux_left_track_13.out net18
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_350_ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_2__A1 net18 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_11.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_3_X cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_12_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_4.ccff_tail net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_0__A0 sb_8__8_.mux_left_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__257
+ VGND VGND VPWR VPWR net257 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__257/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l2_in_3_ net196 sb_8__8_.mux_bottom_track_59.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_92_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mem_left_track_25.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net72 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_26_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_1_ sb_8__8_.mux_bottom_track_11.out
+ net49 cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
X_333_ sb_8__8_.mux_bottom_track_29.out VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_2
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_5.mux_l2_in_1__307 VGND VGND VPWR VPWR net307 sb_8__8_.mux_left_track_5.mux_l2_in_1__307/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_51_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_4__A1 net30 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_0__A0 sb_8__8_.mux_left_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput101 net101 VGND VGND VPWR VPWR chanx_left_out[27] sky130_fd_sc_hd__buf_12
Xoutput134 net134 VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_12
Xoutput123 net123 VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_12
Xoutput112 net112 VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_12
Xoutput156 net156 VGND VGND VPWR VPWR gfpga_pad_io_soc_out_0[2] sky130_fd_sc_hd__buf_12
Xoutput145 net145 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[3] sky130_fd_sc_hd__buf_12
Xoutput167 net167 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_0_ sky130_fd_sc_hd__buf_12
XFILLER_87_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l2_in_3__196 VGND VGND VPWR VPWR net196
+ cby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l2_in_3__196/LO sky130_fd_sc_hd__conb_1
XFILLER_28_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_33.out sky130_fd_sc_hd__clkbuf_2
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_1_ net6 cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net214 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__mux2_8
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_316_ sb_8__8_.mux_left_track_3.out VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput36 chany_bottom_in[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput14 chanx_left_in[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_2
Xinput25 chanx_left_in[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput69 gfpga_pad_io_soc_in_0[2] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput58 chany_bottom_in[5] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_2
Xinput47 chany_bottom_in[22] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_ VGND VGND VPWR
+ VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_1_ sb_8__8_.mux_bottom_track_11.out
+ net49 cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_bottom_track_45.mux_l1_in_1__A1 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_31_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l2_in_3__198 VGND VGND VPWR VPWR net198
+ cby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l2_in_3__198/LO sky130_fd_sc_hd__conb_1
XFILLER_28_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_3__A1 sb_8__8_.mux_left_track_57.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_input52_A chany_bottom_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__8_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net72
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_bottom_track_11.mux_l1_in_1__A0 net163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_4__A0 sb_8__8_.mux_left_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_30_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__8_.mux_left_track_11.mux_l3_in_0_ sb_8__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X sb_8__8_.mem_left_track_11.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_left_track_53.mux_l1_in_0_ net167 net57 sb_8__8_.mem_left_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_0__A0 sb_8__8_.mux_left_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_27.out sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_45_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_45_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_92_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_2_ sb_8__8_.mux_left_track_23.out net12
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_left_track_1.mux_l2_in_0_ sb_8__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mem_bottom_track_23.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__235
+ VGND VGND VPWR VPWR net235 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__235/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_79_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__8_.mux_left_track_53.mux_l1_in_0__A1 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_94_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_1_ sb_8__8_.mux_left_track_7.out net21
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_39_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_bottom_track_9.mux_l1_in_0_ net164 left_width_0_height_0_subtile_1__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_9.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l2_in_3_ net207 sb_8__8_.mux_bottom_track_57.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_11_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_7.ccff_tail net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_13_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l1_in_1_ sb_8__8_.mux_bottom_track_9.out
+ net50 cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_2__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_23_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net241 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_left_track_13.mux_l1_in_1__287 VGND VGND VPWR VPWR net287 sb_8__8_.mux_left_track_13.mux_l1_in_1__287/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_11.mux_l2_in_1_ net286 net174 sb_8__8_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input15_A chanx_left_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_1.mux_l1_in_1_ net169 bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_8__8_.mem_left_track_1.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net178
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_60_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_60_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input7_A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_1_ sb_8__8_.mux_left_track_7.out net21
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.ccff_tail net71 VGND
+ VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_11.mux_l1_in_0__A1 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net212 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l1_in_4_ sb_8__8_.mux_bottom_track_45.out
+ net60 cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_1_prog_clk sb_8__8_.mem_left_track_45.mem_out\[0\]
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_45.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net73 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net75 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_68_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_82_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_0__A1 net22 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_18_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_4__A0 net31 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_37_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l2_in_2_ net33 net31 cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l2_in_3__203 VGND VGND VPWR VPWR net203
+ cby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l2_in_3__203/LO sky130_fd_sc_hd__conb_1
XFILLER_54_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_26_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l1_in_1__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_0_ sb_8__8_.mux_bottom_track_5.out
+ net52 cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
X_332_ sb_8__8_.mux_bottom_track_31.out VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output169_A net169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_9_X cby_8__8_.cby_8__8_.mem_right_ipin_6.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_55.mux_l2_in_0_ net280 sb_8__8_.mux_bottom_track_55.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_bottom_track_55.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_55.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_0__A1 net24 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput102 net102 VGND VGND VPWR VPWR chanx_left_out[28] sky130_fd_sc_hd__buf_12
Xoutput124 net124 VGND VGND VPWR VPWR chany_bottom_out[20] sky130_fd_sc_hd__buf_12
Xoutput113 net113 VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_12
Xoutput146 net146 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir_0[0] sky130_fd_sc_hd__buf_12
Xoutput157 net157 VGND VGND VPWR VPWR gfpga_pad_io_soc_out_0[3] sky130_fd_sc_hd__buf_12
Xoutput168 net168 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_1_ sky130_fd_sc_hd__buf_12
Xoutput135 net135 VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_12
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_17_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mem_left_track_23.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net72 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__221
+ VGND VGND VPWR VPWR net221 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__221/LO
+ sky130_fd_sc_hd__conb_1
X_315_ sb_8__8_.mux_left_track_5.out VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_56_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput26 chanx_left_in[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_2
Xinput37 chany_bottom_in[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_2
Xinput15 chanx_left_in[20] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput48 chany_bottom_in[23] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_2
Xinput59 chany_bottom_in[6] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_0_ sb_8__8_.mux_bottom_track_5.out
+ net52 cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net221 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__247
+ VGND VGND VPWR VPWR net247 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__247/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_24_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net243 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__mux2_4
XFILLER_24_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_58_prog_clk
+ sb_8__8_.mem_bottom_track_53.mem_out\[0\] net175 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_53.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__231
+ VGND VGND VPWR VPWR net231 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__231/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_55.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_55.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_55.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_2__A0 net14 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_78_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input45_A chany_bottom_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__8_.mux_bottom_track_11.mux_l1_in_1__A1 net160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__8_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_4__A1 net30 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net178
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_31_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_ VGND VGND
+ VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_42_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_0__A1 net24 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_7__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_7__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_14_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_14_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_84_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_1_ sb_8__8_.mux_left_track_11.out net19
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_32_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_0_ sb_8__8_.mux_left_track_1.out net24
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_45_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net176 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_39_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_bottom_track_49.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_49.out sky130_fd_sc_hd__buf_4
XFILLER_26_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__8_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l2_in_2_ net44 cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l1_in_0_ sb_8__8_.mux_bottom_track_3.out
+ net53 cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_3__A1 sb_8__8_.mux_left_track_57.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_11.mux_l2_in_0_ sb_8__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_76_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_49.mux_l1_in_0__A0 net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_left_track_1.mux_l1_in_0_ bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ net33 sb_8__8_.mem_left_track_1.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_7_prog_clk sb_8__8_.mem_left_track_13.mem_out\[0\]
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_31_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_0_ sb_8__8_.mux_left_track_1.out net24
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mem_bottom_track_27.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_1__S cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_2_prog_clk sb_8__8_.mem_left_track_43.ccff_tail
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_45.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l1_in_3_ sb_8__8_.mux_bottom_track_33.out
+ net37 cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_2__A1 net48 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__216
+ VGND VGND VPWR VPWR net216 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__216/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_35_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_11.mux_l1_in_1_ net171 net168 sb_8__8_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_3.out sky130_fd_sc_hd__buf_4
XFILLER_73_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_37_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l2_in_1_ net62 cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_26_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_331_ sb_8__8_.mux_bottom_track_33.out VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_46_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input75_A test_enable VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_39_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_39_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput103 net103 VGND VGND VPWR VPWR chanx_left_out[29] sky130_fd_sc_hd__buf_12
Xoutput125 net125 VGND VGND VPWR VPWR chany_bottom_out[21] sky130_fd_sc_hd__buf_12
Xoutput114 net114 VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_12
Xoutput147 net147 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir_0[1] sky130_fd_sc_hd__buf_12
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput158 net158 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_10_
+ sky130_fd_sc_hd__buf_12
Xoutput136 net136 VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_12
Xoutput169 net169 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_2_ sky130_fd_sc_hd__buf_12
XFILLER_87_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l1_in_4__A1 net60 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_ net76 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_6_prog_clk sb_8__8_.mem_bottom_track_21.mem_out\[0\]
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_21.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_11_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_2_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_314_ sb_8__8_.mux_left_track_7.out VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
XFILLER_42_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput27 chanx_left_in[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_2
Xinput16 chanx_left_in[21] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_2
Xclkbuf_3_6__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_6__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xinput38 chany_bottom_in[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_2
Xinput49 chany_bottom_in[24] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_2
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_3__323 VGND VGND VPWR VPWR net323 cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_3__323/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l1_in_2_ sb_8__8_.mux_bottom_track_23.out
+ net42 cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_3_ net316 sb_8__8_.mux_left_track_51.out
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_53_prog_clk
+ sb_8__8_.mem_bottom_track_51.ccff_tail net175 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_53.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_55.mux_l1_in_0_ net14 net161 sb_8__8_.mem_bottom_track_55.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_55.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_input38_A chany_bottom_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_30_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_ VGND VGND
+ VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_63_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_47.mux_l1_in_1__A1 net172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_54_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_54_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_92_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_0_ sb_8__8_.mux_left_track_5.out net22
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mux_bottom_track_57.mux_l1_in_0__A0 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_19_prog_clk cbx_8__8_.cbx_1__8_.ccff_tail net177 VGND VGND VPWR VPWR
+ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_24_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_50_prog_clk
+ cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[2\] net176 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_32_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_44_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net176 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_load_slew178_A net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_4__S cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_39_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_4_ sb_8__8_.mux_left_track_39.out
+ net4 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_1__A0 sb_8__8_.mux_left_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l2_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_2_X cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_8__8_.cby_8__8_.mux_left_ipin_3.out cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_21_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_49.mux_l1_in_0__A1 left_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mem_bottom_track_59.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk sb_8__8_.mem_bottom_track_59.mem_out\[0\]
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_59.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_39_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_22_prog_clk sb_8__8_.mem_left_track_11.ccff_tail
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_82_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_1__A0 sb_8__8_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_9_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_32_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_38_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__8_.mux_bottom_track_15.mux_l1_in_0__A0 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_36_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input20_A chanx_left_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net230 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l1_in_2_ sb_8__8_.mux_bottom_track_21.out
+ net43 cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_42_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_1__D cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l2_in_1__A0 net40 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__317__A sb_8__8_.mux_left_track_1.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_2__A0 sb_8__8_.mux_bottom_track_17.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_11.mux_l1_in_0_ bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ net50 sb_8__8_.mem_left_track_11.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_9_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_9_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_58_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__8_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_26_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_330_ sb_8__8_.mux_bottom_track_35.out VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_5__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_5__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_8__8_.mux_left_track_23.mux_l2_in_0_ net292 sb_8__8_.mux_left_track_23.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_23.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_23.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input68_A gfpga_pad_io_soc_in_0[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_92_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_1__A0 sb_8__8_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput115 net115 VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_12
Xoutput104 net104 VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_12
Xoutput148 net148 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir_0[2] sky130_fd_sc_hd__buf_12
Xoutput126 net126 VGND VGND VPWR VPWR chany_bottom_out[22] sky130_fd_sc_hd__buf_12
Xoutput137 net137 VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_12
Xoutput159 net159 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_11_
+ sky130_fd_sc_hd__buf_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_2__A0 net26 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk sb_8__8_.mem_left_track_19.mem_out\[0\]
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_19.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_51_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_52_prog_clk
+ sb_8__8_.mem_bottom_track_19.ccff_tail net176 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_21.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_4__A0 net4 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_19_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_313_ sb_8__8_.mux_left_track_9.out VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput28 chanx_left_in[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_4
Xinput17 chanx_left_in[22] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput39 chany_bottom_in[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_54_prog_clk
+ cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[2\] net175 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_3.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_output174_A net174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_2__A0 net28 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l1_in_1_ sb_8__8_.mux_bottom_track_11.out
+ net49 cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_bottom_track_3.mux_l1_in_0__A0 net164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_2_ net27 cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_30_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__220
+ VGND VGND VPWR VPWR net220 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__220/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_42_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net225 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__mux2_4
XFILLER_25_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_23_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_23_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_57.mux_l1_in_0__A1 net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net257 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_50_prog_clk
+ cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[1\] net176 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_13.mux_l1_in_1__A1 net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input50_A chany_bottom_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_2__A0 net31 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mem_bottom_track_27.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_35_prog_clk
+ sb_8__8_.mem_bottom_track_27.mem_out\[0\] net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_27.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_39_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_3_ sb_8__8_.mux_left_track_27.out
+ net10 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__8_.mux_bottom_track_23.mux_l1_in_0__A0 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_38_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_13.mux_l2_in_0_ net261 sb_8__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_bottom_track_13.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l1_in_2__A1 net47 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l2_in_2__A0 net58 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_59.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_0_prog_clk sb_8__8_.mem_bottom_track_57.ccff_tail
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_59.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_79_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_1__A1 net19 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__8_.mux_bottom_track_15.mux_l1_in_0__A1 left_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_3__A1 net9 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xclkbuf_3_4__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_4__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_14_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input13_A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_8__8_.cby_8__8_.mux_left_ipin_1.out cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l1_in_1_ sb_8__8_.mux_bottom_track_9.out
+ net50 cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_42_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_3__A1 net11 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_61_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[2\] net175 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__333__A sb_8__8_.mux_bottom_track_29.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input5_A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_26_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_1__A1 net19 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l2_in_3_ net198 net30 cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput116 net116 VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_12
Xoutput105 net105 VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_12
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput149 net149 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir_0[3] sky130_fd_sc_hd__buf_12
Xoutput138 net138 VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_12
Xoutput127 net127 VGND VGND VPWR VPWR chany_bottom_out[23] sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_48_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_48_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_95_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__328__A net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_5_prog_clk sb_8__8_.mem_left_track_17.ccff_tail
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_19.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_51_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_4__A1 net35 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_52_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_312_ sb_8__8_.mux_left_track_11.out VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput18 chanx_left_in[23] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_2
Xinput29 chanx_left_in[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__8_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_58_prog_clk
+ cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[1\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_output167_A net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_3__318 VGND VGND VPWR VPWR net318
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_3__318/LO sky130_fd_sc_hd__conb_1
XFILLER_18_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l1_in_0_ sb_8__8_.mux_bottom_track_5.out
+ net52 cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_19.mux_l2_in_0__264 VGND VGND VPWR VPWR net264 sb_8__8_.mux_bottom_track_19.mux_l2_in_0__264/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l2_in_3_ net194 sb_8__8_.mux_bottom_track_55.out
+ cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_left_track_23.mux_l1_in_0_ net168 net43 sb_8__8_.mem_left_track_23.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_23.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_bottom_track_3.mux_l1_in_0__A1 left_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_1_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_2_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_1__A0 sb_8__8_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_30_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mux_left_track_35.mux_l2_in_0_ sb_8__8_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_35.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_63_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_bottom_track_31.mux_l1_in_0__A0 net161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_6_prog_clk sb_8__8_.mem_left_track_31.mem_out\[0\]
+ net176 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_31.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_65_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_16_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_3__A1 net41 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_36_prog_clk sb_8__8_.mem_bottom_track_3.mem_out\[1\]
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_55_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_11.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_49_prog_clk
+ cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\] net175 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input43_A chany_bottom_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l2_in_3__194 VGND VGND VPWR VPWR net194 cby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l2_in_3__194/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__8_.mem_bottom_track_27.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_35_prog_clk
+ sb_8__8_.mem_bottom_track_25.ccff_tail net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_27.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_4_ net30 net61 cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_39_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.out cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_2_ sb_8__8_.mux_left_track_15.out
+ net17 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__8_.mux_bottom_track_23.mux_l1_in_0__A1 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net73 grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_77_.in net75 VGND
+ VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_38_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_3_ net323 sb_8__8_.mux_left_track_57.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_3__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_3__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_21_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_60_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[2\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_4.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_79_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__213
+ VGND VGND VPWR VPWR net213 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__213/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__8_.mux_left_track_59.mux_l1_in_0__A0 net170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_35.mux_l1_in_1_ net299 net174 sb_8__8_.mem_left_track_35.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_0_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_3__188 VGND VGND VPWR VPWR net188 cbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_3__188/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_clk0 clk0 VGND VGND VPWR VPWR clknet_0_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_12_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_9_X cby_8__8_.cby_8__8_.mem_left_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_left_track_3.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_43_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_bottom_track_5.mux_l3_in_0_ sb_8__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X sb_8__8_.mem_bottom_track_5.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_47_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_25.mux_l2_in_0__293 VGND VGND VPWR VPWR net293 sb_8__8_.mux_left_track_25.mux_l2_in_0__293/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_86_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_bottom_track_1.mux_l2_in_1__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__217
+ VGND VGND VPWR VPWR net217 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__217/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_33_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_3_ net184 sb_8__8_.mux_left_track_45.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net248 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l1_in_0_ sb_8__8_.mux_bottom_track_3.out
+ net53 cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_42_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_bottom_track_13.mux_l1_in_0_ net17 left_width_0_height_0_subtile_0__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_13.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_4_ sb_8__8_.mux_left_track_45.out net30
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_60_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[1\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__8_.mux_left_track_17.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_bottom_track_25.mux_l2_in_0_ net267 sb_8__8_.mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_bottom_track_25.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_26_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_5.mux_l2_in_1_ net277 net21 sb_8__8_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_1_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_23.mux_l2_in_0__266 VGND VGND VPWR VPWR net266 sb_8__8_.mux_bottom_track_23.mux_l2_in_0__266/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_49_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_17_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_64_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_9_X cbx_8__8_.cbx_1__8_.mem_top_ipin_12.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net178
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l2_in_2_ net61 sb_8__8_.mux_bottom_track_31.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput106 net106 VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_12
Xoutput128 net128 VGND VGND VPWR VPWR chany_bottom_out[24] sky130_fd_sc_hd__buf_12
Xoutput139 net139 VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_12
Xoutput117 net117 VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_12
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_31.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_31.out sky130_fd_sc_hd__clkbuf_2
XFILLER_68_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_17_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_17_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_55_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__344__A sb_8__8_.mux_bottom_track_7.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net72
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_311_ sb_8__8_.mux_left_track_13.out VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput19 chanx_left_in[24] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_57_prog_clk
+ cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[0\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_input73_A reset VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net246 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_45_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l2_in_2_ net55 cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__339__A sb_8__8_.mux_bottom_track_17.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_59_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[2\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_7.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_1__A1 net19 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_30_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_left_track_25.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_25.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_25.out sky130_fd_sc_hd__clkbuf_2
XFILLER_34_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__8_.mux_bottom_track_31.mux_l1_in_0__A1 left_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_6_prog_clk sb_8__8_.mem_left_track_29.ccff_tail
+ net176 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_31.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_84_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_35.mux_l1_in_1__273 VGND VGND VPWR VPWR net273 sb_8__8_.mux_bottom_track_35.mux_l1_in_1__273/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_25_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_2__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_2__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_1_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_36_prog_clk sb_8__8_.mem_bottom_track_3.mem_out\[0\]
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_32_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_32_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_4__A0 sb_8__8_.mux_left_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_3_ net189 sb_8__8_.mux_left_track_49.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__8_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_60_prog_clk
+ net1 net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net178
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input36_A chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__8_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_3_ sb_8__8_.mux_bottom_track_31.out
+ net38 cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_1_ sb_8__8_.mux_left_track_9.out
+ net20 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l2_in_2__A0 net58 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_33_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_2_ net14 cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__229
+ VGND VGND VPWR VPWR net229 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__229/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__8_.mux_left_track_19.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_19.out sky130_fd_sc_hd__clkbuf_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_60_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[1\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_left_track_35.mux_l1_in_0_ bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ net37 sb_8__8_.mem_left_track_35.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_left_track_59.mux_l1_in_0__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_9.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_9.out sky130_fd_sc_hd__buf_4
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l2_in_3__202 VGND VGND VPWR VPWR net202
+ cby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l2_in_3__202/LO sky130_fd_sc_hd__conb_1
XFILLER_56_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_2__A0 sb_8__8_.mux_left_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_left_track_47.mux_l2_in_0_ sb_8__8_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_47.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_left_track_3.mux_l1_in_0__A1 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_43_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net178
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_load_slew176_A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_25.mux_l1_in_0__A0 net169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_4_ sb_8__8_.mux_left_track_37.out net5
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_3_X cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_1_prog_clk sb_8__8_.mem_left_track_37.mem_out\[0\]
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_37.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_26_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__347__A sb_8__8_.mux_bottom_track_1.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_34_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.out cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_39_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_2_ net30 sb_8__8_.mux_left_track_27.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_37_prog_clk sb_8__8_.mem_bottom_track_9.mem_out\[1\]
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_43_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_3_ sb_8__8_.mux_left_track_33.out net7
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_3__182 VGND VGND VPWR VPWR net182 cbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_3__182/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_9_X cbx_8__8_.cbx_1__8_.mem_top_ipin_8.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_59_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[0\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_8__8_.mux_bottom_track_5.mux_l1_in_1__A0 net163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_17.mux_l1_in_0__A1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_1__A0 net4 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_54_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_left_track_47.mux_l1_in_1_ net305 net172 sb_8__8_.mem_left_track_47.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_10_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_5.mux_l2_in_0_ sb_8__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_17_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l2_in_1_ net38 cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__239
+ VGND VGND VPWR VPWR net239 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__239/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_40_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput107 net107 VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_12
Xoutput129 net129 VGND VGND VPWR VPWR chany_bottom_out[25] sky130_fd_sc_hd__buf_12
Xoutput118 net118 VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_12
XANTENNA_clkbuf_leaf_35_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_57_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_57_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l1_in_1__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_7__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_79_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_310_ sb_8__8_.mux_left_track_15.out VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_61_prog_clk
+ cby_8__8_.cby_8__8_.mem_left_ipin_2.ccff_tail net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_sb_8__8_.mux_left_track_1.mux_l2_in_1__A1 net172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input66_A gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_53_prog_clk
+ sb_8__8_.mem_bottom_track_45.mem_out\[0\] net175 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_45.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_1__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_1__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_8__8_.mux_bottom_track_25.mux_l1_in_0_ net10 net158 sb_8__8_.mem_bottom_track_25.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_87_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l2_in_1_ cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_2_X cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.out sky130_fd_sc_hd__clkbuf_1
XFILLER_24_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_53.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_53.out sky130_fd_sc_hd__clkbuf_2
Xsb_8__8_.mux_bottom_track_5.mux_l1_in_1_ net163 net160 sb_8__8_.mem_bottom_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_24_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__8_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_33_prog_clk cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.ccff_tail
+ net178 VGND VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_59_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[1\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l1_in_2_ sb_8__8_.mux_bottom_track_13.out
+ net48 cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_29_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_2_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_2_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output172_A net172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_21_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[2\] net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_12.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_36_prog_clk sb_8__8_.mem_bottom_track_1.ccff_tail
+ net177 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_4__A1 net30 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l2_in_3__208 VGND VGND VPWR VPWR net208
+ cby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l2_in_3__208/LO sky130_fd_sc_hd__conb_1
XFILLER_29_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_2_ net28 cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input29_A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net73 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net75 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_77_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_47_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__8_.mux_left_track_33.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_28_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_2_ sb_8__8_.mux_bottom_track_19.out
+ net45 cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_left_track_47.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_47.out sky130_fd_sc_hd__clkbuf_1
XFILLER_7_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_0_ sb_8__8_.mux_left_track_3.out
+ net23 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_4__A1 net32 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_2_X cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_32_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_60_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[0\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_88_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__251
+ VGND VGND VPWR VPWR net251 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__251/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_44_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net175
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_2__A1 net13 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_43_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_3__A1 sb_8__8_.mux_left_track_57.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_3_ sb_8__8_.mux_left_track_25.out net11
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew175 net176 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__buf_12
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_8_prog_clk sb_8__8_.mem_left_track_1.mem_out\[1\]
+ net176 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_0_prog_clk sb_8__8_.mem_left_track_35.ccff_tail
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_37.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_81_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_0__A0 sb_8__8_.mux_left_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net73 net74 net75 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_5_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_1_ net10 cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_37_prog_clk sb_8__8_.mem_bottom_track_9.mem_out\[0\]
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_9.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_44_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_42_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net175
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_2_ sb_8__8_.mux_left_track_21.out net13
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_23.out sky130_fd_sc_hd__clkbuf_2
XFILLER_95_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_0__A0 sb_8__8_.mux_left_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_57_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_0.ccff_tail net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mux_bottom_track_5.mux_l1_in_1__A1 net160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_38_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_54_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mux_left_track_47.mux_l1_in_0_ bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ net60 sb_8__8_.mem_left_track_47.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input11_A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_34_prog_clk
+ sb_8__8_.mem_bottom_track_13.mem_out\[0\] net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_13.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_0__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_0__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_32_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_59.mux_l2_in_0_ sb_8__8_.mux_left_track_59.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_59.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.ccff_head
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_59.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput119 net119 VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_12
XFILLER_31_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput108 net108 VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_12
XFILLER_95_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput90 net90 VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_12
XFILLER_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_ VGND
+ VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_48_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_left_track_7.mux_l3_in_0_ sb_8__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X sb_8__8_.mem_left_track_7.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_26_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_26_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_2_ sb_8__8_.mux_left_track_15.out net17
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_20_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[2\] net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input3_A chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_17.out sky130_fd_sc_hd__buf_4
XFILLER_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_45_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net72 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input59_A chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_53_prog_clk
+ sb_8__8_.mem_bottom_track_35.ccff_tail net175 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_45.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_3__321 VGND VGND VPWR VPWR net321 cbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_3__321/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_0__A0 sb_8__8_.mux_left_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_56_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[2\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_12.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mem_left_track_59.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_1__A0 net10 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_28_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mux_bottom_track_5.mux_l1_in_0_ net165 left_width_0_height_0_subtile_2__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_5.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l2_in_3_ net203 sb_8__8_.mux_bottom_track_49.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_57_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[0\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_78_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l1_in_1_ sb_8__8_.mux_bottom_track_7.out
+ net51 cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l2_in_2__A0 net44 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mux_left_track_41.mux_l1_in_0__A0 net169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_59.mux_l1_in_1_ net312 net174 sb_8__8_.mem_left_track_59.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_59.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_47_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_29_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mux_left_track_5.mux_l1_in_1__A0 net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output165_A net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_left_track_7.mux_l2_in_1_ net313 net172 sb_8__8_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_2_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__246
+ VGND VGND VPWR VPWR net246 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__246/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_80_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_21_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[1\] net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_2_X cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_41_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_41_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_24_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__8_.mux_left_track_33.mux_l1_in_0__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net64 cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_2__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_74_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_28_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_1_ sb_8__8_.mux_bottom_track_7.out
+ net51 cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_8__8_.ccff_tail net71 VGND VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
XFILLER_65_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_4_ net4 net35 cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net227 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l1_in_2__A0 sb_8__8_.mux_bottom_track_17.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_55_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_3.ccff_tail net175 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mux_bottom_track_49.mux_l2_in_0_ sb_8__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_49.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_25_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_15_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input41_A chany_bottom_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_43_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__256
+ VGND VGND VPWR VPWR net256 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__256/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_54_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cby_8__8_.cby_8__8_.mem_right_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mux_bottom_track_51.mux_l2_in_0_ sb_8__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_51.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_2_ sb_8__8_.mux_left_track_13.out net18
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net177 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mem_bottom_track_57.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew176 net72 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__buf_12
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_6_prog_clk sb_8__8_.mem_left_track_1.mem_out\[0\]
+ net176 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_81_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_61_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_51.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_51.out sky130_fd_sc_hd__clkbuf_2
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_36_prog_clk sb_8__8_.mem_bottom_track_7.ccff_tail
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_9.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_57_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_11_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[2\] net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_1_ sb_8__8_.mux_left_track_9.out net20
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_42_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_0__A1 net23 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_51_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[2\] net176 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l2_in_3_ net208 sb_8__8_.mux_bottom_track_53.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_49.mux_l1_in_1_ net276 net27 sb_8__8_.mem_bottom_track_49.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net68 cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR left_width_0_height_0_subtile_2__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_38_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_66_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_2__A1 net17 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_2_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[2\] net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_66_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__8_.mux_bottom_track_51.mux_l1_in_1_ net278 net26 sb_8__8_.mem_bottom_track_51.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_34_prog_clk
+ sb_8__8_.mem_bottom_track_11.ccff_tail net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_13.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l2_in_1__A0 net34 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_bottom_track_33.mux_l1_in_1__A1 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net178
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_3__A1 net37 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
Xoutput109 net109 VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_12
Xoutput91 net91 VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_12
Xoutput80 net80 VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_12
XFILLER_48_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_45.out sky130_fd_sc_hd__clkbuf_2
XFILLER_36_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_1_ sb_8__8_.mux_left_track_9.out net20
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_21_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[1\] net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_1__A1 net50 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_bottom_track_49.mux_l1_in_1__276 VGND VGND VPWR VPWR net276 sb_8__8_.mux_bottom_track_49.mux_l1_in_1__276/LO
+ sky130_fd_sc_hd__conb_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_21_prog_clk sb_8__8_.mem_left_track_7.mem_out\[1\]
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_7.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_45_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net72 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_0__A1 net23 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_48_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[1\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_ VGND VGND
+ VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_41_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_left_track_49.mux_l1_in_1__306 VGND VGND VPWR VPWR net306 sb_8__8_.mux_left_track_49.mux_l1_in_1__306/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_42_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_299_ sb_8__8_.mux_left_track_37.out VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l2_in_2_ net58 cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_56_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_6.ccff_tail net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l1_in_0_ sb_8__8_.mux_bottom_track_1.out
+ net54 cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mux_left_track_41.mux_l1_in_0__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_59.mux_l1_in_0_ net170 net44 sb_8__8_.mem_left_track_59.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_59.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_47_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_32_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__8_.mux_left_track_5.mux_l1_in_1__A1 net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_7.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input71_A isol_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_left_track_7.mux_l2_in_0_ sb_8__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_output158_A net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_9.mux_l1_in_0__A0 net164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_21_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\] net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_8__8_.mem_left_track_57.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net72 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_52_prog_clk
+ sb_8__8_.mem_bottom_track_19.mem_out\[0\] net176 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_19.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_2__A1 net16 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_23_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_left_track_55.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_60_prog_clk sb_8__8_.mem_left_track_55.mem_out\[0\]
+ net72 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_55.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_71_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net178
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_10_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_10_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_58_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_0__A0 sb_8__8_.mux_left_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_44_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_27_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_0_ sb_8__8_.mux_bottom_track_1.out
+ net54 cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_3_ sb_8__8_.mux_bottom_track_25.out
+ net41 cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net244 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__mux2_4
XFILLER_88_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_25_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_52_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_7.mux_l1_in_1_ net169 bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_8__8_.mem_left_track_7.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mem_left_track_43.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net72 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_9_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[2\] net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_4.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__8_.mux_bottom_track_29.mux_l1_in_0__A0 net160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_43_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input34_A chany_bottom_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_0_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_1_ sb_8__8_.mux_left_track_7.out net21
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l1_in_2__A1 net40 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xload_slew177 net178 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__buf_12
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_5_prog_clk sb_8__8_.mem_bottom_track_59.ccff_tail
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_93_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net175
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.ccff_tail net71 VGND
+ VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_42_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_10_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[1\] net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_0_ sb_8__8_.mux_left_track_3.out net23
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_41_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net177 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mem_bottom_track_55.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_53_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[1\] net175 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l2_in_2_ net56 sb_8__8_.mux_bottom_track_35.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_49.mux_l1_in_0_ net158 left_width_0_height_0_subtile_2__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_49.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_2_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[1\] net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__249
+ VGND VGND VPWR VPWR net249 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__249/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_51.mux_l1_in_0_ net159 left_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_51.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_ VGND VGND VPWR VPWR
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
Xoutput81 net81 VGND VGND VPWR VPWR ccff_tail_0 sky130_fd_sc_hd__buf_12
Xoutput92 net92 VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_12
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l2_in_3__A1 net30 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_0_ sb_8__8_.mux_left_track_3.out net23
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_21_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[0\] net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_8__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net177 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_35_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_35_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_22_prog_clk sb_8__8_.mem_left_track_7.mem_out\[0\]
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_10_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_44_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net72 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_38_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__295__A sb_8__8_.mux_left_track_45.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_47_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[0\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_3__316 VGND VGND VPWR VPWR net316
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_3__316/LO sky130_fd_sc_hd__conb_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_ VGND VGND
+ VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
X_298_ sb_8__8_.mux_left_track_39.out VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_18_prog_clk cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.ccff_tail
+ net177 VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dfrtp_2
Xsb_8__8_.mem_left_track_23.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_61_prog_clk sb_8__8_.mem_left_track_23.mem_out\[0\]
+ net72 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_23.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l2_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net211 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_32_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_34_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net216 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input64_A gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_9.mux_l1_in_0__A1 left_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_11_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[2\] net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_7.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_14_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_11.ccff_tail net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xsb_8__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_7_prog_clk sb_8__8_.mem_bottom_track_17.ccff_tail
+ net176 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_19.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_23_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_1__A0 sb_8__8_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_left_track_55.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_60_prog_clk sb_8__8_.mem_left_track_53.ccff_tail
+ net72 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_55.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_83_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_2__A0 sb_8__8_.mux_bottom_track_17.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_50_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_50_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_59_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l2_in_3__192 VGND VGND VPWR VPWR net192 cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l2_in_3__192/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_29_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output170_A net170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_2_ sb_8__8_.mux_bottom_track_13.out
+ net48 cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_17.mux_l2_in_0_ sb_8__8_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_17.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_9_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_3_ net317 sb_8__8_.mux_left_track_53.out
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_3_X cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_3__186 VGND VGND VPWR VPWR net186 cbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_3__186/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_25_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_25_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_64_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_7.mux_l1_in_0_ bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ net52 sb_8__8_.mem_left_track_7.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_9_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[1\] net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__8_.mux_bottom_track_29.mux_l1_in_0__A1 left_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_43_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input27_A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_4__A0 net4 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk
+ sb_8__8_.mem_bottom_track_31.mem_out\[0\] net176 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_31.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_2__S cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_0_ sb_8__8_.mux_left_track_1.out net24
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew178 net179 VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_16
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_left_track_9.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__8_.mem_left_track_41.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net72 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_10_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\] net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_8__8_.mux_bottom_track_7.mux_l2_in_1__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_17.mux_l1_in_1_ net289 net173 sb_8__8_.mem_left_track_17.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_29_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_77_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_4_ sb_8__8_.mux_left_track_41.out
+ net32 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_2__A0 net28 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_49_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[0\] net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1 sb_8__8_.mux_bottom_track_23.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l2_in_1_ net36 cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_45_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net176 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_4__A0 net32 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_1_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[0\] net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_32_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_left_track_19.mux_l2_in_0__290 VGND VGND VPWR VPWR net290 sb_8__8_.mux_left_track_19.mux_l2_in_0__290/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_77_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_4__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_ VGND VGND VPWR VPWR
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_5_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_5_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_2__A0 net27 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xoutput82 net82 VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_12
Xoutput93 net93 VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_12
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_0_clk0_A clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_17_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_14.ccff_tail net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_59_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_0__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_22_prog_clk sb_8__8_.mem_left_track_5.ccff_tail
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_10_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_44_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net72 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_left_track_35.mux_l1_in_1__A1 net174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_37_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l1_in_2_ sb_8__8_.mux_bottom_track_23.out
+ net42 cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net73 grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_86_.in net75 VGND
+ VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_9.out sky130_fd_sc_hd__buf_4
XFILLER_60_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_47_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_11.ccff_tail net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_297_ sb_8__8_.mux_left_track_41.out VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_45_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net176 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_17.mux_l2_in_0__263 VGND VGND VPWR VPWR net263 sb_8__8_.mux_bottom_track_17.mux_l2_in_0__263/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__8_.mux_bottom_track_45.mux_l1_in_0__A0 net164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net177 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_23.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_0_prog_clk sb_8__8_.mem_left_track_21.ccff_tail
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_23.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_51_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net178
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input1_A ccff_head_0_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.out sky130_fd_sc_hd__clkbuf_1
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_2__A0 net14 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input57_A chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_2_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[1\] net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_349_ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_1__A1 net19 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_56_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mem_left_track_39.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_27_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l2_in_2__A0 net57 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output163_A net163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_1__A1 net21 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_1_ sb_8__8_.mux_bottom_track_7.out
+ net51 cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_2_ net26 cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_19_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l2_in_3__200 VGND VGND VPWR VPWR net200
+ cby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l2_in_3__200/LO sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_6_prog_clk sb_8__8_.mem_left_track_29.mem_out\[0\]
+ net176 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_29.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_9_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\] net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_94_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_43_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_4__A1 net35 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_52_prog_clk
+ sb_8__8_.mem_bottom_track_29.ccff_tail net176 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_31.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net226 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__mux2_4
XFILLER_7_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew179 net72 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__buf_12
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_23.mux_l2_in_0__292 VGND VGND VPWR VPWR net292 sb_8__8_.mux_left_track_23.mux_l2_in_0__292/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_3__A1 net10 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_2__A1 net45 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_29_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_29_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_left_track_9.mux_l1_in_0__A1 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_20_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.ccff_tail net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_4_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_1__A1 net21 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_17.mux_l1_in_0_ bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ net47 sb_8__8_.mem_left_track_17.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_3__180 VGND VGND VPWR VPWR net180 cbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_3__180/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_29_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_3_ sb_8__8_.mux_left_track_29.out
+ net9 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_47_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_14.ccff_tail net72 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_31_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_2 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_left_track_29.mux_l2_in_0_ sb_8__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_29.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_14_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_45_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net176 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_4__A1 net34 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_6_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_0.ccff_tail net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_38_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net178
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_53_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_21.mux_l2_in_0__265 VGND VGND VPWR VPWR net265 sb_8__8_.mux_bottom_track_21.mux_l2_in_0__265/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__238
+ VGND VGND VPWR VPWR net238 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__238/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__8_.mux_left_track_31.mux_l2_in_0_ sb_8__8_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_31.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_40_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput94 net94 VGND VGND VPWR VPWR chanx_left_out[20] sky130_fd_sc_hd__buf_12
Xoutput83 net83 VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_12
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_53.mux_l1_in_0__A0 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_3__A1 net7 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_63_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_44_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_44_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_43_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net72 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l1_in_1_ sb_8__8_.mux_bottom_track_11.out
+ net49 cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_296_ sb_8__8_.mux_left_track_43.out VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_1
XFILLER_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_29.mux_l1_in_1_ net295 net171 sb_8__8_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_45_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net176 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__8_.mux_bottom_track_45.mux_l1_in_0__A1 left_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_7.mux_l2_in_1__A1 net172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net229 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_31.mux_l1_in_1_ net297 net172 sb_8__8_.mem_left_track_31.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l2_in_3_ net199 sb_8__8_.mux_bottom_track_57.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_3_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[0\] net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_8__8_.mux_bottom_track_11.mux_l1_in_0__A0 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_348_ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_1
Xsb_8__8_.mux_bottom_track_33.mux_l1_in_1__272 VGND VGND VPWR VPWR net272 sb_8__8_.mux_bottom_track_33.mux_l1_in_1__272/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_bottom_track_1.mux_l3_in_0_ sb_8__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X sb_8__8_.mem_bottom_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l2_in_3__206 VGND VGND VPWR VPWR net206
+ cby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l2_in_3__206/LO sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net178
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_27_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l2_in_2__A1 net32 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_19.mux_l2_in_0_ net264 sb_8__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_bottom_track_19.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_0_ sb_8__8_.mux_bottom_track_1.out
+ net54 cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net252 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_1_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__8_.mux_left_track_39.mux_l1_in_0__A0 net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_bottom_track_21.mux_l2_in_0_ net265 sb_8__8_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_bottom_track_21.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l1_in_4_ sb_8__8_.mux_bottom_track_45.out
+ net60 cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_2__A0 net14 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_4_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_6_prog_clk sb_8__8_.mem_left_track_27.ccff_tail
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_29.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_20_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_3.ccff_tail net178 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_43_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_bottom_track_1.mux_l2_in_1_ net259 net23 sb_8__8_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_85_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_9_X cby_8__8_.cby_8__8_.mem_right_ipin_12.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_43_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_21.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_21.out sky130_fd_sc_hd__buf_4
XFILLER_4_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input32_A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net255 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__mux2_4
XFILLER_63_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_29_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_2_ sb_8__8_.mux_left_track_17.out
+ net16 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mem_left_track_23.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_3 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_3_ net180 sb_8__8_.mux_left_track_47.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mem_left_track_41.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_61_prog_clk sb_8__8_.mem_left_track_41.mem_out\[0\]
+ net72 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_41.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_62_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_50_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_3__A0 sb_8__8_.mux_bottom_track_29.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l1_in_0__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput84 net84 VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_12
XFILLER_95_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput95 net95 VGND VGND VPWR VPWR chanx_left_out[21] sky130_fd_sc_hd__buf_12
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mux_bottom_track_53.mux_l1_in_0__A1 net160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_15.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_15.out sky130_fd_sc_hd__clkbuf_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_5.out sky130_fd_sc_hd__buf_4
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_40_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net73 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net75 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_86_.in
+ sky130_fd_sc_hd__sdfrtp_1
XANTENNA_sb_8__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_3_ net185 sb_8__8_.mux_left_track_53.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
Xclkbuf_leaf_13_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_13_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_43_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_89_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l1_in_0_ sb_8__8_.mux_bottom_track_5.out
+ net52 cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_364_ net79 VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_1
X_295_ sb_8__8_.mux_left_track_45.out VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_1_1__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_left_track_29.mux_l1_in_0_ bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ net40 sb_8__8_.mem_left_track_29.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_53.mux_l2_in_0__279 VGND VGND VPWR VPWR net279 sb_8__8_.mux_bottom_track_53.mux_l2_in_0__279/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_31.mux_l1_in_0_ bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ net39 sb_8__8_.mem_left_track_31.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mux_left_track_53.mux_l2_in_0__309 VGND VGND VPWR VPWR net309 sb_8__8_.mux_left_track_53.mux_l2_in_0__309/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_13.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l2_in_2_ net44 cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_1__A0 net4 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_9_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_6.ccff_tail net176 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_92_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__8_.mux_bottom_track_11.mux_l1_in_0__A1 left_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mux_left_track_43.mux_l2_in_0_ net303 sb_8__8_.mux_left_track_43.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_43.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_43.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_3__A1 net7 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_73_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_347_ sb_8__8_.mux_bottom_track_1.out VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_34_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_43_.in
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net176 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l2_in_2__A0 net44 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net73 grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_32_.in net75 VGND
+ VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_5_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_47.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_4_ sb_8__8_.mux_left_track_41.out net32
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_27_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net178 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input62_A chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_9_X cbx_8__8_.cbx_1__8_.mem_top_ipin_4.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_33_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mem_bottom_track_27.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__8_.mux_left_track_39.mux_l1_in_0__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l1_in_3_ sb_8__8_.mux_bottom_track_33.out
+ net37 cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_42_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_bottom_track_1.mux_l2_in_0_ sb_8__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_85_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__233
+ VGND VGND VPWR VPWR net233 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__233/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_66_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_3_ net190 sb_8__8_.mux_left_track_57.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l1_in_1__A1 net50 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_38_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_38_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_19.mux_l1_in_0_ net13 left_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_19.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net176
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input25_A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_30_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net179 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_1_ sb_8__8_.mux_left_track_11.out
+ net19 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_4 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_2_ net29 sb_8__8_.mux_left_track_35.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_21.mux_l1_in_0_ net12 net164 sb_8__8_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__8_.mem_left_track_41.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_61_prog_clk sb_8__8_.mem_left_track_39.ccff_tail
+ net72 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_41.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_1.mux_l1_in_1_ net161 net158 sb_8__8_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_bottom_track_33.mux_l2_in_0_ sb_8__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_33.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_3__A1 net39 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_43.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_43.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_43.out sky130_fd_sc_hd__dlymetal6s2s_1
Xoutput85 net85 VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_12
Xoutput96 net96 VGND VGND VPWR VPWR chanx_left_out[22] sky130_fd_sc_hd__buf_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_26_prog_clk grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net177 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_2__A1 net10 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
.ends

