magic
tech sky130A
magscale 1 2
timestamp 1625784963
<< obsli1 >>
rect 1104 2159 21896 20689
<< obsm1 >>
rect 198 2128 22802 20868
<< metal2 >>
rect 202 22200 258 23000
rect 662 22200 718 23000
rect 1122 22200 1178 23000
rect 1582 22200 1638 23000
rect 2042 22200 2098 23000
rect 2502 22200 2558 23000
rect 2962 22200 3018 23000
rect 3422 22200 3478 23000
rect 3882 22200 3938 23000
rect 4342 22200 4398 23000
rect 4802 22200 4858 23000
rect 5262 22200 5318 23000
rect 5722 22200 5778 23000
rect 6182 22200 6238 23000
rect 6642 22200 6698 23000
rect 7102 22200 7158 23000
rect 7562 22200 7618 23000
rect 8022 22200 8078 23000
rect 8482 22200 8538 23000
rect 8942 22200 8998 23000
rect 9402 22200 9458 23000
rect 9862 22200 9918 23000
rect 10322 22200 10378 23000
rect 10782 22200 10838 23000
rect 11242 22200 11298 23000
rect 11702 22200 11758 23000
rect 12162 22200 12218 23000
rect 12622 22200 12678 23000
rect 13082 22200 13138 23000
rect 13542 22200 13598 23000
rect 14002 22200 14058 23000
rect 14462 22200 14518 23000
rect 14922 22200 14978 23000
rect 15382 22200 15438 23000
rect 15842 22200 15898 23000
rect 16302 22200 16358 23000
rect 16762 22200 16818 23000
rect 17222 22200 17278 23000
rect 17682 22200 17738 23000
rect 18142 22200 18198 23000
rect 18602 22200 18658 23000
rect 19062 22200 19118 23000
rect 19522 22200 19578 23000
rect 19982 22200 20038 23000
rect 20442 22200 20498 23000
rect 20902 22200 20958 23000
rect 21362 22200 21418 23000
rect 21822 22200 21878 23000
rect 22282 22200 22338 23000
rect 22742 22200 22798 23000
rect 11518 0 11574 800
<< obsm2 >>
rect 314 22144 606 22681
rect 774 22144 1066 22681
rect 1234 22144 1526 22681
rect 1694 22144 1986 22681
rect 2154 22144 2446 22681
rect 2614 22144 2906 22681
rect 3074 22144 3366 22681
rect 3534 22144 3826 22681
rect 3994 22144 4286 22681
rect 4454 22144 4746 22681
rect 4914 22144 5206 22681
rect 5374 22144 5666 22681
rect 5834 22144 6126 22681
rect 6294 22144 6586 22681
rect 6754 22144 7046 22681
rect 7214 22144 7506 22681
rect 7674 22144 7966 22681
rect 8134 22144 8426 22681
rect 8594 22144 8886 22681
rect 9054 22144 9346 22681
rect 9514 22144 9806 22681
rect 9974 22144 10266 22681
rect 10434 22144 10726 22681
rect 10894 22144 11186 22681
rect 11354 22144 11646 22681
rect 11814 22144 12106 22681
rect 12274 22144 12566 22681
rect 12734 22144 13026 22681
rect 13194 22144 13486 22681
rect 13654 22144 13946 22681
rect 14114 22144 14406 22681
rect 14574 22144 14866 22681
rect 15034 22144 15326 22681
rect 15494 22144 15786 22681
rect 15954 22144 16246 22681
rect 16414 22144 16706 22681
rect 16874 22144 17166 22681
rect 17334 22144 17626 22681
rect 17794 22144 18086 22681
rect 18254 22144 18546 22681
rect 18714 22144 19006 22681
rect 19174 22144 19466 22681
rect 19634 22144 19926 22681
rect 20094 22144 20386 22681
rect 20554 22144 20846 22681
rect 21014 22144 21306 22681
rect 21474 22144 21766 22681
rect 21934 22144 22226 22681
rect 22394 22144 22686 22681
rect 204 856 22796 22144
rect 204 167 11462 856
rect 11630 167 22796 856
<< metal3 >>
rect 0 22584 800 22704
rect 0 22176 800 22296
rect 0 21632 800 21752
rect 0 21224 800 21344
rect 0 20680 800 20800
rect 0 20272 800 20392
rect 0 19728 800 19848
rect 0 19320 800 19440
rect 0 18776 800 18896
rect 0 18368 800 18488
rect 0 17960 800 18080
rect 0 17416 800 17536
rect 0 17008 800 17128
rect 0 16464 800 16584
rect 0 16056 800 16176
rect 0 15512 800 15632
rect 0 15104 800 15224
rect 0 14560 800 14680
rect 0 14152 800 14272
rect 0 13744 800 13864
rect 0 13200 800 13320
rect 0 12792 800 12912
rect 0 12248 800 12368
rect 0 11840 800 11960
rect 0 11296 800 11416
rect 22200 11432 23000 11552
rect 0 10888 800 11008
rect 0 10344 800 10464
rect 0 9936 800 10056
rect 0 9392 800 9512
rect 0 8984 800 9104
rect 0 8576 800 8696
rect 0 8032 800 8152
rect 0 7624 800 7744
rect 0 7080 800 7200
rect 0 6672 800 6792
rect 0 6128 800 6248
rect 0 5720 800 5840
rect 0 5176 800 5296
rect 0 4768 800 4888
rect 0 4360 800 4480
rect 0 3816 800 3936
rect 0 3408 800 3528
rect 0 2864 800 2984
rect 0 2456 800 2576
rect 0 1912 800 2032
rect 0 1504 800 1624
rect 0 960 800 1080
rect 0 552 800 672
rect 0 144 800 264
<< obsm3 >>
rect 880 22504 22200 22677
rect 800 22376 22200 22504
rect 880 22096 22200 22376
rect 800 21832 22200 22096
rect 880 21552 22200 21832
rect 800 21424 22200 21552
rect 880 21144 22200 21424
rect 800 20880 22200 21144
rect 880 20600 22200 20880
rect 800 20472 22200 20600
rect 880 20192 22200 20472
rect 800 19928 22200 20192
rect 880 19648 22200 19928
rect 800 19520 22200 19648
rect 880 19240 22200 19520
rect 800 18976 22200 19240
rect 880 18696 22200 18976
rect 800 18568 22200 18696
rect 880 18288 22200 18568
rect 800 18160 22200 18288
rect 880 17880 22200 18160
rect 800 17616 22200 17880
rect 880 17336 22200 17616
rect 800 17208 22200 17336
rect 880 16928 22200 17208
rect 800 16664 22200 16928
rect 880 16384 22200 16664
rect 800 16256 22200 16384
rect 880 15976 22200 16256
rect 800 15712 22200 15976
rect 880 15432 22200 15712
rect 800 15304 22200 15432
rect 880 15024 22200 15304
rect 800 14760 22200 15024
rect 880 14480 22200 14760
rect 800 14352 22200 14480
rect 880 14072 22200 14352
rect 800 13944 22200 14072
rect 880 13664 22200 13944
rect 800 13400 22200 13664
rect 880 13120 22200 13400
rect 800 12992 22200 13120
rect 880 12712 22200 12992
rect 800 12448 22200 12712
rect 880 12168 22200 12448
rect 800 12040 22200 12168
rect 880 11760 22200 12040
rect 800 11632 22200 11760
rect 800 11496 22120 11632
rect 880 11352 22120 11496
rect 880 11216 22200 11352
rect 800 11088 22200 11216
rect 880 10808 22200 11088
rect 800 10544 22200 10808
rect 880 10264 22200 10544
rect 800 10136 22200 10264
rect 880 9856 22200 10136
rect 800 9592 22200 9856
rect 880 9312 22200 9592
rect 800 9184 22200 9312
rect 880 8904 22200 9184
rect 800 8776 22200 8904
rect 880 8496 22200 8776
rect 800 8232 22200 8496
rect 880 7952 22200 8232
rect 800 7824 22200 7952
rect 880 7544 22200 7824
rect 800 7280 22200 7544
rect 880 7000 22200 7280
rect 800 6872 22200 7000
rect 880 6592 22200 6872
rect 800 6328 22200 6592
rect 880 6048 22200 6328
rect 800 5920 22200 6048
rect 880 5640 22200 5920
rect 800 5376 22200 5640
rect 880 5096 22200 5376
rect 800 4968 22200 5096
rect 880 4688 22200 4968
rect 800 4560 22200 4688
rect 880 4280 22200 4560
rect 800 4016 22200 4280
rect 880 3736 22200 4016
rect 800 3608 22200 3736
rect 880 3328 22200 3608
rect 800 3064 22200 3328
rect 880 2784 22200 3064
rect 800 2656 22200 2784
rect 880 2376 22200 2656
rect 800 2112 22200 2376
rect 880 1832 22200 2112
rect 800 1704 22200 1832
rect 880 1424 22200 1704
rect 800 1160 22200 1424
rect 880 880 22200 1160
rect 800 752 22200 880
rect 880 472 22200 752
rect 800 344 22200 472
rect 880 171 22200 344
<< metal4 >>
rect 4409 2128 4729 20720
rect 7875 2128 8195 20720
rect 11340 2128 11660 20720
rect 14805 2128 15125 20720
rect 18271 2128 18591 20720
<< obsm4 >>
rect 8275 2128 11260 20720
rect 11740 2128 14725 20720
rect 15205 2128 18191 20720
<< labels >>
rlabel metal3 s 22200 11432 23000 11552 6 ccff_head
port 1 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 ccff_tail
port 2 nsew signal output
rlabel metal3 s 0 4360 800 4480 6 chanx_left_in[0]
port 3 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[10]
port 4 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[11]
port 5 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 chanx_left_in[12]
port 6 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[13]
port 7 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[14]
port 8 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[15]
port 9 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 chanx_left_in[16]
port 10 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[17]
port 11 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 chanx_left_in[18]
port 12 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 chanx_left_in[19]
port 13 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[1]
port 14 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 chanx_left_in[2]
port 15 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 chanx_left_in[3]
port 16 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 chanx_left_in[4]
port 17 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 chanx_left_in[5]
port 18 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 chanx_left_in[6]
port 19 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 chanx_left_in[7]
port 20 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[8]
port 21 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 chanx_left_in[9]
port 22 nsew signal input
rlabel metal3 s 0 13744 800 13864 6 chanx_left_out[0]
port 23 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 chanx_left_out[10]
port 24 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[11]
port 25 nsew signal output
rlabel metal3 s 0 19320 800 19440 6 chanx_left_out[12]
port 26 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 chanx_left_out[13]
port 27 nsew signal output
rlabel metal3 s 0 20272 800 20392 6 chanx_left_out[14]
port 28 nsew signal output
rlabel metal3 s 0 20680 800 20800 6 chanx_left_out[15]
port 29 nsew signal output
rlabel metal3 s 0 21224 800 21344 6 chanx_left_out[16]
port 30 nsew signal output
rlabel metal3 s 0 21632 800 21752 6 chanx_left_out[17]
port 31 nsew signal output
rlabel metal3 s 0 22176 800 22296 6 chanx_left_out[18]
port 32 nsew signal output
rlabel metal3 s 0 22584 800 22704 6 chanx_left_out[19]
port 33 nsew signal output
rlabel metal3 s 0 14152 800 14272 6 chanx_left_out[1]
port 34 nsew signal output
rlabel metal3 s 0 14560 800 14680 6 chanx_left_out[2]
port 35 nsew signal output
rlabel metal3 s 0 15104 800 15224 6 chanx_left_out[3]
port 36 nsew signal output
rlabel metal3 s 0 15512 800 15632 6 chanx_left_out[4]
port 37 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 chanx_left_out[5]
port 38 nsew signal output
rlabel metal3 s 0 16464 800 16584 6 chanx_left_out[6]
port 39 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 chanx_left_out[7]
port 40 nsew signal output
rlabel metal3 s 0 17416 800 17536 6 chanx_left_out[8]
port 41 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 chanx_left_out[9]
port 42 nsew signal output
rlabel metal2 s 3882 22200 3938 23000 6 chany_top_in[0]
port 43 nsew signal input
rlabel metal2 s 8482 22200 8538 23000 6 chany_top_in[10]
port 44 nsew signal input
rlabel metal2 s 8942 22200 8998 23000 6 chany_top_in[11]
port 45 nsew signal input
rlabel metal2 s 9402 22200 9458 23000 6 chany_top_in[12]
port 46 nsew signal input
rlabel metal2 s 9862 22200 9918 23000 6 chany_top_in[13]
port 47 nsew signal input
rlabel metal2 s 10322 22200 10378 23000 6 chany_top_in[14]
port 48 nsew signal input
rlabel metal2 s 10782 22200 10838 23000 6 chany_top_in[15]
port 49 nsew signal input
rlabel metal2 s 11242 22200 11298 23000 6 chany_top_in[16]
port 50 nsew signal input
rlabel metal2 s 11702 22200 11758 23000 6 chany_top_in[17]
port 51 nsew signal input
rlabel metal2 s 12162 22200 12218 23000 6 chany_top_in[18]
port 52 nsew signal input
rlabel metal2 s 12622 22200 12678 23000 6 chany_top_in[19]
port 53 nsew signal input
rlabel metal2 s 4342 22200 4398 23000 6 chany_top_in[1]
port 54 nsew signal input
rlabel metal2 s 4802 22200 4858 23000 6 chany_top_in[2]
port 55 nsew signal input
rlabel metal2 s 5262 22200 5318 23000 6 chany_top_in[3]
port 56 nsew signal input
rlabel metal2 s 5722 22200 5778 23000 6 chany_top_in[4]
port 57 nsew signal input
rlabel metal2 s 6182 22200 6238 23000 6 chany_top_in[5]
port 58 nsew signal input
rlabel metal2 s 6642 22200 6698 23000 6 chany_top_in[6]
port 59 nsew signal input
rlabel metal2 s 7102 22200 7158 23000 6 chany_top_in[7]
port 60 nsew signal input
rlabel metal2 s 7562 22200 7618 23000 6 chany_top_in[8]
port 61 nsew signal input
rlabel metal2 s 8022 22200 8078 23000 6 chany_top_in[9]
port 62 nsew signal input
rlabel metal2 s 13082 22200 13138 23000 6 chany_top_out[0]
port 63 nsew signal output
rlabel metal2 s 17682 22200 17738 23000 6 chany_top_out[10]
port 64 nsew signal output
rlabel metal2 s 18142 22200 18198 23000 6 chany_top_out[11]
port 65 nsew signal output
rlabel metal2 s 18602 22200 18658 23000 6 chany_top_out[12]
port 66 nsew signal output
rlabel metal2 s 19062 22200 19118 23000 6 chany_top_out[13]
port 67 nsew signal output
rlabel metal2 s 19522 22200 19578 23000 6 chany_top_out[14]
port 68 nsew signal output
rlabel metal2 s 19982 22200 20038 23000 6 chany_top_out[15]
port 69 nsew signal output
rlabel metal2 s 20442 22200 20498 23000 6 chany_top_out[16]
port 70 nsew signal output
rlabel metal2 s 20902 22200 20958 23000 6 chany_top_out[17]
port 71 nsew signal output
rlabel metal2 s 21362 22200 21418 23000 6 chany_top_out[18]
port 72 nsew signal output
rlabel metal2 s 21822 22200 21878 23000 6 chany_top_out[19]
port 73 nsew signal output
rlabel metal2 s 13542 22200 13598 23000 6 chany_top_out[1]
port 74 nsew signal output
rlabel metal2 s 14002 22200 14058 23000 6 chany_top_out[2]
port 75 nsew signal output
rlabel metal2 s 14462 22200 14518 23000 6 chany_top_out[3]
port 76 nsew signal output
rlabel metal2 s 14922 22200 14978 23000 6 chany_top_out[4]
port 77 nsew signal output
rlabel metal2 s 15382 22200 15438 23000 6 chany_top_out[5]
port 78 nsew signal output
rlabel metal2 s 15842 22200 15898 23000 6 chany_top_out[6]
port 79 nsew signal output
rlabel metal2 s 16302 22200 16358 23000 6 chany_top_out[7]
port 80 nsew signal output
rlabel metal2 s 16762 22200 16818 23000 6 chany_top_out[8]
port 81 nsew signal output
rlabel metal2 s 17222 22200 17278 23000 6 chany_top_out[9]
port 82 nsew signal output
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_11_
port 83 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 left_bottom_grid_pin_13_
port 84 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 left_bottom_grid_pin_15_
port 85 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 left_bottom_grid_pin_17_
port 86 nsew signal input
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_1_
port 87 nsew signal input
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_3_
port 88 nsew signal input
rlabel metal3 s 0 960 800 1080 6 left_bottom_grid_pin_5_
port 89 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 left_bottom_grid_pin_7_
port 90 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 left_bottom_grid_pin_9_
port 91 nsew signal input
rlabel metal2 s 22282 22200 22338 23000 6 prog_clk_0_N_in
port 92 nsew signal input
rlabel metal2 s 202 22200 258 23000 6 top_left_grid_pin_42_
port 93 nsew signal input
rlabel metal2 s 662 22200 718 23000 6 top_left_grid_pin_43_
port 94 nsew signal input
rlabel metal2 s 1122 22200 1178 23000 6 top_left_grid_pin_44_
port 95 nsew signal input
rlabel metal2 s 1582 22200 1638 23000 6 top_left_grid_pin_45_
port 96 nsew signal input
rlabel metal2 s 2042 22200 2098 23000 6 top_left_grid_pin_46_
port 97 nsew signal input
rlabel metal2 s 2502 22200 2558 23000 6 top_left_grid_pin_47_
port 98 nsew signal input
rlabel metal2 s 2962 22200 3018 23000 6 top_left_grid_pin_48_
port 99 nsew signal input
rlabel metal2 s 3422 22200 3478 23000 6 top_left_grid_pin_49_
port 100 nsew signal input
rlabel metal2 s 22742 22200 22798 23000 6 top_right_grid_pin_1_
port 101 nsew signal input
rlabel metal4 s 18271 2128 18591 20720 6 VPWR
port 102 nsew power bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VPWR
port 103 nsew power bidirectional
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 104 nsew power bidirectional
rlabel metal4 s 14805 2128 15125 20720 6 VGND
port 105 nsew ground bidirectional
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 106 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 23000 23000
string LEFview TRUE
string GDS_FILE /project/openlane/sb_2__0_/runs/sb_2__0_/results/magic/sb_2__0_.gds
string GDS_END 1078492
string GDS_START 80590
<< end >>

