magic
tech sky130A
magscale 1 2
timestamp 1625785660
<< locali >>
rect 6653 11679 6687 11849
rect 11529 11543 11563 11645
rect 18981 11271 19015 12257
rect 4261 9911 4295 10149
rect 15945 7871 15979 8041
rect 3709 5559 3743 5797
rect 7849 4539 7883 4709
<< viali >>
rect 1869 14569 1903 14603
rect 2237 14569 2271 14603
rect 3617 14569 3651 14603
rect 4445 14569 4479 14603
rect 16313 14569 16347 14603
rect 1501 14501 1535 14535
rect 4905 14501 4939 14535
rect 5917 14501 5951 14535
rect 9873 14501 9907 14535
rect 16037 14501 16071 14535
rect 17509 14501 17543 14535
rect 17693 14501 17727 14535
rect 1961 14433 1995 14467
rect 2329 14433 2363 14467
rect 2697 14433 2731 14467
rect 2789 14433 2823 14467
rect 3065 14433 3099 14467
rect 3525 14433 3559 14467
rect 3893 14433 3927 14467
rect 4353 14433 4387 14467
rect 4629 14433 4663 14467
rect 6101 14433 6135 14467
rect 10057 14433 10091 14467
rect 16129 14433 16163 14467
rect 16589 14433 16623 14467
rect 16957 14433 16991 14467
rect 17233 14433 17267 14467
rect 18153 14433 18187 14467
rect 18429 14433 18463 14467
rect 1685 14297 1719 14331
rect 2973 14297 3007 14331
rect 3249 14297 3283 14331
rect 16405 14297 16439 14331
rect 16773 14297 16807 14331
rect 17969 14297 18003 14331
rect 2513 14229 2547 14263
rect 3341 14229 3375 14263
rect 4077 14229 4111 14263
rect 4169 14229 4203 14263
rect 4721 14229 4755 14263
rect 17417 14229 17451 14263
rect 18337 14229 18371 14263
rect 1869 14025 1903 14059
rect 2789 14025 2823 14059
rect 9781 14025 9815 14059
rect 15393 14025 15427 14059
rect 16405 14025 16439 14059
rect 16773 14025 16807 14059
rect 2145 13957 2179 13991
rect 2513 13957 2547 13991
rect 3065 13957 3099 13991
rect 3341 13957 3375 13991
rect 3893 13957 3927 13991
rect 4169 13957 4203 13991
rect 16589 13957 16623 13991
rect 3525 13889 3559 13923
rect 3801 13889 3835 13923
rect 15853 13889 15887 13923
rect 17049 13889 17083 13923
rect 17877 13889 17911 13923
rect 18245 13889 18279 13923
rect 1409 13821 1443 13855
rect 2329 13821 2363 13855
rect 2697 13821 2731 13855
rect 2973 13821 3007 13855
rect 3249 13821 3283 13855
rect 9597 13821 9631 13855
rect 15577 13821 15611 13855
rect 16221 13821 16255 13855
rect 17141 13821 17175 13855
rect 18429 13821 18463 13855
rect 1593 13753 1627 13787
rect 1961 13753 1995 13787
rect 17325 13753 17359 13787
rect 17693 13753 17727 13787
rect 18061 13753 18095 13787
rect 17601 13685 17635 13719
rect 1777 13481 1811 13515
rect 2421 13481 2455 13515
rect 2973 13481 3007 13515
rect 6101 13481 6135 13515
rect 16405 13481 16439 13515
rect 17141 13481 17175 13515
rect 17325 13481 17359 13515
rect 17969 13481 18003 13515
rect 2697 13413 2731 13447
rect 17509 13413 17543 13447
rect 18429 13413 18463 13447
rect 1501 13345 1535 13379
rect 1961 13345 1995 13379
rect 2145 13345 2179 13379
rect 2605 13345 2639 13379
rect 6285 13345 6319 13379
rect 17785 13345 17819 13379
rect 18061 13345 18095 13379
rect 16129 13277 16163 13311
rect 16589 13277 16623 13311
rect 16773 13277 16807 13311
rect 2329 13209 2363 13243
rect 18245 13209 18279 13243
rect 1593 13141 1627 13175
rect 16865 13141 16899 13175
rect 17601 13141 17635 13175
rect 1961 12937 1995 12971
rect 15485 12937 15519 12971
rect 15669 12937 15703 12971
rect 16313 12937 16347 12971
rect 1685 12869 1719 12903
rect 17601 12869 17635 12903
rect 2513 12801 2547 12835
rect 16037 12801 16071 12835
rect 17049 12801 17083 12835
rect 2697 12733 2731 12767
rect 17325 12733 17359 12767
rect 17785 12733 17819 12767
rect 18429 12733 18463 12767
rect 1501 12665 1535 12699
rect 1869 12665 1903 12699
rect 2237 12665 2271 12699
rect 2881 12665 2915 12699
rect 3157 12665 3191 12699
rect 8861 12665 8895 12699
rect 16405 12665 16439 12699
rect 17233 12665 17267 12699
rect 17877 12665 17911 12699
rect 18061 12665 18095 12699
rect 18245 12665 18279 12699
rect 2329 12597 2363 12631
rect 3341 12597 3375 12631
rect 3617 12597 3651 12631
rect 3801 12597 3835 12631
rect 9137 12597 9171 12631
rect 15853 12597 15887 12631
rect 16773 12597 16807 12631
rect 17509 12597 17543 12631
rect 1593 12393 1627 12427
rect 5549 12393 5583 12427
rect 5733 12393 5767 12427
rect 7941 12393 7975 12427
rect 9873 12393 9907 12427
rect 11161 12393 11195 12427
rect 18337 12393 18371 12427
rect 2145 12325 2179 12359
rect 4353 12325 4387 12359
rect 8493 12325 8527 12359
rect 8677 12325 8711 12359
rect 15393 12325 15427 12359
rect 17417 12325 17451 12359
rect 1501 12257 1535 12291
rect 1869 12257 1903 12291
rect 2881 12257 2915 12291
rect 4169 12257 4203 12291
rect 7021 12257 7055 12291
rect 9505 12257 9539 12291
rect 14841 12257 14875 12291
rect 15301 12257 15335 12291
rect 16221 12257 16255 12291
rect 17969 12257 18003 12291
rect 18429 12257 18463 12291
rect 18981 12257 19015 12291
rect 2697 12189 2731 12223
rect 3525 12189 3559 12223
rect 5181 12189 5215 12223
rect 5365 12189 5399 12223
rect 7205 12189 7239 12223
rect 7297 12189 7331 12223
rect 8217 12189 8251 12223
rect 8769 12189 8803 12223
rect 9229 12189 9263 12223
rect 9413 12189 9447 12223
rect 10333 12189 10367 12223
rect 10609 12189 10643 12223
rect 15025 12189 15059 12223
rect 15577 12189 15611 12223
rect 16773 12189 16807 12223
rect 17141 12189 17175 12223
rect 2329 12121 2363 12155
rect 2605 12121 2639 12155
rect 3709 12121 3743 12155
rect 4997 12121 5031 12155
rect 6009 12121 6043 12155
rect 15853 12121 15887 12155
rect 17785 12121 17819 12155
rect 1961 12053 1995 12087
rect 3065 12053 3099 12087
rect 3341 12053 3375 12087
rect 3985 12053 4019 12087
rect 4537 12053 4571 12087
rect 4813 12053 4847 12087
rect 6193 12053 6227 12087
rect 6377 12053 6411 12087
rect 6561 12053 6595 12087
rect 6837 12053 6871 12087
rect 8033 12053 8067 12087
rect 9965 12053 9999 12087
rect 10241 12053 10275 12087
rect 10793 12053 10827 12087
rect 11253 12053 11287 12087
rect 14565 12053 14599 12087
rect 16037 12053 16071 12087
rect 16405 12053 16439 12087
rect 16865 12053 16899 12087
rect 17509 12053 17543 12087
rect 18061 12053 18095 12087
rect 5457 11849 5491 11883
rect 6653 11849 6687 11883
rect 8033 11849 8067 11883
rect 14289 11849 14323 11883
rect 15025 11849 15059 11883
rect 17233 11849 17267 11883
rect 1685 11781 1719 11815
rect 3157 11781 3191 11815
rect 2237 11713 2271 11747
rect 4813 11713 4847 11747
rect 6469 11713 6503 11747
rect 9689 11781 9723 11815
rect 12081 11781 12115 11815
rect 14657 11781 14691 11815
rect 18153 11781 18187 11815
rect 7297 11713 7331 11747
rect 8125 11713 8159 11747
rect 10425 11713 10459 11747
rect 10793 11713 10827 11747
rect 12265 11713 12299 11747
rect 16773 11713 16807 11747
rect 1777 11645 1811 11679
rect 2973 11645 3007 11679
rect 3709 11645 3743 11679
rect 3985 11645 4019 11679
rect 4997 11645 5031 11679
rect 5641 11645 5675 11679
rect 6009 11645 6043 11679
rect 6653 11645 6687 11679
rect 8309 11645 8343 11679
rect 10977 11645 11011 11679
rect 11529 11645 11563 11679
rect 14841 11645 14875 11679
rect 15117 11645 15151 11679
rect 15945 11645 15979 11679
rect 17049 11645 17083 11679
rect 17509 11645 17543 11679
rect 1501 11577 1535 11611
rect 4537 11577 4571 11611
rect 5825 11577 5859 11611
rect 7113 11577 7147 11611
rect 8565 11577 8599 11611
rect 11069 11577 11103 11611
rect 11713 11577 11747 11611
rect 12449 11577 12483 11611
rect 14473 11577 14507 11611
rect 17877 11577 17911 11611
rect 18429 11577 18463 11611
rect 1961 11509 1995 11543
rect 2329 11509 2363 11543
rect 2421 11509 2455 11543
rect 2789 11509 2823 11543
rect 3249 11509 3283 11543
rect 3525 11509 3559 11543
rect 4077 11509 4111 11543
rect 4261 11509 4295 11543
rect 5273 11509 5307 11543
rect 6285 11509 6319 11543
rect 6745 11509 6779 11543
rect 7205 11509 7239 11543
rect 7665 11509 7699 11543
rect 9781 11509 9815 11543
rect 10149 11509 10183 11543
rect 10241 11509 10275 11543
rect 11437 11509 11471 11543
rect 11529 11509 11563 11543
rect 14013 11509 14047 11543
rect 16313 11509 16347 11543
rect 16497 11509 16531 11543
rect 17417 11509 17451 11543
rect 17785 11509 17819 11543
rect 5181 11305 5215 11339
rect 7205 11305 7239 11339
rect 7573 11305 7607 11339
rect 7665 11305 7699 11339
rect 8585 11305 8619 11339
rect 11253 11305 11287 11339
rect 11713 11305 11747 11339
rect 12265 11305 12299 11339
rect 12909 11305 12943 11339
rect 13461 11305 13495 11339
rect 17969 11305 18003 11339
rect 3893 11237 3927 11271
rect 6592 11237 6626 11271
rect 12173 11237 12207 11271
rect 14105 11237 14139 11271
rect 14473 11237 14507 11271
rect 18981 11237 19015 11271
rect 1501 11169 1535 11203
rect 1869 11169 1903 11203
rect 3442 11169 3476 11203
rect 9321 11169 9355 11203
rect 10618 11169 10652 11203
rect 11345 11169 11379 11203
rect 14841 11169 14875 11203
rect 15373 11169 15407 11203
rect 16773 11169 16807 11203
rect 17049 11169 17083 11203
rect 17417 11169 17451 11203
rect 17877 11169 17911 11203
rect 18337 11169 18371 11203
rect 2145 11101 2179 11135
rect 3709 11101 3743 11135
rect 4169 11101 4203 11135
rect 4813 11101 4847 11135
rect 6837 11101 6871 11135
rect 7757 11101 7791 11135
rect 8125 11101 8159 11135
rect 8309 11101 8343 11135
rect 8493 11101 8527 11135
rect 9137 11101 9171 11135
rect 10885 11101 10919 11135
rect 11069 11101 11103 11135
rect 12357 11101 12391 11135
rect 13001 11101 13035 11135
rect 13553 11101 13587 11135
rect 14657 11101 14691 11135
rect 15117 11101 15151 11135
rect 18153 11101 18187 11135
rect 1685 11033 1719 11067
rect 4353 11033 4387 11067
rect 4445 11033 4479 11067
rect 5457 11033 5491 11067
rect 8953 11033 8987 11067
rect 9505 11033 9539 11067
rect 11805 11033 11839 11067
rect 12633 11033 12667 11067
rect 13277 11033 13311 11067
rect 14013 11033 14047 11067
rect 15025 11033 15059 11067
rect 16589 11033 16623 11067
rect 17233 11033 17267 11067
rect 17509 11033 17543 11067
rect 1961 10965 1995 10999
rect 2329 10965 2363 10999
rect 4721 10965 4755 10999
rect 5089 10965 5123 10999
rect 7021 10965 7055 10999
rect 13829 10965 13863 10999
rect 16497 10965 16531 10999
rect 16865 10965 16899 10999
rect 2329 10761 2363 10795
rect 7941 10761 7975 10795
rect 9505 10761 9539 10795
rect 11989 10761 12023 10795
rect 15117 10761 15151 10795
rect 2237 10693 2271 10727
rect 4077 10693 4111 10727
rect 8953 10693 8987 10727
rect 9137 10693 9171 10727
rect 11437 10693 11471 10727
rect 1685 10625 1719 10659
rect 2973 10625 3007 10659
rect 3893 10625 3927 10659
rect 5733 10625 5767 10659
rect 8493 10625 8527 10659
rect 10149 10625 10183 10659
rect 10885 10625 10919 10659
rect 11713 10625 11747 10659
rect 1869 10557 1903 10591
rect 5457 10557 5491 10591
rect 6469 10557 6503 10591
rect 6725 10557 6759 10591
rect 8309 10557 8343 10591
rect 9965 10557 9999 10591
rect 10701 10557 10735 10591
rect 12265 10557 12299 10591
rect 13737 10557 13771 10591
rect 16589 10557 16623 10591
rect 16957 10557 16991 10591
rect 1777 10489 1811 10523
rect 2697 10489 2731 10523
rect 2789 10489 2823 10523
rect 3709 10489 3743 10523
rect 5190 10489 5224 10523
rect 5917 10489 5951 10523
rect 9873 10489 9907 10523
rect 12532 10489 12566 10523
rect 14004 10489 14038 10523
rect 16344 10489 16378 10523
rect 17202 10489 17236 10523
rect 3249 10421 3283 10455
rect 3617 10421 3651 10455
rect 5825 10421 5859 10455
rect 6285 10421 6319 10455
rect 7849 10421 7883 10455
rect 8401 10421 8435 10455
rect 8769 10421 8803 10455
rect 9321 10421 9355 10455
rect 10333 10421 10367 10455
rect 10793 10421 10827 10455
rect 11253 10421 11287 10455
rect 12081 10421 12115 10455
rect 13645 10421 13679 10455
rect 15209 10421 15243 10455
rect 16681 10421 16715 10455
rect 18337 10421 18371 10455
rect 18521 10421 18555 10455
rect 3249 10217 3283 10251
rect 4353 10217 4387 10251
rect 4813 10217 4847 10251
rect 5641 10217 5675 10251
rect 6009 10217 6043 10251
rect 7021 10217 7055 10251
rect 7573 10217 7607 10251
rect 7941 10217 7975 10251
rect 8309 10217 8343 10251
rect 9781 10217 9815 10251
rect 10149 10217 10183 10251
rect 11713 10217 11747 10251
rect 14105 10217 14139 10251
rect 14749 10217 14783 10251
rect 15577 10217 15611 10251
rect 15945 10217 15979 10251
rect 16589 10217 16623 10251
rect 18153 10217 18187 10251
rect 3341 10149 3375 10183
rect 4261 10149 4295 10183
rect 5549 10149 5583 10183
rect 17417 10149 17451 10183
rect 18245 10149 18279 10183
rect 2533 10081 2567 10115
rect 2789 10081 2823 10115
rect 3985 10081 4019 10115
rect 3157 10013 3191 10047
rect 4169 10013 4203 10047
rect 4721 10081 4755 10115
rect 6653 10081 6687 10115
rect 7481 10081 7515 10115
rect 8769 10081 8803 10115
rect 11354 10081 11388 10115
rect 11621 10081 11655 10115
rect 11897 10081 11931 10115
rect 12164 10081 12198 10115
rect 13737 10081 13771 10115
rect 16497 10081 16531 10115
rect 17325 10081 17359 10115
rect 4905 10013 4939 10047
rect 5733 10013 5767 10047
rect 6377 10013 6411 10047
rect 6561 10013 6595 10047
rect 7665 10013 7699 10047
rect 8401 10013 8435 10047
rect 8493 10013 8527 10047
rect 9137 10013 9171 10047
rect 9597 10013 9631 10047
rect 9689 10013 9723 10047
rect 13461 10013 13495 10047
rect 13645 10013 13679 10047
rect 14841 10013 14875 10047
rect 14933 10013 14967 10047
rect 15301 10013 15335 10047
rect 15485 10013 15519 10047
rect 16681 10013 16715 10047
rect 17509 10013 17543 10047
rect 18337 10013 18371 10047
rect 5181 9945 5215 9979
rect 7113 9945 7147 9979
rect 10241 9945 10275 9979
rect 1409 9877 1443 9911
rect 3709 9877 3743 9911
rect 4261 9877 4295 9911
rect 8953 9877 8987 9911
rect 13277 9877 13311 9911
rect 14381 9877 14415 9911
rect 16129 9877 16163 9911
rect 16957 9877 16991 9911
rect 17785 9877 17819 9911
rect 3065 9673 3099 9707
rect 7849 9673 7883 9707
rect 10793 9673 10827 9707
rect 11253 9673 11287 9707
rect 13737 9673 13771 9707
rect 1777 9605 1811 9639
rect 4169 9605 4203 9639
rect 5733 9605 5767 9639
rect 5825 9605 5859 9639
rect 13277 9605 13311 9639
rect 14565 9605 14599 9639
rect 15485 9605 15519 9639
rect 15945 9605 15979 9639
rect 18521 9605 18555 9639
rect 2329 9537 2363 9571
rect 2513 9537 2547 9571
rect 3525 9537 3559 9571
rect 3617 9537 3651 9571
rect 4813 9537 4847 9571
rect 5089 9537 5123 9571
rect 7941 9537 7975 9571
rect 9413 9537 9447 9571
rect 10885 9537 10919 9571
rect 11805 9537 11839 9571
rect 11897 9537 11931 9571
rect 13093 9537 13127 9571
rect 14381 9537 14415 9571
rect 15209 9537 15243 9571
rect 16405 9537 16439 9571
rect 16497 9537 16531 9571
rect 2145 9469 2179 9503
rect 2605 9469 2639 9503
rect 3433 9469 3467 9503
rect 3893 9469 3927 9503
rect 4629 9469 4663 9503
rect 6009 9469 6043 9503
rect 6285 9469 6319 9503
rect 6469 9469 6503 9503
rect 11437 9469 11471 9503
rect 12265 9469 12299 9503
rect 12817 9469 12851 9503
rect 15025 9469 15059 9503
rect 16313 9469 16347 9503
rect 16957 9469 16991 9503
rect 1501 9401 1535 9435
rect 5365 9401 5399 9435
rect 6714 9401 6748 9435
rect 8186 9401 8220 9435
rect 9680 9401 9714 9435
rect 13645 9401 13679 9435
rect 14933 9401 14967 9435
rect 15669 9401 15703 9435
rect 17224 9401 17258 9435
rect 1961 9333 1995 9367
rect 2973 9333 3007 9367
rect 4077 9333 4111 9367
rect 4537 9333 4571 9367
rect 5273 9333 5307 9367
rect 6101 9333 6135 9367
rect 9321 9333 9355 9367
rect 11161 9333 11195 9367
rect 12081 9333 12115 9367
rect 12449 9333 12483 9367
rect 12909 9333 12943 9367
rect 14105 9333 14139 9367
rect 14197 9333 14231 9367
rect 15761 9333 15795 9367
rect 18337 9333 18371 9367
rect 4629 9129 4663 9163
rect 6377 9129 6411 9163
rect 6837 9129 6871 9163
rect 7205 9129 7239 9163
rect 10701 9129 10735 9163
rect 12081 9129 12115 9163
rect 13001 9129 13035 9163
rect 15761 9129 15795 9163
rect 17785 9129 17819 9163
rect 2890 9061 2924 9095
rect 5264 9061 5298 9095
rect 8585 9061 8619 9095
rect 9496 9061 9530 9095
rect 11069 9061 11103 9095
rect 16098 9061 16132 9095
rect 17693 9061 17727 9095
rect 1501 8993 1535 9027
rect 3341 8993 3375 9027
rect 4261 8993 4295 9027
rect 4905 8993 4939 9027
rect 6745 8993 6779 9027
rect 7665 8993 7699 9027
rect 8677 8993 8711 9027
rect 9229 8993 9263 9027
rect 11161 8993 11195 9027
rect 11897 8993 11931 9027
rect 12541 8993 12575 9027
rect 13369 8993 13403 9027
rect 14013 8993 14047 9027
rect 14648 8993 14682 9027
rect 18521 8993 18555 9027
rect 3157 8925 3191 8959
rect 3617 8925 3651 8959
rect 4077 8925 4111 8959
rect 4169 8925 4203 8959
rect 5004 8925 5038 8959
rect 6653 8925 6687 8959
rect 7389 8925 7423 8959
rect 7573 8925 7607 8959
rect 8861 8925 8895 8959
rect 11253 8925 11287 8959
rect 12357 8925 12391 8959
rect 12449 8925 12483 8959
rect 13461 8925 13495 8959
rect 13645 8925 13679 8959
rect 14381 8925 14415 8959
rect 15853 8925 15887 8959
rect 17877 8925 17911 8959
rect 1685 8857 1719 8891
rect 8033 8857 8067 8891
rect 17325 8857 17359 8891
rect 18337 8857 18371 8891
rect 1777 8789 1811 8823
rect 3433 8789 3467 8823
rect 4721 8789 4755 8823
rect 8217 8789 8251 8823
rect 10609 8789 10643 8823
rect 11621 8789 11655 8823
rect 11805 8789 11839 8823
rect 12909 8789 12943 8823
rect 13921 8789 13955 8823
rect 14197 8789 14231 8823
rect 17233 8789 17267 8823
rect 1501 8585 1535 8619
rect 6193 8585 6227 8619
rect 7849 8585 7883 8619
rect 16405 8585 16439 8619
rect 4353 8517 4387 8551
rect 5825 8517 5859 8551
rect 10149 8517 10183 8551
rect 12173 8517 12207 8551
rect 13185 8517 13219 8551
rect 14013 8517 14047 8551
rect 15393 8517 15427 8551
rect 16957 8517 16991 8551
rect 18337 8517 18371 8551
rect 11529 8449 11563 8483
rect 12081 8449 12115 8483
rect 12449 8449 12483 8483
rect 12633 8449 12667 8483
rect 13829 8449 13863 8483
rect 14657 8449 14691 8483
rect 15301 8449 15335 8483
rect 15853 8449 15887 8483
rect 16037 8449 16071 8483
rect 17509 8449 17543 8483
rect 2614 8381 2648 8415
rect 2881 8381 2915 8415
rect 2973 8381 3007 8415
rect 4445 8381 4479 8415
rect 4712 8381 4746 8415
rect 6101 8381 6135 8415
rect 6469 8381 6503 8415
rect 9146 8381 9180 8415
rect 9413 8381 9447 8415
rect 9781 8381 9815 8415
rect 12725 8381 12759 8415
rect 13553 8381 13587 8415
rect 14841 8381 14875 8415
rect 15117 8381 15151 8415
rect 15761 8381 15795 8415
rect 16221 8381 16255 8415
rect 16773 8381 16807 8415
rect 17417 8381 17451 8415
rect 18521 8381 18555 8415
rect 3240 8313 3274 8347
rect 6736 8313 6770 8347
rect 11262 8313 11296 8347
rect 11897 8313 11931 8347
rect 13645 8313 13679 8347
rect 14381 8313 14415 8347
rect 16589 8313 16623 8347
rect 17325 8313 17359 8347
rect 17969 8313 18003 8347
rect 18153 8313 18187 8347
rect 5917 8245 5951 8279
rect 8033 8245 8067 8279
rect 9597 8245 9631 8279
rect 10057 8245 10091 8279
rect 13093 8245 13127 8279
rect 14473 8245 14507 8279
rect 3065 8041 3099 8075
rect 5457 8041 5491 8075
rect 6101 8041 6135 8075
rect 7849 8041 7883 8075
rect 8401 8041 8435 8075
rect 8769 8041 8803 8075
rect 8953 8041 8987 8075
rect 13737 8041 13771 8075
rect 14197 8041 14231 8075
rect 15945 8041 15979 8075
rect 16405 8041 16439 8075
rect 16773 8041 16807 8075
rect 17325 8041 17359 8075
rect 1501 7973 1535 8007
rect 5089 7973 5123 8007
rect 7941 7973 7975 8007
rect 9137 7973 9171 8007
rect 11437 7973 11471 8007
rect 2237 7905 2271 7939
rect 3525 7905 3559 7939
rect 4261 7905 4295 7939
rect 4353 7905 4387 7939
rect 5825 7905 5859 7939
rect 7225 7905 7259 7939
rect 8585 7905 8619 7939
rect 11897 7905 11931 7939
rect 12624 7905 12658 7939
rect 13829 7905 13863 7939
rect 14013 7905 14047 7939
rect 15597 7905 15631 7939
rect 16313 7905 16347 7939
rect 17233 7905 17267 7939
rect 18061 7905 18095 7939
rect 2329 7837 2363 7871
rect 2421 7837 2455 7871
rect 3157 7837 3191 7871
rect 3249 7837 3283 7871
rect 4445 7837 4479 7871
rect 4905 7837 4939 7871
rect 4997 7837 5031 7871
rect 5733 7837 5767 7871
rect 7481 7837 7515 7871
rect 7665 7837 7699 7871
rect 9321 7837 9355 7871
rect 11621 7837 11655 7871
rect 11805 7837 11839 7871
rect 12357 7837 12391 7871
rect 15853 7837 15887 7871
rect 15945 7837 15979 7871
rect 16221 7837 16255 7871
rect 17509 7837 17543 7871
rect 18153 7837 18187 7871
rect 18245 7837 18279 7871
rect 1685 7769 1719 7803
rect 8309 7769 8343 7803
rect 1869 7701 1903 7735
rect 2697 7701 2731 7735
rect 3709 7701 3743 7735
rect 3893 7701 3927 7735
rect 6009 7701 6043 7735
rect 9505 7701 9539 7735
rect 10149 7701 10183 7735
rect 12265 7701 12299 7735
rect 14473 7701 14507 7735
rect 16865 7701 16899 7735
rect 17693 7701 17727 7735
rect 1593 7497 1627 7531
rect 4169 7497 4203 7531
rect 4813 7497 4847 7531
rect 7573 7497 7607 7531
rect 8677 7497 8711 7531
rect 13185 7497 13219 7531
rect 16681 7497 16715 7531
rect 17785 7497 17819 7531
rect 4537 7429 4571 7463
rect 6469 7429 6503 7463
rect 13093 7429 13127 7463
rect 17693 7429 17727 7463
rect 1961 7361 1995 7395
rect 3157 7361 3191 7395
rect 3617 7361 3651 7395
rect 3709 7361 3743 7395
rect 4261 7361 4295 7395
rect 7021 7361 7055 7395
rect 7941 7361 7975 7395
rect 8125 7361 8159 7395
rect 9229 7361 9263 7395
rect 9597 7361 9631 7395
rect 10425 7361 10459 7395
rect 11713 7361 11747 7395
rect 13737 7361 13771 7395
rect 14473 7361 14507 7395
rect 16129 7361 16163 7395
rect 17141 7361 17175 7395
rect 18337 7361 18371 7395
rect 1409 7293 1443 7327
rect 2053 7293 2087 7327
rect 2145 7293 2179 7327
rect 4721 7293 4755 7327
rect 6193 7293 6227 7327
rect 6837 7293 6871 7327
rect 7757 7293 7791 7327
rect 9045 7293 9079 7327
rect 10701 7293 10735 7327
rect 11345 7293 11379 7327
rect 13553 7293 13587 7327
rect 14197 7293 14231 7327
rect 14740 7293 14774 7327
rect 18245 7293 18279 7327
rect 5926 7225 5960 7259
rect 7481 7225 7515 7259
rect 9781 7225 9815 7259
rect 11958 7225 11992 7259
rect 13645 7225 13679 7259
rect 2513 7157 2547 7191
rect 2605 7157 2639 7191
rect 2973 7157 3007 7191
rect 3065 7157 3099 7191
rect 3801 7157 3835 7191
rect 6929 7157 6963 7191
rect 8217 7157 8251 7191
rect 8585 7157 8619 7191
rect 9137 7157 9171 7191
rect 9873 7157 9907 7191
rect 10241 7157 10275 7191
rect 10609 7157 10643 7191
rect 11069 7157 11103 7191
rect 11253 7157 11287 7191
rect 11529 7157 11563 7191
rect 14013 7157 14047 7191
rect 14381 7157 14415 7191
rect 15853 7157 15887 7191
rect 16221 7157 16255 7191
rect 16313 7157 16347 7191
rect 17233 7157 17267 7191
rect 17325 7157 17359 7191
rect 18153 7157 18187 7191
rect 2973 6953 3007 6987
rect 3341 6953 3375 6987
rect 4261 6953 4295 6987
rect 11529 6953 11563 6987
rect 11621 6953 11655 6987
rect 13461 6953 13495 6987
rect 13829 6953 13863 6987
rect 17325 6953 17359 6987
rect 6653 6885 6687 6919
rect 7113 6885 7147 6919
rect 8033 6885 8067 6919
rect 10609 6885 10643 6919
rect 16098 6885 16132 6919
rect 1768 6817 1802 6851
rect 3433 6817 3467 6851
rect 4353 6817 4387 6851
rect 4905 6817 4939 6851
rect 6213 6817 6247 6851
rect 7021 6817 7055 6851
rect 7941 6817 7975 6851
rect 8493 6817 8527 6851
rect 8769 6817 8803 6851
rect 10261 6817 10295 6851
rect 11161 6817 11195 6851
rect 12734 6817 12768 6851
rect 13185 6817 13219 6851
rect 14648 6817 14682 6851
rect 17601 6817 17635 6851
rect 17785 6817 17819 6851
rect 17969 6817 18003 6851
rect 18153 6817 18187 6851
rect 18337 6817 18371 6851
rect 1501 6749 1535 6783
rect 3617 6749 3651 6783
rect 4445 6749 4479 6783
rect 6469 6749 6503 6783
rect 6929 6749 6963 6783
rect 7757 6749 7791 6783
rect 10517 6749 10551 6783
rect 10977 6749 11011 6783
rect 11069 6749 11103 6783
rect 13001 6749 13035 6783
rect 13921 6749 13955 6783
rect 14105 6749 14139 6783
rect 14381 6749 14415 6783
rect 15853 6749 15887 6783
rect 3893 6681 3927 6715
rect 7481 6681 7515 6715
rect 8401 6681 8435 6715
rect 13369 6681 13403 6715
rect 18521 6681 18555 6715
rect 2881 6613 2915 6647
rect 4813 6613 4847 6647
rect 5089 6613 5123 6647
rect 8677 6613 8711 6647
rect 8953 6613 8987 6647
rect 9137 6613 9171 6647
rect 15761 6613 15795 6647
rect 17233 6613 17267 6647
rect 1777 6409 1811 6443
rect 6469 6409 6503 6443
rect 11529 6409 11563 6443
rect 13921 6409 13955 6443
rect 14841 6409 14875 6443
rect 2789 6341 2823 6375
rect 6745 6341 6779 6375
rect 12357 6341 12391 6375
rect 2237 6273 2271 6307
rect 7481 6273 7515 6307
rect 10149 6273 10183 6307
rect 10977 6273 11011 6307
rect 12909 6273 12943 6307
rect 13369 6273 13403 6307
rect 14105 6273 14139 6307
rect 15485 6273 15519 6307
rect 16221 6273 16255 6307
rect 17509 6273 17543 6307
rect 17693 6273 17727 6307
rect 1501 6205 1535 6239
rect 2421 6205 2455 6239
rect 4261 6205 4295 6239
rect 4353 6205 4387 6239
rect 5825 6205 5859 6239
rect 6009 6205 6043 6239
rect 6653 6205 6687 6239
rect 7849 6205 7883 6239
rect 9597 6205 9631 6239
rect 10333 6205 10367 6239
rect 12081 6205 12115 6239
rect 12817 6205 12851 6239
rect 13461 6205 13495 6239
rect 14381 6205 14415 6239
rect 16129 6205 16163 6239
rect 16589 6205 16623 6239
rect 18337 6205 18371 6239
rect 3994 6137 4028 6171
rect 4598 6137 4632 6171
rect 7297 6137 7331 6171
rect 8116 6137 8150 6171
rect 9873 6137 9907 6171
rect 15301 6137 15335 6171
rect 16037 6137 16071 6171
rect 17969 6137 18003 6171
rect 18521 6137 18555 6171
rect 2329 6069 2363 6103
rect 2881 6069 2915 6103
rect 5733 6069 5767 6103
rect 6193 6069 6227 6103
rect 6929 6069 6963 6103
rect 7389 6069 7423 6103
rect 9229 6069 9263 6103
rect 9413 6069 9447 6103
rect 10241 6069 10275 6103
rect 10701 6069 10735 6103
rect 11069 6069 11103 6103
rect 11161 6069 11195 6103
rect 11805 6069 11839 6103
rect 12265 6069 12299 6103
rect 12725 6069 12759 6103
rect 13553 6069 13587 6103
rect 14289 6069 14323 6103
rect 14749 6069 14783 6103
rect 15209 6069 15243 6103
rect 15669 6069 15703 6103
rect 16773 6069 16807 6103
rect 17049 6069 17083 6103
rect 17417 6069 17451 6103
rect 18061 6069 18095 6103
rect 2329 5865 2363 5899
rect 2881 5865 2915 5899
rect 3249 5865 3283 5899
rect 6009 5865 6043 5899
rect 6377 5865 6411 5899
rect 6561 5865 6595 5899
rect 8033 5865 8067 5899
rect 8861 5865 8895 5899
rect 10977 5865 11011 5899
rect 11437 5865 11471 5899
rect 11805 5865 11839 5899
rect 14105 5865 14139 5899
rect 14749 5865 14783 5899
rect 15117 5865 15151 5899
rect 15945 5865 15979 5899
rect 18153 5865 18187 5899
rect 1501 5797 1535 5831
rect 3709 5797 3743 5831
rect 16764 5797 16798 5831
rect 18521 5797 18555 5831
rect 2421 5729 2455 5763
rect 2237 5661 2271 5695
rect 3341 5661 3375 5695
rect 3525 5661 3559 5695
rect 1777 5593 1811 5627
rect 4261 5729 4295 5763
rect 5181 5729 5215 5763
rect 7674 5729 7708 5763
rect 8401 5729 8435 5763
rect 8493 5729 8527 5763
rect 9393 5729 9427 5763
rect 10885 5729 10919 5763
rect 12521 5729 12555 5763
rect 13737 5729 13771 5763
rect 14657 5729 14691 5763
rect 16037 5729 16071 5763
rect 18337 5729 18371 5763
rect 4353 5661 4387 5695
rect 4445 5661 4479 5695
rect 5273 5661 5307 5695
rect 5457 5661 5491 5695
rect 5733 5661 5767 5695
rect 5917 5661 5951 5695
rect 7941 5661 7975 5695
rect 8585 5661 8619 5695
rect 9137 5661 9171 5695
rect 10701 5661 10735 5695
rect 11897 5661 11931 5695
rect 12081 5661 12115 5695
rect 12265 5661 12299 5695
rect 14473 5661 14507 5695
rect 15577 5661 15611 5695
rect 15853 5661 15887 5695
rect 16497 5661 16531 5695
rect 13645 5593 13679 5627
rect 13921 5593 13955 5627
rect 2789 5525 2823 5559
rect 3709 5525 3743 5559
rect 3893 5525 3927 5559
rect 4813 5525 4847 5559
rect 10517 5525 10551 5559
rect 11345 5525 11379 5559
rect 15209 5525 15243 5559
rect 16405 5525 16439 5559
rect 17877 5525 17911 5559
rect 1501 5321 1535 5355
rect 2329 5321 2363 5355
rect 8401 5321 8435 5355
rect 11713 5321 11747 5355
rect 13185 5321 13219 5355
rect 15117 5321 15151 5355
rect 16497 5321 16531 5355
rect 6009 5253 6043 5287
rect 9229 5253 9263 5287
rect 15393 5253 15427 5287
rect 1777 5185 1811 5219
rect 7389 5185 7423 5219
rect 8125 5185 8159 5219
rect 8953 5185 8987 5219
rect 11161 5185 11195 5219
rect 13093 5185 13127 5219
rect 14841 5185 14875 5219
rect 16129 5185 16163 5219
rect 17785 5185 17819 5219
rect 2421 5117 2455 5151
rect 3893 5117 3927 5151
rect 4445 5117 4479 5151
rect 5917 5117 5951 5151
rect 6193 5117 6227 5151
rect 6653 5117 6687 5151
rect 7113 5117 7147 5151
rect 7941 5117 7975 5151
rect 8861 5117 8895 5151
rect 9413 5117 9447 5151
rect 9689 5117 9723 5151
rect 11437 5117 11471 5151
rect 13369 5117 13403 5151
rect 14574 5117 14608 5151
rect 14933 5117 14967 5151
rect 15209 5117 15243 5151
rect 15853 5117 15887 5151
rect 16313 5117 16347 5151
rect 16589 5117 16623 5151
rect 16957 5117 16991 5151
rect 18153 5117 18187 5151
rect 2688 5049 2722 5083
rect 4077 5049 4111 5083
rect 5650 5049 5684 5083
rect 8769 5049 8803 5083
rect 10894 5049 10928 5083
rect 12826 5049 12860 5083
rect 15945 5049 15979 5083
rect 18337 5049 18371 5083
rect 18521 5049 18555 5083
rect 1869 4981 1903 5015
rect 1961 4981 1995 5015
rect 3801 4981 3835 5015
rect 4261 4981 4295 5015
rect 4537 4981 4571 5015
rect 6469 4981 6503 5015
rect 6745 4981 6779 5015
rect 7205 4981 7239 5015
rect 7573 4981 7607 5015
rect 8033 4981 8067 5015
rect 9505 4981 9539 5015
rect 9781 4981 9815 5015
rect 11253 4981 11287 5015
rect 13461 4981 13495 5015
rect 15485 4981 15519 5015
rect 16773 4981 16807 5015
rect 17141 4981 17175 5015
rect 17509 4981 17543 5015
rect 17601 4981 17635 5015
rect 17969 4981 18003 5015
rect 1777 4777 1811 4811
rect 2237 4777 2271 4811
rect 2973 4777 3007 4811
rect 6193 4777 6227 4811
rect 6653 4777 6687 4811
rect 7021 4777 7055 4811
rect 8125 4777 8159 4811
rect 8493 4777 8527 4811
rect 9597 4777 9631 4811
rect 9965 4777 9999 4811
rect 10057 4777 10091 4811
rect 10793 4777 10827 4811
rect 11529 4777 11563 4811
rect 11989 4777 12023 4811
rect 12817 4777 12851 4811
rect 13369 4777 13403 4811
rect 14197 4777 14231 4811
rect 1593 4709 1627 4743
rect 4997 4709 5031 4743
rect 6561 4709 6595 4743
rect 7849 4709 7883 4743
rect 10701 4709 10735 4743
rect 11621 4709 11655 4743
rect 13737 4709 13771 4743
rect 14933 4709 14967 4743
rect 15292 4709 15326 4743
rect 18337 4709 18371 4743
rect 2145 4641 2179 4675
rect 3433 4641 3467 4675
rect 4077 4641 4111 4675
rect 4353 4641 4387 4675
rect 4905 4641 4939 4675
rect 5549 4641 5583 4675
rect 5825 4641 5859 4675
rect 6101 4641 6135 4675
rect 7389 4641 7423 4675
rect 2329 4573 2363 4607
rect 3065 4573 3099 4607
rect 3249 4573 3283 4607
rect 5181 4573 5215 4607
rect 6745 4573 6779 4607
rect 7481 4573 7515 4607
rect 7573 4573 7607 4607
rect 8585 4641 8619 4675
rect 9321 4641 9355 4675
rect 9413 4641 9447 4675
rect 12449 4641 12483 4675
rect 13277 4641 13311 4675
rect 14565 4641 14599 4675
rect 14749 4641 14783 4675
rect 16589 4641 16623 4675
rect 16865 4641 16899 4675
rect 17509 4641 17543 4675
rect 17969 4641 18003 4675
rect 18521 4641 18555 4675
rect 8309 4573 8343 4607
rect 10241 4573 10275 4607
rect 10609 4573 10643 4607
rect 11437 4573 11471 4607
rect 12173 4573 12207 4607
rect 12357 4573 12391 4607
rect 13553 4573 13587 4607
rect 15025 4573 15059 4607
rect 17601 4573 17635 4607
rect 17785 4573 17819 4607
rect 2605 4505 2639 4539
rect 3893 4505 3927 4539
rect 4169 4505 4203 4539
rect 5641 4505 5675 4539
rect 7849 4505 7883 4539
rect 9137 4505 9171 4539
rect 14381 4505 14415 4539
rect 17049 4505 17083 4539
rect 1501 4437 1535 4471
rect 3617 4437 3651 4471
rect 4537 4437 4571 4471
rect 5365 4437 5399 4471
rect 5917 4437 5951 4471
rect 8953 4437 8987 4471
rect 11161 4437 11195 4471
rect 12909 4437 12943 4471
rect 16405 4437 16439 4471
rect 16773 4437 16807 4471
rect 17141 4437 17175 4471
rect 18153 4437 18187 4471
rect 6285 4233 6319 4267
rect 8309 4233 8343 4267
rect 16497 4233 16531 4267
rect 2513 4165 2547 4199
rect 5365 4165 5399 4199
rect 6745 4165 6779 4199
rect 11897 4165 11931 4199
rect 13553 4165 13587 4199
rect 2145 4097 2179 4131
rect 5181 4097 5215 4131
rect 5825 4097 5859 4131
rect 5917 4097 5951 4131
rect 6929 4097 6963 4131
rect 9781 4097 9815 4131
rect 11069 4097 11103 4131
rect 11161 4097 11195 4131
rect 11529 4097 11563 4131
rect 12357 4097 12391 4131
rect 12541 4097 12575 4131
rect 12817 4097 12851 4131
rect 14105 4097 14139 4131
rect 16313 4097 16347 4131
rect 17417 4097 17451 4131
rect 17601 4097 17635 4131
rect 18153 4097 18187 4131
rect 1593 4029 1627 4063
rect 2973 4029 3007 4063
rect 3240 4029 3274 4063
rect 6653 4029 6687 4063
rect 7196 4029 7230 4063
rect 9525 4029 9559 4063
rect 10057 4029 10091 4063
rect 10333 4029 10367 4063
rect 10517 4029 10551 4063
rect 10977 4029 11011 4063
rect 12265 4029 12299 4063
rect 13093 4029 13127 4063
rect 13921 4029 13955 4063
rect 14565 4029 14599 4063
rect 14841 4029 14875 4063
rect 16057 4029 16091 4063
rect 16589 4029 16623 4063
rect 17325 4029 17359 4063
rect 17969 4029 18003 4063
rect 1961 3961 1995 3995
rect 2329 3961 2363 3995
rect 2697 3961 2731 3995
rect 14013 3961 14047 3995
rect 18337 3961 18371 3995
rect 18521 3961 18555 3995
rect 1501 3893 1535 3927
rect 1869 3893 1903 3927
rect 4353 3893 4387 3927
rect 4537 3893 4571 3927
rect 4905 3893 4939 3927
rect 4997 3893 5031 3927
rect 5733 3893 5767 3927
rect 6469 3893 6503 3927
rect 8401 3893 8435 3927
rect 9873 3893 9907 3927
rect 10149 3893 10183 3927
rect 10609 3893 10643 3927
rect 11805 3893 11839 3927
rect 13001 3893 13035 3927
rect 13461 3893 13495 3927
rect 14381 3893 14415 3927
rect 14657 3893 14691 3927
rect 14933 3893 14967 3927
rect 16773 3893 16807 3927
rect 16957 3893 16991 3927
rect 1409 3689 1443 3723
rect 7481 3689 7515 3723
rect 8585 3689 8619 3723
rect 9137 3689 9171 3723
rect 10885 3689 10919 3723
rect 13829 3689 13863 3723
rect 15853 3689 15887 3723
rect 16313 3689 16347 3723
rect 16681 3689 16715 3723
rect 16773 3689 16807 3723
rect 17509 3689 17543 3723
rect 2544 3621 2578 3655
rect 4077 3621 4111 3655
rect 4874 3621 4908 3655
rect 8677 3621 8711 3655
rect 11222 3621 11256 3655
rect 12716 3621 12750 3655
rect 14933 3621 14967 3655
rect 17969 3621 18003 3655
rect 18337 3621 18371 3655
rect 2789 3553 2823 3587
rect 3341 3553 3375 3587
rect 4261 3553 4295 3587
rect 4445 3553 4479 3587
rect 6357 3553 6391 3587
rect 7757 3553 7791 3587
rect 8033 3553 8067 3587
rect 10261 3553 10295 3587
rect 14105 3553 14139 3587
rect 14565 3553 14599 3587
rect 15025 3553 15059 3587
rect 15945 3553 15979 3587
rect 17325 3553 17359 3587
rect 17601 3553 17635 3587
rect 18153 3553 18187 3587
rect 3065 3485 3099 3519
rect 3249 3485 3283 3519
rect 4629 3485 4663 3519
rect 6101 3485 6135 3519
rect 8861 3485 8895 3519
rect 10517 3485 10551 3519
rect 10984 3485 11018 3519
rect 12449 3485 12483 3519
rect 14749 3485 14783 3519
rect 16129 3485 16163 3519
rect 16865 3485 16899 3519
rect 12357 3417 12391 3451
rect 14381 3417 14415 3451
rect 15393 3417 15427 3451
rect 18521 3417 18555 3451
rect 3709 3349 3743 3383
rect 3985 3349 4019 3383
rect 6009 3349 6043 3383
rect 7573 3349 7607 3383
rect 7849 3349 7883 3383
rect 8217 3349 8251 3383
rect 13921 3349 13955 3383
rect 15485 3349 15519 3383
rect 17141 3349 17175 3383
rect 17785 3349 17819 3383
rect 1869 3145 1903 3179
rect 2237 3145 2271 3179
rect 4077 3145 4111 3179
rect 12541 3145 12575 3179
rect 15301 3145 15335 3179
rect 1409 3077 1443 3111
rect 17049 3077 17083 3111
rect 2513 3009 2547 3043
rect 4537 3009 4571 3043
rect 4629 3009 4663 3043
rect 4905 3009 4939 3043
rect 5733 3009 5767 3043
rect 6561 3009 6595 3043
rect 7573 3009 7607 3043
rect 8309 3009 8343 3043
rect 8493 3009 8527 3043
rect 9597 3009 9631 3043
rect 10517 3009 10551 3043
rect 11253 3009 11287 3043
rect 11805 3009 11839 3043
rect 13093 3009 13127 3043
rect 15761 3009 15795 3043
rect 15945 3009 15979 3043
rect 1961 2941 1995 2975
rect 2329 2941 2363 2975
rect 2697 2941 2731 2975
rect 2881 2941 2915 2975
rect 3433 2941 3467 2975
rect 3801 2941 3835 2975
rect 4445 2941 4479 2975
rect 6193 2941 6227 2975
rect 6745 2941 6779 2975
rect 7113 2941 7147 2975
rect 12081 2941 12115 2975
rect 13645 2941 13679 2975
rect 14105 2941 14139 2975
rect 14381 2941 14415 2975
rect 14749 2941 14783 2975
rect 15117 2941 15151 2975
rect 15669 2941 15703 2975
rect 16313 2941 16347 2975
rect 16773 2941 16807 2975
rect 17233 2941 17267 2975
rect 17601 2941 17635 2975
rect 17969 2941 18003 2975
rect 18337 2941 18371 2975
rect 1593 2873 1627 2907
rect 3065 2873 3099 2907
rect 5457 2873 5491 2907
rect 5917 2873 5951 2907
rect 7297 2873 7331 2907
rect 8585 2873 8619 2907
rect 9413 2873 9447 2907
rect 11069 2873 11103 2907
rect 11989 2873 12023 2907
rect 12909 2873 12943 2907
rect 13829 2873 13863 2907
rect 17785 2873 17819 2907
rect 18153 2873 18187 2907
rect 3341 2805 3375 2839
rect 3709 2805 3743 2839
rect 5089 2805 5123 2839
rect 5549 2805 5583 2839
rect 6837 2805 6871 2839
rect 7665 2805 7699 2839
rect 7757 2805 7791 2839
rect 8125 2805 8159 2839
rect 8953 2805 8987 2839
rect 9045 2805 9079 2839
rect 9505 2805 9539 2839
rect 9873 2805 9907 2839
rect 10241 2805 10275 2839
rect 10333 2805 10367 2839
rect 10701 2805 10735 2839
rect 11161 2805 11195 2839
rect 12449 2805 12483 2839
rect 13001 2805 13035 2839
rect 13461 2805 13495 2839
rect 13921 2805 13955 2839
rect 14197 2805 14231 2839
rect 14565 2805 14599 2839
rect 14933 2805 14967 2839
rect 16129 2805 16163 2839
rect 16405 2805 16439 2839
rect 16589 2805 16623 2839
rect 17325 2805 17359 2839
rect 18429 2805 18463 2839
rect 2605 2601 2639 2635
rect 2973 2601 3007 2635
rect 4445 2601 4479 2635
rect 4813 2601 4847 2635
rect 5733 2601 5767 2635
rect 7481 2601 7515 2635
rect 7849 2601 7883 2635
rect 8309 2601 8343 2635
rect 8769 2601 8803 2635
rect 9321 2601 9355 2635
rect 11621 2601 11655 2635
rect 12265 2601 12299 2635
rect 12633 2601 12667 2635
rect 15301 2601 15335 2635
rect 16313 2601 16347 2635
rect 18153 2601 18187 2635
rect 1961 2533 1995 2567
rect 3617 2533 3651 2567
rect 4905 2533 4939 2567
rect 5457 2533 5491 2567
rect 9781 2533 9815 2567
rect 11437 2533 11471 2567
rect 12909 2533 12943 2567
rect 13277 2533 13311 2567
rect 14105 2533 14139 2567
rect 15025 2533 15059 2567
rect 15945 2533 15979 2567
rect 16497 2533 16531 2567
rect 16865 2533 16899 2567
rect 17325 2533 17359 2567
rect 17785 2533 17819 2567
rect 18337 2533 18371 2567
rect 1593 2465 1627 2499
rect 2329 2465 2363 2499
rect 2697 2465 2731 2499
rect 3249 2465 3283 2499
rect 4169 2465 4203 2499
rect 6009 2465 6043 2499
rect 6377 2465 6411 2499
rect 6929 2465 6963 2499
rect 7205 2465 7239 2499
rect 8677 2465 8711 2499
rect 9873 2465 9907 2499
rect 10609 2465 10643 2499
rect 12173 2465 12207 2499
rect 13461 2465 13495 2499
rect 13645 2465 13679 2499
rect 14749 2465 14783 2499
rect 15485 2465 15519 2499
rect 16129 2465 16163 2499
rect 17969 2465 18003 2499
rect 1777 2397 1811 2431
rect 4997 2397 5031 2431
rect 7941 2397 7975 2431
rect 8125 2397 8159 2431
rect 8953 2397 8987 2431
rect 10057 2397 10091 2431
rect 10701 2397 10735 2431
rect 10793 2397 10827 2431
rect 11989 2397 12023 2431
rect 1409 2329 1443 2363
rect 2145 2329 2179 2363
rect 3065 2329 3099 2363
rect 3433 2329 3467 2363
rect 3985 2329 4019 2363
rect 5825 2329 5859 2363
rect 6193 2329 6227 2363
rect 6745 2329 6779 2363
rect 7389 2329 7423 2363
rect 9413 2329 9447 2363
rect 10241 2329 10275 2363
rect 11253 2329 11287 2363
rect 12725 2329 12759 2363
rect 13093 2329 13127 2363
rect 13921 2329 13955 2363
rect 14565 2329 14599 2363
rect 14841 2329 14875 2363
rect 15761 2329 15795 2363
rect 16681 2329 16715 2363
rect 17049 2329 17083 2363
rect 17601 2329 17635 2363
rect 18521 2329 18555 2363
rect 5365 2261 5399 2295
rect 6653 2261 6687 2295
rect 11161 2261 11195 2295
rect 14289 2261 14323 2295
rect 15577 2261 15611 2295
rect 17417 2261 17451 2295
<< metal1 >>
rect 1486 14764 1492 14816
rect 1544 14804 1550 14816
rect 2958 14804 2964 14816
rect 1544 14776 2964 14804
rect 1544 14764 1550 14776
rect 2958 14764 2964 14776
rect 3016 14764 3022 14816
rect 11882 14764 11888 14816
rect 11940 14804 11946 14816
rect 17494 14804 17500 14816
rect 11940 14776 17500 14804
rect 11940 14764 11946 14776
rect 17494 14764 17500 14776
rect 17552 14764 17558 14816
rect 1104 14714 18860 14736
rect 1104 14662 6912 14714
rect 6964 14662 6976 14714
rect 7028 14662 7040 14714
rect 7092 14662 7104 14714
rect 7156 14662 12843 14714
rect 12895 14662 12907 14714
rect 12959 14662 12971 14714
rect 13023 14662 13035 14714
rect 13087 14662 18860 14714
rect 1104 14640 18860 14662
rect 1854 14600 1860 14612
rect 1815 14572 1860 14600
rect 1854 14560 1860 14572
rect 1912 14560 1918 14612
rect 2222 14600 2228 14612
rect 2183 14572 2228 14600
rect 2222 14560 2228 14572
rect 2280 14560 2286 14612
rect 2774 14560 2780 14612
rect 2832 14600 2838 14612
rect 3605 14603 3663 14609
rect 3605 14600 3617 14603
rect 2832 14572 3617 14600
rect 2832 14560 2838 14572
rect 3605 14569 3617 14572
rect 3651 14569 3663 14603
rect 4430 14600 4436 14612
rect 4343 14572 4436 14600
rect 3605 14563 3663 14569
rect 4430 14560 4436 14572
rect 4488 14600 4494 14612
rect 14458 14600 14464 14612
rect 4488 14572 14464 14600
rect 4488 14560 4494 14572
rect 14458 14560 14464 14572
rect 14516 14560 14522 14612
rect 16301 14603 16359 14609
rect 16301 14569 16313 14603
rect 16347 14600 16359 14603
rect 17862 14600 17868 14612
rect 16347 14572 17868 14600
rect 16347 14569 16359 14572
rect 16301 14563 16359 14569
rect 17862 14560 17868 14572
rect 17920 14560 17926 14612
rect 1486 14532 1492 14544
rect 1447 14504 1492 14532
rect 1486 14492 1492 14504
rect 1544 14492 1550 14544
rect 2038 14492 2044 14544
rect 2096 14532 2102 14544
rect 3326 14532 3332 14544
rect 2096 14504 3332 14532
rect 2096 14492 2102 14504
rect 1949 14467 2007 14473
rect 1949 14433 1961 14467
rect 1995 14433 2007 14467
rect 2314 14464 2320 14476
rect 2275 14436 2320 14464
rect 1949 14427 2007 14433
rect 1964 14396 1992 14427
rect 2314 14424 2320 14436
rect 2372 14424 2378 14476
rect 2682 14464 2688 14476
rect 2643 14436 2688 14464
rect 2682 14424 2688 14436
rect 2740 14424 2746 14476
rect 2792 14473 2820 14504
rect 3326 14492 3332 14504
rect 3384 14492 3390 14544
rect 4154 14492 4160 14544
rect 4212 14532 4218 14544
rect 4893 14535 4951 14541
rect 4893 14532 4905 14535
rect 4212 14504 4905 14532
rect 4212 14492 4218 14504
rect 2777 14467 2835 14473
rect 2777 14433 2789 14467
rect 2823 14433 2835 14467
rect 3050 14464 3056 14476
rect 3011 14436 3056 14464
rect 2777 14427 2835 14433
rect 3050 14424 3056 14436
rect 3108 14424 3114 14476
rect 3510 14464 3516 14476
rect 3471 14436 3516 14464
rect 3510 14424 3516 14436
rect 3568 14424 3574 14476
rect 3878 14464 3884 14476
rect 3839 14436 3884 14464
rect 3878 14424 3884 14436
rect 3936 14424 3942 14476
rect 4246 14424 4252 14476
rect 4304 14464 4310 14476
rect 4632 14473 4660 14504
rect 4893 14501 4905 14504
rect 4939 14501 4951 14535
rect 5902 14532 5908 14544
rect 5863 14504 5908 14532
rect 4893 14495 4951 14501
rect 5902 14492 5908 14504
rect 5960 14492 5966 14544
rect 9858 14532 9864 14544
rect 9819 14504 9864 14532
rect 9858 14492 9864 14504
rect 9916 14492 9922 14544
rect 16025 14535 16083 14541
rect 16025 14501 16037 14535
rect 16071 14532 16083 14535
rect 17494 14532 17500 14544
rect 16071 14504 17356 14532
rect 17455 14504 17500 14532
rect 16071 14501 16083 14504
rect 16025 14495 16083 14501
rect 4341 14467 4399 14473
rect 4341 14464 4353 14467
rect 4304 14436 4353 14464
rect 4304 14424 4310 14436
rect 4341 14433 4353 14436
rect 4387 14433 4399 14467
rect 4341 14427 4399 14433
rect 4617 14467 4675 14473
rect 4617 14433 4629 14467
rect 4663 14433 4675 14467
rect 6086 14464 6092 14476
rect 6047 14436 6092 14464
rect 4617 14427 4675 14433
rect 6086 14424 6092 14436
rect 6144 14424 6150 14476
rect 9766 14424 9772 14476
rect 9824 14464 9830 14476
rect 10045 14467 10103 14473
rect 10045 14464 10057 14467
rect 9824 14436 10057 14464
rect 9824 14424 9830 14436
rect 10045 14433 10057 14436
rect 10091 14433 10103 14467
rect 16114 14464 16120 14476
rect 16075 14436 16120 14464
rect 10045 14427 10103 14433
rect 16114 14424 16120 14436
rect 16172 14424 16178 14476
rect 16482 14424 16488 14476
rect 16540 14464 16546 14476
rect 16577 14467 16635 14473
rect 16577 14464 16589 14467
rect 16540 14436 16589 14464
rect 16540 14424 16546 14436
rect 16577 14433 16589 14436
rect 16623 14433 16635 14467
rect 16942 14464 16948 14476
rect 16903 14436 16948 14464
rect 16577 14427 16635 14433
rect 16942 14424 16948 14436
rect 17000 14424 17006 14476
rect 17221 14467 17279 14473
rect 17221 14433 17233 14467
rect 17267 14433 17279 14467
rect 17328 14464 17356 14504
rect 17494 14492 17500 14504
rect 17552 14492 17558 14544
rect 17678 14532 17684 14544
rect 17639 14504 17684 14532
rect 17678 14492 17684 14504
rect 17736 14492 17742 14544
rect 18138 14464 18144 14476
rect 17328 14436 17632 14464
rect 18099 14436 18144 14464
rect 17221 14427 17279 14433
rect 2498 14396 2504 14408
rect 1964 14368 2504 14396
rect 2498 14356 2504 14368
rect 2556 14356 2562 14408
rect 17236 14396 17264 14427
rect 2976 14368 17264 14396
rect 17604 14396 17632 14436
rect 18138 14424 18144 14436
rect 18196 14424 18202 14476
rect 18414 14464 18420 14476
rect 18375 14436 18420 14464
rect 18414 14424 18420 14436
rect 18472 14424 18478 14476
rect 18432 14396 18460 14424
rect 17604 14368 18460 14396
rect 1673 14331 1731 14337
rect 1673 14297 1685 14331
rect 1719 14328 1731 14331
rect 2866 14328 2872 14340
rect 1719 14300 2872 14328
rect 1719 14297 1731 14300
rect 1673 14291 1731 14297
rect 2866 14288 2872 14300
rect 2924 14288 2930 14340
rect 2976 14337 3004 14368
rect 2961 14331 3019 14337
rect 2961 14297 2973 14331
rect 3007 14297 3019 14331
rect 2961 14291 3019 14297
rect 3237 14331 3295 14337
rect 3237 14297 3249 14331
rect 3283 14328 3295 14331
rect 9582 14328 9588 14340
rect 3283 14300 9588 14328
rect 3283 14297 3295 14300
rect 3237 14291 3295 14297
rect 9582 14288 9588 14300
rect 9640 14328 9646 14340
rect 9640 14300 12434 14328
rect 9640 14288 9646 14300
rect 2038 14220 2044 14272
rect 2096 14260 2102 14272
rect 2501 14263 2559 14269
rect 2501 14260 2513 14263
rect 2096 14232 2513 14260
rect 2096 14220 2102 14232
rect 2501 14229 2513 14232
rect 2547 14229 2559 14263
rect 2501 14223 2559 14229
rect 3329 14263 3387 14269
rect 3329 14229 3341 14263
rect 3375 14260 3387 14263
rect 3418 14260 3424 14272
rect 3375 14232 3424 14260
rect 3375 14229 3387 14232
rect 3329 14223 3387 14229
rect 3418 14220 3424 14232
rect 3476 14220 3482 14272
rect 3786 14220 3792 14272
rect 3844 14260 3850 14272
rect 4065 14263 4123 14269
rect 4065 14260 4077 14263
rect 3844 14232 4077 14260
rect 3844 14220 3850 14232
rect 4065 14229 4077 14232
rect 4111 14229 4123 14263
rect 4065 14223 4123 14229
rect 4157 14263 4215 14269
rect 4157 14229 4169 14263
rect 4203 14260 4215 14263
rect 4246 14260 4252 14272
rect 4203 14232 4252 14260
rect 4203 14229 4215 14232
rect 4157 14223 4215 14229
rect 4246 14220 4252 14232
rect 4304 14220 4310 14272
rect 4338 14220 4344 14272
rect 4396 14260 4402 14272
rect 4709 14263 4767 14269
rect 4709 14260 4721 14263
rect 4396 14232 4721 14260
rect 4396 14220 4402 14232
rect 4709 14229 4721 14232
rect 4755 14229 4767 14263
rect 12406 14260 12434 14300
rect 15378 14288 15384 14340
rect 15436 14328 15442 14340
rect 16393 14331 16451 14337
rect 16393 14328 16405 14331
rect 15436 14300 16405 14328
rect 15436 14288 15442 14300
rect 16393 14297 16405 14300
rect 16439 14297 16451 14331
rect 16393 14291 16451 14297
rect 16574 14288 16580 14340
rect 16632 14328 16638 14340
rect 16761 14331 16819 14337
rect 16761 14328 16773 14331
rect 16632 14300 16773 14328
rect 16632 14288 16638 14300
rect 16761 14297 16773 14300
rect 16807 14297 16819 14331
rect 17494 14328 17500 14340
rect 16761 14291 16819 14297
rect 16868 14300 17500 14328
rect 16868 14260 16896 14300
rect 17494 14288 17500 14300
rect 17552 14288 17558 14340
rect 17957 14331 18015 14337
rect 17957 14297 17969 14331
rect 18003 14328 18015 14331
rect 18506 14328 18512 14340
rect 18003 14300 18512 14328
rect 18003 14297 18015 14300
rect 17957 14291 18015 14297
rect 18506 14288 18512 14300
rect 18564 14288 18570 14340
rect 17402 14260 17408 14272
rect 12406 14232 16896 14260
rect 17363 14232 17408 14260
rect 4709 14223 4767 14229
rect 17402 14220 17408 14232
rect 17460 14220 17466 14272
rect 18322 14260 18328 14272
rect 18283 14232 18328 14260
rect 18322 14220 18328 14232
rect 18380 14220 18386 14272
rect 1104 14170 18860 14192
rect 1104 14118 3947 14170
rect 3999 14118 4011 14170
rect 4063 14118 4075 14170
rect 4127 14118 4139 14170
rect 4191 14118 9878 14170
rect 9930 14118 9942 14170
rect 9994 14118 10006 14170
rect 10058 14118 10070 14170
rect 10122 14118 15808 14170
rect 15860 14118 15872 14170
rect 15924 14118 15936 14170
rect 15988 14118 16000 14170
rect 16052 14118 18860 14170
rect 1104 14096 18860 14118
rect 1854 14056 1860 14068
rect 1815 14028 1860 14056
rect 1854 14016 1860 14028
rect 1912 14016 1918 14068
rect 2314 14016 2320 14068
rect 2372 14056 2378 14068
rect 2777 14059 2835 14065
rect 2777 14056 2789 14059
rect 2372 14028 2789 14056
rect 2372 14016 2378 14028
rect 2777 14025 2789 14028
rect 2823 14025 2835 14059
rect 2777 14019 2835 14025
rect 2866 14016 2872 14068
rect 2924 14056 2930 14068
rect 9766 14056 9772 14068
rect 2924 14028 6914 14056
rect 9727 14028 9772 14056
rect 2924 14016 2930 14028
rect 2130 13988 2136 14000
rect 2091 13960 2136 13988
rect 2130 13948 2136 13960
rect 2188 13948 2194 14000
rect 2498 13988 2504 14000
rect 2459 13960 2504 13988
rect 2498 13948 2504 13960
rect 2556 13948 2562 14000
rect 3053 13991 3111 13997
rect 3053 13957 3065 13991
rect 3099 13957 3111 13991
rect 3326 13988 3332 14000
rect 3287 13960 3332 13988
rect 3053 13951 3111 13957
rect 3068 13920 3096 13951
rect 3326 13948 3332 13960
rect 3384 13948 3390 14000
rect 3694 13948 3700 14000
rect 3752 13988 3758 14000
rect 3881 13991 3939 13997
rect 3881 13988 3893 13991
rect 3752 13960 3893 13988
rect 3752 13948 3758 13960
rect 3881 13957 3893 13960
rect 3927 13957 3939 13991
rect 3881 13951 3939 13957
rect 4157 13991 4215 13997
rect 4157 13957 4169 13991
rect 4203 13988 4215 13991
rect 4430 13988 4436 14000
rect 4203 13960 4436 13988
rect 4203 13957 4215 13960
rect 4157 13951 4215 13957
rect 2332 13892 3096 13920
rect 1394 13852 1400 13864
rect 1355 13824 1400 13852
rect 1394 13812 1400 13824
rect 1452 13812 1458 13864
rect 2332 13861 2360 13892
rect 3142 13880 3148 13932
rect 3200 13920 3206 13932
rect 3513 13923 3571 13929
rect 3513 13920 3525 13923
rect 3200 13892 3525 13920
rect 3200 13880 3206 13892
rect 3513 13889 3525 13892
rect 3559 13889 3571 13923
rect 3513 13883 3571 13889
rect 3602 13880 3608 13932
rect 3660 13920 3666 13932
rect 3789 13923 3847 13929
rect 3789 13920 3801 13923
rect 3660 13892 3801 13920
rect 3660 13880 3666 13892
rect 3789 13889 3801 13892
rect 3835 13889 3847 13923
rect 3789 13883 3847 13889
rect 2317 13855 2375 13861
rect 2317 13821 2329 13855
rect 2363 13821 2375 13855
rect 2317 13815 2375 13821
rect 2685 13855 2743 13861
rect 2685 13821 2697 13855
rect 2731 13852 2743 13855
rect 2961 13855 3019 13861
rect 2731 13824 2912 13852
rect 2731 13821 2743 13824
rect 2685 13815 2743 13821
rect 1578 13784 1584 13796
rect 1539 13756 1584 13784
rect 1578 13744 1584 13756
rect 1636 13744 1642 13796
rect 1946 13784 1952 13796
rect 1907 13756 1952 13784
rect 1946 13744 1952 13756
rect 2004 13744 2010 13796
rect 2884 13716 2912 13824
rect 2961 13821 2973 13855
rect 3007 13821 3019 13855
rect 2961 13815 3019 13821
rect 3237 13855 3295 13861
rect 3237 13821 3249 13855
rect 3283 13852 3295 13855
rect 4172 13852 4200 13951
rect 4430 13948 4436 13960
rect 4488 13948 4494 14000
rect 6886 13988 6914 14028
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 13906 14016 13912 14068
rect 13964 14056 13970 14068
rect 15010 14056 15016 14068
rect 13964 14028 15016 14056
rect 13964 14016 13970 14028
rect 15010 14016 15016 14028
rect 15068 14056 15074 14068
rect 15381 14059 15439 14065
rect 15381 14056 15393 14059
rect 15068 14028 15393 14056
rect 15068 14016 15074 14028
rect 15381 14025 15393 14028
rect 15427 14025 15439 14059
rect 15381 14019 15439 14025
rect 16393 14059 16451 14065
rect 16393 14025 16405 14059
rect 16439 14056 16451 14059
rect 16482 14056 16488 14068
rect 16439 14028 16488 14056
rect 16439 14025 16451 14028
rect 16393 14019 16451 14025
rect 15286 13988 15292 14000
rect 6886 13960 15292 13988
rect 15286 13948 15292 13960
rect 15344 13948 15350 14000
rect 9582 13852 9588 13864
rect 3283 13824 4200 13852
rect 9543 13824 9588 13852
rect 3283 13821 3295 13824
rect 3237 13815 3295 13821
rect 2976 13784 3004 13815
rect 9582 13812 9588 13824
rect 9640 13812 9646 13864
rect 15396 13852 15424 14019
rect 16482 14016 16488 14028
rect 16540 14016 16546 14068
rect 16761 14059 16819 14065
rect 16761 14025 16773 14059
rect 16807 14056 16819 14059
rect 18138 14056 18144 14068
rect 16807 14028 18144 14056
rect 16807 14025 16819 14028
rect 16761 14019 16819 14025
rect 18138 14016 18144 14028
rect 18196 14016 18202 14068
rect 16577 13991 16635 13997
rect 16577 13957 16589 13991
rect 16623 13988 16635 13991
rect 16942 13988 16948 14000
rect 16623 13960 16948 13988
rect 16623 13957 16635 13960
rect 16577 13951 16635 13957
rect 16942 13948 16948 13960
rect 17000 13948 17006 14000
rect 17218 13948 17224 14000
rect 17276 13988 17282 14000
rect 17770 13988 17776 14000
rect 17276 13960 17776 13988
rect 17276 13948 17282 13960
rect 17770 13948 17776 13960
rect 17828 13948 17834 14000
rect 15841 13923 15899 13929
rect 15841 13889 15853 13923
rect 15887 13920 15899 13923
rect 16114 13920 16120 13932
rect 15887 13892 16120 13920
rect 15887 13889 15899 13892
rect 15841 13883 15899 13889
rect 16114 13880 16120 13892
rect 16172 13880 16178 13932
rect 17037 13923 17095 13929
rect 17037 13889 17049 13923
rect 17083 13920 17095 13923
rect 17083 13892 17632 13920
rect 17083 13889 17095 13892
rect 17037 13883 17095 13889
rect 15565 13855 15623 13861
rect 15565 13852 15577 13855
rect 15396 13824 15577 13852
rect 15565 13821 15577 13824
rect 15611 13821 15623 13855
rect 16206 13852 16212 13864
rect 16167 13824 16212 13852
rect 15565 13815 15623 13821
rect 16206 13812 16212 13824
rect 16264 13852 16270 13864
rect 17126 13852 17132 13864
rect 16264 13824 16988 13852
rect 17087 13824 17132 13852
rect 16264 13812 16270 13824
rect 3786 13784 3792 13796
rect 2976 13756 3792 13784
rect 3786 13744 3792 13756
rect 3844 13744 3850 13796
rect 16960 13784 16988 13824
rect 17126 13812 17132 13824
rect 17184 13812 17190 13864
rect 17604 13852 17632 13892
rect 17678 13880 17684 13932
rect 17736 13920 17742 13932
rect 17865 13923 17923 13929
rect 17865 13920 17877 13923
rect 17736 13892 17877 13920
rect 17736 13880 17742 13892
rect 17865 13889 17877 13892
rect 17911 13889 17923 13923
rect 17865 13883 17923 13889
rect 17954 13880 17960 13932
rect 18012 13920 18018 13932
rect 18233 13923 18291 13929
rect 18233 13920 18245 13923
rect 18012 13892 18245 13920
rect 18012 13880 18018 13892
rect 18233 13889 18245 13892
rect 18279 13889 18291 13923
rect 18233 13883 18291 13889
rect 18414 13852 18420 13864
rect 17236 13824 17540 13852
rect 17604 13824 18420 13852
rect 17236 13784 17264 13824
rect 16960 13756 17264 13784
rect 17310 13744 17316 13796
rect 17368 13784 17374 13796
rect 17512 13784 17540 13824
rect 18414 13812 18420 13824
rect 18472 13812 18478 13864
rect 17681 13787 17739 13793
rect 17681 13784 17693 13787
rect 17368 13756 17413 13784
rect 17512 13756 17693 13784
rect 17368 13744 17374 13756
rect 17681 13753 17693 13756
rect 17727 13753 17739 13787
rect 17681 13747 17739 13753
rect 17770 13744 17776 13796
rect 17828 13784 17834 13796
rect 18049 13787 18107 13793
rect 18049 13784 18061 13787
rect 17828 13756 18061 13784
rect 17828 13744 17834 13756
rect 18049 13753 18061 13756
rect 18095 13753 18107 13787
rect 18049 13747 18107 13753
rect 3418 13716 3424 13728
rect 2884 13688 3424 13716
rect 3418 13676 3424 13688
rect 3476 13676 3482 13728
rect 16298 13676 16304 13728
rect 16356 13716 16362 13728
rect 17589 13719 17647 13725
rect 17589 13716 17601 13719
rect 16356 13688 17601 13716
rect 16356 13676 16362 13688
rect 17589 13685 17601 13688
rect 17635 13685 17647 13719
rect 17589 13679 17647 13685
rect 1104 13626 18860 13648
rect 1104 13574 6912 13626
rect 6964 13574 6976 13626
rect 7028 13574 7040 13626
rect 7092 13574 7104 13626
rect 7156 13574 12843 13626
rect 12895 13574 12907 13626
rect 12959 13574 12971 13626
rect 13023 13574 13035 13626
rect 13087 13574 18860 13626
rect 1104 13552 18860 13574
rect 1578 13472 1584 13524
rect 1636 13512 1642 13524
rect 1765 13515 1823 13521
rect 1765 13512 1777 13515
rect 1636 13484 1777 13512
rect 1636 13472 1642 13484
rect 1765 13481 1777 13484
rect 1811 13481 1823 13515
rect 1765 13475 1823 13481
rect 1946 13472 1952 13524
rect 2004 13512 2010 13524
rect 2409 13515 2467 13521
rect 2409 13512 2421 13515
rect 2004 13484 2421 13512
rect 2004 13472 2010 13484
rect 2409 13481 2421 13484
rect 2455 13481 2467 13515
rect 2958 13512 2964 13524
rect 2919 13484 2964 13512
rect 2409 13475 2467 13481
rect 2958 13472 2964 13484
rect 3016 13472 3022 13524
rect 6086 13512 6092 13524
rect 6047 13484 6092 13512
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 14274 13472 14280 13524
rect 14332 13512 14338 13524
rect 16390 13512 16396 13524
rect 14332 13484 16396 13512
rect 14332 13472 14338 13484
rect 16390 13472 16396 13484
rect 16448 13472 16454 13524
rect 17129 13515 17187 13521
rect 17129 13481 17141 13515
rect 17175 13512 17187 13515
rect 17218 13512 17224 13524
rect 17175 13484 17224 13512
rect 17175 13481 17187 13484
rect 17129 13475 17187 13481
rect 17218 13472 17224 13484
rect 17276 13472 17282 13524
rect 17313 13515 17371 13521
rect 17313 13481 17325 13515
rect 17359 13512 17371 13515
rect 17586 13512 17592 13524
rect 17359 13484 17592 13512
rect 17359 13481 17371 13484
rect 17313 13475 17371 13481
rect 17586 13472 17592 13484
rect 17644 13472 17650 13524
rect 17770 13472 17776 13524
rect 17828 13512 17834 13524
rect 17957 13515 18015 13521
rect 17957 13512 17969 13515
rect 17828 13484 17969 13512
rect 17828 13472 17834 13484
rect 17957 13481 17969 13484
rect 18003 13512 18015 13515
rect 18230 13512 18236 13524
rect 18003 13484 18236 13512
rect 18003 13481 18015 13484
rect 17957 13475 18015 13481
rect 18230 13472 18236 13484
rect 18288 13472 18294 13524
rect 2685 13447 2743 13453
rect 2685 13444 2697 13447
rect 1504 13416 2697 13444
rect 1504 13388 1532 13416
rect 2685 13413 2697 13416
rect 2731 13413 2743 13447
rect 2685 13407 2743 13413
rect 3786 13404 3792 13456
rect 3844 13444 3850 13456
rect 17497 13447 17555 13453
rect 3844 13416 6914 13444
rect 3844 13404 3850 13416
rect 1486 13376 1492 13388
rect 1447 13348 1492 13376
rect 1486 13336 1492 13348
rect 1544 13336 1550 13388
rect 1949 13379 2007 13385
rect 1949 13345 1961 13379
rect 1995 13376 2007 13379
rect 2038 13376 2044 13388
rect 1995 13348 2044 13376
rect 1995 13345 2007 13348
rect 1949 13339 2007 13345
rect 2038 13336 2044 13348
rect 2096 13336 2102 13388
rect 2133 13379 2191 13385
rect 2133 13345 2145 13379
rect 2179 13376 2191 13379
rect 2593 13379 2651 13385
rect 2593 13376 2605 13379
rect 2179 13348 2605 13376
rect 2179 13345 2191 13348
rect 2133 13339 2191 13345
rect 2593 13345 2605 13348
rect 2639 13376 2651 13379
rect 4246 13376 4252 13388
rect 2639 13348 4252 13376
rect 2639 13345 2651 13348
rect 2593 13339 2651 13345
rect 4246 13336 4252 13348
rect 4304 13336 4310 13388
rect 6178 13336 6184 13388
rect 6236 13376 6242 13388
rect 6273 13379 6331 13385
rect 6273 13376 6285 13379
rect 6236 13348 6285 13376
rect 6236 13336 6242 13348
rect 6273 13345 6285 13348
rect 6319 13345 6331 13379
rect 6886 13376 6914 13416
rect 17497 13413 17509 13447
rect 17543 13444 17555 13447
rect 18414 13444 18420 13456
rect 17543 13416 18420 13444
rect 17543 13413 17555 13416
rect 17497 13407 17555 13413
rect 18414 13404 18420 13416
rect 18472 13404 18478 13456
rect 17773 13379 17831 13385
rect 17773 13376 17785 13379
rect 6886 13348 17785 13376
rect 6273 13339 6331 13345
rect 17773 13345 17785 13348
rect 17819 13345 17831 13379
rect 18046 13376 18052 13388
rect 18007 13348 18052 13376
rect 17773 13339 17831 13345
rect 18046 13336 18052 13348
rect 18104 13336 18110 13388
rect 16117 13311 16175 13317
rect 16117 13308 16129 13311
rect 6886 13280 16129 13308
rect 2317 13243 2375 13249
rect 2317 13209 2329 13243
rect 2363 13240 2375 13243
rect 6886 13240 6914 13280
rect 16117 13277 16129 13280
rect 16163 13308 16175 13311
rect 16390 13308 16396 13320
rect 16163 13280 16396 13308
rect 16163 13277 16175 13280
rect 16117 13271 16175 13277
rect 16390 13268 16396 13280
rect 16448 13268 16454 13320
rect 16577 13311 16635 13317
rect 16577 13277 16589 13311
rect 16623 13308 16635 13311
rect 16666 13308 16672 13320
rect 16623 13280 16672 13308
rect 16623 13277 16635 13280
rect 16577 13271 16635 13277
rect 16666 13268 16672 13280
rect 16724 13268 16730 13320
rect 16761 13311 16819 13317
rect 16761 13277 16773 13311
rect 16807 13308 16819 13311
rect 18064 13308 18092 13336
rect 16807 13280 18092 13308
rect 16807 13277 16819 13280
rect 16761 13271 16819 13277
rect 2363 13212 6914 13240
rect 2363 13209 2375 13212
rect 2317 13203 2375 13209
rect 16942 13200 16948 13252
rect 17000 13240 17006 13252
rect 18233 13243 18291 13249
rect 18233 13240 18245 13243
rect 17000 13212 18245 13240
rect 17000 13200 17006 13212
rect 18233 13209 18245 13212
rect 18279 13209 18291 13243
rect 18233 13203 18291 13209
rect 1581 13175 1639 13181
rect 1581 13141 1593 13175
rect 1627 13172 1639 13175
rect 7834 13172 7840 13184
rect 1627 13144 7840 13172
rect 1627 13141 1639 13144
rect 1581 13135 1639 13141
rect 7834 13132 7840 13144
rect 7892 13132 7898 13184
rect 16853 13175 16911 13181
rect 16853 13141 16865 13175
rect 16899 13172 16911 13175
rect 17310 13172 17316 13184
rect 16899 13144 17316 13172
rect 16899 13141 16911 13144
rect 16853 13135 16911 13141
rect 17310 13132 17316 13144
rect 17368 13132 17374 13184
rect 17586 13172 17592 13184
rect 17547 13144 17592 13172
rect 17586 13132 17592 13144
rect 17644 13132 17650 13184
rect 1104 13082 18860 13104
rect 1104 13030 3947 13082
rect 3999 13030 4011 13082
rect 4063 13030 4075 13082
rect 4127 13030 4139 13082
rect 4191 13030 9878 13082
rect 9930 13030 9942 13082
rect 9994 13030 10006 13082
rect 10058 13030 10070 13082
rect 10122 13030 15808 13082
rect 15860 13030 15872 13082
rect 15924 13030 15936 13082
rect 15988 13030 16000 13082
rect 16052 13030 18860 13082
rect 1104 13008 18860 13030
rect 1949 12971 2007 12977
rect 1949 12937 1961 12971
rect 1995 12968 2007 12971
rect 8478 12968 8484 12980
rect 1995 12940 8484 12968
rect 1995 12937 2007 12940
rect 1949 12931 2007 12937
rect 8478 12928 8484 12940
rect 8536 12928 8542 12980
rect 15286 12928 15292 12980
rect 15344 12968 15350 12980
rect 15473 12971 15531 12977
rect 15473 12968 15485 12971
rect 15344 12940 15485 12968
rect 15344 12928 15350 12940
rect 15473 12937 15485 12940
rect 15519 12968 15531 12971
rect 15562 12968 15568 12980
rect 15519 12940 15568 12968
rect 15519 12937 15531 12940
rect 15473 12931 15531 12937
rect 15562 12928 15568 12940
rect 15620 12968 15626 12980
rect 15657 12971 15715 12977
rect 15657 12968 15669 12971
rect 15620 12940 15669 12968
rect 15620 12928 15626 12940
rect 15657 12937 15669 12940
rect 15703 12937 15715 12971
rect 16298 12968 16304 12980
rect 16259 12940 16304 12968
rect 15657 12931 15715 12937
rect 16298 12928 16304 12940
rect 16356 12928 16362 12980
rect 16850 12928 16856 12980
rect 16908 12968 16914 12980
rect 18322 12968 18328 12980
rect 16908 12940 18328 12968
rect 16908 12928 16914 12940
rect 18322 12928 18328 12940
rect 18380 12928 18386 12980
rect 1673 12903 1731 12909
rect 1673 12869 1685 12903
rect 1719 12900 1731 12903
rect 5074 12900 5080 12912
rect 1719 12872 5080 12900
rect 1719 12869 1731 12872
rect 1673 12863 1731 12869
rect 5074 12860 5080 12872
rect 5132 12860 5138 12912
rect 9766 12860 9772 12912
rect 9824 12900 9830 12912
rect 10226 12900 10232 12912
rect 9824 12872 10232 12900
rect 9824 12860 9830 12872
rect 10226 12860 10232 12872
rect 10284 12900 10290 12912
rect 11514 12900 11520 12912
rect 10284 12872 11520 12900
rect 10284 12860 10290 12872
rect 11514 12860 11520 12872
rect 11572 12900 11578 12912
rect 12434 12900 12440 12912
rect 11572 12872 12440 12900
rect 11572 12860 11578 12872
rect 12434 12860 12440 12872
rect 12492 12900 12498 12912
rect 16316 12900 16344 12928
rect 12492 12872 16344 12900
rect 12492 12860 12498 12872
rect 17310 12860 17316 12912
rect 17368 12900 17374 12912
rect 17589 12903 17647 12909
rect 17589 12900 17601 12903
rect 17368 12872 17601 12900
rect 17368 12860 17374 12872
rect 17589 12869 17601 12872
rect 17635 12869 17647 12903
rect 17589 12863 17647 12869
rect 2501 12835 2559 12841
rect 2501 12832 2513 12835
rect 1504 12804 2513 12832
rect 1394 12656 1400 12708
rect 1452 12696 1458 12708
rect 1504 12705 1532 12804
rect 2501 12801 2513 12804
rect 2547 12801 2559 12835
rect 2501 12795 2559 12801
rect 15286 12792 15292 12844
rect 15344 12832 15350 12844
rect 16025 12835 16083 12841
rect 16025 12832 16037 12835
rect 15344 12804 16037 12832
rect 15344 12792 15350 12804
rect 16025 12801 16037 12804
rect 16071 12801 16083 12835
rect 16025 12795 16083 12801
rect 17037 12835 17095 12841
rect 17037 12801 17049 12835
rect 17083 12832 17095 12835
rect 17083 12804 18092 12832
rect 17083 12801 17095 12804
rect 17037 12795 17095 12801
rect 2685 12767 2743 12773
rect 2685 12764 2697 12767
rect 1872 12736 2697 12764
rect 1872 12708 1900 12736
rect 2685 12733 2697 12736
rect 2731 12733 2743 12767
rect 2685 12727 2743 12733
rect 3418 12724 3424 12776
rect 3476 12764 3482 12776
rect 17313 12767 17371 12773
rect 17313 12764 17325 12767
rect 3476 12736 17325 12764
rect 3476 12724 3482 12736
rect 17313 12733 17325 12736
rect 17359 12733 17371 12767
rect 17313 12727 17371 12733
rect 17494 12724 17500 12776
rect 17552 12764 17558 12776
rect 17773 12767 17831 12773
rect 17773 12764 17785 12767
rect 17552 12736 17785 12764
rect 17552 12724 17558 12736
rect 17773 12733 17785 12736
rect 17819 12733 17831 12767
rect 17773 12727 17831 12733
rect 18064 12708 18092 12804
rect 18414 12764 18420 12776
rect 18327 12736 18420 12764
rect 1489 12699 1547 12705
rect 1489 12696 1501 12699
rect 1452 12668 1501 12696
rect 1452 12656 1458 12668
rect 1489 12665 1501 12668
rect 1535 12665 1547 12699
rect 1854 12696 1860 12708
rect 1815 12668 1860 12696
rect 1489 12659 1547 12665
rect 1854 12656 1860 12668
rect 1912 12656 1918 12708
rect 2222 12696 2228 12708
rect 2183 12668 2228 12696
rect 2222 12656 2228 12668
rect 2280 12696 2286 12708
rect 2869 12699 2927 12705
rect 2869 12696 2881 12699
rect 2280 12668 2881 12696
rect 2280 12656 2286 12668
rect 2869 12665 2881 12668
rect 2915 12665 2927 12699
rect 2869 12659 2927 12665
rect 2958 12656 2964 12708
rect 3016 12696 3022 12708
rect 3145 12699 3203 12705
rect 3145 12696 3157 12699
rect 3016 12668 3157 12696
rect 3016 12656 3022 12668
rect 3145 12665 3157 12668
rect 3191 12696 3203 12699
rect 8110 12696 8116 12708
rect 3191 12668 8116 12696
rect 3191 12665 3203 12668
rect 3145 12659 3203 12665
rect 8110 12656 8116 12668
rect 8168 12656 8174 12708
rect 8849 12699 8907 12705
rect 8849 12665 8861 12699
rect 8895 12696 8907 12699
rect 10318 12696 10324 12708
rect 8895 12668 10324 12696
rect 8895 12665 8907 12668
rect 8849 12659 8907 12665
rect 10318 12656 10324 12668
rect 10376 12656 10382 12708
rect 14550 12656 14556 12708
rect 14608 12696 14614 12708
rect 16393 12699 16451 12705
rect 16393 12696 16405 12699
rect 14608 12668 16405 12696
rect 14608 12656 14614 12668
rect 16393 12665 16405 12668
rect 16439 12665 16451 12699
rect 16393 12659 16451 12665
rect 17221 12699 17279 12705
rect 17221 12665 17233 12699
rect 17267 12696 17279 12699
rect 17862 12696 17868 12708
rect 17267 12668 17724 12696
rect 17823 12668 17868 12696
rect 17267 12665 17279 12668
rect 17221 12659 17279 12665
rect 2130 12588 2136 12640
rect 2188 12628 2194 12640
rect 2317 12631 2375 12637
rect 2317 12628 2329 12631
rect 2188 12600 2329 12628
rect 2188 12588 2194 12600
rect 2317 12597 2329 12600
rect 2363 12597 2375 12631
rect 2317 12591 2375 12597
rect 3329 12631 3387 12637
rect 3329 12597 3341 12631
rect 3375 12628 3387 12631
rect 3602 12628 3608 12640
rect 3375 12600 3608 12628
rect 3375 12597 3387 12600
rect 3329 12591 3387 12597
rect 3602 12588 3608 12600
rect 3660 12588 3666 12640
rect 3789 12631 3847 12637
rect 3789 12597 3801 12631
rect 3835 12628 3847 12631
rect 4798 12628 4804 12640
rect 3835 12600 4804 12628
rect 3835 12597 3847 12600
rect 3789 12591 3847 12597
rect 4798 12588 4804 12600
rect 4856 12588 4862 12640
rect 9030 12588 9036 12640
rect 9088 12628 9094 12640
rect 9125 12631 9183 12637
rect 9125 12628 9137 12631
rect 9088 12600 9137 12628
rect 9088 12588 9094 12600
rect 9125 12597 9137 12600
rect 9171 12628 9183 12631
rect 10778 12628 10784 12640
rect 9171 12600 10784 12628
rect 9171 12597 9183 12600
rect 9125 12591 9183 12597
rect 10778 12588 10784 12600
rect 10836 12588 10842 12640
rect 14826 12588 14832 12640
rect 14884 12628 14890 12640
rect 15841 12631 15899 12637
rect 15841 12628 15853 12631
rect 14884 12600 15853 12628
rect 14884 12588 14890 12600
rect 15841 12597 15853 12600
rect 15887 12628 15899 12631
rect 16482 12628 16488 12640
rect 15887 12600 16488 12628
rect 15887 12597 15899 12600
rect 15841 12591 15899 12597
rect 16482 12588 16488 12600
rect 16540 12588 16546 12640
rect 16758 12628 16764 12640
rect 16719 12600 16764 12628
rect 16758 12588 16764 12600
rect 16816 12588 16822 12640
rect 17494 12628 17500 12640
rect 17455 12600 17500 12628
rect 17494 12588 17500 12600
rect 17552 12588 17558 12640
rect 17696 12628 17724 12668
rect 17862 12656 17868 12668
rect 17920 12656 17926 12708
rect 18046 12696 18052 12708
rect 18007 12668 18052 12696
rect 18046 12656 18052 12668
rect 18104 12656 18110 12708
rect 18138 12656 18144 12708
rect 18196 12696 18202 12708
rect 18233 12699 18291 12705
rect 18233 12696 18245 12699
rect 18196 12668 18245 12696
rect 18196 12656 18202 12668
rect 18233 12665 18245 12668
rect 18279 12665 18291 12699
rect 18233 12659 18291 12665
rect 18340 12628 18368 12736
rect 18414 12724 18420 12736
rect 18472 12724 18478 12776
rect 17696 12600 18368 12628
rect 1104 12538 18860 12560
rect 1104 12486 6912 12538
rect 6964 12486 6976 12538
rect 7028 12486 7040 12538
rect 7092 12486 7104 12538
rect 7156 12486 12843 12538
rect 12895 12486 12907 12538
rect 12959 12486 12971 12538
rect 13023 12486 13035 12538
rect 13087 12486 18860 12538
rect 1104 12464 18860 12486
rect 1581 12427 1639 12433
rect 1581 12393 1593 12427
rect 1627 12424 1639 12427
rect 5258 12424 5264 12436
rect 1627 12396 5264 12424
rect 1627 12393 1639 12396
rect 1581 12387 1639 12393
rect 5258 12384 5264 12396
rect 5316 12384 5322 12436
rect 5537 12427 5595 12433
rect 5537 12393 5549 12427
rect 5583 12424 5595 12427
rect 5721 12427 5779 12433
rect 5721 12424 5733 12427
rect 5583 12396 5733 12424
rect 5583 12393 5595 12396
rect 5537 12387 5595 12393
rect 5721 12393 5733 12396
rect 5767 12424 5779 12427
rect 5902 12424 5908 12436
rect 5767 12396 5908 12424
rect 5767 12393 5779 12396
rect 5721 12387 5779 12393
rect 5902 12384 5908 12396
rect 5960 12384 5966 12436
rect 7929 12427 7987 12433
rect 7929 12393 7941 12427
rect 7975 12424 7987 12427
rect 9766 12424 9772 12436
rect 7975 12396 9772 12424
rect 7975 12393 7987 12396
rect 7929 12387 7987 12393
rect 9766 12384 9772 12396
rect 9824 12384 9830 12436
rect 9861 12427 9919 12433
rect 9861 12393 9873 12427
rect 9907 12424 9919 12427
rect 10686 12424 10692 12436
rect 9907 12396 10692 12424
rect 9907 12393 9919 12396
rect 9861 12387 9919 12393
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 11149 12427 11207 12433
rect 11149 12393 11161 12427
rect 11195 12424 11207 12427
rect 12158 12424 12164 12436
rect 11195 12396 12164 12424
rect 11195 12393 11207 12396
rect 11149 12387 11207 12393
rect 12158 12384 12164 12396
rect 12216 12384 12222 12436
rect 16942 12424 16948 12436
rect 12406 12396 16948 12424
rect 1670 12316 1676 12368
rect 1728 12356 1734 12368
rect 2133 12359 2191 12365
rect 2133 12356 2145 12359
rect 1728 12328 2145 12356
rect 1728 12316 1734 12328
rect 2133 12325 2145 12328
rect 2179 12325 2191 12359
rect 2133 12319 2191 12325
rect 3602 12316 3608 12368
rect 3660 12356 3666 12368
rect 4341 12359 4399 12365
rect 4341 12356 4353 12359
rect 3660 12328 4353 12356
rect 3660 12316 3666 12328
rect 4341 12325 4353 12328
rect 4387 12356 4399 12359
rect 8481 12359 8539 12365
rect 8481 12356 8493 12359
rect 4387 12328 8493 12356
rect 4387 12325 4399 12328
rect 4341 12319 4399 12325
rect 8481 12325 8493 12328
rect 8527 12356 8539 12359
rect 8665 12359 8723 12365
rect 8665 12356 8677 12359
rect 8527 12328 8677 12356
rect 8527 12325 8539 12328
rect 8481 12319 8539 12325
rect 8665 12325 8677 12328
rect 8711 12356 8723 12359
rect 12250 12356 12256 12368
rect 8711 12328 12256 12356
rect 8711 12325 8723 12328
rect 8665 12319 8723 12325
rect 12250 12316 12256 12328
rect 12308 12316 12314 12368
rect 1486 12288 1492 12300
rect 1447 12260 1492 12288
rect 1486 12248 1492 12260
rect 1544 12248 1550 12300
rect 1762 12248 1768 12300
rect 1820 12288 1826 12300
rect 1857 12291 1915 12297
rect 1857 12288 1869 12291
rect 1820 12260 1869 12288
rect 1820 12248 1826 12260
rect 1857 12257 1869 12260
rect 1903 12288 1915 12291
rect 2869 12291 2927 12297
rect 2869 12288 2881 12291
rect 1903 12260 2881 12288
rect 1903 12257 1915 12260
rect 1857 12251 1915 12257
rect 2869 12257 2881 12260
rect 2915 12257 2927 12291
rect 2869 12251 2927 12257
rect 4157 12291 4215 12297
rect 4157 12257 4169 12291
rect 4203 12288 4215 12291
rect 6178 12288 6184 12300
rect 4203 12260 6184 12288
rect 4203 12257 4215 12260
rect 4157 12251 4215 12257
rect 6178 12248 6184 12260
rect 6236 12248 6242 12300
rect 7009 12291 7067 12297
rect 7009 12257 7021 12291
rect 7055 12288 7067 12291
rect 7742 12288 7748 12300
rect 7055 12260 7748 12288
rect 7055 12257 7067 12260
rect 7009 12251 7067 12257
rect 7742 12248 7748 12260
rect 7800 12248 7806 12300
rect 9493 12291 9551 12297
rect 9493 12257 9505 12291
rect 9539 12288 9551 12291
rect 11790 12288 11796 12300
rect 9539 12260 11796 12288
rect 9539 12257 9551 12260
rect 9493 12251 9551 12257
rect 11790 12248 11796 12260
rect 11848 12248 11854 12300
rect 11882 12248 11888 12300
rect 11940 12288 11946 12300
rect 12406 12288 12434 12396
rect 16942 12384 16948 12396
rect 17000 12384 17006 12436
rect 17034 12384 17040 12436
rect 17092 12424 17098 12436
rect 18325 12427 18383 12433
rect 18325 12424 18337 12427
rect 17092 12396 18337 12424
rect 17092 12384 17098 12396
rect 18325 12393 18337 12396
rect 18371 12393 18383 12427
rect 18325 12387 18383 12393
rect 15378 12356 15384 12368
rect 15339 12328 15384 12356
rect 15378 12316 15384 12328
rect 15436 12316 15442 12368
rect 16666 12356 16672 12368
rect 15488 12328 16672 12356
rect 11940 12260 12434 12288
rect 11940 12248 11946 12260
rect 13906 12248 13912 12300
rect 13964 12288 13970 12300
rect 14826 12288 14832 12300
rect 13964 12260 14832 12288
rect 13964 12248 13970 12260
rect 14826 12248 14832 12260
rect 14884 12248 14890 12300
rect 15286 12288 15292 12300
rect 15247 12260 15292 12288
rect 15286 12248 15292 12260
rect 15344 12248 15350 12300
rect 1504 12220 1532 12248
rect 2685 12223 2743 12229
rect 2685 12220 2697 12223
rect 1504 12192 2697 12220
rect 2685 12189 2697 12192
rect 2731 12189 2743 12223
rect 2685 12183 2743 12189
rect 3513 12223 3571 12229
rect 3513 12189 3525 12223
rect 3559 12220 3571 12223
rect 4522 12220 4528 12232
rect 3559 12192 4528 12220
rect 3559 12189 3571 12192
rect 3513 12183 3571 12189
rect 4522 12180 4528 12192
rect 4580 12180 4586 12232
rect 4614 12180 4620 12232
rect 4672 12220 4678 12232
rect 5169 12223 5227 12229
rect 5169 12220 5181 12223
rect 4672 12192 5181 12220
rect 4672 12180 4678 12192
rect 5169 12189 5181 12192
rect 5215 12220 5227 12223
rect 5350 12220 5356 12232
rect 5215 12192 5356 12220
rect 5215 12189 5227 12192
rect 5169 12183 5227 12189
rect 5350 12180 5356 12192
rect 5408 12180 5414 12232
rect 5626 12180 5632 12232
rect 5684 12220 5690 12232
rect 7193 12223 7251 12229
rect 7193 12220 7205 12223
rect 5684 12192 7205 12220
rect 5684 12180 5690 12192
rect 7193 12189 7205 12192
rect 7239 12220 7251 12223
rect 7285 12223 7343 12229
rect 7285 12220 7297 12223
rect 7239 12192 7297 12220
rect 7239 12189 7251 12192
rect 7193 12183 7251 12189
rect 7285 12189 7297 12192
rect 7331 12189 7343 12223
rect 7285 12183 7343 12189
rect 7834 12180 7840 12232
rect 7892 12220 7898 12232
rect 8205 12223 8263 12229
rect 8205 12220 8217 12223
rect 7892 12192 8217 12220
rect 7892 12180 7898 12192
rect 8205 12189 8217 12192
rect 8251 12220 8263 12223
rect 8757 12223 8815 12229
rect 8757 12220 8769 12223
rect 8251 12192 8769 12220
rect 8251 12189 8263 12192
rect 8205 12183 8263 12189
rect 8757 12189 8769 12192
rect 8803 12220 8815 12223
rect 9030 12220 9036 12232
rect 8803 12192 9036 12220
rect 8803 12189 8815 12192
rect 8757 12183 8815 12189
rect 9030 12180 9036 12192
rect 9088 12180 9094 12232
rect 9217 12223 9275 12229
rect 9217 12189 9229 12223
rect 9263 12189 9275 12223
rect 9398 12220 9404 12232
rect 9359 12192 9404 12220
rect 9217 12183 9275 12189
rect 1854 12112 1860 12164
rect 1912 12152 1918 12164
rect 2317 12155 2375 12161
rect 2317 12152 2329 12155
rect 1912 12124 2329 12152
rect 1912 12112 1918 12124
rect 2317 12121 2329 12124
rect 2363 12121 2375 12155
rect 2317 12115 2375 12121
rect 2593 12155 2651 12161
rect 2593 12121 2605 12155
rect 2639 12152 2651 12155
rect 2774 12152 2780 12164
rect 2639 12124 2780 12152
rect 2639 12121 2651 12124
rect 2593 12115 2651 12121
rect 2774 12112 2780 12124
rect 2832 12112 2838 12164
rect 2866 12112 2872 12164
rect 2924 12152 2930 12164
rect 3697 12155 3755 12161
rect 3697 12152 3709 12155
rect 2924 12124 3709 12152
rect 2924 12112 2930 12124
rect 3697 12121 3709 12124
rect 3743 12152 3755 12155
rect 4985 12155 5043 12161
rect 3743 12124 4936 12152
rect 3743 12121 3755 12124
rect 3697 12115 3755 12121
rect 1949 12087 2007 12093
rect 1949 12053 1961 12087
rect 1995 12084 2007 12087
rect 2038 12084 2044 12096
rect 1995 12056 2044 12084
rect 1995 12053 2007 12056
rect 1949 12047 2007 12053
rect 2038 12044 2044 12056
rect 2096 12044 2102 12096
rect 3050 12084 3056 12096
rect 3011 12056 3056 12084
rect 3050 12044 3056 12056
rect 3108 12044 3114 12096
rect 3329 12087 3387 12093
rect 3329 12053 3341 12087
rect 3375 12084 3387 12087
rect 3602 12084 3608 12096
rect 3375 12056 3608 12084
rect 3375 12053 3387 12056
rect 3329 12047 3387 12053
rect 3602 12044 3608 12056
rect 3660 12044 3666 12096
rect 3973 12087 4031 12093
rect 3973 12053 3985 12087
rect 4019 12084 4031 12087
rect 4246 12084 4252 12096
rect 4019 12056 4252 12084
rect 4019 12053 4031 12056
rect 3973 12047 4031 12053
rect 4246 12044 4252 12056
rect 4304 12044 4310 12096
rect 4525 12087 4583 12093
rect 4525 12053 4537 12087
rect 4571 12084 4583 12087
rect 4798 12084 4804 12096
rect 4571 12056 4804 12084
rect 4571 12053 4583 12056
rect 4525 12047 4583 12053
rect 4798 12044 4804 12056
rect 4856 12044 4862 12096
rect 4908 12084 4936 12124
rect 4985 12121 4997 12155
rect 5031 12152 5043 12155
rect 5997 12155 6055 12161
rect 5997 12152 6009 12155
rect 5031 12124 6009 12152
rect 5031 12121 5043 12124
rect 4985 12115 5043 12121
rect 5997 12121 6009 12124
rect 6043 12152 6055 12155
rect 9232 12152 9260 12183
rect 9398 12180 9404 12192
rect 9456 12180 9462 12232
rect 9674 12180 9680 12232
rect 9732 12220 9738 12232
rect 10321 12223 10379 12229
rect 10321 12220 10333 12223
rect 9732 12192 10333 12220
rect 9732 12180 9738 12192
rect 10321 12189 10333 12192
rect 10367 12220 10379 12223
rect 10410 12220 10416 12232
rect 10367 12192 10416 12220
rect 10367 12189 10379 12192
rect 10321 12183 10379 12189
rect 10410 12180 10416 12192
rect 10468 12180 10474 12232
rect 10594 12220 10600 12232
rect 10555 12192 10600 12220
rect 10594 12180 10600 12192
rect 10652 12180 10658 12232
rect 11146 12180 11152 12232
rect 11204 12220 11210 12232
rect 13814 12220 13820 12232
rect 11204 12192 13820 12220
rect 11204 12180 11210 12192
rect 13814 12180 13820 12192
rect 13872 12220 13878 12232
rect 15013 12223 15071 12229
rect 15013 12220 15025 12223
rect 13872 12192 15025 12220
rect 13872 12180 13878 12192
rect 15013 12189 15025 12192
rect 15059 12220 15071 12223
rect 15488 12220 15516 12328
rect 16666 12316 16672 12328
rect 16724 12316 16730 12368
rect 17405 12359 17463 12365
rect 17405 12325 17417 12359
rect 17451 12356 17463 12359
rect 17451 12328 18460 12356
rect 17451 12325 17463 12328
rect 17405 12319 17463 12325
rect 15654 12248 15660 12300
rect 15712 12288 15718 12300
rect 16209 12291 16267 12297
rect 16209 12288 16221 12291
rect 15712 12260 16221 12288
rect 15712 12248 15718 12260
rect 16209 12257 16221 12260
rect 16255 12257 16267 12291
rect 16209 12251 16267 12257
rect 17218 12248 17224 12300
rect 17276 12288 17282 12300
rect 18432 12297 18460 12328
rect 17957 12291 18015 12297
rect 17957 12288 17969 12291
rect 17276 12260 17969 12288
rect 17276 12248 17282 12260
rect 17957 12257 17969 12260
rect 18003 12257 18015 12291
rect 17957 12251 18015 12257
rect 18417 12291 18475 12297
rect 18417 12257 18429 12291
rect 18463 12288 18475 12291
rect 18969 12291 19027 12297
rect 18969 12288 18981 12291
rect 18463 12260 18981 12288
rect 18463 12257 18475 12260
rect 18417 12251 18475 12257
rect 18969 12257 18981 12260
rect 19015 12257 19027 12291
rect 18969 12251 19027 12257
rect 15059 12192 15516 12220
rect 15565 12223 15623 12229
rect 15059 12189 15071 12192
rect 15013 12183 15071 12189
rect 15565 12189 15577 12223
rect 15611 12220 15623 12223
rect 16574 12220 16580 12232
rect 15611 12192 16580 12220
rect 15611 12189 15623 12192
rect 15565 12183 15623 12189
rect 9582 12152 9588 12164
rect 6043 12124 8156 12152
rect 9232 12124 9588 12152
rect 6043 12121 6055 12124
rect 5997 12115 6055 12121
rect 5718 12084 5724 12096
rect 4908 12056 5724 12084
rect 5718 12044 5724 12056
rect 5776 12044 5782 12096
rect 6178 12084 6184 12096
rect 6139 12056 6184 12084
rect 6178 12044 6184 12056
rect 6236 12044 6242 12096
rect 6365 12087 6423 12093
rect 6365 12053 6377 12087
rect 6411 12084 6423 12087
rect 6454 12084 6460 12096
rect 6411 12056 6460 12084
rect 6411 12053 6423 12056
rect 6365 12047 6423 12053
rect 6454 12044 6460 12056
rect 6512 12044 6518 12096
rect 6546 12044 6552 12096
rect 6604 12084 6610 12096
rect 6825 12087 6883 12093
rect 6604 12056 6649 12084
rect 6604 12044 6610 12056
rect 6825 12053 6837 12087
rect 6871 12084 6883 12087
rect 7834 12084 7840 12096
rect 6871 12056 7840 12084
rect 6871 12053 6883 12056
rect 6825 12047 6883 12053
rect 7834 12044 7840 12056
rect 7892 12044 7898 12096
rect 8018 12084 8024 12096
rect 7979 12056 8024 12084
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 8128 12084 8156 12124
rect 9582 12112 9588 12124
rect 9640 12112 9646 12164
rect 9692 12124 12434 12152
rect 9692 12084 9720 12124
rect 8128 12056 9720 12084
rect 9766 12044 9772 12096
rect 9824 12084 9830 12096
rect 9953 12087 10011 12093
rect 9953 12084 9965 12087
rect 9824 12056 9965 12084
rect 9824 12044 9830 12056
rect 9953 12053 9965 12056
rect 9999 12053 10011 12087
rect 10226 12084 10232 12096
rect 10187 12056 10232 12084
rect 9953 12047 10011 12053
rect 10226 12044 10232 12056
rect 10284 12044 10290 12096
rect 10778 12084 10784 12096
rect 10739 12056 10784 12084
rect 10778 12044 10784 12056
rect 10836 12044 10842 12096
rect 11146 12044 11152 12096
rect 11204 12084 11210 12096
rect 11241 12087 11299 12093
rect 11241 12084 11253 12087
rect 11204 12056 11253 12084
rect 11204 12044 11210 12056
rect 11241 12053 11253 12056
rect 11287 12053 11299 12087
rect 11241 12047 11299 12053
rect 11330 12044 11336 12096
rect 11388 12084 11394 12096
rect 11974 12084 11980 12096
rect 11388 12056 11980 12084
rect 11388 12044 11394 12056
rect 11974 12044 11980 12056
rect 12032 12044 12038 12096
rect 12406 12084 12434 12124
rect 13170 12112 13176 12164
rect 13228 12152 13234 12164
rect 15580 12152 15608 12183
rect 16574 12180 16580 12192
rect 16632 12180 16638 12232
rect 16761 12223 16819 12229
rect 16761 12189 16773 12223
rect 16807 12220 16819 12223
rect 17129 12223 17187 12229
rect 16807 12192 17080 12220
rect 16807 12189 16819 12192
rect 16761 12183 16819 12189
rect 13228 12124 15608 12152
rect 15841 12155 15899 12161
rect 13228 12112 13234 12124
rect 15841 12121 15853 12155
rect 15887 12152 15899 12155
rect 16942 12152 16948 12164
rect 15887 12124 16948 12152
rect 15887 12121 15899 12124
rect 15841 12115 15899 12121
rect 16942 12112 16948 12124
rect 17000 12112 17006 12164
rect 17052 12152 17080 12192
rect 17129 12189 17141 12223
rect 17175 12220 17187 12223
rect 17494 12220 17500 12232
rect 17175 12192 17500 12220
rect 17175 12189 17187 12192
rect 17129 12183 17187 12189
rect 17494 12180 17500 12192
rect 17552 12180 17558 12232
rect 17773 12155 17831 12161
rect 17052 12124 17632 12152
rect 13262 12084 13268 12096
rect 12406 12056 13268 12084
rect 13262 12044 13268 12056
rect 13320 12044 13326 12096
rect 14458 12044 14464 12096
rect 14516 12084 14522 12096
rect 14553 12087 14611 12093
rect 14553 12084 14565 12087
rect 14516 12056 14565 12084
rect 14516 12044 14522 12056
rect 14553 12053 14565 12056
rect 14599 12084 14611 12087
rect 14734 12084 14740 12096
rect 14599 12056 14740 12084
rect 14599 12053 14611 12056
rect 14553 12047 14611 12053
rect 14734 12044 14740 12056
rect 14792 12044 14798 12096
rect 16025 12087 16083 12093
rect 16025 12053 16037 12087
rect 16071 12084 16083 12087
rect 16114 12084 16120 12096
rect 16071 12056 16120 12084
rect 16071 12053 16083 12056
rect 16025 12047 16083 12053
rect 16114 12044 16120 12056
rect 16172 12044 16178 12096
rect 16390 12084 16396 12096
rect 16351 12056 16396 12084
rect 16390 12044 16396 12056
rect 16448 12044 16454 12096
rect 16853 12087 16911 12093
rect 16853 12053 16865 12087
rect 16899 12084 16911 12087
rect 17034 12084 17040 12096
rect 16899 12056 17040 12084
rect 16899 12053 16911 12056
rect 16853 12047 16911 12053
rect 17034 12044 17040 12056
rect 17092 12044 17098 12096
rect 17402 12044 17408 12096
rect 17460 12084 17466 12096
rect 17497 12087 17555 12093
rect 17497 12084 17509 12087
rect 17460 12056 17509 12084
rect 17460 12044 17466 12056
rect 17497 12053 17509 12056
rect 17543 12053 17555 12087
rect 17604 12084 17632 12124
rect 17773 12121 17785 12155
rect 17819 12152 17831 12155
rect 18414 12152 18420 12164
rect 17819 12124 18420 12152
rect 17819 12121 17831 12124
rect 17773 12115 17831 12121
rect 18414 12112 18420 12124
rect 18472 12112 18478 12164
rect 17862 12084 17868 12096
rect 17604 12056 17868 12084
rect 17497 12047 17555 12053
rect 17862 12044 17868 12056
rect 17920 12044 17926 12096
rect 18046 12084 18052 12096
rect 18007 12056 18052 12084
rect 18046 12044 18052 12056
rect 18104 12044 18110 12096
rect 1104 11994 18860 12016
rect 1104 11942 3947 11994
rect 3999 11942 4011 11994
rect 4063 11942 4075 11994
rect 4127 11942 4139 11994
rect 4191 11942 9878 11994
rect 9930 11942 9942 11994
rect 9994 11942 10006 11994
rect 10058 11942 10070 11994
rect 10122 11942 15808 11994
rect 15860 11942 15872 11994
rect 15924 11942 15936 11994
rect 15988 11942 16000 11994
rect 16052 11942 18860 11994
rect 1104 11920 18860 11942
rect 3510 11880 3516 11892
rect 2746 11852 3516 11880
rect 1673 11815 1731 11821
rect 1673 11781 1685 11815
rect 1719 11812 1731 11815
rect 2746 11812 2774 11852
rect 3510 11840 3516 11852
rect 3568 11840 3574 11892
rect 5445 11883 5503 11889
rect 5445 11849 5457 11883
rect 5491 11880 5503 11883
rect 5534 11880 5540 11892
rect 5491 11852 5540 11880
rect 5491 11849 5503 11852
rect 5445 11843 5503 11849
rect 5534 11840 5540 11852
rect 5592 11880 5598 11892
rect 6546 11880 6552 11892
rect 5592 11852 6552 11880
rect 5592 11840 5598 11852
rect 6546 11840 6552 11852
rect 6604 11840 6610 11892
rect 6641 11883 6699 11889
rect 6641 11849 6653 11883
rect 6687 11880 6699 11883
rect 8021 11883 8079 11889
rect 8021 11880 8033 11883
rect 6687 11852 8033 11880
rect 6687 11849 6699 11852
rect 6641 11843 6699 11849
rect 8021 11849 8033 11852
rect 8067 11880 8079 11883
rect 8110 11880 8116 11892
rect 8067 11852 8116 11880
rect 8067 11849 8079 11852
rect 8021 11843 8079 11849
rect 8110 11840 8116 11852
rect 8168 11840 8174 11892
rect 8662 11880 8668 11892
rect 8220 11852 8668 11880
rect 1719 11784 2774 11812
rect 3145 11815 3203 11821
rect 1719 11781 1731 11784
rect 1673 11775 1731 11781
rect 3145 11781 3157 11815
rect 3191 11812 3203 11815
rect 8220 11812 8248 11852
rect 8662 11840 8668 11852
rect 8720 11880 8726 11892
rect 8720 11852 9996 11880
rect 8720 11840 8726 11852
rect 9968 11824 9996 11852
rect 10318 11840 10324 11892
rect 10376 11880 10382 11892
rect 10778 11880 10784 11892
rect 10376 11852 10784 11880
rect 10376 11840 10382 11852
rect 10778 11840 10784 11852
rect 10836 11880 10842 11892
rect 14274 11880 14280 11892
rect 10836 11852 14280 11880
rect 10836 11840 10842 11852
rect 14274 11840 14280 11852
rect 14332 11840 14338 11892
rect 14366 11840 14372 11892
rect 14424 11880 14430 11892
rect 15010 11880 15016 11892
rect 14424 11852 14688 11880
rect 14971 11852 15016 11880
rect 14424 11840 14430 11852
rect 3191 11784 8248 11812
rect 3191 11781 3203 11784
rect 3145 11775 3203 11781
rect 9582 11772 9588 11824
rect 9640 11812 9646 11824
rect 9677 11815 9735 11821
rect 9677 11812 9689 11815
rect 9640 11784 9689 11812
rect 9640 11772 9646 11784
rect 9677 11781 9689 11784
rect 9723 11781 9735 11815
rect 9677 11775 9735 11781
rect 9950 11772 9956 11824
rect 10008 11772 10014 11824
rect 12066 11812 12072 11824
rect 11979 11784 12072 11812
rect 12066 11772 12072 11784
rect 12124 11812 12130 11824
rect 14660 11821 14688 11852
rect 15010 11840 15016 11852
rect 15068 11840 15074 11892
rect 15102 11840 15108 11892
rect 15160 11880 15166 11892
rect 16390 11880 16396 11892
rect 15160 11852 16396 11880
rect 15160 11840 15166 11852
rect 16390 11840 16396 11852
rect 16448 11840 16454 11892
rect 16850 11880 16856 11892
rect 16500 11852 16856 11880
rect 14645 11815 14703 11821
rect 12124 11784 14504 11812
rect 12124 11772 12130 11784
rect 2222 11744 2228 11756
rect 2183 11716 2228 11744
rect 2222 11704 2228 11716
rect 2280 11704 2286 11756
rect 2590 11744 2596 11756
rect 2503 11716 2596 11744
rect 1670 11636 1676 11688
rect 1728 11676 1734 11688
rect 1765 11679 1823 11685
rect 1765 11676 1777 11679
rect 1728 11648 1777 11676
rect 1728 11636 1734 11648
rect 1765 11645 1777 11648
rect 1811 11645 1823 11679
rect 1765 11639 1823 11645
rect 2130 11636 2136 11688
rect 2188 11676 2194 11688
rect 2516 11676 2544 11716
rect 2590 11704 2596 11716
rect 2648 11744 2654 11756
rect 4801 11747 4859 11753
rect 2648 11716 4016 11744
rect 2648 11704 2654 11716
rect 3988 11688 4016 11716
rect 4801 11713 4813 11747
rect 4847 11744 4859 11747
rect 4847 11716 6040 11744
rect 4847 11713 4859 11716
rect 4801 11707 4859 11713
rect 2774 11676 2780 11688
rect 2188 11648 2544 11676
rect 2188 11636 2194 11648
rect 2746 11636 2780 11676
rect 2832 11636 2838 11688
rect 2961 11679 3019 11685
rect 2961 11645 2973 11679
rect 3007 11676 3019 11679
rect 3050 11676 3056 11688
rect 3007 11648 3056 11676
rect 3007 11645 3019 11648
rect 2961 11639 3019 11645
rect 3050 11636 3056 11648
rect 3108 11636 3114 11688
rect 3510 11636 3516 11688
rect 3568 11676 3574 11688
rect 3697 11679 3755 11685
rect 3697 11676 3709 11679
rect 3568 11648 3709 11676
rect 3568 11636 3574 11648
rect 3697 11645 3709 11648
rect 3743 11645 3755 11679
rect 3970 11676 3976 11688
rect 3931 11648 3976 11676
rect 3697 11639 3755 11645
rect 3970 11636 3976 11648
rect 4028 11636 4034 11688
rect 4246 11636 4252 11688
rect 4304 11676 4310 11688
rect 4982 11676 4988 11688
rect 4304 11648 4988 11676
rect 4304 11636 4310 11648
rect 4982 11636 4988 11648
rect 5040 11676 5046 11688
rect 5442 11676 5448 11688
rect 5040 11648 5448 11676
rect 5040 11636 5046 11648
rect 5442 11636 5448 11648
rect 5500 11636 5506 11688
rect 5626 11676 5632 11688
rect 5587 11648 5632 11676
rect 5626 11636 5632 11648
rect 5684 11636 5690 11688
rect 6012 11685 6040 11716
rect 6086 11704 6092 11756
rect 6144 11744 6150 11756
rect 6457 11747 6515 11753
rect 6457 11744 6469 11747
rect 6144 11716 6469 11744
rect 6144 11704 6150 11716
rect 6457 11713 6469 11716
rect 6503 11713 6515 11747
rect 6457 11707 6515 11713
rect 6546 11704 6552 11756
rect 6604 11744 6610 11756
rect 7285 11747 7343 11753
rect 7285 11744 7297 11747
rect 6604 11716 7297 11744
rect 6604 11704 6610 11716
rect 7285 11713 7297 11716
rect 7331 11713 7343 11747
rect 7285 11707 7343 11713
rect 7742 11704 7748 11756
rect 7800 11744 7806 11756
rect 8113 11747 8171 11753
rect 8113 11744 8125 11747
rect 7800 11716 8125 11744
rect 7800 11704 7806 11716
rect 5997 11679 6055 11685
rect 5997 11645 6009 11679
rect 6043 11676 6055 11679
rect 6638 11676 6644 11688
rect 6043 11648 6644 11676
rect 6043 11645 6055 11648
rect 5997 11639 6055 11645
rect 6638 11636 6644 11648
rect 6696 11636 6702 11688
rect 7374 11676 7380 11688
rect 6840 11648 7380 11676
rect 1394 11568 1400 11620
rect 1452 11608 1458 11620
rect 1489 11611 1547 11617
rect 1489 11608 1501 11611
rect 1452 11580 1501 11608
rect 1452 11568 1458 11580
rect 1489 11577 1501 11580
rect 1535 11608 1547 11611
rect 2746 11608 2774 11636
rect 1535 11580 2774 11608
rect 4525 11611 4583 11617
rect 1535 11577 1547 11580
rect 1489 11571 1547 11577
rect 4525 11577 4537 11611
rect 4571 11608 4583 11611
rect 5350 11608 5356 11620
rect 4571 11580 5356 11608
rect 4571 11577 4583 11580
rect 4525 11571 4583 11577
rect 5350 11568 5356 11580
rect 5408 11568 5414 11620
rect 1946 11540 1952 11552
rect 1907 11512 1952 11540
rect 1946 11500 1952 11512
rect 2004 11500 2010 11552
rect 2314 11540 2320 11552
rect 2275 11512 2320 11540
rect 2314 11500 2320 11512
rect 2372 11500 2378 11552
rect 2406 11500 2412 11552
rect 2464 11540 2470 11552
rect 2464 11512 2509 11540
rect 2464 11500 2470 11512
rect 2774 11500 2780 11552
rect 2832 11540 2838 11552
rect 3234 11540 3240 11552
rect 2832 11512 2877 11540
rect 3195 11512 3240 11540
rect 2832 11500 2838 11512
rect 3234 11500 3240 11512
rect 3292 11500 3298 11552
rect 3418 11500 3424 11552
rect 3476 11540 3482 11552
rect 3513 11543 3571 11549
rect 3513 11540 3525 11543
rect 3476 11512 3525 11540
rect 3476 11500 3482 11512
rect 3513 11509 3525 11512
rect 3559 11509 3571 11543
rect 3513 11503 3571 11509
rect 3602 11500 3608 11552
rect 3660 11540 3666 11552
rect 4065 11543 4123 11549
rect 4065 11540 4077 11543
rect 3660 11512 4077 11540
rect 3660 11500 3666 11512
rect 4065 11509 4077 11512
rect 4111 11509 4123 11543
rect 4246 11540 4252 11552
rect 4207 11512 4252 11540
rect 4065 11503 4123 11509
rect 4246 11500 4252 11512
rect 4304 11500 4310 11552
rect 5261 11543 5319 11549
rect 5261 11509 5273 11543
rect 5307 11540 5319 11543
rect 5644 11540 5672 11636
rect 5718 11568 5724 11620
rect 5776 11608 5782 11620
rect 5813 11611 5871 11617
rect 5813 11608 5825 11611
rect 5776 11580 5825 11608
rect 5776 11568 5782 11580
rect 5813 11577 5825 11580
rect 5859 11608 5871 11611
rect 6454 11608 6460 11620
rect 5859 11580 6460 11608
rect 5859 11577 5871 11580
rect 5813 11571 5871 11577
rect 6454 11568 6460 11580
rect 6512 11608 6518 11620
rect 6840 11608 6868 11648
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 6512 11580 6868 11608
rect 7101 11611 7159 11617
rect 6512 11568 6518 11580
rect 7101 11577 7113 11611
rect 7147 11608 7159 11611
rect 7282 11608 7288 11620
rect 7147 11580 7288 11608
rect 7147 11577 7159 11580
rect 7101 11571 7159 11577
rect 7282 11568 7288 11580
rect 7340 11568 7346 11620
rect 6270 11540 6276 11552
rect 5307 11512 5672 11540
rect 6231 11512 6276 11540
rect 5307 11509 5319 11512
rect 5261 11503 5319 11509
rect 6270 11500 6276 11512
rect 6328 11500 6334 11552
rect 6730 11540 6736 11552
rect 6691 11512 6736 11540
rect 6730 11500 6736 11512
rect 6788 11500 6794 11552
rect 7193 11543 7251 11549
rect 7193 11509 7205 11543
rect 7239 11540 7251 11543
rect 7466 11540 7472 11552
rect 7239 11512 7472 11540
rect 7239 11509 7251 11512
rect 7193 11503 7251 11509
rect 7466 11500 7472 11512
rect 7524 11500 7530 11552
rect 7558 11500 7564 11552
rect 7616 11540 7622 11552
rect 7653 11543 7711 11549
rect 7653 11540 7665 11543
rect 7616 11512 7665 11540
rect 7616 11500 7622 11512
rect 7653 11509 7665 11512
rect 7699 11509 7711 11543
rect 7944 11540 7972 11716
rect 8113 11713 8125 11716
rect 8159 11713 8171 11747
rect 8113 11707 8171 11713
rect 9306 11704 9312 11756
rect 9364 11744 9370 11756
rect 9490 11744 9496 11756
rect 9364 11716 9496 11744
rect 9364 11704 9370 11716
rect 9490 11704 9496 11716
rect 9548 11704 9554 11756
rect 10413 11747 10471 11753
rect 10413 11713 10425 11747
rect 10459 11744 10471 11747
rect 10594 11744 10600 11756
rect 10459 11716 10600 11744
rect 10459 11713 10471 11716
rect 10413 11707 10471 11713
rect 10594 11704 10600 11716
rect 10652 11744 10658 11756
rect 10781 11747 10839 11753
rect 10781 11744 10793 11747
rect 10652 11716 10793 11744
rect 10652 11704 10658 11716
rect 10781 11713 10793 11716
rect 10827 11713 10839 11747
rect 10781 11707 10839 11713
rect 12253 11747 12311 11753
rect 12253 11713 12265 11747
rect 12299 11744 12311 11747
rect 12434 11744 12440 11756
rect 12299 11716 12440 11744
rect 12299 11713 12311 11716
rect 12253 11707 12311 11713
rect 12434 11704 12440 11716
rect 12492 11704 12498 11756
rect 14476 11744 14504 11784
rect 14645 11781 14657 11815
rect 14691 11812 14703 11815
rect 16500 11812 16528 11852
rect 16850 11840 16856 11852
rect 16908 11840 16914 11892
rect 17218 11880 17224 11892
rect 17179 11852 17224 11880
rect 17218 11840 17224 11852
rect 17276 11840 17282 11892
rect 14691 11784 16528 11812
rect 14691 11781 14703 11784
rect 14645 11775 14703 11781
rect 16666 11772 16672 11824
rect 16724 11812 16730 11824
rect 17126 11812 17132 11824
rect 16724 11784 17132 11812
rect 16724 11772 16730 11784
rect 17126 11772 17132 11784
rect 17184 11812 17190 11824
rect 18141 11815 18199 11821
rect 18141 11812 18153 11815
rect 17184 11784 18153 11812
rect 17184 11772 17190 11784
rect 18141 11781 18153 11784
rect 18187 11781 18199 11815
rect 18141 11775 18199 11781
rect 14476 11716 14872 11744
rect 8294 11676 8300 11688
rect 8255 11648 8300 11676
rect 8294 11636 8300 11648
rect 8352 11636 8358 11688
rect 14844 11685 14872 11716
rect 15470 11704 15476 11756
rect 15528 11744 15534 11756
rect 16574 11744 16580 11756
rect 15528 11716 16580 11744
rect 15528 11704 15534 11716
rect 16574 11704 16580 11716
rect 16632 11704 16638 11756
rect 16761 11747 16819 11753
rect 16761 11713 16773 11747
rect 16807 11744 16819 11747
rect 16807 11716 17908 11744
rect 16807 11713 16819 11716
rect 16761 11707 16819 11713
rect 10965 11679 11023 11685
rect 10965 11676 10977 11679
rect 8404 11648 10977 11676
rect 8018 11568 8024 11620
rect 8076 11608 8082 11620
rect 8404 11608 8432 11648
rect 10965 11645 10977 11648
rect 11011 11676 11023 11679
rect 11517 11679 11575 11685
rect 11517 11676 11529 11679
rect 11011 11648 11529 11676
rect 11011 11645 11023 11648
rect 10965 11639 11023 11645
rect 11517 11645 11529 11648
rect 11563 11645 11575 11679
rect 11517 11639 11575 11645
rect 14829 11679 14887 11685
rect 14829 11645 14841 11679
rect 14875 11676 14887 11679
rect 14918 11676 14924 11688
rect 14875 11648 14924 11676
rect 14875 11645 14887 11648
rect 14829 11639 14887 11645
rect 14918 11636 14924 11648
rect 14976 11636 14982 11688
rect 15010 11636 15016 11688
rect 15068 11676 15074 11688
rect 15105 11679 15163 11685
rect 15105 11676 15117 11679
rect 15068 11648 15117 11676
rect 15068 11636 15074 11648
rect 15105 11645 15117 11648
rect 15151 11645 15163 11679
rect 15105 11639 15163 11645
rect 15933 11679 15991 11685
rect 15933 11645 15945 11679
rect 15979 11676 15991 11679
rect 16206 11676 16212 11688
rect 15979 11648 16212 11676
rect 15979 11645 15991 11648
rect 15933 11639 15991 11645
rect 16206 11636 16212 11648
rect 16264 11636 16270 11688
rect 17034 11676 17040 11688
rect 16995 11648 17040 11676
rect 17034 11636 17040 11648
rect 17092 11636 17098 11688
rect 17494 11676 17500 11688
rect 17455 11648 17500 11676
rect 17494 11636 17500 11648
rect 17552 11636 17558 11688
rect 8076 11580 8432 11608
rect 8553 11611 8611 11617
rect 8076 11568 8082 11580
rect 8553 11577 8565 11611
rect 8599 11608 8611 11611
rect 8754 11608 8760 11620
rect 8599 11580 8760 11608
rect 8599 11577 8611 11580
rect 8553 11571 8611 11577
rect 8754 11568 8760 11580
rect 8812 11568 8818 11620
rect 9490 11568 9496 11620
rect 9548 11608 9554 11620
rect 11057 11611 11115 11617
rect 9548 11580 10456 11608
rect 9548 11568 9554 11580
rect 8110 11540 8116 11552
rect 7944 11512 8116 11540
rect 7653 11503 7711 11509
rect 8110 11500 8116 11512
rect 8168 11540 8174 11552
rect 9306 11540 9312 11552
rect 8168 11512 9312 11540
rect 8168 11500 8174 11512
rect 9306 11500 9312 11512
rect 9364 11500 9370 11552
rect 9766 11540 9772 11552
rect 9727 11512 9772 11540
rect 9766 11500 9772 11512
rect 9824 11500 9830 11552
rect 9858 11500 9864 11552
rect 9916 11540 9922 11552
rect 10134 11540 10140 11552
rect 9916 11512 10140 11540
rect 9916 11500 9922 11512
rect 10134 11500 10140 11512
rect 10192 11500 10198 11552
rect 10226 11500 10232 11552
rect 10284 11540 10290 11552
rect 10428 11540 10456 11580
rect 11057 11577 11069 11611
rect 11103 11608 11115 11611
rect 11701 11611 11759 11617
rect 11701 11608 11713 11611
rect 11103 11580 11713 11608
rect 11103 11577 11115 11580
rect 11057 11571 11115 11577
rect 11701 11577 11713 11580
rect 11747 11577 11759 11611
rect 11701 11571 11759 11577
rect 12158 11568 12164 11620
rect 12216 11608 12222 11620
rect 12437 11611 12495 11617
rect 12437 11608 12449 11611
rect 12216 11580 12449 11608
rect 12216 11568 12222 11580
rect 12437 11577 12449 11580
rect 12483 11608 12495 11611
rect 14461 11611 14519 11617
rect 14461 11608 14473 11611
rect 12483 11580 14473 11608
rect 12483 11577 12495 11580
rect 12437 11571 12495 11577
rect 14461 11577 14473 11580
rect 14507 11608 14519 11611
rect 15286 11608 15292 11620
rect 14507 11580 15292 11608
rect 14507 11577 14519 11580
rect 14461 11571 14519 11577
rect 15286 11568 15292 11580
rect 15344 11568 15350 11620
rect 17880 11617 17908 11716
rect 17865 11611 17923 11617
rect 17865 11577 17877 11611
rect 17911 11608 17923 11611
rect 18138 11608 18144 11620
rect 17911 11580 18144 11608
rect 17911 11577 17923 11580
rect 17865 11571 17923 11577
rect 18138 11568 18144 11580
rect 18196 11568 18202 11620
rect 18414 11608 18420 11620
rect 18375 11580 18420 11608
rect 18414 11568 18420 11580
rect 18472 11568 18478 11620
rect 11238 11540 11244 11552
rect 10284 11512 10329 11540
rect 10428 11512 11244 11540
rect 10284 11500 10290 11512
rect 11238 11500 11244 11512
rect 11296 11500 11302 11552
rect 11422 11540 11428 11552
rect 11383 11512 11428 11540
rect 11422 11500 11428 11512
rect 11480 11500 11486 11552
rect 11517 11543 11575 11549
rect 11517 11509 11529 11543
rect 11563 11540 11575 11543
rect 12066 11540 12072 11552
rect 11563 11512 12072 11540
rect 11563 11509 11575 11512
rect 11517 11503 11575 11509
rect 12066 11500 12072 11512
rect 12124 11500 12130 11552
rect 13262 11500 13268 11552
rect 13320 11540 13326 11552
rect 14001 11543 14059 11549
rect 14001 11540 14013 11543
rect 13320 11512 14013 11540
rect 13320 11500 13326 11512
rect 14001 11509 14013 11512
rect 14047 11509 14059 11543
rect 14001 11503 14059 11509
rect 16301 11543 16359 11549
rect 16301 11509 16313 11543
rect 16347 11540 16359 11543
rect 16390 11540 16396 11552
rect 16347 11512 16396 11540
rect 16347 11509 16359 11512
rect 16301 11503 16359 11509
rect 16390 11500 16396 11512
rect 16448 11500 16454 11552
rect 16485 11543 16543 11549
rect 16485 11509 16497 11543
rect 16531 11540 16543 11543
rect 16758 11540 16764 11552
rect 16531 11512 16764 11540
rect 16531 11509 16543 11512
rect 16485 11503 16543 11509
rect 16758 11500 16764 11512
rect 16816 11500 16822 11552
rect 16850 11500 16856 11552
rect 16908 11540 16914 11552
rect 17405 11543 17463 11549
rect 17405 11540 17417 11543
rect 16908 11512 17417 11540
rect 16908 11500 16914 11512
rect 17405 11509 17417 11512
rect 17451 11509 17463 11543
rect 17405 11503 17463 11509
rect 17494 11500 17500 11552
rect 17552 11540 17558 11552
rect 17773 11543 17831 11549
rect 17773 11540 17785 11543
rect 17552 11512 17785 11540
rect 17552 11500 17558 11512
rect 17773 11509 17785 11512
rect 17819 11509 17831 11543
rect 17773 11503 17831 11509
rect 1104 11450 18860 11472
rect 1104 11398 6912 11450
rect 6964 11398 6976 11450
rect 7028 11398 7040 11450
rect 7092 11398 7104 11450
rect 7156 11398 12843 11450
rect 12895 11398 12907 11450
rect 12959 11398 12971 11450
rect 13023 11398 13035 11450
rect 13087 11398 18860 11450
rect 1104 11376 18860 11398
rect 4522 11296 4528 11348
rect 4580 11336 4586 11348
rect 5169 11339 5227 11345
rect 5169 11336 5181 11339
rect 4580 11308 5181 11336
rect 4580 11296 4586 11308
rect 5169 11305 5181 11308
rect 5215 11336 5227 11339
rect 6086 11336 6092 11348
rect 5215 11308 6092 11336
rect 5215 11305 5227 11308
rect 5169 11299 5227 11305
rect 6086 11296 6092 11308
rect 6144 11296 6150 11348
rect 7193 11339 7251 11345
rect 7193 11305 7205 11339
rect 7239 11336 7251 11339
rect 7282 11336 7288 11348
rect 7239 11308 7288 11336
rect 7239 11305 7251 11308
rect 7193 11299 7251 11305
rect 7282 11296 7288 11308
rect 7340 11296 7346 11348
rect 7558 11336 7564 11348
rect 7519 11308 7564 11336
rect 7558 11296 7564 11308
rect 7616 11296 7622 11348
rect 7653 11339 7711 11345
rect 7653 11305 7665 11339
rect 7699 11336 7711 11339
rect 8018 11336 8024 11348
rect 7699 11308 8024 11336
rect 7699 11305 7711 11308
rect 7653 11299 7711 11305
rect 8018 11296 8024 11308
rect 8076 11296 8082 11348
rect 8573 11339 8631 11345
rect 8573 11305 8585 11339
rect 8619 11336 8631 11339
rect 9766 11336 9772 11348
rect 8619 11308 9772 11336
rect 8619 11305 8631 11308
rect 8573 11299 8631 11305
rect 9766 11296 9772 11308
rect 9824 11296 9830 11348
rect 10134 11296 10140 11348
rect 10192 11336 10198 11348
rect 10962 11336 10968 11348
rect 10192 11308 10968 11336
rect 10192 11296 10198 11308
rect 10962 11296 10968 11308
rect 11020 11296 11026 11348
rect 11054 11296 11060 11348
rect 11112 11336 11118 11348
rect 11241 11339 11299 11345
rect 11241 11336 11253 11339
rect 11112 11308 11253 11336
rect 11112 11296 11118 11308
rect 11241 11305 11253 11308
rect 11287 11305 11299 11339
rect 11241 11299 11299 11305
rect 11701 11339 11759 11345
rect 11701 11305 11713 11339
rect 11747 11336 11759 11339
rect 12253 11339 12311 11345
rect 12253 11336 12265 11339
rect 11747 11308 12265 11336
rect 11747 11305 11759 11308
rect 11701 11299 11759 11305
rect 12253 11305 12265 11308
rect 12299 11305 12311 11339
rect 12253 11299 12311 11305
rect 12897 11339 12955 11345
rect 12897 11305 12909 11339
rect 12943 11336 12955 11339
rect 13170 11336 13176 11348
rect 12943 11308 13176 11336
rect 12943 11305 12955 11308
rect 12897 11299 12955 11305
rect 13170 11296 13176 11308
rect 13228 11336 13234 11348
rect 13354 11336 13360 11348
rect 13228 11308 13360 11336
rect 13228 11296 13234 11308
rect 13354 11296 13360 11308
rect 13412 11296 13418 11348
rect 13449 11339 13507 11345
rect 13449 11305 13461 11339
rect 13495 11336 13507 11339
rect 13814 11336 13820 11348
rect 13495 11308 13820 11336
rect 13495 11305 13507 11308
rect 13449 11299 13507 11305
rect 13814 11296 13820 11308
rect 13872 11296 13878 11348
rect 14918 11296 14924 11348
rect 14976 11336 14982 11348
rect 17678 11336 17684 11348
rect 14976 11308 17684 11336
rect 14976 11296 14982 11308
rect 17678 11296 17684 11308
rect 17736 11336 17742 11348
rect 17957 11339 18015 11345
rect 17957 11336 17969 11339
rect 17736 11308 17969 11336
rect 17736 11296 17742 11308
rect 17957 11305 17969 11308
rect 18003 11305 18015 11339
rect 17957 11299 18015 11305
rect 3326 11228 3332 11280
rect 3384 11268 3390 11280
rect 3881 11271 3939 11277
rect 3881 11268 3893 11271
rect 3384 11240 3893 11268
rect 3384 11228 3390 11240
rect 3881 11237 3893 11240
rect 3927 11237 3939 11271
rect 3881 11231 3939 11237
rect 6580 11271 6638 11277
rect 6580 11237 6592 11271
rect 6626 11268 6638 11271
rect 6626 11240 7788 11268
rect 6626 11237 6638 11240
rect 6580 11231 6638 11237
rect 1486 11200 1492 11212
rect 1447 11172 1492 11200
rect 1486 11160 1492 11172
rect 1544 11160 1550 11212
rect 1854 11200 1860 11212
rect 1815 11172 1860 11200
rect 1854 11160 1860 11172
rect 1912 11160 1918 11212
rect 3142 11160 3148 11212
rect 3200 11200 3206 11212
rect 3430 11203 3488 11209
rect 3430 11200 3442 11203
rect 3200 11172 3442 11200
rect 3200 11160 3206 11172
rect 3430 11169 3442 11172
rect 3476 11169 3488 11203
rect 3430 11163 3488 11169
rect 4816 11172 7512 11200
rect 1504 11132 1532 11160
rect 2133 11135 2191 11141
rect 2133 11132 2145 11135
rect 1504 11104 2145 11132
rect 2133 11101 2145 11104
rect 2179 11101 2191 11135
rect 2133 11095 2191 11101
rect 3697 11135 3755 11141
rect 3697 11101 3709 11135
rect 3743 11132 3755 11135
rect 3786 11132 3792 11144
rect 3743 11104 3792 11132
rect 3743 11101 3755 11104
rect 3697 11095 3755 11101
rect 3786 11092 3792 11104
rect 3844 11092 3850 11144
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11132 4215 11135
rect 4522 11132 4528 11144
rect 4203 11104 4528 11132
rect 4203 11101 4215 11104
rect 4157 11095 4215 11101
rect 4522 11092 4528 11104
rect 4580 11092 4586 11144
rect 4706 11092 4712 11144
rect 4764 11132 4770 11144
rect 4816 11141 4844 11172
rect 4801 11135 4859 11141
rect 4801 11132 4813 11135
rect 4764 11104 4813 11132
rect 4764 11092 4770 11104
rect 4801 11101 4813 11104
rect 4847 11101 4859 11135
rect 4801 11095 4859 11101
rect 6822 11092 6828 11144
rect 6880 11132 6886 11144
rect 6880 11104 6925 11132
rect 6880 11092 6886 11104
rect 1578 11024 1584 11076
rect 1636 11064 1642 11076
rect 1673 11067 1731 11073
rect 1673 11064 1685 11067
rect 1636 11036 1685 11064
rect 1636 11024 1642 11036
rect 1673 11033 1685 11036
rect 1719 11033 1731 11067
rect 4338 11064 4344 11076
rect 4299 11036 4344 11064
rect 1673 11027 1731 11033
rect 4338 11024 4344 11036
rect 4396 11024 4402 11076
rect 4430 11024 4436 11076
rect 4488 11064 4494 11076
rect 5445 11067 5503 11073
rect 4488 11036 4533 11064
rect 4488 11024 4494 11036
rect 5445 11033 5457 11067
rect 5491 11064 5503 11067
rect 5718 11064 5724 11076
rect 5491 11036 5724 11064
rect 5491 11033 5503 11036
rect 5445 11027 5503 11033
rect 5718 11024 5724 11036
rect 5776 11024 5782 11076
rect 7484 11064 7512 11172
rect 7558 11092 7564 11144
rect 7616 11132 7622 11144
rect 7760 11141 7788 11240
rect 8202 11228 8208 11280
rect 8260 11228 8266 11280
rect 8754 11228 8760 11280
rect 8812 11268 8818 11280
rect 8812 11240 9674 11268
rect 8812 11228 8818 11240
rect 8220 11200 8248 11228
rect 9306 11200 9312 11212
rect 8220 11172 8340 11200
rect 9267 11172 9312 11200
rect 7745 11135 7803 11141
rect 7745 11132 7757 11135
rect 7616 11104 7757 11132
rect 7616 11092 7622 11104
rect 7745 11101 7757 11104
rect 7791 11101 7803 11135
rect 7745 11095 7803 11101
rect 8113 11135 8171 11141
rect 8113 11101 8125 11135
rect 8159 11132 8171 11135
rect 8202 11132 8208 11144
rect 8159 11104 8208 11132
rect 8159 11101 8171 11104
rect 8113 11095 8171 11101
rect 8202 11092 8208 11104
rect 8260 11092 8266 11144
rect 8312 11141 8340 11172
rect 9306 11160 9312 11172
rect 9364 11160 9370 11212
rect 9646 11200 9674 11240
rect 9876 11240 11192 11268
rect 9876 11200 9904 11240
rect 9646 11172 9904 11200
rect 8297 11135 8355 11141
rect 8297 11101 8309 11135
rect 8343 11101 8355 11135
rect 8478 11132 8484 11144
rect 8439 11104 8484 11132
rect 8297 11095 8355 11101
rect 8478 11092 8484 11104
rect 8536 11092 8542 11144
rect 9122 11132 9128 11144
rect 9083 11104 9128 11132
rect 9122 11092 9128 11104
rect 9180 11092 9186 11144
rect 9214 11092 9220 11144
rect 9272 11132 9278 11144
rect 9766 11132 9772 11144
rect 9272 11104 9772 11132
rect 9272 11092 9278 11104
rect 9766 11092 9772 11104
rect 9824 11092 9830 11144
rect 8754 11064 8760 11076
rect 7484 11036 8760 11064
rect 8754 11024 8760 11036
rect 8812 11024 8818 11076
rect 8941 11067 8999 11073
rect 8941 11033 8953 11067
rect 8987 11064 8999 11067
rect 9398 11064 9404 11076
rect 8987 11036 9404 11064
rect 8987 11033 8999 11036
rect 8941 11027 8999 11033
rect 9398 11024 9404 11036
rect 9456 11024 9462 11076
rect 9493 11067 9551 11073
rect 9493 11033 9505 11067
rect 9539 11064 9551 11067
rect 9876 11064 9904 11172
rect 10594 11160 10600 11212
rect 10652 11209 10658 11212
rect 10652 11200 10664 11209
rect 10652 11172 11100 11200
rect 10652 11163 10664 11172
rect 10652 11160 10658 11163
rect 11072 11141 11100 11172
rect 10873 11135 10931 11141
rect 10873 11101 10885 11135
rect 10919 11101 10931 11135
rect 10873 11095 10931 11101
rect 11057 11135 11115 11141
rect 11057 11101 11069 11135
rect 11103 11101 11115 11135
rect 11164 11132 11192 11240
rect 11422 11228 11428 11280
rect 11480 11268 11486 11280
rect 12161 11271 12219 11277
rect 12161 11268 12173 11271
rect 11480 11240 12173 11268
rect 11480 11228 11486 11240
rect 12161 11237 12173 11240
rect 12207 11237 12219 11271
rect 12161 11231 12219 11237
rect 12618 11228 12624 11280
rect 12676 11268 12682 11280
rect 14093 11271 14151 11277
rect 14093 11268 14105 11271
rect 12676 11240 14105 11268
rect 12676 11228 12682 11240
rect 14093 11237 14105 11240
rect 14139 11268 14151 11271
rect 14461 11271 14519 11277
rect 14461 11268 14473 11271
rect 14139 11240 14473 11268
rect 14139 11237 14151 11240
rect 14093 11231 14151 11237
rect 14461 11237 14473 11240
rect 14507 11268 14519 11271
rect 14550 11268 14556 11280
rect 14507 11240 14556 11268
rect 14507 11237 14519 11240
rect 14461 11231 14519 11237
rect 14550 11228 14556 11240
rect 14608 11268 14614 11280
rect 17770 11268 17776 11280
rect 14608 11240 17776 11268
rect 14608 11228 14614 11240
rect 17770 11228 17776 11240
rect 17828 11228 17834 11280
rect 18966 11268 18972 11280
rect 18927 11240 18972 11268
rect 18966 11228 18972 11240
rect 19024 11228 19030 11280
rect 11330 11200 11336 11212
rect 11291 11172 11336 11200
rect 11330 11160 11336 11172
rect 11388 11160 11394 11212
rect 12066 11160 12072 11212
rect 12124 11200 12130 11212
rect 14829 11203 14887 11209
rect 14829 11200 14841 11203
rect 12124 11172 14841 11200
rect 12124 11160 12130 11172
rect 14829 11169 14841 11172
rect 14875 11169 14887 11203
rect 14829 11163 14887 11169
rect 15194 11160 15200 11212
rect 15252 11200 15258 11212
rect 15361 11203 15419 11209
rect 15361 11200 15373 11203
rect 15252 11172 15373 11200
rect 15252 11160 15258 11172
rect 15361 11169 15373 11172
rect 15407 11169 15419 11203
rect 15361 11163 15419 11169
rect 16482 11160 16488 11212
rect 16540 11160 16546 11212
rect 16758 11200 16764 11212
rect 16719 11172 16764 11200
rect 16758 11160 16764 11172
rect 16816 11160 16822 11212
rect 17034 11200 17040 11212
rect 16995 11172 17040 11200
rect 17034 11160 17040 11172
rect 17092 11160 17098 11212
rect 17402 11200 17408 11212
rect 17363 11172 17408 11200
rect 17402 11160 17408 11172
rect 17460 11160 17466 11212
rect 17865 11203 17923 11209
rect 17865 11169 17877 11203
rect 17911 11200 17923 11203
rect 18325 11203 18383 11209
rect 18325 11200 18337 11203
rect 17911 11172 18337 11200
rect 17911 11169 17923 11172
rect 17865 11163 17923 11169
rect 18325 11169 18337 11172
rect 18371 11169 18383 11203
rect 18325 11163 18383 11169
rect 12345 11135 12403 11141
rect 12345 11132 12357 11135
rect 11164 11104 12357 11132
rect 11057 11095 11115 11101
rect 12345 11101 12357 11104
rect 12391 11101 12403 11135
rect 12345 11095 12403 11101
rect 9539 11036 9904 11064
rect 10888 11064 10916 11095
rect 12526 11092 12532 11144
rect 12584 11132 12590 11144
rect 12989 11135 13047 11141
rect 12989 11132 13001 11135
rect 12584 11104 13001 11132
rect 12584 11092 12590 11104
rect 12989 11101 13001 11104
rect 13035 11132 13047 11135
rect 13541 11135 13599 11141
rect 13541 11132 13553 11135
rect 13035 11104 13553 11132
rect 13035 11101 13047 11104
rect 12989 11095 13047 11101
rect 13541 11101 13553 11104
rect 13587 11132 13599 11135
rect 13906 11132 13912 11144
rect 13587 11104 13912 11132
rect 13587 11101 13599 11104
rect 13541 11095 13599 11101
rect 13906 11092 13912 11104
rect 13964 11092 13970 11144
rect 14182 11092 14188 11144
rect 14240 11132 14246 11144
rect 14645 11135 14703 11141
rect 14645 11132 14657 11135
rect 14240 11104 14657 11132
rect 14240 11092 14246 11104
rect 14645 11101 14657 11104
rect 14691 11101 14703 11135
rect 14645 11095 14703 11101
rect 15105 11135 15163 11141
rect 15105 11101 15117 11135
rect 15151 11101 15163 11135
rect 16500 11132 16528 11160
rect 18138 11132 18144 11144
rect 16500 11104 17264 11132
rect 18099 11104 18144 11132
rect 15105 11095 15163 11101
rect 11606 11064 11612 11076
rect 10888 11036 11612 11064
rect 9539 11033 9551 11036
rect 9493 11027 9551 11033
rect 11606 11024 11612 11036
rect 11664 11024 11670 11076
rect 11790 11064 11796 11076
rect 11751 11036 11796 11064
rect 11790 11024 11796 11036
rect 11848 11024 11854 11076
rect 12621 11067 12679 11073
rect 12621 11064 12633 11067
rect 12544 11036 12633 11064
rect 1946 10996 1952 11008
rect 1907 10968 1952 10996
rect 1946 10956 1952 10968
rect 2004 10956 2010 11008
rect 2222 10956 2228 11008
rect 2280 10996 2286 11008
rect 2317 10999 2375 11005
rect 2317 10996 2329 10999
rect 2280 10968 2329 10996
rect 2280 10956 2286 10968
rect 2317 10965 2329 10968
rect 2363 10996 2375 10999
rect 2682 10996 2688 11008
rect 2363 10968 2688 10996
rect 2363 10965 2375 10968
rect 2317 10959 2375 10965
rect 2682 10956 2688 10968
rect 2740 10956 2746 11008
rect 4709 10999 4767 11005
rect 4709 10965 4721 10999
rect 4755 10996 4767 10999
rect 4798 10996 4804 11008
rect 4755 10968 4804 10996
rect 4755 10965 4767 10968
rect 4709 10959 4767 10965
rect 4798 10956 4804 10968
rect 4856 10956 4862 11008
rect 5074 10996 5080 11008
rect 5035 10968 5080 10996
rect 5074 10956 5080 10968
rect 5132 10956 5138 11008
rect 6454 10956 6460 11008
rect 6512 10996 6518 11008
rect 6822 10996 6828 11008
rect 6512 10968 6828 10996
rect 6512 10956 6518 10968
rect 6822 10956 6828 10968
rect 6880 10956 6886 11008
rect 7009 10999 7067 11005
rect 7009 10965 7021 10999
rect 7055 10996 7067 10999
rect 7282 10996 7288 11008
rect 7055 10968 7288 10996
rect 7055 10965 7067 10968
rect 7009 10959 7067 10965
rect 7282 10956 7288 10968
rect 7340 10956 7346 11008
rect 7834 10956 7840 11008
rect 7892 10996 7898 11008
rect 11422 10996 11428 11008
rect 7892 10968 11428 10996
rect 7892 10956 7898 10968
rect 11422 10956 11428 10968
rect 11480 10956 11486 11008
rect 11698 10956 11704 11008
rect 11756 10996 11762 11008
rect 12342 10996 12348 11008
rect 11756 10968 12348 10996
rect 11756 10956 11762 10968
rect 12342 10956 12348 10968
rect 12400 10996 12406 11008
rect 12544 10996 12572 11036
rect 12621 11033 12633 11036
rect 12667 11033 12679 11067
rect 13262 11064 13268 11076
rect 13223 11036 13268 11064
rect 12621 11027 12679 11033
rect 13262 11024 13268 11036
rect 13320 11024 13326 11076
rect 13446 11024 13452 11076
rect 13504 11064 13510 11076
rect 14001 11067 14059 11073
rect 14001 11064 14013 11067
rect 13504 11036 14013 11064
rect 13504 11024 13510 11036
rect 14001 11033 14013 11036
rect 14047 11064 14059 11067
rect 15010 11064 15016 11076
rect 14047 11036 14872 11064
rect 14971 11036 15016 11064
rect 14047 11033 14059 11036
rect 14001 11027 14059 11033
rect 12400 10968 12572 10996
rect 13817 10999 13875 11005
rect 12400 10956 12406 10968
rect 13817 10965 13829 10999
rect 13863 10996 13875 10999
rect 14090 10996 14096 11008
rect 13863 10968 14096 10996
rect 13863 10965 13875 10968
rect 13817 10959 13875 10965
rect 14090 10956 14096 10968
rect 14148 10956 14154 11008
rect 14844 10996 14872 11036
rect 15010 11024 15016 11036
rect 15068 11064 15074 11076
rect 15120 11064 15148 11095
rect 16390 11064 16396 11076
rect 15068 11036 15148 11064
rect 16040 11036 16396 11064
rect 15068 11024 15074 11036
rect 16040 10996 16068 11036
rect 16390 11024 16396 11036
rect 16448 11024 16454 11076
rect 16577 11067 16635 11073
rect 16577 11033 16589 11067
rect 16623 11064 16635 11067
rect 16666 11064 16672 11076
rect 16623 11036 16672 11064
rect 16623 11033 16635 11036
rect 16577 11027 16635 11033
rect 16666 11024 16672 11036
rect 16724 11024 16730 11076
rect 17236 11073 17264 11104
rect 18138 11092 18144 11104
rect 18196 11092 18202 11144
rect 17221 11067 17279 11073
rect 17221 11033 17233 11067
rect 17267 11033 17279 11067
rect 17221 11027 17279 11033
rect 17497 11067 17555 11073
rect 17497 11033 17509 11067
rect 17543 11064 17555 11067
rect 17678 11064 17684 11076
rect 17543 11036 17684 11064
rect 17543 11033 17555 11036
rect 17497 11027 17555 11033
rect 17678 11024 17684 11036
rect 17736 11024 17742 11076
rect 16482 10996 16488 11008
rect 14844 10968 16068 10996
rect 16443 10968 16488 10996
rect 16482 10956 16488 10968
rect 16540 10956 16546 11008
rect 16850 10956 16856 11008
rect 16908 10996 16914 11008
rect 16908 10968 16953 10996
rect 16908 10956 16914 10968
rect 1104 10906 18860 10928
rect 1104 10854 3947 10906
rect 3999 10854 4011 10906
rect 4063 10854 4075 10906
rect 4127 10854 4139 10906
rect 4191 10854 9878 10906
rect 9930 10854 9942 10906
rect 9994 10854 10006 10906
rect 10058 10854 10070 10906
rect 10122 10854 15808 10906
rect 15860 10854 15872 10906
rect 15924 10854 15936 10906
rect 15988 10854 16000 10906
rect 16052 10854 18860 10906
rect 1104 10832 18860 10854
rect 2314 10792 2320 10804
rect 2275 10764 2320 10792
rect 2314 10752 2320 10764
rect 2372 10752 2378 10804
rect 2498 10752 2504 10804
rect 2556 10792 2562 10804
rect 5994 10792 6000 10804
rect 2556 10764 6000 10792
rect 2556 10752 2562 10764
rect 5994 10752 6000 10764
rect 6052 10792 6058 10804
rect 6178 10792 6184 10804
rect 6052 10764 6184 10792
rect 6052 10752 6058 10764
rect 6178 10752 6184 10764
rect 6236 10752 6242 10804
rect 6288 10764 7420 10792
rect 2225 10727 2283 10733
rect 2225 10693 2237 10727
rect 2271 10724 2283 10727
rect 2406 10724 2412 10736
rect 2271 10696 2412 10724
rect 2271 10693 2283 10696
rect 2225 10687 2283 10693
rect 2406 10684 2412 10696
rect 2464 10684 2470 10736
rect 4065 10727 4123 10733
rect 4065 10724 4077 10727
rect 3896 10696 4077 10724
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 2961 10659 3019 10665
rect 2961 10656 2973 10659
rect 1719 10628 2973 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 2961 10625 2973 10628
rect 3007 10656 3019 10659
rect 3142 10656 3148 10668
rect 3007 10628 3148 10656
rect 3007 10625 3019 10628
rect 2961 10619 3019 10625
rect 3142 10616 3148 10628
rect 3200 10656 3206 10668
rect 3896 10665 3924 10696
rect 4065 10693 4077 10696
rect 4111 10693 4123 10727
rect 4065 10687 4123 10693
rect 5442 10684 5448 10736
rect 5500 10724 5506 10736
rect 6288 10724 6316 10764
rect 5500 10696 6316 10724
rect 7392 10724 7420 10764
rect 7466 10752 7472 10804
rect 7524 10792 7530 10804
rect 7929 10795 7987 10801
rect 7929 10792 7941 10795
rect 7524 10764 7941 10792
rect 7524 10752 7530 10764
rect 7929 10761 7941 10764
rect 7975 10761 7987 10795
rect 7929 10755 7987 10761
rect 8478 10752 8484 10804
rect 8536 10792 8542 10804
rect 9493 10795 9551 10801
rect 9493 10792 9505 10795
rect 8536 10764 9505 10792
rect 8536 10752 8542 10764
rect 9493 10761 9505 10764
rect 9539 10761 9551 10795
rect 9493 10755 9551 10761
rect 9674 10752 9680 10804
rect 9732 10792 9738 10804
rect 10318 10792 10324 10804
rect 9732 10764 10324 10792
rect 9732 10752 9738 10764
rect 10318 10752 10324 10764
rect 10376 10752 10382 10804
rect 11974 10792 11980 10804
rect 11935 10764 11980 10792
rect 11974 10752 11980 10764
rect 12032 10752 12038 10804
rect 14366 10792 14372 10804
rect 12268 10764 14372 10792
rect 7392 10696 8616 10724
rect 5500 10684 5506 10696
rect 3881 10659 3939 10665
rect 3881 10656 3893 10659
rect 3200 10628 3893 10656
rect 3200 10616 3206 10628
rect 3881 10625 3893 10628
rect 3927 10625 3939 10659
rect 5718 10656 5724 10668
rect 5631 10628 5724 10656
rect 3881 10619 3939 10625
rect 5718 10616 5724 10628
rect 5776 10656 5782 10668
rect 5776 10628 6592 10656
rect 5776 10616 5782 10628
rect 6564 10600 6592 10628
rect 7558 10616 7564 10668
rect 7616 10656 7622 10668
rect 8481 10659 8539 10665
rect 8481 10656 8493 10659
rect 7616 10628 8493 10656
rect 7616 10616 7622 10628
rect 8481 10625 8493 10628
rect 8527 10625 8539 10659
rect 8588 10656 8616 10696
rect 8662 10684 8668 10736
rect 8720 10724 8726 10736
rect 8941 10727 8999 10733
rect 8941 10724 8953 10727
rect 8720 10696 8953 10724
rect 8720 10684 8726 10696
rect 8941 10693 8953 10696
rect 8987 10693 8999 10727
rect 9122 10724 9128 10736
rect 9083 10696 9128 10724
rect 8941 10687 8999 10693
rect 9122 10684 9128 10696
rect 9180 10684 9186 10736
rect 11330 10724 11336 10736
rect 9646 10696 11336 10724
rect 9214 10656 9220 10668
rect 8588 10628 9220 10656
rect 8481 10619 8539 10625
rect 9214 10616 9220 10628
rect 9272 10616 9278 10668
rect 1857 10591 1915 10597
rect 1857 10557 1869 10591
rect 1903 10588 1915 10591
rect 3234 10588 3240 10600
rect 1903 10560 3240 10588
rect 1903 10557 1915 10560
rect 1857 10551 1915 10557
rect 3234 10548 3240 10560
rect 3292 10548 3298 10600
rect 3786 10548 3792 10600
rect 3844 10588 3850 10600
rect 5442 10588 5448 10600
rect 3844 10560 5448 10588
rect 3844 10548 3850 10560
rect 5442 10548 5448 10560
rect 5500 10548 5506 10600
rect 6178 10588 6184 10600
rect 5828 10560 6184 10588
rect 1765 10523 1823 10529
rect 1765 10489 1777 10523
rect 1811 10520 1823 10523
rect 2498 10520 2504 10532
rect 1811 10492 2504 10520
rect 1811 10489 1823 10492
rect 1765 10483 1823 10489
rect 2498 10480 2504 10492
rect 2556 10480 2562 10532
rect 2590 10480 2596 10532
rect 2648 10520 2654 10532
rect 2685 10523 2743 10529
rect 2685 10520 2697 10523
rect 2648 10492 2697 10520
rect 2648 10480 2654 10492
rect 2685 10489 2697 10492
rect 2731 10489 2743 10523
rect 2685 10483 2743 10489
rect 2777 10523 2835 10529
rect 2777 10489 2789 10523
rect 2823 10520 2835 10523
rect 2866 10520 2872 10532
rect 2823 10492 2872 10520
rect 2823 10489 2835 10492
rect 2777 10483 2835 10489
rect 2866 10480 2872 10492
rect 2924 10480 2930 10532
rect 3697 10523 3755 10529
rect 3697 10489 3709 10523
rect 3743 10520 3755 10523
rect 4246 10520 4252 10532
rect 3743 10492 4252 10520
rect 3743 10489 3755 10492
rect 3697 10483 3755 10489
rect 4246 10480 4252 10492
rect 4304 10480 4310 10532
rect 4890 10480 4896 10532
rect 4948 10520 4954 10532
rect 5178 10523 5236 10529
rect 5178 10520 5190 10523
rect 4948 10492 5190 10520
rect 4948 10480 4954 10492
rect 5178 10489 5190 10492
rect 5224 10489 5236 10523
rect 5828 10520 5856 10560
rect 6178 10548 6184 10560
rect 6236 10548 6242 10600
rect 6454 10588 6460 10600
rect 6415 10560 6460 10588
rect 6454 10548 6460 10560
rect 6512 10548 6518 10600
rect 6546 10548 6552 10600
rect 6604 10588 6610 10600
rect 6713 10591 6771 10597
rect 6713 10588 6725 10591
rect 6604 10560 6725 10588
rect 6604 10548 6610 10560
rect 6713 10557 6725 10560
rect 6759 10557 6771 10591
rect 6713 10551 6771 10557
rect 8202 10548 8208 10600
rect 8260 10588 8266 10600
rect 8297 10591 8355 10597
rect 8297 10588 8309 10591
rect 8260 10560 8309 10588
rect 8260 10548 8266 10560
rect 8297 10557 8309 10560
rect 8343 10588 8355 10591
rect 8386 10588 8392 10600
rect 8343 10560 8392 10588
rect 8343 10557 8355 10560
rect 8297 10551 8355 10557
rect 8386 10548 8392 10560
rect 8444 10588 8450 10600
rect 9646 10588 9674 10696
rect 11330 10684 11336 10696
rect 11388 10684 11394 10736
rect 11422 10684 11428 10736
rect 11480 10724 11486 10736
rect 12268 10724 12296 10764
rect 14366 10752 14372 10764
rect 14424 10752 14430 10804
rect 15105 10795 15163 10801
rect 15105 10761 15117 10795
rect 15151 10792 15163 10795
rect 15194 10792 15200 10804
rect 15151 10764 15200 10792
rect 15151 10761 15163 10764
rect 15105 10755 15163 10761
rect 15194 10752 15200 10764
rect 15252 10752 15258 10804
rect 16942 10752 16948 10804
rect 17000 10792 17006 10804
rect 17218 10792 17224 10804
rect 17000 10764 17224 10792
rect 17000 10752 17006 10764
rect 17218 10752 17224 10764
rect 17276 10752 17282 10804
rect 11480 10696 12296 10724
rect 11480 10684 11486 10696
rect 10134 10656 10140 10668
rect 10095 10628 10140 10656
rect 10134 10616 10140 10628
rect 10192 10656 10198 10668
rect 10594 10656 10600 10668
rect 10192 10628 10600 10656
rect 10192 10616 10198 10628
rect 10594 10616 10600 10628
rect 10652 10616 10658 10668
rect 10778 10616 10784 10668
rect 10836 10656 10842 10668
rect 10873 10659 10931 10665
rect 10873 10656 10885 10659
rect 10836 10628 10885 10656
rect 10836 10616 10842 10628
rect 10873 10625 10885 10628
rect 10919 10625 10931 10659
rect 10873 10619 10931 10625
rect 11054 10616 11060 10668
rect 11112 10656 11118 10668
rect 11698 10656 11704 10668
rect 11112 10628 11704 10656
rect 11112 10616 11118 10628
rect 11698 10616 11704 10628
rect 11756 10616 11762 10668
rect 8444 10560 9674 10588
rect 9953 10591 10011 10597
rect 8444 10548 8450 10560
rect 9953 10557 9965 10591
rect 9999 10588 10011 10591
rect 10318 10588 10324 10600
rect 9999 10560 10324 10588
rect 9999 10557 10011 10560
rect 9953 10551 10011 10557
rect 10318 10548 10324 10560
rect 10376 10548 10382 10600
rect 10689 10591 10747 10597
rect 10689 10557 10701 10591
rect 10735 10588 10747 10591
rect 11146 10588 11152 10600
rect 10735 10560 11152 10588
rect 10735 10557 10747 10560
rect 10689 10551 10747 10557
rect 11146 10548 11152 10560
rect 11204 10548 11210 10600
rect 11606 10548 11612 10600
rect 11664 10588 11670 10600
rect 12253 10591 12311 10597
rect 12253 10588 12265 10591
rect 11664 10560 12265 10588
rect 11664 10548 11670 10560
rect 12253 10557 12265 10560
rect 12299 10557 12311 10591
rect 12253 10551 12311 10557
rect 13725 10591 13783 10597
rect 13725 10557 13737 10591
rect 13771 10588 13783 10591
rect 15010 10588 15016 10600
rect 13771 10560 15016 10588
rect 13771 10557 13783 10560
rect 13725 10551 13783 10557
rect 15010 10548 15016 10560
rect 15068 10548 15074 10600
rect 16577 10591 16635 10597
rect 16577 10557 16589 10591
rect 16623 10588 16635 10591
rect 16942 10588 16948 10600
rect 16623 10560 16948 10588
rect 16623 10557 16635 10560
rect 16577 10551 16635 10557
rect 16942 10548 16948 10560
rect 17000 10548 17006 10600
rect 5178 10483 5236 10489
rect 5644 10492 5856 10520
rect 5905 10523 5963 10529
rect 3234 10452 3240 10464
rect 3195 10424 3240 10452
rect 3234 10412 3240 10424
rect 3292 10412 3298 10464
rect 3510 10412 3516 10464
rect 3568 10452 3574 10464
rect 3605 10455 3663 10461
rect 3605 10452 3617 10455
rect 3568 10424 3617 10452
rect 3568 10412 3574 10424
rect 3605 10421 3617 10424
rect 3651 10452 3663 10455
rect 5644 10452 5672 10492
rect 5905 10489 5917 10523
rect 5951 10520 5963 10523
rect 9674 10520 9680 10532
rect 5951 10492 6684 10520
rect 5951 10489 5963 10492
rect 5905 10483 5963 10489
rect 5810 10452 5816 10464
rect 3651 10424 5672 10452
rect 5771 10424 5816 10452
rect 3651 10421 3663 10424
rect 3605 10415 3663 10421
rect 5810 10412 5816 10424
rect 5868 10412 5874 10464
rect 6270 10452 6276 10464
rect 6231 10424 6276 10452
rect 6270 10412 6276 10424
rect 6328 10412 6334 10464
rect 6656 10452 6684 10492
rect 8404 10492 9680 10520
rect 7742 10452 7748 10464
rect 6656 10424 7748 10452
rect 7742 10412 7748 10424
rect 7800 10412 7806 10464
rect 7834 10412 7840 10464
rect 7892 10452 7898 10464
rect 8404 10461 8432 10492
rect 9674 10480 9680 10492
rect 9732 10480 9738 10532
rect 9858 10520 9864 10532
rect 9819 10492 9864 10520
rect 9858 10480 9864 10492
rect 9916 10480 9922 10532
rect 12526 10529 12532 10532
rect 12520 10520 12532 10529
rect 12487 10492 12532 10520
rect 12520 10483 12532 10492
rect 12526 10480 12532 10483
rect 12584 10480 12590 10532
rect 13992 10523 14050 10529
rect 13992 10520 14004 10523
rect 13648 10492 14004 10520
rect 8389 10455 8447 10461
rect 7892 10424 7937 10452
rect 7892 10412 7898 10424
rect 8389 10421 8401 10455
rect 8435 10421 8447 10455
rect 8754 10452 8760 10464
rect 8715 10424 8760 10452
rect 8389 10415 8447 10421
rect 8754 10412 8760 10424
rect 8812 10412 8818 10464
rect 9306 10452 9312 10464
rect 9267 10424 9312 10452
rect 9306 10412 9312 10424
rect 9364 10452 9370 10464
rect 10042 10452 10048 10464
rect 9364 10424 10048 10452
rect 9364 10412 9370 10424
rect 10042 10412 10048 10424
rect 10100 10412 10106 10464
rect 10321 10455 10379 10461
rect 10321 10421 10333 10455
rect 10367 10452 10379 10455
rect 10410 10452 10416 10464
rect 10367 10424 10416 10452
rect 10367 10421 10379 10424
rect 10321 10415 10379 10421
rect 10410 10412 10416 10424
rect 10468 10412 10474 10464
rect 10502 10412 10508 10464
rect 10560 10452 10566 10464
rect 10781 10455 10839 10461
rect 10781 10452 10793 10455
rect 10560 10424 10793 10452
rect 10560 10412 10566 10424
rect 10781 10421 10793 10424
rect 10827 10421 10839 10455
rect 10781 10415 10839 10421
rect 11241 10455 11299 10461
rect 11241 10421 11253 10455
rect 11287 10452 11299 10455
rect 11330 10452 11336 10464
rect 11287 10424 11336 10452
rect 11287 10421 11299 10424
rect 11241 10415 11299 10421
rect 11330 10412 11336 10424
rect 11388 10452 11394 10464
rect 11790 10452 11796 10464
rect 11388 10424 11796 10452
rect 11388 10412 11394 10424
rect 11790 10412 11796 10424
rect 11848 10412 11854 10464
rect 11974 10412 11980 10464
rect 12032 10452 12038 10464
rect 12069 10455 12127 10461
rect 12069 10452 12081 10455
rect 12032 10424 12081 10452
rect 12032 10412 12038 10424
rect 12069 10421 12081 10424
rect 12115 10452 12127 10455
rect 12250 10452 12256 10464
rect 12115 10424 12256 10452
rect 12115 10421 12127 10424
rect 12069 10415 12127 10421
rect 12250 10412 12256 10424
rect 12308 10412 12314 10464
rect 13648 10461 13676 10492
rect 13992 10489 14004 10492
rect 14038 10520 14050 10523
rect 14918 10520 14924 10532
rect 14038 10492 14924 10520
rect 14038 10489 14050 10492
rect 13992 10483 14050 10489
rect 14918 10480 14924 10492
rect 14976 10480 14982 10532
rect 15470 10480 15476 10532
rect 15528 10520 15534 10532
rect 16390 10529 16396 10532
rect 16332 10523 16396 10529
rect 15528 10492 15976 10520
rect 15528 10480 15534 10492
rect 13633 10455 13691 10461
rect 13633 10421 13645 10455
rect 13679 10421 13691 10455
rect 13633 10415 13691 10421
rect 15197 10455 15255 10461
rect 15197 10421 15209 10455
rect 15243 10452 15255 10455
rect 15654 10452 15660 10464
rect 15243 10424 15660 10452
rect 15243 10421 15255 10424
rect 15197 10415 15255 10421
rect 15654 10412 15660 10424
rect 15712 10412 15718 10464
rect 15948 10452 15976 10492
rect 16332 10489 16344 10523
rect 16378 10489 16396 10523
rect 16332 10483 16396 10489
rect 16390 10480 16396 10483
rect 16448 10480 16454 10532
rect 16482 10480 16488 10532
rect 16540 10520 16546 10532
rect 17190 10523 17248 10529
rect 17190 10520 17202 10523
rect 16540 10492 17202 10520
rect 16540 10480 16546 10492
rect 17190 10489 17202 10492
rect 17236 10489 17248 10523
rect 17190 10483 17248 10489
rect 16669 10455 16727 10461
rect 16669 10452 16681 10455
rect 15948 10424 16681 10452
rect 16669 10421 16681 10424
rect 16715 10452 16727 10455
rect 17034 10452 17040 10464
rect 16715 10424 17040 10452
rect 16715 10421 16727 10424
rect 16669 10415 16727 10421
rect 17034 10412 17040 10424
rect 17092 10412 17098 10464
rect 17862 10412 17868 10464
rect 17920 10452 17926 10464
rect 18325 10455 18383 10461
rect 18325 10452 18337 10455
rect 17920 10424 18337 10452
rect 17920 10412 17926 10424
rect 18325 10421 18337 10424
rect 18371 10421 18383 10455
rect 18506 10452 18512 10464
rect 18467 10424 18512 10452
rect 18325 10415 18383 10421
rect 18506 10412 18512 10424
rect 18564 10412 18570 10464
rect 1104 10362 18860 10384
rect 1104 10310 6912 10362
rect 6964 10310 6976 10362
rect 7028 10310 7040 10362
rect 7092 10310 7104 10362
rect 7156 10310 12843 10362
rect 12895 10310 12907 10362
rect 12959 10310 12971 10362
rect 13023 10310 13035 10362
rect 13087 10310 18860 10362
rect 1104 10288 18860 10310
rect 3237 10251 3295 10257
rect 3237 10217 3249 10251
rect 3283 10248 3295 10251
rect 4341 10251 4399 10257
rect 4341 10248 4353 10251
rect 3283 10220 4353 10248
rect 3283 10217 3295 10220
rect 3237 10211 3295 10217
rect 4341 10217 4353 10220
rect 4387 10217 4399 10251
rect 4798 10248 4804 10260
rect 4759 10220 4804 10248
rect 4341 10211 4399 10217
rect 4798 10208 4804 10220
rect 4856 10208 4862 10260
rect 5074 10208 5080 10260
rect 5132 10248 5138 10260
rect 5629 10251 5687 10257
rect 5629 10248 5641 10251
rect 5132 10220 5641 10248
rect 5132 10208 5138 10220
rect 5629 10217 5641 10220
rect 5675 10217 5687 10251
rect 5629 10211 5687 10217
rect 5902 10208 5908 10260
rect 5960 10248 5966 10260
rect 5997 10251 6055 10257
rect 5997 10248 6009 10251
rect 5960 10220 6009 10248
rect 5960 10208 5966 10220
rect 5997 10217 6009 10220
rect 6043 10217 6055 10251
rect 5997 10211 6055 10217
rect 6362 10208 6368 10260
rect 6420 10248 6426 10260
rect 6546 10248 6552 10260
rect 6420 10220 6552 10248
rect 6420 10208 6426 10220
rect 6546 10208 6552 10220
rect 6604 10208 6610 10260
rect 7009 10251 7067 10257
rect 7009 10217 7021 10251
rect 7055 10248 7067 10251
rect 7561 10251 7619 10257
rect 7561 10248 7573 10251
rect 7055 10220 7573 10248
rect 7055 10217 7067 10220
rect 7009 10211 7067 10217
rect 7561 10217 7573 10220
rect 7607 10217 7619 10251
rect 7561 10211 7619 10217
rect 7742 10208 7748 10260
rect 7800 10248 7806 10260
rect 7929 10251 7987 10257
rect 7929 10248 7941 10251
rect 7800 10220 7941 10248
rect 7800 10208 7806 10220
rect 7929 10217 7941 10220
rect 7975 10217 7987 10251
rect 7929 10211 7987 10217
rect 8297 10251 8355 10257
rect 8297 10217 8309 10251
rect 8343 10248 8355 10251
rect 8662 10248 8668 10260
rect 8343 10220 8668 10248
rect 8343 10217 8355 10220
rect 8297 10211 8355 10217
rect 8662 10208 8668 10220
rect 8720 10208 8726 10260
rect 9766 10248 9772 10260
rect 9727 10220 9772 10248
rect 9766 10208 9772 10220
rect 9824 10208 9830 10260
rect 10137 10251 10195 10257
rect 10137 10217 10149 10251
rect 10183 10248 10195 10251
rect 10226 10248 10232 10260
rect 10183 10220 10232 10248
rect 10183 10217 10195 10220
rect 10137 10211 10195 10217
rect 10226 10208 10232 10220
rect 10284 10208 10290 10260
rect 10410 10208 10416 10260
rect 10468 10248 10474 10260
rect 11698 10248 11704 10260
rect 10468 10220 11704 10248
rect 10468 10208 10474 10220
rect 11698 10208 11704 10220
rect 11756 10208 11762 10260
rect 13538 10248 13544 10260
rect 12360 10220 13544 10248
rect 3329 10183 3387 10189
rect 3329 10149 3341 10183
rect 3375 10180 3387 10183
rect 4249 10183 4307 10189
rect 4249 10180 4261 10183
rect 3375 10152 4261 10180
rect 3375 10149 3387 10152
rect 3329 10143 3387 10149
rect 4249 10149 4261 10152
rect 4295 10149 4307 10183
rect 5534 10180 5540 10192
rect 5495 10152 5540 10180
rect 4249 10143 4307 10149
rect 5534 10140 5540 10152
rect 5592 10140 5598 10192
rect 6086 10140 6092 10192
rect 6144 10180 6150 10192
rect 12360 10180 12388 10220
rect 13538 10208 13544 10220
rect 13596 10208 13602 10260
rect 14093 10251 14151 10257
rect 14093 10217 14105 10251
rect 14139 10248 14151 10251
rect 14737 10251 14795 10257
rect 14737 10248 14749 10251
rect 14139 10220 14749 10248
rect 14139 10217 14151 10220
rect 14093 10211 14151 10217
rect 14737 10217 14749 10220
rect 14783 10217 14795 10251
rect 14737 10211 14795 10217
rect 15286 10208 15292 10260
rect 15344 10248 15350 10260
rect 15565 10251 15623 10257
rect 15565 10248 15577 10251
rect 15344 10220 15577 10248
rect 15344 10208 15350 10220
rect 15565 10217 15577 10220
rect 15611 10217 15623 10251
rect 15565 10211 15623 10217
rect 15933 10251 15991 10257
rect 15933 10217 15945 10251
rect 15979 10248 15991 10251
rect 16577 10251 16635 10257
rect 16577 10248 16589 10251
rect 15979 10220 16589 10248
rect 15979 10217 15991 10220
rect 15933 10211 15991 10217
rect 16577 10217 16589 10220
rect 16623 10217 16635 10251
rect 16577 10211 16635 10217
rect 17034 10208 17040 10260
rect 17092 10248 17098 10260
rect 18141 10251 18199 10257
rect 18141 10248 18153 10251
rect 17092 10220 18153 10248
rect 17092 10208 17098 10220
rect 18141 10217 18153 10220
rect 18187 10217 18199 10251
rect 18141 10211 18199 10217
rect 6144 10152 10548 10180
rect 6144 10140 6150 10152
rect 2521 10115 2579 10121
rect 2521 10081 2533 10115
rect 2567 10112 2579 10115
rect 2682 10112 2688 10124
rect 2567 10084 2688 10112
rect 2567 10081 2579 10084
rect 2521 10075 2579 10081
rect 2682 10072 2688 10084
rect 2740 10072 2746 10124
rect 2777 10115 2835 10121
rect 2777 10081 2789 10115
rect 2823 10112 2835 10115
rect 3694 10112 3700 10124
rect 2823 10084 3700 10112
rect 2823 10081 2835 10084
rect 2777 10075 2835 10081
rect 3694 10072 3700 10084
rect 3752 10072 3758 10124
rect 3786 10072 3792 10124
rect 3844 10112 3850 10124
rect 3973 10115 4031 10121
rect 3973 10112 3985 10115
rect 3844 10084 3985 10112
rect 3844 10072 3850 10084
rect 3973 10081 3985 10084
rect 4019 10112 4031 10115
rect 4430 10112 4436 10124
rect 4019 10084 4436 10112
rect 4019 10081 4031 10084
rect 3973 10075 4031 10081
rect 4430 10072 4436 10084
rect 4488 10072 4494 10124
rect 4709 10115 4767 10121
rect 4709 10081 4721 10115
rect 4755 10112 4767 10115
rect 5626 10112 5632 10124
rect 4755 10084 5632 10112
rect 4755 10081 4767 10084
rect 4709 10075 4767 10081
rect 5626 10072 5632 10084
rect 5684 10112 5690 10124
rect 6638 10112 6644 10124
rect 5684 10084 6644 10112
rect 5684 10072 5690 10084
rect 6638 10072 6644 10084
rect 6696 10072 6702 10124
rect 7469 10115 7527 10121
rect 7469 10081 7481 10115
rect 7515 10112 7527 10115
rect 7515 10084 8607 10112
rect 7515 10081 7527 10084
rect 7469 10075 7527 10081
rect 3142 10044 3148 10056
rect 3103 10016 3148 10044
rect 3142 10004 3148 10016
rect 3200 10004 3206 10056
rect 4154 10044 4160 10056
rect 4115 10016 4160 10044
rect 4154 10004 4160 10016
rect 4212 10044 4218 10056
rect 4890 10044 4896 10056
rect 4212 10016 4752 10044
rect 4851 10016 4896 10044
rect 4212 10004 4218 10016
rect 4724 9988 4752 10016
rect 4890 10004 4896 10016
rect 4948 10004 4954 10056
rect 5534 10004 5540 10056
rect 5592 10044 5598 10056
rect 5721 10047 5779 10053
rect 5721 10044 5733 10047
rect 5592 10016 5733 10044
rect 5592 10004 5598 10016
rect 5721 10013 5733 10016
rect 5767 10013 5779 10047
rect 6362 10044 6368 10056
rect 6323 10016 6368 10044
rect 5721 10007 5779 10013
rect 6362 10004 6368 10016
rect 6420 10004 6426 10056
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10044 6607 10047
rect 6914 10044 6920 10056
rect 6595 10016 6920 10044
rect 6595 10013 6607 10016
rect 6549 10007 6607 10013
rect 6914 10004 6920 10016
rect 6972 10004 6978 10056
rect 4706 9936 4712 9988
rect 4764 9936 4770 9988
rect 5169 9979 5227 9985
rect 5169 9976 5181 9979
rect 4816 9948 5181 9976
rect 1394 9908 1400 9920
rect 1355 9880 1400 9908
rect 1394 9868 1400 9880
rect 1452 9868 1458 9920
rect 2130 9868 2136 9920
rect 2188 9908 2194 9920
rect 2958 9908 2964 9920
rect 2188 9880 2964 9908
rect 2188 9868 2194 9880
rect 2958 9868 2964 9880
rect 3016 9868 3022 9920
rect 3510 9868 3516 9920
rect 3568 9908 3574 9920
rect 3697 9911 3755 9917
rect 3697 9908 3709 9911
rect 3568 9880 3709 9908
rect 3568 9868 3574 9880
rect 3697 9877 3709 9880
rect 3743 9877 3755 9911
rect 3697 9871 3755 9877
rect 4249 9911 4307 9917
rect 4249 9877 4261 9911
rect 4295 9908 4307 9911
rect 4816 9908 4844 9948
rect 5169 9945 5181 9948
rect 5215 9945 5227 9979
rect 5169 9939 5227 9945
rect 5810 9936 5816 9988
rect 5868 9976 5874 9988
rect 7101 9979 7159 9985
rect 7101 9976 7113 9979
rect 5868 9948 7113 9976
rect 5868 9936 5874 9948
rect 7101 9945 7113 9948
rect 7147 9945 7159 9979
rect 7101 9939 7159 9945
rect 4295 9880 4844 9908
rect 4295 9877 4307 9880
rect 4249 9871 4307 9877
rect 5074 9868 5080 9920
rect 5132 9908 5138 9920
rect 7484 9908 7512 10075
rect 7558 10004 7564 10056
rect 7616 10044 7622 10056
rect 7653 10047 7711 10053
rect 7653 10044 7665 10047
rect 7616 10016 7665 10044
rect 7616 10004 7622 10016
rect 7653 10013 7665 10016
rect 7699 10013 7711 10047
rect 7653 10007 7711 10013
rect 7668 9976 7696 10007
rect 8018 10004 8024 10056
rect 8076 10044 8082 10056
rect 8389 10047 8447 10053
rect 8389 10044 8401 10047
rect 8076 10016 8401 10044
rect 8076 10004 8082 10016
rect 8389 10013 8401 10016
rect 8435 10013 8447 10047
rect 8389 10007 8447 10013
rect 8481 10047 8539 10053
rect 8481 10013 8493 10047
rect 8527 10013 8539 10047
rect 8579 10044 8607 10084
rect 8754 10072 8760 10124
rect 8812 10112 8818 10124
rect 8812 10084 8857 10112
rect 8812 10072 8818 10084
rect 9490 10072 9496 10124
rect 9548 10112 9554 10124
rect 10410 10112 10416 10124
rect 9548 10084 10416 10112
rect 9548 10072 9554 10084
rect 10410 10072 10416 10084
rect 10468 10072 10474 10124
rect 10520 10112 10548 10152
rect 10704 10152 12388 10180
rect 10704 10112 10732 10152
rect 17126 10140 17132 10192
rect 17184 10180 17190 10192
rect 17405 10183 17463 10189
rect 17405 10180 17417 10183
rect 17184 10152 17417 10180
rect 17184 10140 17190 10152
rect 17405 10149 17417 10152
rect 17451 10149 17463 10183
rect 17405 10143 17463 10149
rect 17494 10140 17500 10192
rect 17552 10140 17558 10192
rect 18230 10180 18236 10192
rect 18191 10152 18236 10180
rect 18230 10140 18236 10152
rect 18288 10140 18294 10192
rect 10520 10084 10732 10112
rect 10778 10072 10784 10124
rect 10836 10112 10842 10124
rect 11342 10115 11400 10121
rect 11342 10112 11354 10115
rect 10836 10084 11354 10112
rect 10836 10072 10842 10084
rect 11342 10081 11354 10084
rect 11388 10081 11400 10115
rect 11606 10112 11612 10124
rect 11567 10084 11612 10112
rect 11342 10075 11400 10081
rect 11606 10072 11612 10084
rect 11664 10112 11670 10124
rect 11885 10115 11943 10121
rect 11885 10112 11897 10115
rect 11664 10084 11897 10112
rect 11664 10072 11670 10084
rect 11885 10081 11897 10084
rect 11931 10081 11943 10115
rect 11885 10075 11943 10081
rect 12152 10115 12210 10121
rect 12152 10081 12164 10115
rect 12198 10112 12210 10115
rect 12618 10112 12624 10124
rect 12198 10084 12624 10112
rect 12198 10081 12210 10084
rect 12152 10075 12210 10081
rect 12618 10072 12624 10084
rect 12676 10072 12682 10124
rect 13725 10115 13783 10121
rect 13725 10081 13737 10115
rect 13771 10112 13783 10115
rect 14550 10112 14556 10124
rect 13771 10084 14556 10112
rect 13771 10081 13783 10084
rect 13725 10075 13783 10081
rect 14550 10072 14556 10084
rect 14608 10072 14614 10124
rect 14642 10072 14648 10124
rect 14700 10112 14706 10124
rect 16114 10112 16120 10124
rect 14700 10084 16120 10112
rect 14700 10072 14706 10084
rect 16114 10072 16120 10084
rect 16172 10112 16178 10124
rect 16485 10115 16543 10121
rect 16485 10112 16497 10115
rect 16172 10084 16497 10112
rect 16172 10072 16178 10084
rect 16485 10081 16497 10084
rect 16531 10081 16543 10115
rect 16485 10075 16543 10081
rect 16574 10072 16580 10124
rect 16632 10112 16638 10124
rect 17034 10112 17040 10124
rect 16632 10084 17040 10112
rect 16632 10072 16638 10084
rect 17034 10072 17040 10084
rect 17092 10072 17098 10124
rect 17313 10115 17371 10121
rect 17313 10081 17325 10115
rect 17359 10112 17371 10115
rect 17512 10112 17540 10140
rect 17770 10112 17776 10124
rect 17359 10084 17776 10112
rect 17359 10081 17371 10084
rect 17313 10075 17371 10081
rect 17770 10072 17776 10084
rect 17828 10072 17834 10124
rect 9125 10047 9183 10053
rect 9125 10044 9137 10047
rect 8579 10016 9137 10044
rect 8481 10007 8539 10013
rect 9125 10013 9137 10016
rect 9171 10044 9183 10047
rect 9306 10044 9312 10056
rect 9171 10016 9312 10044
rect 9171 10013 9183 10016
rect 9125 10007 9183 10013
rect 8496 9976 8524 10007
rect 9306 10004 9312 10016
rect 9364 10004 9370 10056
rect 9585 10047 9643 10053
rect 9585 10013 9597 10047
rect 9631 10013 9643 10047
rect 9585 10007 9643 10013
rect 9677 10047 9735 10053
rect 9677 10013 9689 10047
rect 9723 10044 9735 10047
rect 10502 10044 10508 10056
rect 9723 10016 10508 10044
rect 9723 10013 9735 10016
rect 9677 10007 9735 10013
rect 7668 9948 8524 9976
rect 9600 9976 9628 10007
rect 10502 10004 10508 10016
rect 10560 10004 10566 10056
rect 13449 10047 13507 10053
rect 13449 10044 13461 10047
rect 13280 10016 13461 10044
rect 9766 9976 9772 9988
rect 9600 9948 9772 9976
rect 9766 9936 9772 9948
rect 9824 9936 9830 9988
rect 10134 9936 10140 9988
rect 10192 9976 10198 9988
rect 10229 9979 10287 9985
rect 10229 9976 10241 9979
rect 10192 9948 10241 9976
rect 10192 9936 10198 9948
rect 10229 9945 10241 9948
rect 10275 9945 10287 9979
rect 10229 9939 10287 9945
rect 5132 9880 7512 9908
rect 5132 9868 5138 9880
rect 8294 9868 8300 9920
rect 8352 9908 8358 9920
rect 8941 9911 8999 9917
rect 8941 9908 8953 9911
rect 8352 9880 8953 9908
rect 8352 9868 8358 9880
rect 8941 9877 8953 9880
rect 8987 9908 8999 9911
rect 9122 9908 9128 9920
rect 8987 9880 9128 9908
rect 8987 9877 8999 9880
rect 8941 9871 8999 9877
rect 9122 9868 9128 9880
rect 9180 9868 9186 9920
rect 9214 9868 9220 9920
rect 9272 9908 9278 9920
rect 12250 9908 12256 9920
rect 9272 9880 12256 9908
rect 9272 9868 9278 9880
rect 12250 9868 12256 9880
rect 12308 9868 12314 9920
rect 12526 9868 12532 9920
rect 12584 9908 12590 9920
rect 13280 9917 13308 10016
rect 13449 10013 13461 10016
rect 13495 10013 13507 10047
rect 13630 10044 13636 10056
rect 13591 10016 13636 10044
rect 13449 10007 13507 10013
rect 13630 10004 13636 10016
rect 13688 10004 13694 10056
rect 13814 10004 13820 10056
rect 13872 10044 13878 10056
rect 14829 10047 14887 10053
rect 14829 10044 14841 10047
rect 13872 10016 14841 10044
rect 13872 10004 13878 10016
rect 14829 10013 14841 10016
rect 14875 10013 14887 10047
rect 14829 10007 14887 10013
rect 14918 10004 14924 10056
rect 14976 10044 14982 10056
rect 14976 10016 15021 10044
rect 14976 10004 14982 10016
rect 15194 10004 15200 10056
rect 15252 10044 15258 10056
rect 15289 10047 15347 10053
rect 15289 10044 15301 10047
rect 15252 10016 15301 10044
rect 15252 10004 15258 10016
rect 15289 10013 15301 10016
rect 15335 10013 15347 10047
rect 15289 10007 15347 10013
rect 15473 10047 15531 10053
rect 15473 10013 15485 10047
rect 15519 10013 15531 10047
rect 15473 10007 15531 10013
rect 16669 10047 16727 10053
rect 16669 10013 16681 10047
rect 16715 10044 16727 10047
rect 17497 10047 17555 10053
rect 17497 10044 17509 10047
rect 16715 10016 17509 10044
rect 16715 10013 16727 10016
rect 16669 10007 16727 10013
rect 17497 10013 17509 10016
rect 17543 10044 17555 10047
rect 18138 10044 18144 10056
rect 17543 10016 18144 10044
rect 17543 10013 17555 10016
rect 17497 10007 17555 10013
rect 14182 9936 14188 9988
rect 14240 9976 14246 9988
rect 15488 9976 15516 10007
rect 14240 9948 15516 9976
rect 14240 9936 14246 9948
rect 16482 9936 16488 9988
rect 16540 9976 16546 9988
rect 16684 9976 16712 10007
rect 18138 10004 18144 10016
rect 18196 10044 18202 10056
rect 18325 10047 18383 10053
rect 18325 10044 18337 10047
rect 18196 10016 18337 10044
rect 18196 10004 18202 10016
rect 18325 10013 18337 10016
rect 18371 10013 18383 10047
rect 18325 10007 18383 10013
rect 16540 9948 16712 9976
rect 16540 9936 16546 9948
rect 17402 9936 17408 9988
rect 17460 9976 17466 9988
rect 18230 9976 18236 9988
rect 17460 9948 18236 9976
rect 17460 9936 17466 9948
rect 18230 9936 18236 9948
rect 18288 9936 18294 9988
rect 13265 9911 13323 9917
rect 13265 9908 13277 9911
rect 12584 9880 13277 9908
rect 12584 9868 12590 9880
rect 13265 9877 13277 9880
rect 13311 9877 13323 9911
rect 13265 9871 13323 9877
rect 14369 9911 14427 9917
rect 14369 9877 14381 9911
rect 14415 9908 14427 9911
rect 14458 9908 14464 9920
rect 14415 9880 14464 9908
rect 14415 9877 14427 9880
rect 14369 9871 14427 9877
rect 14458 9868 14464 9880
rect 14516 9868 14522 9920
rect 16114 9908 16120 9920
rect 16075 9880 16120 9908
rect 16114 9868 16120 9880
rect 16172 9868 16178 9920
rect 16574 9868 16580 9920
rect 16632 9908 16638 9920
rect 16945 9911 17003 9917
rect 16945 9908 16957 9911
rect 16632 9880 16957 9908
rect 16632 9868 16638 9880
rect 16945 9877 16957 9880
rect 16991 9877 17003 9911
rect 17770 9908 17776 9920
rect 17731 9880 17776 9908
rect 16945 9871 17003 9877
rect 17770 9868 17776 9880
rect 17828 9868 17834 9920
rect 1104 9818 18860 9840
rect 1104 9766 3947 9818
rect 3999 9766 4011 9818
rect 4063 9766 4075 9818
rect 4127 9766 4139 9818
rect 4191 9766 9878 9818
rect 9930 9766 9942 9818
rect 9994 9766 10006 9818
rect 10058 9766 10070 9818
rect 10122 9766 15808 9818
rect 15860 9766 15872 9818
rect 15924 9766 15936 9818
rect 15988 9766 16000 9818
rect 16052 9766 18860 9818
rect 1104 9744 18860 9766
rect 1394 9664 1400 9716
rect 1452 9704 1458 9716
rect 2866 9704 2872 9716
rect 1452 9676 2872 9704
rect 1452 9664 1458 9676
rect 1765 9639 1823 9645
rect 1765 9605 1777 9639
rect 1811 9636 1823 9639
rect 2222 9636 2228 9648
rect 1811 9608 2228 9636
rect 1811 9605 1823 9608
rect 1765 9599 1823 9605
rect 2222 9596 2228 9608
rect 2280 9596 2286 9648
rect 2332 9577 2360 9676
rect 2866 9664 2872 9676
rect 2924 9664 2930 9716
rect 3053 9707 3111 9713
rect 3053 9673 3065 9707
rect 3099 9673 3111 9707
rect 4890 9704 4896 9716
rect 3053 9667 3111 9673
rect 4816 9676 4896 9704
rect 2317 9571 2375 9577
rect 2317 9537 2329 9571
rect 2363 9537 2375 9571
rect 2317 9531 2375 9537
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9568 2559 9571
rect 3068 9568 3096 9667
rect 4157 9639 4215 9645
rect 2547 9540 3096 9568
rect 3160 9608 3648 9636
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 2130 9500 2136 9512
rect 2091 9472 2136 9500
rect 2130 9460 2136 9472
rect 2188 9460 2194 9512
rect 2593 9503 2651 9509
rect 2593 9469 2605 9503
rect 2639 9500 2651 9503
rect 2774 9500 2780 9512
rect 2639 9472 2780 9500
rect 2639 9469 2651 9472
rect 2593 9463 2651 9469
rect 2774 9460 2780 9472
rect 2832 9460 2838 9512
rect 3160 9500 3188 9608
rect 3510 9568 3516 9580
rect 3471 9540 3516 9568
rect 3510 9528 3516 9540
rect 3568 9528 3574 9580
rect 3620 9577 3648 9608
rect 4157 9605 4169 9639
rect 4203 9636 4215 9639
rect 4246 9636 4252 9648
rect 4203 9608 4252 9636
rect 4203 9605 4215 9608
rect 4157 9599 4215 9605
rect 4246 9596 4252 9608
rect 4304 9596 4310 9648
rect 3605 9571 3663 9577
rect 3605 9537 3617 9571
rect 3651 9537 3663 9571
rect 4430 9568 4436 9580
rect 3605 9531 3663 9537
rect 3712 9540 4436 9568
rect 2884 9472 3188 9500
rect 1394 9392 1400 9444
rect 1452 9432 1458 9444
rect 1489 9435 1547 9441
rect 1489 9432 1501 9435
rect 1452 9404 1501 9432
rect 1452 9392 1458 9404
rect 1489 9401 1501 9404
rect 1535 9401 1547 9435
rect 1489 9395 1547 9401
rect 2682 9392 2688 9444
rect 2740 9432 2746 9444
rect 2884 9432 2912 9472
rect 3234 9460 3240 9512
rect 3292 9500 3298 9512
rect 3421 9503 3479 9509
rect 3421 9500 3433 9503
rect 3292 9472 3433 9500
rect 3292 9460 3298 9472
rect 3421 9469 3433 9472
rect 3467 9469 3479 9503
rect 3421 9463 3479 9469
rect 2740 9404 2912 9432
rect 2740 9392 2746 9404
rect 3142 9392 3148 9444
rect 3200 9432 3206 9444
rect 3712 9432 3740 9540
rect 4430 9528 4436 9540
rect 4488 9528 4494 9580
rect 4816 9577 4844 9676
rect 4890 9664 4896 9676
rect 4948 9664 4954 9716
rect 5442 9664 5448 9716
rect 5500 9704 5506 9716
rect 5500 9676 5856 9704
rect 5500 9664 5506 9676
rect 5828 9645 5856 9676
rect 6454 9664 6460 9716
rect 6512 9704 6518 9716
rect 6512 9676 7420 9704
rect 6512 9664 6518 9676
rect 5721 9639 5779 9645
rect 5721 9605 5733 9639
rect 5767 9605 5779 9639
rect 5721 9599 5779 9605
rect 5813 9639 5871 9645
rect 5813 9605 5825 9639
rect 5859 9636 5871 9639
rect 7392 9636 7420 9676
rect 7558 9664 7564 9716
rect 7616 9704 7622 9716
rect 7837 9707 7895 9713
rect 7837 9704 7849 9707
rect 7616 9676 7849 9704
rect 7616 9664 7622 9676
rect 7837 9673 7849 9676
rect 7883 9673 7895 9707
rect 8294 9704 8300 9716
rect 7837 9667 7895 9673
rect 7944 9676 8300 9704
rect 7944 9636 7972 9676
rect 8294 9664 8300 9676
rect 8352 9664 8358 9716
rect 9766 9664 9772 9716
rect 9824 9704 9830 9716
rect 10778 9704 10784 9716
rect 9824 9676 10784 9704
rect 9824 9664 9830 9676
rect 10778 9664 10784 9676
rect 10836 9664 10842 9716
rect 11241 9707 11299 9713
rect 11241 9673 11253 9707
rect 11287 9704 11299 9707
rect 11606 9704 11612 9716
rect 11287 9676 11612 9704
rect 11287 9673 11299 9676
rect 11241 9667 11299 9673
rect 11606 9664 11612 9676
rect 11664 9664 11670 9716
rect 11790 9664 11796 9716
rect 11848 9704 11854 9716
rect 11848 9676 12296 9704
rect 11848 9664 11854 9676
rect 12268 9648 12296 9676
rect 12342 9664 12348 9716
rect 12400 9704 12406 9716
rect 12400 9676 13584 9704
rect 12400 9664 12406 9676
rect 5859 9608 5893 9636
rect 7392 9608 7972 9636
rect 5859 9605 5871 9608
rect 5813 9599 5871 9605
rect 4801 9571 4859 9577
rect 4801 9537 4813 9571
rect 4847 9537 4859 9571
rect 5074 9568 5080 9580
rect 5035 9540 5080 9568
rect 4801 9531 4859 9537
rect 3878 9500 3884 9512
rect 3791 9472 3884 9500
rect 3878 9460 3884 9472
rect 3936 9500 3942 9512
rect 4338 9500 4344 9512
rect 3936 9472 4344 9500
rect 3936 9460 3942 9472
rect 4338 9460 4344 9472
rect 4396 9460 4402 9512
rect 4617 9503 4675 9509
rect 4617 9469 4629 9503
rect 4663 9500 4675 9503
rect 4663 9472 4752 9500
rect 4663 9469 4675 9472
rect 4617 9463 4675 9469
rect 4724 9432 4752 9472
rect 4816 9444 4844 9531
rect 5074 9528 5080 9540
rect 5132 9528 5138 9580
rect 5258 9528 5264 9580
rect 5316 9568 5322 9580
rect 5626 9568 5632 9580
rect 5316 9540 5632 9568
rect 5316 9528 5322 9540
rect 5626 9528 5632 9540
rect 5684 9528 5690 9580
rect 5736 9568 5764 9599
rect 5736 9540 6592 9568
rect 5534 9500 5540 9512
rect 5276 9472 5540 9500
rect 3200 9404 3740 9432
rect 4080 9404 4752 9432
rect 3200 9392 3206 9404
rect 1854 9324 1860 9376
rect 1912 9364 1918 9376
rect 1949 9367 2007 9373
rect 1949 9364 1961 9367
rect 1912 9336 1961 9364
rect 1912 9324 1918 9336
rect 1949 9333 1961 9336
rect 1995 9333 2007 9367
rect 1949 9327 2007 9333
rect 2961 9367 3019 9373
rect 2961 9333 2973 9367
rect 3007 9364 3019 9367
rect 3694 9364 3700 9376
rect 3007 9336 3700 9364
rect 3007 9333 3019 9336
rect 2961 9327 3019 9333
rect 3694 9324 3700 9336
rect 3752 9324 3758 9376
rect 4080 9373 4108 9404
rect 4065 9367 4123 9373
rect 4065 9333 4077 9367
rect 4111 9333 4123 9367
rect 4065 9327 4123 9333
rect 4525 9367 4583 9373
rect 4525 9333 4537 9367
rect 4571 9364 4583 9367
rect 4614 9364 4620 9376
rect 4571 9336 4620 9364
rect 4571 9333 4583 9336
rect 4525 9327 4583 9333
rect 4614 9324 4620 9336
rect 4672 9324 4678 9376
rect 4724 9364 4752 9404
rect 4798 9392 4804 9444
rect 4856 9392 4862 9444
rect 5276 9432 5304 9472
rect 5534 9460 5540 9472
rect 5592 9460 5598 9512
rect 5810 9460 5816 9512
rect 5868 9500 5874 9512
rect 5997 9503 6055 9509
rect 5997 9500 6009 9503
rect 5868 9472 6009 9500
rect 5868 9460 5874 9472
rect 5997 9469 6009 9472
rect 6043 9469 6055 9503
rect 5997 9463 6055 9469
rect 6086 9460 6092 9512
rect 6144 9500 6150 9512
rect 6273 9503 6331 9509
rect 6273 9500 6285 9503
rect 6144 9472 6285 9500
rect 6144 9460 6150 9472
rect 6273 9469 6285 9472
rect 6319 9469 6331 9503
rect 6454 9500 6460 9512
rect 6415 9472 6460 9500
rect 6273 9463 6331 9469
rect 6454 9460 6460 9472
rect 6512 9460 6518 9512
rect 6564 9500 6592 9540
rect 7466 9528 7472 9580
rect 7524 9568 7530 9580
rect 7944 9577 7972 9608
rect 10428 9608 12204 9636
rect 7929 9571 7987 9577
rect 7524 9540 7880 9568
rect 7524 9528 7530 9540
rect 7742 9500 7748 9512
rect 6564 9472 7748 9500
rect 7742 9460 7748 9472
rect 7800 9460 7806 9512
rect 7852 9500 7880 9540
rect 7929 9537 7941 9571
rect 7975 9568 7987 9571
rect 7975 9540 8009 9568
rect 7975 9537 7987 9540
rect 7929 9531 7987 9537
rect 9122 9528 9128 9580
rect 9180 9568 9186 9580
rect 9401 9571 9459 9577
rect 9401 9568 9413 9571
rect 9180 9540 9413 9568
rect 9180 9528 9186 9540
rect 9401 9537 9413 9540
rect 9447 9537 9459 9571
rect 9401 9531 9459 9537
rect 7852 9472 8340 9500
rect 5092 9404 5304 9432
rect 5353 9435 5411 9441
rect 5092 9364 5120 9404
rect 5353 9401 5365 9435
rect 5399 9432 5411 9435
rect 6178 9432 6184 9444
rect 5399 9404 6184 9432
rect 5399 9401 5411 9404
rect 5353 9395 5411 9401
rect 6178 9392 6184 9404
rect 6236 9392 6242 9444
rect 6362 9392 6368 9444
rect 6420 9432 6426 9444
rect 6702 9435 6760 9441
rect 6702 9432 6714 9435
rect 6420 9404 6714 9432
rect 6420 9392 6426 9404
rect 6702 9401 6714 9404
rect 6748 9401 6760 9435
rect 6702 9395 6760 9401
rect 7282 9392 7288 9444
rect 7340 9432 7346 9444
rect 7834 9432 7840 9444
rect 7340 9404 7840 9432
rect 7340 9392 7346 9404
rect 7834 9392 7840 9404
rect 7892 9432 7898 9444
rect 8174 9435 8232 9441
rect 8174 9432 8186 9435
rect 7892 9404 8186 9432
rect 7892 9392 7898 9404
rect 8174 9401 8186 9404
rect 8220 9401 8232 9435
rect 8312 9432 8340 9472
rect 8570 9460 8576 9512
rect 8628 9500 8634 9512
rect 9214 9500 9220 9512
rect 8628 9472 9220 9500
rect 8628 9460 8634 9472
rect 9214 9460 9220 9472
rect 9272 9500 9278 9512
rect 10428 9500 10456 9608
rect 10686 9528 10692 9580
rect 10744 9568 10750 9580
rect 10873 9571 10931 9577
rect 10873 9568 10885 9571
rect 10744 9540 10885 9568
rect 10744 9528 10750 9540
rect 10873 9537 10885 9540
rect 10919 9537 10931 9571
rect 11790 9568 11796 9580
rect 11751 9540 11796 9568
rect 10873 9531 10931 9537
rect 11790 9528 11796 9540
rect 11848 9528 11854 9580
rect 11882 9528 11888 9580
rect 11940 9568 11946 9580
rect 11940 9540 11985 9568
rect 11940 9528 11946 9540
rect 9272 9472 10456 9500
rect 11425 9503 11483 9509
rect 9272 9460 9278 9472
rect 11425 9469 11437 9503
rect 11471 9500 11483 9503
rect 12066 9500 12072 9512
rect 11471 9472 12072 9500
rect 11471 9469 11483 9472
rect 11425 9463 11483 9469
rect 12066 9460 12072 9472
rect 12124 9460 12130 9512
rect 12176 9500 12204 9608
rect 12250 9596 12256 9648
rect 12308 9596 12314 9648
rect 13265 9639 13323 9645
rect 13265 9636 13277 9639
rect 12360 9608 13277 9636
rect 12360 9580 12388 9608
rect 13265 9605 13277 9608
rect 13311 9636 13323 9639
rect 13354 9636 13360 9648
rect 13311 9608 13360 9636
rect 13311 9605 13323 9608
rect 13265 9599 13323 9605
rect 13354 9596 13360 9608
rect 13412 9596 13418 9648
rect 13556 9636 13584 9676
rect 13630 9664 13636 9716
rect 13688 9704 13694 9716
rect 13725 9707 13783 9713
rect 13725 9704 13737 9707
rect 13688 9676 13737 9704
rect 13688 9664 13694 9676
rect 13725 9673 13737 9676
rect 13771 9673 13783 9707
rect 13725 9667 13783 9673
rect 14090 9664 14096 9716
rect 14148 9704 14154 9716
rect 15286 9704 15292 9716
rect 14148 9676 15292 9704
rect 14148 9664 14154 9676
rect 15286 9664 15292 9676
rect 15344 9664 15350 9716
rect 16390 9664 16396 9716
rect 16448 9704 16454 9716
rect 17862 9704 17868 9716
rect 16448 9676 17868 9704
rect 16448 9664 16454 9676
rect 14274 9636 14280 9648
rect 13556 9608 14280 9636
rect 14274 9596 14280 9608
rect 14332 9596 14338 9648
rect 14550 9636 14556 9648
rect 14511 9608 14556 9636
rect 14550 9596 14556 9608
rect 14608 9596 14614 9648
rect 14918 9596 14924 9648
rect 14976 9636 14982 9648
rect 15470 9636 15476 9648
rect 14976 9608 15332 9636
rect 15431 9608 15476 9636
rect 14976 9596 14982 9608
rect 12342 9528 12348 9580
rect 12400 9528 12406 9580
rect 12618 9528 12624 9580
rect 12676 9568 12682 9580
rect 13081 9571 13139 9577
rect 13081 9568 13093 9571
rect 12676 9540 13093 9568
rect 12676 9528 12682 9540
rect 13081 9537 13093 9540
rect 13127 9568 13139 9571
rect 14369 9571 14427 9577
rect 14369 9568 14381 9571
rect 13127 9540 14381 9568
rect 13127 9537 13139 9540
rect 13081 9531 13139 9537
rect 14369 9537 14381 9540
rect 14415 9568 14427 9571
rect 15194 9568 15200 9580
rect 14415 9540 15200 9568
rect 14415 9537 14427 9540
rect 14369 9531 14427 9537
rect 15194 9528 15200 9540
rect 15252 9528 15258 9580
rect 15304 9568 15332 9608
rect 15470 9596 15476 9608
rect 15528 9596 15534 9648
rect 15933 9639 15991 9645
rect 15933 9605 15945 9639
rect 15979 9605 15991 9639
rect 15933 9599 15991 9605
rect 15948 9568 15976 9599
rect 15304 9540 15976 9568
rect 16114 9528 16120 9580
rect 16172 9568 16178 9580
rect 16500 9577 16528 9676
rect 17862 9664 17868 9676
rect 17920 9664 17926 9716
rect 18506 9636 18512 9648
rect 18467 9608 18512 9636
rect 18506 9596 18512 9608
rect 18564 9596 18570 9648
rect 16393 9571 16451 9577
rect 16393 9568 16405 9571
rect 16172 9540 16405 9568
rect 16172 9528 16178 9540
rect 16393 9537 16405 9540
rect 16439 9537 16451 9571
rect 16393 9531 16451 9537
rect 16485 9571 16543 9577
rect 16485 9537 16497 9571
rect 16531 9537 16543 9571
rect 16485 9531 16543 9537
rect 12253 9503 12311 9509
rect 12253 9500 12265 9503
rect 12176 9472 12265 9500
rect 12253 9469 12265 9472
rect 12299 9500 12311 9503
rect 12805 9503 12863 9509
rect 12805 9500 12817 9503
rect 12299 9472 12817 9500
rect 12299 9469 12311 9472
rect 12253 9463 12311 9469
rect 12805 9469 12817 9472
rect 12851 9500 12863 9503
rect 14090 9500 14096 9512
rect 12851 9472 14096 9500
rect 12851 9469 12863 9472
rect 12805 9463 12863 9469
rect 14090 9460 14096 9472
rect 14148 9460 14154 9512
rect 14274 9460 14280 9512
rect 14332 9500 14338 9512
rect 15013 9503 15071 9509
rect 15013 9500 15025 9503
rect 14332 9472 15025 9500
rect 14332 9460 14338 9472
rect 15013 9469 15025 9472
rect 15059 9500 15071 9503
rect 15102 9500 15108 9512
rect 15059 9472 15108 9500
rect 15059 9469 15071 9472
rect 15013 9463 15071 9469
rect 15102 9460 15108 9472
rect 15160 9460 15166 9512
rect 15378 9460 15384 9512
rect 15436 9500 15442 9512
rect 16206 9500 16212 9512
rect 15436 9472 16212 9500
rect 15436 9460 15442 9472
rect 16206 9460 16212 9472
rect 16264 9460 16270 9512
rect 16301 9503 16359 9509
rect 16301 9469 16313 9503
rect 16347 9500 16359 9503
rect 16574 9500 16580 9512
rect 16347 9472 16580 9500
rect 16347 9469 16359 9472
rect 16301 9463 16359 9469
rect 16574 9460 16580 9472
rect 16632 9460 16638 9512
rect 16942 9500 16948 9512
rect 16903 9472 16948 9500
rect 16942 9460 16948 9472
rect 17000 9460 17006 9512
rect 9668 9435 9726 9441
rect 8312 9404 9444 9432
rect 8174 9395 8232 9401
rect 5258 9364 5264 9376
rect 4724 9336 5120 9364
rect 5219 9336 5264 9364
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 5810 9324 5816 9376
rect 5868 9364 5874 9376
rect 6089 9367 6147 9373
rect 6089 9364 6101 9367
rect 5868 9336 6101 9364
rect 5868 9324 5874 9336
rect 6089 9333 6101 9336
rect 6135 9364 6147 9367
rect 8662 9364 8668 9376
rect 6135 9336 8668 9364
rect 6135 9333 6147 9336
rect 6089 9327 6147 9333
rect 8662 9324 8668 9336
rect 8720 9324 8726 9376
rect 8846 9324 8852 9376
rect 8904 9364 8910 9376
rect 9309 9367 9367 9373
rect 9309 9364 9321 9367
rect 8904 9336 9321 9364
rect 8904 9324 8910 9336
rect 9309 9333 9321 9336
rect 9355 9333 9367 9367
rect 9416 9364 9444 9404
rect 9668 9401 9680 9435
rect 9714 9432 9726 9435
rect 10410 9432 10416 9444
rect 9714 9404 10416 9432
rect 9714 9401 9726 9404
rect 9668 9395 9726 9401
rect 10410 9392 10416 9404
rect 10468 9392 10474 9444
rect 13633 9435 13691 9441
rect 10980 9404 11293 9432
rect 10980 9364 11008 9404
rect 11146 9364 11152 9376
rect 9416 9336 11008 9364
rect 11107 9336 11152 9364
rect 9309 9327 9367 9333
rect 11146 9324 11152 9336
rect 11204 9324 11210 9376
rect 11265 9364 11293 9404
rect 13633 9401 13645 9435
rect 13679 9432 13691 9435
rect 14921 9435 14979 9441
rect 14921 9432 14933 9435
rect 13679 9404 14933 9432
rect 13679 9401 13691 9404
rect 13633 9395 13691 9401
rect 14921 9401 14933 9404
rect 14967 9401 14979 9435
rect 14921 9395 14979 9401
rect 15657 9435 15715 9441
rect 15657 9401 15669 9435
rect 15703 9432 15715 9435
rect 16666 9432 16672 9444
rect 15703 9404 16672 9432
rect 15703 9401 15715 9404
rect 15657 9395 15715 9401
rect 16666 9392 16672 9404
rect 16724 9392 16730 9444
rect 17218 9441 17224 9444
rect 17212 9432 17224 9441
rect 17179 9404 17224 9432
rect 17212 9395 17224 9404
rect 17218 9392 17224 9395
rect 17276 9392 17282 9444
rect 12069 9367 12127 9373
rect 12069 9364 12081 9367
rect 11265 9336 12081 9364
rect 12069 9333 12081 9336
rect 12115 9364 12127 9367
rect 12342 9364 12348 9376
rect 12115 9336 12348 9364
rect 12115 9333 12127 9336
rect 12069 9327 12127 9333
rect 12342 9324 12348 9336
rect 12400 9324 12406 9376
rect 12437 9367 12495 9373
rect 12437 9333 12449 9367
rect 12483 9364 12495 9367
rect 12710 9364 12716 9376
rect 12483 9336 12716 9364
rect 12483 9333 12495 9336
rect 12437 9327 12495 9333
rect 12710 9324 12716 9336
rect 12768 9324 12774 9376
rect 12897 9367 12955 9373
rect 12897 9333 12909 9367
rect 12943 9364 12955 9367
rect 13170 9364 13176 9376
rect 12943 9336 13176 9364
rect 12943 9333 12955 9336
rect 12897 9327 12955 9333
rect 13170 9324 13176 9336
rect 13228 9324 13234 9376
rect 13354 9324 13360 9376
rect 13412 9364 13418 9376
rect 13998 9364 14004 9376
rect 13412 9336 14004 9364
rect 13412 9324 13418 9336
rect 13998 9324 14004 9336
rect 14056 9364 14062 9376
rect 14093 9367 14151 9373
rect 14093 9364 14105 9367
rect 14056 9336 14105 9364
rect 14056 9324 14062 9336
rect 14093 9333 14105 9336
rect 14139 9333 14151 9367
rect 14093 9327 14151 9333
rect 14185 9367 14243 9373
rect 14185 9333 14197 9367
rect 14231 9364 14243 9367
rect 14366 9364 14372 9376
rect 14231 9336 14372 9364
rect 14231 9333 14243 9336
rect 14185 9327 14243 9333
rect 14366 9324 14372 9336
rect 14424 9324 14430 9376
rect 15746 9364 15752 9376
rect 15707 9336 15752 9364
rect 15746 9324 15752 9336
rect 15804 9324 15810 9376
rect 18322 9364 18328 9376
rect 18283 9336 18328 9364
rect 18322 9324 18328 9336
rect 18380 9324 18386 9376
rect 1104 9274 18860 9296
rect 1104 9222 6912 9274
rect 6964 9222 6976 9274
rect 7028 9222 7040 9274
rect 7092 9222 7104 9274
rect 7156 9222 12843 9274
rect 12895 9222 12907 9274
rect 12959 9222 12971 9274
rect 13023 9222 13035 9274
rect 13087 9222 18860 9274
rect 1104 9200 18860 9222
rect 1394 9120 1400 9172
rect 1452 9160 1458 9172
rect 3326 9160 3332 9172
rect 1452 9132 3332 9160
rect 1452 9120 1458 9132
rect 3326 9120 3332 9132
rect 3384 9120 3390 9172
rect 4522 9160 4528 9172
rect 3528 9132 4528 9160
rect 2866 9052 2872 9104
rect 2924 9101 2930 9104
rect 2924 9092 2936 9101
rect 3418 9092 3424 9104
rect 2924 9064 2969 9092
rect 3160 9064 3424 9092
rect 2924 9055 2936 9064
rect 2924 9052 2930 9055
rect 1486 9024 1492 9036
rect 1447 8996 1492 9024
rect 1486 8984 1492 8996
rect 1544 9024 1550 9036
rect 3160 9024 3188 9064
rect 3418 9052 3424 9064
rect 3476 9052 3482 9104
rect 3326 9024 3332 9036
rect 1544 8996 3188 9024
rect 3239 8996 3332 9024
rect 1544 8984 1550 8996
rect 3326 8984 3332 8996
rect 3384 9024 3390 9036
rect 3528 9024 3556 9132
rect 4522 9120 4528 9132
rect 4580 9120 4586 9172
rect 4617 9163 4675 9169
rect 4617 9129 4629 9163
rect 4663 9129 4675 9163
rect 5442 9160 5448 9172
rect 4617 9123 4675 9129
rect 5092 9132 5448 9160
rect 4154 9052 4160 9104
rect 4212 9092 4218 9104
rect 4632 9092 4660 9123
rect 5092 9092 5120 9132
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 6362 9160 6368 9172
rect 6323 9132 6368 9160
rect 6362 9120 6368 9132
rect 6420 9120 6426 9172
rect 6730 9120 6736 9172
rect 6788 9160 6794 9172
rect 6825 9163 6883 9169
rect 6825 9160 6837 9163
rect 6788 9132 6837 9160
rect 6788 9120 6794 9132
rect 6825 9129 6837 9132
rect 6871 9129 6883 9163
rect 6825 9123 6883 9129
rect 7193 9163 7251 9169
rect 7193 9129 7205 9163
rect 7239 9160 7251 9163
rect 9398 9160 9404 9172
rect 7239 9132 9404 9160
rect 7239 9129 7251 9132
rect 7193 9123 7251 9129
rect 9398 9120 9404 9132
rect 9456 9120 9462 9172
rect 10318 9120 10324 9172
rect 10376 9160 10382 9172
rect 10689 9163 10747 9169
rect 10689 9160 10701 9163
rect 10376 9132 10701 9160
rect 10376 9120 10382 9132
rect 10689 9129 10701 9132
rect 10735 9129 10747 9163
rect 12066 9160 12072 9172
rect 12027 9132 12072 9160
rect 10689 9123 10747 9129
rect 12066 9120 12072 9132
rect 12124 9120 12130 9172
rect 12342 9120 12348 9172
rect 12400 9160 12406 9172
rect 12989 9163 13047 9169
rect 12400 9132 12940 9160
rect 12400 9120 12406 9132
rect 4212 9064 4660 9092
rect 4816 9064 5120 9092
rect 4212 9052 4218 9064
rect 4246 9024 4252 9036
rect 3384 8996 3556 9024
rect 4207 8996 4252 9024
rect 3384 8984 3390 8996
rect 4246 8984 4252 8996
rect 4304 8984 4310 9036
rect 4816 9024 4844 9064
rect 4448 8996 4844 9024
rect 4893 9027 4951 9033
rect 4448 8968 4476 8996
rect 4893 8993 4905 9027
rect 4939 8993 4951 9027
rect 4893 8987 4951 8993
rect 3145 8959 3203 8965
rect 3145 8925 3157 8959
rect 3191 8925 3203 8959
rect 3145 8919 3203 8925
rect 1673 8891 1731 8897
rect 1673 8857 1685 8891
rect 1719 8888 1731 8891
rect 3160 8888 3188 8919
rect 3418 8916 3424 8968
rect 3476 8956 3482 8968
rect 3605 8959 3663 8965
rect 3605 8956 3617 8959
rect 3476 8928 3617 8956
rect 3476 8916 3482 8928
rect 3605 8925 3617 8928
rect 3651 8925 3663 8959
rect 4062 8956 4068 8968
rect 4023 8928 4068 8956
rect 3605 8919 3663 8925
rect 4062 8916 4068 8928
rect 4120 8916 4126 8968
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8956 4215 8959
rect 4338 8956 4344 8968
rect 4203 8928 4344 8956
rect 4203 8925 4215 8928
rect 4157 8919 4215 8925
rect 4338 8916 4344 8928
rect 4396 8916 4402 8968
rect 4430 8916 4436 8968
rect 4488 8916 4494 8968
rect 4448 8888 4476 8916
rect 4908 8888 4936 8987
rect 4992 8959 5050 8965
rect 4992 8925 5004 8959
rect 5038 8956 5050 8959
rect 5092 8956 5120 9064
rect 5252 9095 5310 9101
rect 5252 9061 5264 9095
rect 5298 9092 5310 9095
rect 5902 9092 5908 9104
rect 5298 9064 5908 9092
rect 5298 9061 5310 9064
rect 5252 9055 5310 9061
rect 5902 9052 5908 9064
rect 5960 9052 5966 9104
rect 6086 9052 6092 9104
rect 6144 9092 6150 9104
rect 8386 9092 8392 9104
rect 6144 9064 8392 9092
rect 6144 9052 6150 9064
rect 8386 9052 8392 9064
rect 8444 9052 8450 9104
rect 8478 9052 8484 9104
rect 8536 9092 8542 9104
rect 8573 9095 8631 9101
rect 8573 9092 8585 9095
rect 8536 9064 8585 9092
rect 8536 9052 8542 9064
rect 8573 9061 8585 9064
rect 8619 9061 8631 9095
rect 8573 9055 8631 9061
rect 9484 9095 9542 9101
rect 9484 9061 9496 9095
rect 9530 9092 9542 9095
rect 9582 9092 9588 9104
rect 9530 9064 9588 9092
rect 9530 9061 9542 9064
rect 9484 9055 9542 9061
rect 9582 9052 9588 9064
rect 9640 9052 9646 9104
rect 11057 9095 11115 9101
rect 11057 9061 11069 9095
rect 11103 9092 11115 9095
rect 11238 9092 11244 9104
rect 11103 9064 11244 9092
rect 11103 9061 11115 9064
rect 11057 9055 11115 9061
rect 11238 9052 11244 9064
rect 11296 9092 11302 9104
rect 12158 9092 12164 9104
rect 11296 9064 12164 9092
rect 11296 9052 11302 9064
rect 12158 9052 12164 9064
rect 12216 9052 12222 9104
rect 12618 9092 12624 9104
rect 12406 9064 12624 9092
rect 6270 8984 6276 9036
rect 6328 9024 6334 9036
rect 6733 9027 6791 9033
rect 6733 9024 6745 9027
rect 6328 8996 6745 9024
rect 6328 8984 6334 8996
rect 6733 8993 6745 8996
rect 6779 8993 6791 9027
rect 7282 9024 7288 9036
rect 6733 8987 6791 8993
rect 7208 8996 7288 9024
rect 5038 8928 5120 8956
rect 6641 8959 6699 8965
rect 5038 8925 5050 8928
rect 4992 8919 5050 8925
rect 6641 8925 6653 8959
rect 6687 8956 6699 8959
rect 7208 8956 7236 8996
rect 7282 8984 7288 8996
rect 7340 8984 7346 9036
rect 7653 9027 7711 9033
rect 7653 8993 7665 9027
rect 7699 9024 7711 9027
rect 8202 9024 8208 9036
rect 7699 8996 8208 9024
rect 7699 8993 7711 8996
rect 7653 8987 7711 8993
rect 8202 8984 8208 8996
rect 8260 8984 8266 9036
rect 8665 9027 8723 9033
rect 8665 8993 8677 9027
rect 8711 9024 8723 9027
rect 8938 9024 8944 9036
rect 8711 8996 8944 9024
rect 8711 8993 8723 8996
rect 8665 8987 8723 8993
rect 8938 8984 8944 8996
rect 8996 8984 9002 9036
rect 9122 8984 9128 9036
rect 9180 9024 9186 9036
rect 9217 9027 9275 9033
rect 9217 9024 9229 9027
rect 9180 8996 9229 9024
rect 9180 8984 9186 8996
rect 9217 8993 9229 8996
rect 9263 9024 9275 9027
rect 9306 9024 9312 9036
rect 9263 8996 9312 9024
rect 9263 8993 9275 8996
rect 9217 8987 9275 8993
rect 9306 8984 9312 8996
rect 9364 8984 9370 9036
rect 10686 8984 10692 9036
rect 10744 9024 10750 9036
rect 11149 9027 11207 9033
rect 11149 9024 11161 9027
rect 10744 8996 11161 9024
rect 10744 8984 10750 8996
rect 11149 8993 11161 8996
rect 11195 9024 11207 9027
rect 11885 9027 11943 9033
rect 11195 8996 11836 9024
rect 11195 8993 11207 8996
rect 11149 8987 11207 8993
rect 7374 8956 7380 8968
rect 6687 8928 7236 8956
rect 7335 8928 7380 8956
rect 6687 8925 6699 8928
rect 6641 8919 6699 8925
rect 7374 8916 7380 8928
rect 7432 8916 7438 8968
rect 7466 8916 7472 8968
rect 7524 8956 7530 8968
rect 7561 8959 7619 8965
rect 7561 8956 7573 8959
rect 7524 8928 7573 8956
rect 7524 8916 7530 8928
rect 7561 8925 7573 8928
rect 7607 8925 7619 8959
rect 8846 8956 8852 8968
rect 8807 8928 8852 8956
rect 7561 8919 7619 8925
rect 8846 8916 8852 8928
rect 8904 8916 8910 8968
rect 11241 8959 11299 8965
rect 11241 8925 11253 8959
rect 11287 8925 11299 8959
rect 11241 8919 11299 8925
rect 1719 8860 2176 8888
rect 3160 8860 4476 8888
rect 4540 8860 4936 8888
rect 8021 8891 8079 8897
rect 1719 8857 1731 8860
rect 1673 8851 1731 8857
rect 1762 8820 1768 8832
rect 1723 8792 1768 8820
rect 1762 8780 1768 8792
rect 1820 8780 1826 8832
rect 2148 8820 2176 8860
rect 3142 8820 3148 8832
rect 2148 8792 3148 8820
rect 3142 8780 3148 8792
rect 3200 8780 3206 8832
rect 3234 8780 3240 8832
rect 3292 8820 3298 8832
rect 3421 8823 3479 8829
rect 3421 8820 3433 8823
rect 3292 8792 3433 8820
rect 3292 8780 3298 8792
rect 3421 8789 3433 8792
rect 3467 8789 3479 8823
rect 3421 8783 3479 8789
rect 3510 8780 3516 8832
rect 3568 8820 3574 8832
rect 4540 8820 4568 8860
rect 8021 8857 8033 8891
rect 8067 8888 8079 8891
rect 9122 8888 9128 8900
rect 8067 8860 9128 8888
rect 8067 8857 8079 8860
rect 8021 8851 8079 8857
rect 9122 8848 9128 8860
rect 9180 8848 9186 8900
rect 10152 8860 10732 8888
rect 3568 8792 4568 8820
rect 3568 8780 3574 8792
rect 4614 8780 4620 8832
rect 4672 8820 4678 8832
rect 4709 8823 4767 8829
rect 4709 8820 4721 8823
rect 4672 8792 4721 8820
rect 4672 8780 4678 8792
rect 4709 8789 4721 8792
rect 4755 8789 4767 8823
rect 4709 8783 4767 8789
rect 6362 8780 6368 8832
rect 6420 8820 6426 8832
rect 6546 8820 6552 8832
rect 6420 8792 6552 8820
rect 6420 8780 6426 8792
rect 6546 8780 6552 8792
rect 6604 8780 6610 8832
rect 8202 8820 8208 8832
rect 8163 8792 8208 8820
rect 8202 8780 8208 8792
rect 8260 8780 8266 8832
rect 8938 8780 8944 8832
rect 8996 8820 9002 8832
rect 10152 8820 10180 8860
rect 8996 8792 10180 8820
rect 8996 8780 9002 8792
rect 10226 8780 10232 8832
rect 10284 8820 10290 8832
rect 10597 8823 10655 8829
rect 10597 8820 10609 8823
rect 10284 8792 10609 8820
rect 10284 8780 10290 8792
rect 10597 8789 10609 8792
rect 10643 8789 10655 8823
rect 10704 8820 10732 8860
rect 10778 8848 10784 8900
rect 10836 8888 10842 8900
rect 11256 8888 11284 8919
rect 11698 8916 11704 8968
rect 11756 8956 11762 8968
rect 11808 8956 11836 8996
rect 11885 8993 11897 9027
rect 11931 9024 11943 9027
rect 12250 9024 12256 9036
rect 11931 8996 12256 9024
rect 11931 8993 11943 8996
rect 11885 8987 11943 8993
rect 12250 8984 12256 8996
rect 12308 8984 12314 9036
rect 12406 9024 12434 9064
rect 12618 9052 12624 9064
rect 12676 9052 12682 9104
rect 12912 9092 12940 9132
rect 12989 9129 13001 9163
rect 13035 9160 13047 9163
rect 13170 9160 13176 9172
rect 13035 9132 13176 9160
rect 13035 9129 13047 9132
rect 12989 9123 13047 9129
rect 13170 9120 13176 9132
rect 13228 9120 13234 9172
rect 14642 9160 14648 9172
rect 14292 9132 14648 9160
rect 14292 9092 14320 9132
rect 14642 9120 14648 9132
rect 14700 9120 14706 9172
rect 15194 9120 15200 9172
rect 15252 9160 15258 9172
rect 15749 9163 15807 9169
rect 15749 9160 15761 9163
rect 15252 9132 15761 9160
rect 15252 9120 15258 9132
rect 15749 9129 15761 9132
rect 15795 9129 15807 9163
rect 16942 9160 16948 9172
rect 15749 9123 15807 9129
rect 15856 9132 16948 9160
rect 15856 9104 15884 9132
rect 16942 9120 16948 9132
rect 17000 9120 17006 9172
rect 17770 9160 17776 9172
rect 17731 9132 17776 9160
rect 17770 9120 17776 9132
rect 17828 9120 17834 9172
rect 12912 9064 14320 9092
rect 14366 9052 14372 9104
rect 14424 9092 14430 9104
rect 15010 9092 15016 9104
rect 14424 9064 15016 9092
rect 14424 9052 14430 9064
rect 15010 9052 15016 9064
rect 15068 9092 15074 9104
rect 15838 9092 15844 9104
rect 15068 9064 15844 9092
rect 15068 9052 15074 9064
rect 15838 9052 15844 9064
rect 15896 9052 15902 9104
rect 15930 9052 15936 9104
rect 15988 9092 15994 9104
rect 16086 9095 16144 9101
rect 16086 9092 16098 9095
rect 15988 9064 16098 9092
rect 15988 9052 15994 9064
rect 16086 9061 16098 9064
rect 16132 9061 16144 9095
rect 17678 9092 17684 9104
rect 17639 9064 17684 9092
rect 16086 9055 16144 9061
rect 17678 9052 17684 9064
rect 17736 9052 17742 9104
rect 12360 8996 12434 9024
rect 12529 9027 12587 9033
rect 12360 8965 12388 8996
rect 12529 8993 12541 9027
rect 12575 9024 12587 9027
rect 12575 8996 13308 9024
rect 12575 8993 12587 8996
rect 12529 8987 12587 8993
rect 13280 8968 13308 8996
rect 13354 8984 13360 9036
rect 13412 9024 13418 9036
rect 13722 9024 13728 9036
rect 13412 8996 13728 9024
rect 13412 8984 13418 8996
rect 13722 8984 13728 8996
rect 13780 8984 13786 9036
rect 13998 9024 14004 9036
rect 13959 8996 14004 9024
rect 13998 8984 14004 8996
rect 14056 8984 14062 9036
rect 14642 9033 14648 9036
rect 14636 9024 14648 9033
rect 14108 8996 14648 9024
rect 12345 8959 12403 8965
rect 11756 8928 12296 8956
rect 11756 8916 11762 8928
rect 12158 8888 12164 8900
rect 10836 8860 11284 8888
rect 11532 8860 12164 8888
rect 10836 8848 10842 8860
rect 11532 8820 11560 8860
rect 12158 8848 12164 8860
rect 12216 8848 12222 8900
rect 12268 8888 12296 8928
rect 12345 8925 12357 8959
rect 12391 8925 12403 8959
rect 12345 8919 12403 8925
rect 12437 8959 12495 8965
rect 12437 8925 12449 8959
rect 12483 8956 12495 8959
rect 13170 8956 13176 8968
rect 12483 8928 13176 8956
rect 12483 8925 12495 8928
rect 12437 8919 12495 8925
rect 13170 8916 13176 8928
rect 13228 8916 13234 8968
rect 13262 8916 13268 8968
rect 13320 8916 13326 8968
rect 13449 8959 13507 8965
rect 13449 8925 13461 8959
rect 13495 8925 13507 8959
rect 13449 8919 13507 8925
rect 13633 8959 13691 8965
rect 13633 8925 13645 8959
rect 13679 8956 13691 8959
rect 14108 8956 14136 8996
rect 14636 8987 14648 8996
rect 14700 9024 14706 9036
rect 14700 8996 14736 9024
rect 14642 8984 14648 8987
rect 14700 8984 14706 8996
rect 15102 8984 15108 9036
rect 15160 9024 15166 9036
rect 16850 9024 16856 9036
rect 15160 8996 16856 9024
rect 15160 8984 15166 8996
rect 16850 8984 16856 8996
rect 16908 8984 16914 9036
rect 18506 9024 18512 9036
rect 18467 8996 18512 9024
rect 18506 8984 18512 8996
rect 18564 8984 18570 9036
rect 13679 8928 14136 8956
rect 13679 8925 13691 8928
rect 13633 8919 13691 8925
rect 12268 8860 13308 8888
rect 10704 8792 11560 8820
rect 11609 8823 11667 8829
rect 10597 8783 10655 8789
rect 11609 8789 11621 8823
rect 11655 8820 11667 8823
rect 11790 8820 11796 8832
rect 11655 8792 11796 8820
rect 11655 8789 11667 8792
rect 11609 8783 11667 8789
rect 11790 8780 11796 8792
rect 11848 8780 11854 8832
rect 12618 8780 12624 8832
rect 12676 8820 12682 8832
rect 12897 8823 12955 8829
rect 12897 8820 12909 8823
rect 12676 8792 12909 8820
rect 12676 8780 12682 8792
rect 12897 8789 12909 8792
rect 12943 8789 12955 8823
rect 13280 8820 13308 8860
rect 13354 8848 13360 8900
rect 13412 8888 13418 8900
rect 13464 8888 13492 8919
rect 14182 8916 14188 8968
rect 14240 8916 14246 8968
rect 14366 8956 14372 8968
rect 14327 8928 14372 8956
rect 14366 8916 14372 8928
rect 14424 8916 14430 8968
rect 15838 8956 15844 8968
rect 15799 8928 15844 8956
rect 15838 8916 15844 8928
rect 15896 8916 15902 8968
rect 17034 8916 17040 8968
rect 17092 8956 17098 8968
rect 17862 8956 17868 8968
rect 17092 8928 17632 8956
rect 17823 8928 17868 8956
rect 17092 8916 17098 8928
rect 14200 8888 14228 8916
rect 17313 8891 17371 8897
rect 17313 8888 17325 8891
rect 13412 8860 13492 8888
rect 13648 8860 14228 8888
rect 16776 8860 17325 8888
rect 13412 8848 13418 8860
rect 13648 8832 13676 8860
rect 13630 8820 13636 8832
rect 13280 8792 13636 8820
rect 12897 8783 12955 8789
rect 13630 8780 13636 8792
rect 13688 8780 13694 8832
rect 13906 8820 13912 8832
rect 13867 8792 13912 8820
rect 13906 8780 13912 8792
rect 13964 8780 13970 8832
rect 14185 8823 14243 8829
rect 14185 8789 14197 8823
rect 14231 8820 14243 8823
rect 15654 8820 15660 8832
rect 14231 8792 15660 8820
rect 14231 8789 14243 8792
rect 14185 8783 14243 8789
rect 15654 8780 15660 8792
rect 15712 8780 15718 8832
rect 16206 8780 16212 8832
rect 16264 8820 16270 8832
rect 16776 8820 16804 8860
rect 17313 8857 17325 8860
rect 17359 8857 17371 8891
rect 17604 8888 17632 8928
rect 17862 8916 17868 8928
rect 17920 8916 17926 8968
rect 18325 8891 18383 8897
rect 18325 8888 18337 8891
rect 17604 8860 18337 8888
rect 17313 8851 17371 8857
rect 18325 8857 18337 8860
rect 18371 8857 18383 8891
rect 18325 8851 18383 8857
rect 17218 8820 17224 8832
rect 16264 8792 16804 8820
rect 17179 8792 17224 8820
rect 16264 8780 16270 8792
rect 17218 8780 17224 8792
rect 17276 8780 17282 8832
rect 17494 8780 17500 8832
rect 17552 8820 17558 8832
rect 17862 8820 17868 8832
rect 17552 8792 17868 8820
rect 17552 8780 17558 8792
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 1104 8730 18860 8752
rect 1104 8678 3947 8730
rect 3999 8678 4011 8730
rect 4063 8678 4075 8730
rect 4127 8678 4139 8730
rect 4191 8678 9878 8730
rect 9930 8678 9942 8730
rect 9994 8678 10006 8730
rect 10058 8678 10070 8730
rect 10122 8678 15808 8730
rect 15860 8678 15872 8730
rect 15924 8678 15936 8730
rect 15988 8678 16000 8730
rect 16052 8678 18860 8730
rect 1104 8656 18860 8678
rect 1489 8619 1547 8625
rect 1489 8585 1501 8619
rect 1535 8616 1547 8619
rect 2682 8616 2688 8628
rect 1535 8588 2688 8616
rect 1535 8585 1547 8588
rect 1489 8579 1547 8585
rect 2682 8576 2688 8588
rect 2740 8576 2746 8628
rect 3694 8576 3700 8628
rect 3752 8616 3758 8628
rect 6181 8619 6239 8625
rect 6181 8616 6193 8619
rect 3752 8588 6193 8616
rect 3752 8576 3758 8588
rect 6181 8585 6193 8588
rect 6227 8585 6239 8619
rect 7837 8619 7895 8625
rect 6181 8579 6239 8585
rect 6472 8588 7788 8616
rect 4341 8551 4399 8557
rect 4341 8517 4353 8551
rect 4387 8517 4399 8551
rect 4341 8511 4399 8517
rect 5813 8551 5871 8557
rect 5813 8517 5825 8551
rect 5859 8548 5871 8551
rect 5902 8548 5908 8560
rect 5859 8520 5908 8548
rect 5859 8517 5871 8520
rect 5813 8511 5871 8517
rect 4356 8480 4384 8511
rect 5902 8508 5908 8520
rect 5960 8508 5966 8560
rect 6472 8548 6500 8588
rect 6012 8520 6500 8548
rect 7760 8548 7788 8588
rect 7837 8585 7849 8619
rect 7883 8616 7895 8619
rect 10410 8616 10416 8628
rect 7883 8588 10416 8616
rect 7883 8585 7895 8588
rect 7837 8579 7895 8585
rect 10410 8576 10416 8588
rect 10468 8576 10474 8628
rect 10502 8576 10508 8628
rect 10560 8616 10566 8628
rect 16393 8619 16451 8625
rect 10560 8588 16160 8616
rect 10560 8576 10566 8588
rect 8294 8548 8300 8560
rect 7760 8520 8300 8548
rect 4356 8452 4568 8480
rect 1762 8372 1768 8424
rect 1820 8412 1826 8424
rect 2590 8412 2596 8424
rect 2648 8421 2654 8424
rect 1820 8384 2596 8412
rect 1820 8372 1826 8384
rect 2590 8372 2596 8384
rect 2648 8375 2660 8421
rect 2869 8415 2927 8421
rect 2869 8381 2881 8415
rect 2915 8412 2927 8415
rect 2961 8415 3019 8421
rect 2961 8412 2973 8415
rect 2915 8384 2973 8412
rect 2915 8381 2927 8384
rect 2869 8375 2927 8381
rect 2961 8381 2973 8384
rect 3007 8412 3019 8415
rect 4430 8412 4436 8424
rect 3007 8384 4436 8412
rect 3007 8381 3019 8384
rect 2961 8375 3019 8381
rect 2648 8372 2654 8375
rect 4430 8372 4436 8384
rect 4488 8372 4494 8424
rect 4540 8412 4568 8452
rect 4700 8415 4758 8421
rect 4700 8412 4712 8415
rect 4540 8384 4712 8412
rect 4700 8381 4712 8384
rect 4746 8412 4758 8415
rect 5074 8412 5080 8424
rect 4746 8384 5080 8412
rect 4746 8381 4758 8384
rect 4700 8375 4758 8381
rect 5074 8372 5080 8384
rect 5132 8372 5138 8424
rect 2682 8304 2688 8356
rect 2740 8344 2746 8356
rect 2774 8344 2780 8356
rect 2740 8316 2780 8344
rect 2740 8304 2746 8316
rect 2774 8304 2780 8316
rect 2832 8344 2838 8356
rect 3228 8347 3286 8353
rect 3228 8344 3240 8347
rect 2832 8316 3240 8344
rect 2832 8304 2838 8316
rect 3228 8313 3240 8316
rect 3274 8344 3286 8347
rect 3602 8344 3608 8356
rect 3274 8316 3608 8344
rect 3274 8313 3286 8316
rect 3228 8307 3286 8313
rect 3602 8304 3608 8316
rect 3660 8304 3666 8356
rect 3786 8304 3792 8356
rect 3844 8344 3850 8356
rect 6012 8344 6040 8520
rect 8294 8508 8300 8520
rect 8352 8508 8358 8560
rect 9490 8508 9496 8560
rect 9548 8508 9554 8560
rect 10137 8551 10195 8557
rect 10137 8517 10149 8551
rect 10183 8548 10195 8551
rect 10318 8548 10324 8560
rect 10183 8520 10324 8548
rect 10183 8517 10195 8520
rect 10137 8511 10195 8517
rect 10318 8508 10324 8520
rect 10376 8508 10382 8560
rect 12158 8548 12164 8560
rect 12119 8520 12164 8548
rect 12158 8508 12164 8520
rect 12216 8508 12222 8560
rect 12526 8548 12532 8560
rect 12452 8520 12532 8548
rect 9508 8480 9536 8508
rect 10502 8480 10508 8492
rect 6104 8452 6592 8480
rect 9508 8452 10508 8480
rect 6104 8421 6132 8452
rect 6089 8415 6147 8421
rect 6089 8381 6101 8415
rect 6135 8381 6147 8415
rect 6089 8375 6147 8381
rect 6457 8415 6515 8421
rect 6457 8381 6469 8415
rect 6503 8381 6515 8415
rect 6564 8412 6592 8452
rect 10502 8440 10508 8452
rect 10560 8440 10566 8492
rect 11517 8483 11575 8489
rect 11517 8449 11529 8483
rect 11563 8480 11575 8483
rect 11606 8480 11612 8492
rect 11563 8452 11612 8480
rect 11563 8449 11575 8452
rect 11517 8443 11575 8449
rect 11606 8440 11612 8452
rect 11664 8440 11670 8492
rect 11698 8440 11704 8492
rect 11756 8480 11762 8492
rect 12452 8489 12480 8520
rect 12526 8508 12532 8520
rect 12584 8508 12590 8560
rect 13170 8548 13176 8560
rect 13131 8520 13176 8548
rect 13170 8508 13176 8520
rect 13228 8508 13234 8560
rect 13262 8508 13268 8560
rect 13320 8548 13326 8560
rect 14001 8551 14059 8557
rect 14001 8548 14013 8551
rect 13320 8520 14013 8548
rect 13320 8508 13326 8520
rect 14001 8517 14013 8520
rect 14047 8517 14059 8551
rect 14001 8511 14059 8517
rect 14826 8508 14832 8560
rect 14884 8548 14890 8560
rect 15381 8551 15439 8557
rect 15381 8548 15393 8551
rect 14884 8520 15393 8548
rect 14884 8508 14890 8520
rect 15381 8517 15393 8520
rect 15427 8517 15439 8551
rect 15381 8511 15439 8517
rect 12069 8483 12127 8489
rect 12069 8480 12081 8483
rect 11756 8452 12081 8480
rect 11756 8440 11762 8452
rect 12069 8449 12081 8452
rect 12115 8449 12127 8483
rect 12069 8443 12127 8449
rect 12437 8483 12495 8489
rect 12437 8449 12449 8483
rect 12483 8449 12495 8483
rect 12618 8480 12624 8492
rect 12579 8452 12624 8480
rect 12437 8443 12495 8449
rect 12618 8440 12624 8452
rect 12676 8440 12682 8492
rect 13722 8440 13728 8492
rect 13780 8480 13786 8492
rect 13817 8483 13875 8489
rect 13817 8480 13829 8483
rect 13780 8452 13829 8480
rect 13780 8440 13786 8452
rect 13817 8449 13829 8452
rect 13863 8480 13875 8483
rect 14642 8480 14648 8492
rect 13863 8452 14648 8480
rect 13863 8449 13875 8452
rect 13817 8443 13875 8449
rect 14642 8440 14648 8452
rect 14700 8440 14706 8492
rect 15286 8480 15292 8492
rect 15247 8452 15292 8480
rect 15286 8440 15292 8452
rect 15344 8440 15350 8492
rect 15841 8483 15899 8489
rect 15841 8480 15853 8483
rect 15580 8452 15853 8480
rect 8754 8412 8760 8424
rect 6564 8384 8760 8412
rect 6457 8375 6515 8381
rect 3844 8316 6040 8344
rect 6472 8344 6500 8375
rect 8754 8372 8760 8384
rect 8812 8372 8818 8424
rect 8846 8372 8852 8424
rect 8904 8412 8910 8424
rect 9134 8415 9192 8421
rect 9134 8412 9146 8415
rect 8904 8384 9146 8412
rect 8904 8372 8910 8384
rect 9134 8381 9146 8384
rect 9180 8381 9192 8415
rect 9134 8375 9192 8381
rect 9306 8372 9312 8424
rect 9364 8412 9370 8424
rect 9401 8415 9459 8421
rect 9401 8412 9413 8415
rect 9364 8384 9413 8412
rect 9364 8372 9370 8384
rect 9401 8381 9413 8384
rect 9447 8381 9459 8415
rect 9401 8375 9459 8381
rect 9490 8372 9496 8424
rect 9548 8372 9554 8424
rect 9769 8415 9827 8421
rect 9769 8381 9781 8415
rect 9815 8412 9827 8415
rect 10686 8412 10692 8424
rect 9815 8384 10692 8412
rect 9815 8381 9827 8384
rect 9769 8375 9827 8381
rect 10686 8372 10692 8384
rect 10744 8412 10750 8424
rect 11790 8412 11796 8424
rect 10744 8384 11796 8412
rect 10744 8372 10750 8384
rect 11790 8372 11796 8384
rect 11848 8412 11854 8424
rect 12342 8412 12348 8424
rect 11848 8384 12348 8412
rect 11848 8372 11854 8384
rect 12342 8372 12348 8384
rect 12400 8372 12406 8424
rect 12710 8412 12716 8424
rect 12671 8384 12716 8412
rect 12710 8372 12716 8384
rect 12768 8372 12774 8424
rect 13446 8372 13452 8424
rect 13504 8412 13510 8424
rect 13541 8415 13599 8421
rect 13541 8412 13553 8415
rect 13504 8384 13553 8412
rect 13504 8372 13510 8384
rect 13541 8381 13553 8384
rect 13587 8381 13599 8415
rect 14829 8415 14887 8421
rect 14829 8412 14841 8415
rect 13541 8375 13599 8381
rect 13648 8384 14841 8412
rect 6546 8344 6552 8356
rect 6472 8316 6552 8344
rect 3844 8304 3850 8316
rect 6546 8304 6552 8316
rect 6604 8304 6610 8356
rect 6724 8347 6782 8353
rect 6724 8344 6736 8347
rect 6656 8316 6736 8344
rect 2038 8236 2044 8288
rect 2096 8276 2102 8288
rect 4062 8276 4068 8288
rect 2096 8248 4068 8276
rect 2096 8236 2102 8248
rect 4062 8236 4068 8248
rect 4120 8236 4126 8288
rect 4154 8236 4160 8288
rect 4212 8276 4218 8288
rect 5350 8276 5356 8288
rect 4212 8248 5356 8276
rect 4212 8236 4218 8248
rect 5350 8236 5356 8248
rect 5408 8236 5414 8288
rect 5718 8236 5724 8288
rect 5776 8276 5782 8288
rect 5905 8279 5963 8285
rect 5905 8276 5917 8279
rect 5776 8248 5917 8276
rect 5776 8236 5782 8248
rect 5905 8245 5917 8248
rect 5951 8245 5963 8279
rect 5905 8239 5963 8245
rect 6086 8236 6092 8288
rect 6144 8276 6150 8288
rect 6656 8276 6684 8316
rect 6724 8313 6736 8316
rect 6770 8344 6782 8347
rect 7374 8344 7380 8356
rect 6770 8316 7380 8344
rect 6770 8313 6782 8316
rect 6724 8307 6782 8313
rect 7374 8304 7380 8316
rect 7432 8344 7438 8356
rect 7432 8316 8156 8344
rect 7432 8304 7438 8316
rect 6144 8248 6684 8276
rect 6144 8236 6150 8248
rect 7834 8236 7840 8288
rect 7892 8276 7898 8288
rect 8021 8279 8079 8285
rect 8021 8276 8033 8279
rect 7892 8248 8033 8276
rect 7892 8236 7898 8248
rect 8021 8245 8033 8248
rect 8067 8245 8079 8279
rect 8128 8276 8156 8316
rect 8294 8304 8300 8356
rect 8352 8344 8358 8356
rect 9508 8344 9536 8372
rect 8352 8316 9536 8344
rect 8352 8304 8358 8316
rect 10226 8304 10232 8356
rect 10284 8344 10290 8356
rect 11250 8347 11308 8353
rect 11250 8344 11262 8347
rect 10284 8316 11262 8344
rect 10284 8304 10290 8316
rect 11250 8313 11262 8316
rect 11296 8313 11308 8347
rect 11882 8344 11888 8356
rect 11843 8316 11888 8344
rect 11250 8307 11308 8313
rect 11882 8304 11888 8316
rect 11940 8304 11946 8356
rect 12158 8304 12164 8356
rect 12216 8344 12222 8356
rect 13648 8353 13676 8384
rect 14829 8381 14841 8384
rect 14875 8381 14887 8415
rect 15102 8412 15108 8424
rect 15063 8384 15108 8412
rect 14829 8375 14887 8381
rect 13633 8347 13691 8353
rect 13633 8344 13645 8347
rect 12216 8316 13645 8344
rect 12216 8304 12222 8316
rect 13633 8313 13645 8316
rect 13679 8313 13691 8347
rect 13814 8344 13820 8356
rect 13633 8307 13691 8313
rect 13740 8316 13820 8344
rect 9306 8276 9312 8288
rect 8128 8248 9312 8276
rect 8021 8239 8079 8245
rect 9306 8236 9312 8248
rect 9364 8236 9370 8288
rect 9585 8279 9643 8285
rect 9585 8245 9597 8279
rect 9631 8276 9643 8279
rect 9674 8276 9680 8288
rect 9631 8248 9680 8276
rect 9631 8245 9643 8248
rect 9585 8239 9643 8245
rect 9674 8236 9680 8248
rect 9732 8276 9738 8288
rect 10045 8279 10103 8285
rect 10045 8276 10057 8279
rect 9732 8248 10057 8276
rect 9732 8236 9738 8248
rect 10045 8245 10057 8248
rect 10091 8276 10103 8279
rect 10778 8276 10784 8288
rect 10091 8248 10784 8276
rect 10091 8245 10103 8248
rect 10045 8239 10103 8245
rect 10778 8236 10784 8248
rect 10836 8276 10842 8288
rect 11900 8276 11928 8304
rect 10836 8248 11928 8276
rect 13081 8279 13139 8285
rect 10836 8236 10842 8248
rect 13081 8245 13093 8279
rect 13127 8276 13139 8279
rect 13740 8276 13768 8316
rect 13814 8304 13820 8316
rect 13872 8304 13878 8356
rect 13998 8304 14004 8356
rect 14056 8344 14062 8356
rect 14274 8344 14280 8356
rect 14056 8316 14280 8344
rect 14056 8304 14062 8316
rect 14274 8304 14280 8316
rect 14332 8344 14338 8356
rect 14369 8347 14427 8353
rect 14369 8344 14381 8347
rect 14332 8316 14381 8344
rect 14332 8304 14338 8316
rect 14369 8313 14381 8316
rect 14415 8313 14427 8347
rect 14369 8307 14427 8313
rect 13127 8248 13768 8276
rect 14461 8279 14519 8285
rect 13127 8245 13139 8248
rect 13081 8239 13139 8245
rect 14461 8245 14473 8279
rect 14507 8276 14519 8279
rect 14550 8276 14556 8288
rect 14507 8248 14556 8276
rect 14507 8245 14519 8248
rect 14461 8239 14519 8245
rect 14550 8236 14556 8248
rect 14608 8236 14614 8288
rect 14844 8276 14872 8375
rect 15102 8372 15108 8384
rect 15160 8372 15166 8424
rect 14918 8304 14924 8356
rect 14976 8344 14982 8356
rect 15580 8344 15608 8452
rect 15841 8449 15853 8452
rect 15887 8449 15899 8483
rect 16022 8480 16028 8492
rect 15983 8452 16028 8480
rect 15841 8443 15899 8449
rect 16022 8440 16028 8452
rect 16080 8440 16086 8492
rect 15749 8415 15807 8421
rect 15749 8381 15761 8415
rect 15795 8412 15807 8415
rect 15930 8412 15936 8424
rect 15795 8384 15936 8412
rect 15795 8381 15807 8384
rect 15749 8375 15807 8381
rect 15930 8372 15936 8384
rect 15988 8372 15994 8424
rect 16132 8412 16160 8588
rect 16393 8585 16405 8619
rect 16439 8616 16451 8619
rect 17494 8616 17500 8628
rect 16439 8588 17500 8616
rect 16439 8585 16451 8588
rect 16393 8579 16451 8585
rect 17494 8576 17500 8588
rect 17552 8576 17558 8628
rect 16666 8508 16672 8560
rect 16724 8548 16730 8560
rect 16945 8551 17003 8557
rect 16945 8548 16957 8551
rect 16724 8520 16957 8548
rect 16724 8508 16730 8520
rect 16945 8517 16957 8520
rect 16991 8517 17003 8551
rect 16945 8511 17003 8517
rect 17034 8508 17040 8560
rect 17092 8548 17098 8560
rect 18325 8551 18383 8557
rect 18325 8548 18337 8551
rect 17092 8520 18337 8548
rect 17092 8508 17098 8520
rect 18325 8517 18337 8520
rect 18371 8517 18383 8551
rect 18325 8511 18383 8517
rect 17218 8440 17224 8492
rect 17276 8480 17282 8492
rect 17497 8483 17555 8489
rect 17497 8480 17509 8483
rect 17276 8452 17509 8480
rect 17276 8440 17282 8452
rect 17497 8449 17509 8452
rect 17543 8449 17555 8483
rect 17497 8443 17555 8449
rect 16209 8415 16267 8421
rect 16209 8412 16221 8415
rect 16132 8384 16221 8412
rect 16209 8381 16221 8384
rect 16255 8381 16267 8415
rect 16209 8375 16267 8381
rect 16482 8372 16488 8424
rect 16540 8412 16546 8424
rect 16761 8415 16819 8421
rect 16761 8412 16773 8415
rect 16540 8384 16773 8412
rect 16540 8372 16546 8384
rect 16761 8381 16773 8384
rect 16807 8381 16819 8415
rect 17405 8415 17463 8421
rect 17405 8412 17417 8415
rect 16761 8375 16819 8381
rect 16868 8384 17417 8412
rect 14976 8316 15608 8344
rect 14976 8304 14982 8316
rect 15654 8304 15660 8356
rect 15712 8344 15718 8356
rect 16577 8347 16635 8353
rect 16577 8344 16589 8347
rect 15712 8316 16589 8344
rect 15712 8304 15718 8316
rect 16577 8313 16589 8316
rect 16623 8313 16635 8347
rect 16868 8344 16896 8384
rect 17405 8381 17417 8384
rect 17451 8381 17463 8415
rect 17405 8375 17463 8381
rect 18509 8415 18567 8421
rect 18509 8381 18521 8415
rect 18555 8412 18567 8415
rect 18598 8412 18604 8424
rect 18555 8384 18604 8412
rect 18555 8381 18567 8384
rect 18509 8375 18567 8381
rect 18598 8372 18604 8384
rect 18656 8372 18662 8424
rect 16577 8307 16635 8313
rect 16684 8316 16896 8344
rect 16684 8276 16712 8316
rect 16942 8304 16948 8356
rect 17000 8344 17006 8356
rect 17313 8347 17371 8353
rect 17313 8344 17325 8347
rect 17000 8316 17325 8344
rect 17000 8304 17006 8316
rect 17313 8313 17325 8316
rect 17359 8313 17371 8347
rect 17954 8344 17960 8356
rect 17915 8316 17960 8344
rect 17313 8307 17371 8313
rect 17954 8304 17960 8316
rect 18012 8304 18018 8356
rect 18138 8344 18144 8356
rect 18099 8316 18144 8344
rect 18138 8304 18144 8316
rect 18196 8304 18202 8356
rect 14844 8248 16712 8276
rect 17218 8236 17224 8288
rect 17276 8276 17282 8288
rect 17402 8276 17408 8288
rect 17276 8248 17408 8276
rect 17276 8236 17282 8248
rect 17402 8236 17408 8248
rect 17460 8236 17466 8288
rect 1104 8186 18860 8208
rect 1104 8134 6912 8186
rect 6964 8134 6976 8186
rect 7028 8134 7040 8186
rect 7092 8134 7104 8186
rect 7156 8134 12843 8186
rect 12895 8134 12907 8186
rect 12959 8134 12971 8186
rect 13023 8134 13035 8186
rect 13087 8134 18860 8186
rect 1104 8112 18860 8134
rect 3053 8075 3111 8081
rect 3053 8041 3065 8075
rect 3099 8072 3111 8075
rect 3510 8072 3516 8084
rect 3099 8044 3516 8072
rect 3099 8041 3111 8044
rect 3053 8035 3111 8041
rect 3510 8032 3516 8044
rect 3568 8032 3574 8084
rect 4062 8032 4068 8084
rect 4120 8072 4126 8084
rect 5166 8072 5172 8084
rect 4120 8044 5172 8072
rect 4120 8032 4126 8044
rect 5166 8032 5172 8044
rect 5224 8032 5230 8084
rect 5258 8032 5264 8084
rect 5316 8072 5322 8084
rect 5445 8075 5503 8081
rect 5445 8072 5457 8075
rect 5316 8044 5457 8072
rect 5316 8032 5322 8044
rect 5445 8041 5457 8044
rect 5491 8041 5503 8075
rect 5445 8035 5503 8041
rect 5810 8032 5816 8084
rect 5868 8032 5874 8084
rect 6086 8072 6092 8084
rect 6047 8044 6092 8072
rect 6086 8032 6092 8044
rect 6144 8032 6150 8084
rect 7558 8032 7564 8084
rect 7616 8072 7622 8084
rect 7837 8075 7895 8081
rect 7837 8072 7849 8075
rect 7616 8044 7849 8072
rect 7616 8032 7622 8044
rect 7837 8041 7849 8044
rect 7883 8041 7895 8075
rect 8386 8072 8392 8084
rect 8347 8044 8392 8072
rect 7837 8035 7895 8041
rect 8386 8032 8392 8044
rect 8444 8032 8450 8084
rect 8757 8075 8815 8081
rect 8757 8041 8769 8075
rect 8803 8072 8815 8075
rect 8938 8072 8944 8084
rect 8803 8044 8944 8072
rect 8803 8041 8815 8044
rect 8757 8035 8815 8041
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 12526 8072 12532 8084
rect 9646 8044 12532 8072
rect 1486 8004 1492 8016
rect 1447 7976 1492 8004
rect 1486 7964 1492 7976
rect 1544 8004 1550 8016
rect 3694 8004 3700 8016
rect 1544 7976 3700 8004
rect 1544 7964 1550 7976
rect 3694 7964 3700 7976
rect 3752 7964 3758 8016
rect 5077 8007 5135 8013
rect 3804 7976 4936 8004
rect 2225 7939 2283 7945
rect 2225 7905 2237 7939
rect 2271 7936 2283 7939
rect 2682 7936 2688 7948
rect 2271 7908 2688 7936
rect 2271 7905 2283 7908
rect 2225 7899 2283 7905
rect 2682 7896 2688 7908
rect 2740 7896 2746 7948
rect 3513 7939 3571 7945
rect 3513 7905 3525 7939
rect 3559 7905 3571 7939
rect 3513 7899 3571 7905
rect 2314 7868 2320 7880
rect 2275 7840 2320 7868
rect 2314 7828 2320 7840
rect 2372 7828 2378 7880
rect 2409 7871 2467 7877
rect 2409 7837 2421 7871
rect 2455 7837 2467 7871
rect 3142 7868 3148 7880
rect 3103 7840 3148 7868
rect 2409 7831 2467 7837
rect 1670 7800 1676 7812
rect 1631 7772 1676 7800
rect 1670 7760 1676 7772
rect 1728 7760 1734 7812
rect 2424 7800 2452 7831
rect 3142 7828 3148 7840
rect 3200 7828 3206 7880
rect 3237 7871 3295 7877
rect 3237 7837 3249 7871
rect 3283 7837 3295 7871
rect 3528 7868 3556 7899
rect 3602 7896 3608 7948
rect 3660 7936 3666 7948
rect 3804 7936 3832 7976
rect 3660 7908 3832 7936
rect 3660 7896 3666 7908
rect 3970 7896 3976 7948
rect 4028 7936 4034 7948
rect 4249 7939 4307 7945
rect 4249 7936 4261 7939
rect 4028 7908 4261 7936
rect 4028 7896 4034 7908
rect 4249 7905 4261 7908
rect 4295 7905 4307 7939
rect 4249 7899 4307 7905
rect 4341 7939 4399 7945
rect 4341 7905 4353 7939
rect 4387 7936 4399 7939
rect 4387 7908 4568 7936
rect 4387 7905 4399 7908
rect 4341 7899 4399 7905
rect 4154 7868 4160 7880
rect 3528 7840 4160 7868
rect 3237 7831 3295 7837
rect 2590 7800 2596 7812
rect 2424 7772 2596 7800
rect 2590 7760 2596 7772
rect 2648 7800 2654 7812
rect 3252 7800 3280 7831
rect 4154 7828 4160 7840
rect 4212 7828 4218 7880
rect 4433 7871 4491 7877
rect 4433 7868 4445 7871
rect 4356 7840 4445 7868
rect 2648 7772 4200 7800
rect 2648 7760 2654 7772
rect 1857 7735 1915 7741
rect 1857 7701 1869 7735
rect 1903 7732 1915 7735
rect 2038 7732 2044 7744
rect 1903 7704 2044 7732
rect 1903 7701 1915 7704
rect 1857 7695 1915 7701
rect 2038 7692 2044 7704
rect 2096 7692 2102 7744
rect 2130 7692 2136 7744
rect 2188 7732 2194 7744
rect 2685 7735 2743 7741
rect 2685 7732 2697 7735
rect 2188 7704 2697 7732
rect 2188 7692 2194 7704
rect 2685 7701 2697 7704
rect 2731 7701 2743 7735
rect 3694 7732 3700 7744
rect 3655 7704 3700 7732
rect 2685 7695 2743 7701
rect 3694 7692 3700 7704
rect 3752 7692 3758 7744
rect 3786 7692 3792 7744
rect 3844 7732 3850 7744
rect 3881 7735 3939 7741
rect 3881 7732 3893 7735
rect 3844 7704 3893 7732
rect 3844 7692 3850 7704
rect 3881 7701 3893 7704
rect 3927 7701 3939 7735
rect 4172 7732 4200 7772
rect 4356 7732 4384 7840
rect 4433 7837 4445 7840
rect 4479 7837 4491 7871
rect 4433 7831 4491 7837
rect 4172 7704 4384 7732
rect 4540 7732 4568 7908
rect 4908 7877 4936 7976
rect 5077 7973 5089 8007
rect 5123 8004 5135 8007
rect 5828 8004 5856 8032
rect 5123 7976 5856 8004
rect 5123 7973 5135 7976
rect 5077 7967 5135 7973
rect 5902 7964 5908 8016
rect 5960 8004 5966 8016
rect 5960 7976 7696 8004
rect 5960 7964 5966 7976
rect 5813 7939 5871 7945
rect 5813 7905 5825 7939
rect 5859 7936 5871 7939
rect 5994 7936 6000 7948
rect 5859 7908 6000 7936
rect 5859 7905 5871 7908
rect 5813 7899 5871 7905
rect 5994 7896 6000 7908
rect 6052 7896 6058 7948
rect 7213 7939 7271 7945
rect 7213 7905 7225 7939
rect 7259 7936 7271 7939
rect 7259 7908 7604 7936
rect 7259 7905 7271 7908
rect 7213 7899 7271 7905
rect 4893 7871 4951 7877
rect 4893 7837 4905 7871
rect 4939 7837 4951 7871
rect 4893 7831 4951 7837
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7868 5043 7871
rect 5074 7868 5080 7880
rect 5031 7840 5080 7868
rect 5031 7837 5043 7840
rect 4985 7831 5043 7837
rect 4908 7800 4936 7831
rect 5074 7828 5080 7840
rect 5132 7868 5138 7880
rect 5626 7868 5632 7880
rect 5132 7840 5632 7868
rect 5132 7828 5138 7840
rect 5626 7828 5632 7840
rect 5684 7828 5690 7880
rect 5721 7871 5779 7877
rect 5721 7837 5733 7871
rect 5767 7868 5779 7871
rect 6454 7868 6460 7880
rect 5767 7840 6460 7868
rect 5767 7837 5779 7840
rect 5721 7831 5779 7837
rect 6454 7828 6460 7840
rect 6512 7828 6518 7880
rect 7469 7871 7527 7877
rect 7469 7837 7481 7871
rect 7515 7837 7527 7871
rect 7469 7831 7527 7837
rect 6270 7800 6276 7812
rect 4908 7772 6276 7800
rect 6270 7760 6276 7772
rect 6328 7760 6334 7812
rect 4890 7732 4896 7744
rect 4540 7704 4896 7732
rect 3881 7695 3939 7701
rect 4890 7692 4896 7704
rect 4948 7692 4954 7744
rect 5994 7732 6000 7744
rect 5955 7704 6000 7732
rect 5994 7692 6000 7704
rect 6052 7692 6058 7744
rect 6546 7692 6552 7744
rect 6604 7732 6610 7744
rect 7484 7732 7512 7831
rect 7576 7800 7604 7908
rect 7668 7877 7696 7976
rect 7742 7964 7748 8016
rect 7800 8004 7806 8016
rect 7929 8007 7987 8013
rect 7929 8004 7941 8007
rect 7800 7976 7941 8004
rect 7800 7964 7806 7976
rect 7929 7973 7941 7976
rect 7975 7973 7987 8007
rect 7929 7967 7987 7973
rect 8846 7964 8852 8016
rect 8904 8004 8910 8016
rect 9125 8007 9183 8013
rect 9125 8004 9137 8007
rect 8904 7976 9137 8004
rect 8904 7964 8910 7976
rect 9125 7973 9137 7976
rect 9171 8004 9183 8007
rect 9646 8004 9674 8044
rect 12526 8032 12532 8044
rect 12584 8072 12590 8084
rect 13722 8072 13728 8084
rect 12584 8044 13216 8072
rect 13683 8044 13728 8072
rect 12584 8032 12590 8044
rect 9171 7976 9674 8004
rect 11425 8007 11483 8013
rect 9171 7973 9183 7976
rect 9125 7967 9183 7973
rect 11425 7973 11437 8007
rect 11471 8004 11483 8007
rect 13188 8004 13216 8044
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 14185 8075 14243 8081
rect 14185 8041 14197 8075
rect 14231 8041 14243 8075
rect 14185 8035 14243 8041
rect 14200 8004 14228 8035
rect 14366 8032 14372 8084
rect 14424 8072 14430 8084
rect 15933 8075 15991 8081
rect 15933 8072 15945 8075
rect 14424 8044 15945 8072
rect 14424 8032 14430 8044
rect 15933 8041 15945 8044
rect 15979 8041 15991 8075
rect 15933 8035 15991 8041
rect 16206 8032 16212 8084
rect 16264 8072 16270 8084
rect 16393 8075 16451 8081
rect 16393 8072 16405 8075
rect 16264 8044 16405 8072
rect 16264 8032 16270 8044
rect 16393 8041 16405 8044
rect 16439 8041 16451 8075
rect 16393 8035 16451 8041
rect 16761 8075 16819 8081
rect 16761 8041 16773 8075
rect 16807 8072 16819 8075
rect 17313 8075 17371 8081
rect 17313 8072 17325 8075
rect 16807 8044 17325 8072
rect 16807 8041 16819 8044
rect 16761 8035 16819 8041
rect 17313 8041 17325 8044
rect 17359 8041 17371 8075
rect 17313 8035 17371 8041
rect 17954 8004 17960 8016
rect 11471 7976 13124 8004
rect 13188 7976 13952 8004
rect 14200 7976 17960 8004
rect 11471 7973 11483 7976
rect 11425 7967 11483 7973
rect 8110 7936 8116 7948
rect 7760 7908 8116 7936
rect 7760 7880 7788 7908
rect 8110 7896 8116 7908
rect 8168 7896 8174 7948
rect 8573 7939 8631 7945
rect 8573 7905 8585 7939
rect 8619 7936 8631 7939
rect 8619 7908 10180 7936
rect 8619 7905 8631 7908
rect 8573 7899 8631 7905
rect 7653 7871 7711 7877
rect 7653 7837 7665 7871
rect 7699 7837 7711 7871
rect 7653 7831 7711 7837
rect 7742 7828 7748 7880
rect 7800 7828 7806 7880
rect 7926 7828 7932 7880
rect 7984 7868 7990 7880
rect 9309 7871 9367 7877
rect 9309 7868 9321 7871
rect 7984 7840 9321 7868
rect 7984 7828 7990 7840
rect 9309 7837 9321 7840
rect 9355 7868 9367 7871
rect 9858 7868 9864 7880
rect 9355 7840 9864 7868
rect 9355 7837 9367 7840
rect 9309 7831 9367 7837
rect 9858 7828 9864 7840
rect 9916 7828 9922 7880
rect 7834 7800 7840 7812
rect 7576 7772 7840 7800
rect 7834 7760 7840 7772
rect 7892 7760 7898 7812
rect 6604 7704 7512 7732
rect 6604 7692 6610 7704
rect 7558 7692 7564 7744
rect 7616 7732 7622 7744
rect 7944 7732 7972 7828
rect 8297 7803 8355 7809
rect 8297 7769 8309 7803
rect 8343 7800 8355 7803
rect 9582 7800 9588 7812
rect 8343 7772 9588 7800
rect 8343 7769 8355 7772
rect 8297 7763 8355 7769
rect 9582 7760 9588 7772
rect 9640 7760 9646 7812
rect 7616 7704 7972 7732
rect 7616 7692 7622 7704
rect 8018 7692 8024 7744
rect 8076 7732 8082 7744
rect 9493 7735 9551 7741
rect 9493 7732 9505 7735
rect 8076 7704 9505 7732
rect 8076 7692 8082 7704
rect 9493 7701 9505 7704
rect 9539 7732 9551 7735
rect 9674 7732 9680 7744
rect 9539 7704 9680 7732
rect 9539 7701 9551 7704
rect 9493 7695 9551 7701
rect 9674 7692 9680 7704
rect 9732 7692 9738 7744
rect 10152 7741 10180 7908
rect 11514 7896 11520 7948
rect 11572 7936 11578 7948
rect 11885 7939 11943 7945
rect 11885 7936 11897 7939
rect 11572 7908 11897 7936
rect 11572 7896 11578 7908
rect 11885 7905 11897 7908
rect 11931 7905 11943 7939
rect 12612 7939 12670 7945
rect 12612 7936 12624 7939
rect 11885 7899 11943 7905
rect 11992 7908 12624 7936
rect 11609 7871 11667 7877
rect 11609 7837 11621 7871
rect 11655 7837 11667 7871
rect 11790 7868 11796 7880
rect 11751 7840 11796 7868
rect 11609 7831 11667 7837
rect 10594 7760 10600 7812
rect 10652 7800 10658 7812
rect 11146 7800 11152 7812
rect 10652 7772 11152 7800
rect 10652 7760 10658 7772
rect 11146 7760 11152 7772
rect 11204 7760 11210 7812
rect 11624 7800 11652 7831
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 11992 7800 12020 7908
rect 12612 7905 12624 7908
rect 12658 7936 12670 7939
rect 12894 7936 12900 7948
rect 12658 7908 12900 7936
rect 12658 7905 12670 7908
rect 12612 7899 12670 7905
rect 12894 7896 12900 7908
rect 12952 7896 12958 7948
rect 13096 7936 13124 7976
rect 13924 7948 13952 7976
rect 17954 7964 17960 7976
rect 18012 7964 18018 8016
rect 13814 7936 13820 7948
rect 13096 7908 13400 7936
rect 13775 7908 13820 7936
rect 12066 7828 12072 7880
rect 12124 7868 12130 7880
rect 12345 7871 12403 7877
rect 12345 7868 12357 7871
rect 12124 7840 12357 7868
rect 12124 7828 12130 7840
rect 12345 7837 12357 7840
rect 12391 7837 12403 7871
rect 13372 7868 13400 7908
rect 13814 7896 13820 7908
rect 13872 7896 13878 7948
rect 13906 7896 13912 7948
rect 13964 7936 13970 7948
rect 14001 7939 14059 7945
rect 14001 7936 14013 7939
rect 13964 7908 14013 7936
rect 13964 7896 13970 7908
rect 14001 7905 14013 7908
rect 14047 7905 14059 7939
rect 15286 7936 15292 7948
rect 14001 7899 14059 7905
rect 14108 7908 15292 7936
rect 14108 7868 14136 7908
rect 15286 7896 15292 7908
rect 15344 7896 15350 7948
rect 15585 7939 15643 7945
rect 15585 7905 15597 7939
rect 15631 7936 15643 7939
rect 15631 7908 16252 7936
rect 15631 7905 15643 7908
rect 15585 7899 15643 7905
rect 16224 7880 16252 7908
rect 16298 7896 16304 7948
rect 16356 7936 16362 7948
rect 16356 7908 16401 7936
rect 16356 7896 16362 7908
rect 16666 7896 16672 7948
rect 16724 7936 16730 7948
rect 17221 7939 17279 7945
rect 17221 7936 17233 7939
rect 16724 7908 17233 7936
rect 16724 7896 16730 7908
rect 17221 7905 17233 7908
rect 17267 7905 17279 7939
rect 17221 7899 17279 7905
rect 17770 7896 17776 7948
rect 17828 7936 17834 7948
rect 18049 7939 18107 7945
rect 18049 7936 18061 7939
rect 17828 7908 18061 7936
rect 17828 7896 17834 7908
rect 18049 7905 18061 7908
rect 18095 7905 18107 7939
rect 18049 7899 18107 7905
rect 13372 7840 14136 7868
rect 15841 7871 15899 7877
rect 12345 7831 12403 7837
rect 15841 7837 15853 7871
rect 15887 7868 15899 7871
rect 15933 7871 15991 7877
rect 15933 7868 15945 7871
rect 15887 7840 15945 7868
rect 15887 7837 15899 7840
rect 15841 7831 15899 7837
rect 15933 7837 15945 7840
rect 15979 7837 15991 7871
rect 16206 7868 16212 7880
rect 16167 7840 16212 7868
rect 15933 7831 15991 7837
rect 16206 7828 16212 7840
rect 16264 7828 16270 7880
rect 17497 7871 17555 7877
rect 17497 7837 17509 7871
rect 17543 7837 17555 7871
rect 17497 7831 17555 7837
rect 17512 7800 17540 7831
rect 17678 7828 17684 7880
rect 17736 7868 17742 7880
rect 18141 7871 18199 7877
rect 18141 7868 18153 7871
rect 17736 7840 18153 7868
rect 17736 7828 17742 7840
rect 18141 7837 18153 7840
rect 18187 7837 18199 7871
rect 18141 7831 18199 7837
rect 18233 7871 18291 7877
rect 18233 7837 18245 7871
rect 18279 7837 18291 7871
rect 18233 7831 18291 7837
rect 18248 7800 18276 7831
rect 11624 7772 12020 7800
rect 16224 7772 18276 7800
rect 10137 7735 10195 7741
rect 10137 7701 10149 7735
rect 10183 7732 10195 7735
rect 11330 7732 11336 7744
rect 10183 7704 11336 7732
rect 10183 7701 10195 7704
rect 10137 7695 10195 7701
rect 11330 7692 11336 7704
rect 11388 7692 11394 7744
rect 12253 7735 12311 7741
rect 12253 7701 12265 7735
rect 12299 7732 12311 7735
rect 14274 7732 14280 7744
rect 12299 7704 14280 7732
rect 12299 7701 12311 7704
rect 12253 7695 12311 7701
rect 14274 7692 14280 7704
rect 14332 7692 14338 7744
rect 14461 7735 14519 7741
rect 14461 7701 14473 7735
rect 14507 7732 14519 7735
rect 14734 7732 14740 7744
rect 14507 7704 14740 7732
rect 14507 7701 14519 7704
rect 14461 7695 14519 7701
rect 14734 7692 14740 7704
rect 14792 7732 14798 7744
rect 16224 7732 16252 7772
rect 16850 7732 16856 7744
rect 14792 7704 16252 7732
rect 16811 7704 16856 7732
rect 14792 7692 14798 7704
rect 16850 7692 16856 7704
rect 16908 7692 16914 7744
rect 16942 7692 16948 7744
rect 17000 7732 17006 7744
rect 17681 7735 17739 7741
rect 17681 7732 17693 7735
rect 17000 7704 17693 7732
rect 17000 7692 17006 7704
rect 17681 7701 17693 7704
rect 17727 7701 17739 7735
rect 17681 7695 17739 7701
rect 1104 7642 18860 7664
rect 1104 7590 3947 7642
rect 3999 7590 4011 7642
rect 4063 7590 4075 7642
rect 4127 7590 4139 7642
rect 4191 7590 9878 7642
rect 9930 7590 9942 7642
rect 9994 7590 10006 7642
rect 10058 7590 10070 7642
rect 10122 7590 15808 7642
rect 15860 7590 15872 7642
rect 15924 7590 15936 7642
rect 15988 7590 16000 7642
rect 16052 7590 18860 7642
rect 1104 7568 18860 7590
rect 1581 7531 1639 7537
rect 1581 7497 1593 7531
rect 1627 7528 1639 7531
rect 1946 7528 1952 7540
rect 1627 7500 1952 7528
rect 1627 7497 1639 7500
rect 1581 7491 1639 7497
rect 1946 7488 1952 7500
rect 2004 7528 2010 7540
rect 3142 7528 3148 7540
rect 2004 7500 3148 7528
rect 2004 7488 2010 7500
rect 3142 7488 3148 7500
rect 3200 7488 3206 7540
rect 4157 7531 4215 7537
rect 4157 7497 4169 7531
rect 4203 7528 4215 7531
rect 4246 7528 4252 7540
rect 4203 7500 4252 7528
rect 4203 7497 4215 7500
rect 4157 7491 4215 7497
rect 4246 7488 4252 7500
rect 4304 7488 4310 7540
rect 4798 7528 4804 7540
rect 4759 7500 4804 7528
rect 4798 7488 4804 7500
rect 4856 7488 4862 7540
rect 5810 7488 5816 7540
rect 5868 7528 5874 7540
rect 7561 7531 7619 7537
rect 7561 7528 7573 7531
rect 5868 7500 7573 7528
rect 5868 7488 5874 7500
rect 7561 7497 7573 7500
rect 7607 7497 7619 7531
rect 7561 7491 7619 7497
rect 8478 7488 8484 7540
rect 8536 7528 8542 7540
rect 8665 7531 8723 7537
rect 8665 7528 8677 7531
rect 8536 7500 8677 7528
rect 8536 7488 8542 7500
rect 8665 7497 8677 7500
rect 8711 7497 8723 7531
rect 8665 7491 8723 7497
rect 11882 7488 11888 7540
rect 11940 7528 11946 7540
rect 13173 7531 13231 7537
rect 13173 7528 13185 7531
rect 11940 7500 13185 7528
rect 11940 7488 11946 7500
rect 13173 7497 13185 7500
rect 13219 7497 13231 7531
rect 16666 7528 16672 7540
rect 16627 7500 16672 7528
rect 13173 7491 13231 7497
rect 16666 7488 16672 7500
rect 16724 7488 16730 7540
rect 17770 7528 17776 7540
rect 17731 7500 17776 7528
rect 17770 7488 17776 7500
rect 17828 7488 17834 7540
rect 2498 7420 2504 7472
rect 2556 7460 2562 7472
rect 4525 7463 4583 7469
rect 4525 7460 4537 7463
rect 2556 7432 4537 7460
rect 2556 7420 2562 7432
rect 4525 7429 4537 7432
rect 4571 7429 4583 7463
rect 4525 7423 4583 7429
rect 6178 7420 6184 7472
rect 6236 7460 6242 7472
rect 6457 7463 6515 7469
rect 6457 7460 6469 7463
rect 6236 7432 6469 7460
rect 6236 7420 6242 7432
rect 6457 7429 6469 7432
rect 6503 7429 6515 7463
rect 6457 7423 6515 7429
rect 7944 7432 9260 7460
rect 1949 7395 2007 7401
rect 1949 7361 1961 7395
rect 1995 7392 2007 7395
rect 2774 7392 2780 7404
rect 1995 7364 2780 7392
rect 1995 7361 2007 7364
rect 1949 7355 2007 7361
rect 2774 7352 2780 7364
rect 2832 7352 2838 7404
rect 3142 7392 3148 7404
rect 3103 7364 3148 7392
rect 3142 7352 3148 7364
rect 3200 7352 3206 7404
rect 3602 7392 3608 7404
rect 3563 7364 3608 7392
rect 3602 7352 3608 7364
rect 3660 7352 3666 7404
rect 3697 7395 3755 7401
rect 3697 7361 3709 7395
rect 3743 7392 3755 7395
rect 3786 7392 3792 7404
rect 3743 7364 3792 7392
rect 3743 7361 3755 7364
rect 3697 7355 3755 7361
rect 3786 7352 3792 7364
rect 3844 7352 3850 7404
rect 3970 7352 3976 7404
rect 4028 7392 4034 7404
rect 4249 7395 4307 7401
rect 4249 7392 4261 7395
rect 4028 7364 4261 7392
rect 4028 7352 4034 7364
rect 4249 7361 4261 7364
rect 4295 7361 4307 7395
rect 4249 7355 4307 7361
rect 6270 7352 6276 7404
rect 6328 7392 6334 7404
rect 7009 7395 7067 7401
rect 7009 7392 7021 7395
rect 6328 7364 7021 7392
rect 6328 7352 6334 7364
rect 7009 7361 7021 7364
rect 7055 7361 7067 7395
rect 7009 7355 7067 7361
rect 7834 7352 7840 7404
rect 7892 7392 7898 7404
rect 7944 7401 7972 7432
rect 7929 7395 7987 7401
rect 7929 7392 7941 7395
rect 7892 7364 7941 7392
rect 7892 7352 7898 7364
rect 7929 7361 7941 7364
rect 7975 7361 7987 7395
rect 7929 7355 7987 7361
rect 8113 7395 8171 7401
rect 8113 7361 8125 7395
rect 8159 7392 8171 7395
rect 8202 7392 8208 7404
rect 8159 7364 8208 7392
rect 8159 7361 8171 7364
rect 8113 7355 8171 7361
rect 8202 7352 8208 7364
rect 8260 7352 8266 7404
rect 8662 7392 8668 7404
rect 8312 7364 8668 7392
rect 1394 7324 1400 7336
rect 1355 7296 1400 7324
rect 1394 7284 1400 7296
rect 1452 7284 1458 7336
rect 2038 7324 2044 7336
rect 1999 7296 2044 7324
rect 2038 7284 2044 7296
rect 2096 7284 2102 7336
rect 2130 7284 2136 7336
rect 2188 7324 2194 7336
rect 4062 7324 4068 7336
rect 2188 7296 2233 7324
rect 2332 7296 4068 7324
rect 2188 7284 2194 7296
rect 1412 7256 1440 7284
rect 2332 7256 2360 7296
rect 4062 7284 4068 7296
rect 4120 7284 4126 7336
rect 4154 7284 4160 7336
rect 4212 7324 4218 7336
rect 4709 7327 4767 7333
rect 4709 7324 4721 7327
rect 4212 7296 4721 7324
rect 4212 7284 4218 7296
rect 4709 7293 4721 7296
rect 4755 7324 4767 7327
rect 4982 7324 4988 7336
rect 4755 7296 4988 7324
rect 4755 7293 4767 7296
rect 4709 7287 4767 7293
rect 4982 7284 4988 7296
rect 5040 7284 5046 7336
rect 6181 7327 6239 7333
rect 6181 7293 6193 7327
rect 6227 7293 6239 7327
rect 6181 7287 6239 7293
rect 4338 7256 4344 7268
rect 1412 7228 2360 7256
rect 2516 7228 4344 7256
rect 2516 7197 2544 7228
rect 4338 7216 4344 7228
rect 4396 7216 4402 7268
rect 4890 7216 4896 7268
rect 4948 7256 4954 7268
rect 5442 7256 5448 7268
rect 4948 7228 5448 7256
rect 4948 7216 4954 7228
rect 5442 7216 5448 7228
rect 5500 7216 5506 7268
rect 5534 7216 5540 7268
rect 5592 7256 5598 7268
rect 5914 7259 5972 7265
rect 5914 7256 5926 7259
rect 5592 7228 5926 7256
rect 5592 7216 5598 7228
rect 5914 7225 5926 7228
rect 5960 7225 5972 7259
rect 6196 7256 6224 7287
rect 6454 7284 6460 7336
rect 6512 7324 6518 7336
rect 6825 7327 6883 7333
rect 6825 7324 6837 7327
rect 6512 7296 6837 7324
rect 6512 7284 6518 7296
rect 6825 7293 6837 7296
rect 6871 7293 6883 7327
rect 6825 7287 6883 7293
rect 7374 7284 7380 7336
rect 7432 7324 7438 7336
rect 7558 7324 7564 7336
rect 7432 7296 7564 7324
rect 7432 7284 7438 7296
rect 7558 7284 7564 7296
rect 7616 7284 7622 7336
rect 7745 7327 7803 7333
rect 7745 7293 7757 7327
rect 7791 7324 7803 7327
rect 8312 7324 8340 7364
rect 8662 7352 8668 7364
rect 8720 7352 8726 7404
rect 9232 7401 9260 7432
rect 9674 7420 9680 7472
rect 9732 7460 9738 7472
rect 11422 7460 11428 7472
rect 9732 7432 11428 7460
rect 9732 7420 9738 7432
rect 11422 7420 11428 7432
rect 11480 7420 11486 7472
rect 12894 7420 12900 7472
rect 12952 7460 12958 7472
rect 13081 7463 13139 7469
rect 13081 7460 13093 7463
rect 12952 7432 13093 7460
rect 12952 7420 12958 7432
rect 13081 7429 13093 7432
rect 13127 7429 13139 7463
rect 13081 7423 13139 7429
rect 13538 7420 13544 7472
rect 13596 7420 13602 7472
rect 17678 7460 17684 7472
rect 17639 7432 17684 7460
rect 17678 7420 17684 7432
rect 17736 7420 17742 7472
rect 9217 7395 9275 7401
rect 9217 7361 9229 7395
rect 9263 7361 9275 7395
rect 9217 7355 9275 7361
rect 9306 7352 9312 7404
rect 9364 7392 9370 7404
rect 9585 7395 9643 7401
rect 9585 7392 9597 7395
rect 9364 7364 9597 7392
rect 9364 7352 9370 7364
rect 9585 7361 9597 7364
rect 9631 7361 9643 7395
rect 10410 7392 10416 7404
rect 10371 7364 10416 7392
rect 9585 7355 9643 7361
rect 10410 7352 10416 7364
rect 10468 7352 10474 7404
rect 11606 7352 11612 7404
rect 11664 7392 11670 7404
rect 11701 7395 11759 7401
rect 11701 7392 11713 7395
rect 11664 7364 11713 7392
rect 11664 7352 11670 7364
rect 11701 7361 11713 7364
rect 11747 7361 11759 7395
rect 11701 7355 11759 7361
rect 9033 7327 9091 7333
rect 9033 7324 9045 7327
rect 7791 7296 8340 7324
rect 8404 7296 9045 7324
rect 7791 7293 7803 7296
rect 7745 7287 7803 7293
rect 6730 7256 6736 7268
rect 6196 7228 6736 7256
rect 5914 7219 5972 7225
rect 6730 7216 6736 7228
rect 6788 7216 6794 7268
rect 7469 7259 7527 7265
rect 7469 7225 7481 7259
rect 7515 7256 7527 7259
rect 8404 7256 8432 7296
rect 9033 7293 9045 7296
rect 9079 7293 9091 7327
rect 9033 7287 9091 7293
rect 9122 7284 9128 7336
rect 9180 7324 9186 7336
rect 10689 7327 10747 7333
rect 10689 7324 10701 7327
rect 9180 7296 10701 7324
rect 9180 7284 9186 7296
rect 10689 7293 10701 7296
rect 10735 7293 10747 7327
rect 11330 7324 11336 7336
rect 11291 7296 11336 7324
rect 10689 7287 10747 7293
rect 11330 7284 11336 7296
rect 11388 7284 11394 7336
rect 13556 7333 13584 7420
rect 13722 7392 13728 7404
rect 13683 7364 13728 7392
rect 13722 7352 13728 7364
rect 13780 7352 13786 7404
rect 14366 7352 14372 7404
rect 14424 7392 14430 7404
rect 14461 7395 14519 7401
rect 14461 7392 14473 7395
rect 14424 7364 14473 7392
rect 14424 7352 14430 7364
rect 14461 7361 14473 7364
rect 14507 7361 14519 7395
rect 14461 7355 14519 7361
rect 16117 7395 16175 7401
rect 16117 7361 16129 7395
rect 16163 7392 16175 7395
rect 16206 7392 16212 7404
rect 16163 7364 16212 7392
rect 16163 7361 16175 7364
rect 16117 7355 16175 7361
rect 16206 7352 16212 7364
rect 16264 7392 16270 7404
rect 17129 7395 17187 7401
rect 17129 7392 17141 7395
rect 16264 7364 17141 7392
rect 16264 7352 16270 7364
rect 17129 7361 17141 7364
rect 17175 7392 17187 7395
rect 18322 7392 18328 7404
rect 17175 7364 18328 7392
rect 17175 7361 17187 7364
rect 17129 7355 17187 7361
rect 18322 7352 18328 7364
rect 18380 7352 18386 7404
rect 13541 7327 13599 7333
rect 11808 7296 12112 7324
rect 9769 7259 9827 7265
rect 9769 7256 9781 7259
rect 7515 7228 8432 7256
rect 8588 7228 9781 7256
rect 7515 7225 7527 7228
rect 7469 7219 7527 7225
rect 2501 7191 2559 7197
rect 2501 7157 2513 7191
rect 2547 7157 2559 7191
rect 2501 7151 2559 7157
rect 2590 7148 2596 7200
rect 2648 7188 2654 7200
rect 2958 7188 2964 7200
rect 2648 7160 2693 7188
rect 2919 7160 2964 7188
rect 2648 7148 2654 7160
rect 2958 7148 2964 7160
rect 3016 7148 3022 7200
rect 3050 7148 3056 7200
rect 3108 7188 3114 7200
rect 3789 7191 3847 7197
rect 3108 7160 3153 7188
rect 3108 7148 3114 7160
rect 3789 7157 3801 7191
rect 3835 7188 3847 7191
rect 4706 7188 4712 7200
rect 3835 7160 4712 7188
rect 3835 7157 3847 7160
rect 3789 7151 3847 7157
rect 4706 7148 4712 7160
rect 4764 7148 4770 7200
rect 6454 7148 6460 7200
rect 6512 7188 6518 7200
rect 6917 7191 6975 7197
rect 6917 7188 6929 7191
rect 6512 7160 6929 7188
rect 6512 7148 6518 7160
rect 6917 7157 6929 7160
rect 6963 7188 6975 7191
rect 7742 7188 7748 7200
rect 6963 7160 7748 7188
rect 6963 7157 6975 7160
rect 6917 7151 6975 7157
rect 7742 7148 7748 7160
rect 7800 7148 7806 7200
rect 8018 7148 8024 7200
rect 8076 7188 8082 7200
rect 8588 7197 8616 7228
rect 9769 7225 9781 7228
rect 9815 7225 9827 7259
rect 11808 7256 11836 7296
rect 9769 7219 9827 7225
rect 11072 7228 11836 7256
rect 8205 7191 8263 7197
rect 8205 7188 8217 7191
rect 8076 7160 8217 7188
rect 8076 7148 8082 7160
rect 8205 7157 8217 7160
rect 8251 7157 8263 7191
rect 8205 7151 8263 7157
rect 8573 7191 8631 7197
rect 8573 7157 8585 7191
rect 8619 7157 8631 7191
rect 8573 7151 8631 7157
rect 8662 7148 8668 7200
rect 8720 7188 8726 7200
rect 9125 7191 9183 7197
rect 9125 7188 9137 7191
rect 8720 7160 9137 7188
rect 8720 7148 8726 7160
rect 9125 7157 9137 7160
rect 9171 7188 9183 7191
rect 9674 7188 9680 7200
rect 9171 7160 9680 7188
rect 9171 7157 9183 7160
rect 9125 7151 9183 7157
rect 9674 7148 9680 7160
rect 9732 7148 9738 7200
rect 9858 7188 9864 7200
rect 9819 7160 9864 7188
rect 9858 7148 9864 7160
rect 9916 7148 9922 7200
rect 11072 7197 11100 7228
rect 11882 7216 11888 7268
rect 11940 7265 11946 7268
rect 11940 7259 12004 7265
rect 11940 7225 11958 7259
rect 11992 7225 12004 7259
rect 12084 7256 12112 7296
rect 13541 7293 13553 7327
rect 13587 7293 13599 7327
rect 13541 7287 13599 7293
rect 14090 7284 14096 7336
rect 14148 7324 14154 7336
rect 14734 7333 14740 7336
rect 14185 7327 14243 7333
rect 14185 7324 14197 7327
rect 14148 7296 14197 7324
rect 14148 7284 14154 7296
rect 14185 7293 14197 7296
rect 14231 7293 14243 7327
rect 14728 7324 14740 7333
rect 14695 7296 14740 7324
rect 14185 7287 14243 7293
rect 14728 7287 14740 7296
rect 14734 7284 14740 7287
rect 14792 7284 14798 7336
rect 15654 7284 15660 7336
rect 15712 7324 15718 7336
rect 18233 7327 18291 7333
rect 18233 7324 18245 7327
rect 15712 7296 18245 7324
rect 15712 7284 15718 7296
rect 18233 7293 18245 7296
rect 18279 7293 18291 7327
rect 18233 7287 18291 7293
rect 13633 7259 13691 7265
rect 12084 7228 13400 7256
rect 11940 7219 12004 7225
rect 11940 7216 11946 7219
rect 10229 7191 10287 7197
rect 10229 7157 10241 7191
rect 10275 7188 10287 7191
rect 10597 7191 10655 7197
rect 10597 7188 10609 7191
rect 10275 7160 10609 7188
rect 10275 7157 10287 7160
rect 10229 7151 10287 7157
rect 10597 7157 10609 7160
rect 10643 7157 10655 7191
rect 10597 7151 10655 7157
rect 11057 7191 11115 7197
rect 11057 7157 11069 7191
rect 11103 7157 11115 7191
rect 11057 7151 11115 7157
rect 11241 7191 11299 7197
rect 11241 7157 11253 7191
rect 11287 7188 11299 7191
rect 11330 7188 11336 7200
rect 11287 7160 11336 7188
rect 11287 7157 11299 7160
rect 11241 7151 11299 7157
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 11517 7191 11575 7197
rect 11517 7157 11529 7191
rect 11563 7188 11575 7191
rect 12250 7188 12256 7200
rect 11563 7160 12256 7188
rect 11563 7157 11575 7160
rect 11517 7151 11575 7157
rect 12250 7148 12256 7160
rect 12308 7188 12314 7200
rect 13262 7188 13268 7200
rect 12308 7160 13268 7188
rect 12308 7148 12314 7160
rect 13262 7148 13268 7160
rect 13320 7148 13326 7200
rect 13372 7188 13400 7228
rect 13633 7225 13645 7259
rect 13679 7256 13691 7259
rect 14550 7256 14556 7268
rect 13679 7228 14556 7256
rect 13679 7225 13691 7228
rect 13633 7219 13691 7225
rect 14550 7216 14556 7228
rect 14608 7216 14614 7268
rect 15286 7216 15292 7268
rect 15344 7256 15350 7268
rect 15562 7256 15568 7268
rect 15344 7228 15568 7256
rect 15344 7216 15350 7228
rect 15562 7216 15568 7228
rect 15620 7216 15626 7268
rect 18322 7256 18328 7268
rect 15672 7228 18328 7256
rect 13814 7188 13820 7200
rect 13372 7160 13820 7188
rect 13814 7148 13820 7160
rect 13872 7148 13878 7200
rect 13998 7188 14004 7200
rect 13959 7160 14004 7188
rect 13998 7148 14004 7160
rect 14056 7148 14062 7200
rect 14369 7191 14427 7197
rect 14369 7157 14381 7191
rect 14415 7188 14427 7191
rect 15672 7188 15700 7228
rect 18322 7216 18328 7228
rect 18380 7216 18386 7268
rect 15838 7188 15844 7200
rect 14415 7160 15700 7188
rect 15799 7160 15844 7188
rect 14415 7157 14427 7160
rect 14369 7151 14427 7157
rect 15838 7148 15844 7160
rect 15896 7148 15902 7200
rect 16022 7148 16028 7200
rect 16080 7188 16086 7200
rect 16209 7191 16267 7197
rect 16209 7188 16221 7191
rect 16080 7160 16221 7188
rect 16080 7148 16086 7160
rect 16209 7157 16221 7160
rect 16255 7157 16267 7191
rect 16209 7151 16267 7157
rect 16298 7148 16304 7200
rect 16356 7188 16362 7200
rect 16356 7160 16401 7188
rect 16356 7148 16362 7160
rect 17126 7148 17132 7200
rect 17184 7188 17190 7200
rect 17221 7191 17279 7197
rect 17221 7188 17233 7191
rect 17184 7160 17233 7188
rect 17184 7148 17190 7160
rect 17221 7157 17233 7160
rect 17267 7157 17279 7191
rect 17221 7151 17279 7157
rect 17313 7191 17371 7197
rect 17313 7157 17325 7191
rect 17359 7188 17371 7191
rect 17402 7188 17408 7200
rect 17359 7160 17408 7188
rect 17359 7157 17371 7160
rect 17313 7151 17371 7157
rect 17402 7148 17408 7160
rect 17460 7148 17466 7200
rect 18138 7188 18144 7200
rect 18099 7160 18144 7188
rect 18138 7148 18144 7160
rect 18196 7148 18202 7200
rect 1104 7098 18860 7120
rect 1104 7046 6912 7098
rect 6964 7046 6976 7098
rect 7028 7046 7040 7098
rect 7092 7046 7104 7098
rect 7156 7046 12843 7098
rect 12895 7046 12907 7098
rect 12959 7046 12971 7098
rect 13023 7046 13035 7098
rect 13087 7046 18860 7098
rect 1104 7024 18860 7046
rect 2958 6984 2964 6996
rect 2919 6956 2964 6984
rect 2958 6944 2964 6956
rect 3016 6944 3022 6996
rect 3329 6987 3387 6993
rect 3329 6953 3341 6987
rect 3375 6984 3387 6987
rect 3970 6984 3976 6996
rect 3375 6956 3976 6984
rect 3375 6953 3387 6956
rect 3329 6947 3387 6953
rect 3970 6944 3976 6956
rect 4028 6944 4034 6996
rect 4249 6987 4307 6993
rect 4249 6953 4261 6987
rect 4295 6984 4307 6987
rect 4890 6984 4896 6996
rect 4295 6956 4896 6984
rect 4295 6953 4307 6956
rect 4249 6947 4307 6953
rect 4890 6944 4896 6956
rect 4948 6944 4954 6996
rect 5166 6944 5172 6996
rect 5224 6984 5230 6996
rect 11330 6984 11336 6996
rect 5224 6956 11336 6984
rect 5224 6944 5230 6956
rect 11330 6944 11336 6956
rect 11388 6944 11394 6996
rect 11514 6984 11520 6996
rect 11475 6956 11520 6984
rect 11514 6944 11520 6956
rect 11572 6944 11578 6996
rect 11609 6987 11667 6993
rect 11609 6953 11621 6987
rect 11655 6953 11667 6987
rect 11609 6947 11667 6953
rect 4062 6876 4068 6928
rect 4120 6916 4126 6928
rect 6641 6919 6699 6925
rect 6641 6916 6653 6919
rect 4120 6888 6653 6916
rect 4120 6876 4126 6888
rect 6641 6885 6653 6888
rect 6687 6885 6699 6919
rect 6641 6879 6699 6885
rect 7101 6919 7159 6925
rect 7101 6885 7113 6919
rect 7147 6916 7159 6919
rect 7374 6916 7380 6928
rect 7147 6888 7380 6916
rect 7147 6885 7159 6888
rect 7101 6879 7159 6885
rect 7374 6876 7380 6888
rect 7432 6876 7438 6928
rect 7742 6876 7748 6928
rect 7800 6916 7806 6928
rect 8021 6919 8079 6925
rect 8021 6916 8033 6919
rect 7800 6888 8033 6916
rect 7800 6876 7806 6888
rect 8021 6885 8033 6888
rect 8067 6916 8079 6919
rect 8202 6916 8208 6928
rect 8067 6888 8208 6916
rect 8067 6885 8079 6888
rect 8021 6879 8079 6885
rect 8202 6876 8208 6888
rect 8260 6876 8266 6928
rect 8938 6876 8944 6928
rect 8996 6916 9002 6928
rect 9674 6916 9680 6928
rect 8996 6888 9680 6916
rect 8996 6876 9002 6888
rect 9674 6876 9680 6888
rect 9732 6916 9738 6928
rect 10597 6919 10655 6925
rect 10597 6916 10609 6919
rect 9732 6888 10609 6916
rect 9732 6876 9738 6888
rect 10597 6885 10609 6888
rect 10643 6885 10655 6919
rect 11624 6916 11652 6947
rect 12066 6944 12072 6996
rect 12124 6984 12130 6996
rect 13449 6987 13507 6993
rect 12124 6956 13400 6984
rect 12124 6944 12130 6956
rect 11790 6916 11796 6928
rect 10597 6879 10655 6885
rect 10980 6888 11796 6916
rect 1756 6851 1814 6857
rect 1756 6817 1768 6851
rect 1802 6848 1814 6851
rect 3421 6851 3479 6857
rect 1802 6820 2774 6848
rect 1802 6817 1814 6820
rect 1756 6811 1814 6817
rect 1489 6783 1547 6789
rect 1489 6749 1501 6783
rect 1535 6749 1547 6783
rect 2746 6780 2774 6820
rect 3421 6817 3433 6851
rect 3467 6848 3479 6851
rect 4154 6848 4160 6860
rect 3467 6820 4160 6848
rect 3467 6817 3479 6820
rect 3421 6811 3479 6817
rect 4154 6808 4160 6820
rect 4212 6808 4218 6860
rect 4341 6851 4399 6857
rect 4341 6817 4353 6851
rect 4387 6848 4399 6851
rect 4893 6851 4951 6857
rect 4387 6820 4568 6848
rect 4387 6817 4399 6820
rect 4341 6811 4399 6817
rect 3234 6780 3240 6792
rect 2746 6752 3240 6780
rect 1489 6743 1547 6749
rect 1504 6644 1532 6743
rect 3234 6740 3240 6752
rect 3292 6780 3298 6792
rect 3605 6783 3663 6789
rect 3605 6780 3617 6783
rect 3292 6752 3617 6780
rect 3292 6740 3298 6752
rect 3605 6749 3617 6752
rect 3651 6780 3663 6783
rect 4433 6783 4491 6789
rect 4433 6780 4445 6783
rect 3651 6752 4445 6780
rect 3651 6749 3663 6752
rect 3605 6743 3663 6749
rect 4433 6749 4445 6752
rect 4479 6749 4491 6783
rect 4433 6743 4491 6749
rect 3050 6672 3056 6724
rect 3108 6712 3114 6724
rect 3881 6715 3939 6721
rect 3881 6712 3893 6715
rect 3108 6684 3893 6712
rect 3108 6672 3114 6684
rect 3881 6681 3893 6684
rect 3927 6681 3939 6715
rect 4540 6712 4568 6820
rect 4893 6817 4905 6851
rect 4939 6848 4951 6851
rect 5810 6848 5816 6860
rect 4939 6820 5816 6848
rect 4939 6817 4951 6820
rect 4893 6811 4951 6817
rect 5810 6808 5816 6820
rect 5868 6808 5874 6860
rect 6201 6851 6259 6857
rect 6201 6817 6213 6851
rect 6247 6848 6259 6851
rect 6546 6848 6552 6860
rect 6247 6820 6552 6848
rect 6247 6817 6259 6820
rect 6201 6811 6259 6817
rect 6546 6808 6552 6820
rect 6604 6808 6610 6860
rect 7009 6851 7067 6857
rect 7009 6848 7021 6851
rect 6840 6820 7021 6848
rect 6457 6783 6515 6789
rect 6457 6749 6469 6783
rect 6503 6780 6515 6783
rect 6730 6780 6736 6792
rect 6503 6752 6736 6780
rect 6503 6749 6515 6752
rect 6457 6743 6515 6749
rect 6730 6740 6736 6752
rect 6788 6740 6794 6792
rect 4540 6684 5580 6712
rect 3881 6675 3939 6681
rect 2130 6644 2136 6656
rect 1504 6616 2136 6644
rect 2130 6604 2136 6616
rect 2188 6604 2194 6656
rect 2869 6647 2927 6653
rect 2869 6613 2881 6647
rect 2915 6644 2927 6647
rect 2958 6644 2964 6656
rect 2915 6616 2964 6644
rect 2915 6613 2927 6616
rect 2869 6607 2927 6613
rect 2958 6604 2964 6616
rect 3016 6644 3022 6656
rect 3142 6644 3148 6656
rect 3016 6616 3148 6644
rect 3016 6604 3022 6616
rect 3142 6604 3148 6616
rect 3200 6604 3206 6656
rect 3786 6604 3792 6656
rect 3844 6644 3850 6656
rect 4801 6647 4859 6653
rect 4801 6644 4813 6647
rect 3844 6616 4813 6644
rect 3844 6604 3850 6616
rect 4801 6613 4813 6616
rect 4847 6613 4859 6647
rect 4801 6607 4859 6613
rect 5077 6647 5135 6653
rect 5077 6613 5089 6647
rect 5123 6644 5135 6647
rect 5442 6644 5448 6656
rect 5123 6616 5448 6644
rect 5123 6613 5135 6616
rect 5077 6607 5135 6613
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 5552 6644 5580 6684
rect 6270 6644 6276 6656
rect 5552 6616 6276 6644
rect 6270 6604 6276 6616
rect 6328 6644 6334 6656
rect 6840 6644 6868 6820
rect 7009 6817 7021 6820
rect 7055 6848 7067 6851
rect 7190 6848 7196 6860
rect 7055 6820 7196 6848
rect 7055 6817 7067 6820
rect 7009 6811 7067 6817
rect 7190 6808 7196 6820
rect 7248 6808 7254 6860
rect 7558 6808 7564 6860
rect 7616 6848 7622 6860
rect 7929 6851 7987 6857
rect 7929 6848 7941 6851
rect 7616 6820 7941 6848
rect 7616 6808 7622 6820
rect 7929 6817 7941 6820
rect 7975 6817 7987 6851
rect 7929 6811 7987 6817
rect 6917 6783 6975 6789
rect 6917 6749 6929 6783
rect 6963 6749 6975 6783
rect 7745 6783 7803 6789
rect 7745 6780 7757 6783
rect 6917 6743 6975 6749
rect 7300 6752 7757 6780
rect 6932 6712 6960 6743
rect 7300 6712 7328 6752
rect 7745 6749 7757 6752
rect 7791 6780 7803 6783
rect 7834 6780 7840 6792
rect 7791 6752 7840 6780
rect 7791 6749 7803 6752
rect 7745 6743 7803 6749
rect 7834 6740 7840 6752
rect 7892 6740 7898 6792
rect 7944 6780 7972 6811
rect 8386 6808 8392 6860
rect 8444 6848 8450 6860
rect 8481 6851 8539 6857
rect 8481 6848 8493 6851
rect 8444 6820 8493 6848
rect 8444 6808 8450 6820
rect 8481 6817 8493 6820
rect 8527 6817 8539 6851
rect 8754 6848 8760 6860
rect 8715 6820 8760 6848
rect 8481 6811 8539 6817
rect 8754 6808 8760 6820
rect 8812 6808 8818 6860
rect 9858 6848 9864 6860
rect 9048 6820 9864 6848
rect 8938 6780 8944 6792
rect 7944 6752 8944 6780
rect 8938 6740 8944 6752
rect 8996 6740 9002 6792
rect 7466 6712 7472 6724
rect 6932 6684 7328 6712
rect 7427 6684 7472 6712
rect 7466 6672 7472 6684
rect 7524 6672 7530 6724
rect 8389 6715 8447 6721
rect 8389 6681 8401 6715
rect 8435 6712 8447 6715
rect 9048 6712 9076 6820
rect 9858 6808 9864 6820
rect 9916 6808 9922 6860
rect 10249 6851 10307 6857
rect 10249 6817 10261 6851
rect 10295 6848 10307 6851
rect 10410 6848 10416 6860
rect 10295 6820 10416 6848
rect 10295 6817 10307 6820
rect 10249 6811 10307 6817
rect 10410 6808 10416 6820
rect 10468 6808 10474 6860
rect 10980 6789 11008 6888
rect 11790 6876 11796 6888
rect 11848 6916 11854 6928
rect 13372 6916 13400 6956
rect 13449 6953 13461 6987
rect 13495 6984 13507 6987
rect 13538 6984 13544 6996
rect 13495 6956 13544 6984
rect 13495 6953 13507 6956
rect 13449 6947 13507 6953
rect 13538 6944 13544 6956
rect 13596 6944 13602 6996
rect 13817 6987 13875 6993
rect 13817 6953 13829 6987
rect 13863 6984 13875 6987
rect 13906 6984 13912 6996
rect 13863 6956 13912 6984
rect 13863 6953 13875 6956
rect 13817 6947 13875 6953
rect 13906 6944 13912 6956
rect 13964 6984 13970 6996
rect 16482 6984 16488 6996
rect 13964 6956 16488 6984
rect 13964 6944 13970 6956
rect 16482 6944 16488 6956
rect 16540 6944 16546 6996
rect 16758 6944 16764 6996
rect 16816 6984 16822 6996
rect 17313 6987 17371 6993
rect 17313 6984 17325 6987
rect 16816 6956 17325 6984
rect 16816 6944 16822 6956
rect 17313 6953 17325 6956
rect 17359 6984 17371 6987
rect 17402 6984 17408 6996
rect 17359 6956 17408 6984
rect 17359 6953 17371 6956
rect 17313 6947 17371 6953
rect 17402 6944 17408 6956
rect 17460 6944 17466 6996
rect 15654 6916 15660 6928
rect 11848 6888 13308 6916
rect 13372 6888 15660 6916
rect 11848 6876 11854 6888
rect 11146 6848 11152 6860
rect 11107 6820 11152 6848
rect 11146 6808 11152 6820
rect 11204 6808 11210 6860
rect 12158 6808 12164 6860
rect 12216 6848 12222 6860
rect 12710 6848 12716 6860
rect 12768 6857 12774 6860
rect 12216 6820 12716 6848
rect 12216 6808 12222 6820
rect 12710 6808 12716 6820
rect 12768 6848 12780 6857
rect 13173 6851 13231 6857
rect 12768 6820 12813 6848
rect 12768 6811 12780 6820
rect 13173 6817 13185 6851
rect 13219 6817 13231 6851
rect 13280 6848 13308 6888
rect 15654 6876 15660 6888
rect 15712 6876 15718 6928
rect 15838 6876 15844 6928
rect 15896 6916 15902 6928
rect 16086 6919 16144 6925
rect 16086 6916 16098 6919
rect 15896 6888 16098 6916
rect 15896 6876 15902 6888
rect 16086 6885 16098 6888
rect 16132 6916 16144 6919
rect 16206 6916 16212 6928
rect 16132 6888 16212 6916
rect 16132 6885 16144 6888
rect 16086 6879 16144 6885
rect 16206 6876 16212 6888
rect 16264 6876 16270 6928
rect 13722 6848 13728 6860
rect 13280 6820 13728 6848
rect 13173 6811 13231 6817
rect 12768 6808 12774 6811
rect 10505 6783 10563 6789
rect 10505 6749 10517 6783
rect 10551 6749 10563 6783
rect 10505 6743 10563 6749
rect 10965 6783 11023 6789
rect 10965 6749 10977 6783
rect 11011 6749 11023 6783
rect 10965 6743 11023 6749
rect 11057 6783 11115 6789
rect 11057 6749 11069 6783
rect 11103 6780 11115 6783
rect 11514 6780 11520 6792
rect 11103 6752 11520 6780
rect 11103 6749 11115 6752
rect 11057 6743 11115 6749
rect 8435 6684 9076 6712
rect 10520 6712 10548 6743
rect 11514 6740 11520 6752
rect 11572 6740 11578 6792
rect 11606 6740 11612 6792
rect 11664 6780 11670 6792
rect 11974 6780 11980 6792
rect 11664 6752 11980 6780
rect 11664 6740 11670 6752
rect 11974 6740 11980 6752
rect 12032 6740 12038 6792
rect 12989 6783 13047 6789
rect 12989 6749 13001 6783
rect 13035 6780 13047 6783
rect 13078 6780 13084 6792
rect 13035 6752 13084 6780
rect 13035 6749 13047 6752
rect 12989 6743 13047 6749
rect 13078 6740 13084 6752
rect 13136 6740 13142 6792
rect 11422 6712 11428 6724
rect 10520 6684 11428 6712
rect 8435 6681 8447 6684
rect 8389 6675 8447 6681
rect 11422 6672 11428 6684
rect 11480 6672 11486 6724
rect 6328 6616 6868 6644
rect 8665 6647 8723 6653
rect 6328 6604 6334 6616
rect 8665 6613 8677 6647
rect 8711 6644 8723 6647
rect 8754 6644 8760 6656
rect 8711 6616 8760 6644
rect 8711 6613 8723 6616
rect 8665 6607 8723 6613
rect 8754 6604 8760 6616
rect 8812 6604 8818 6656
rect 8846 6604 8852 6656
rect 8904 6644 8910 6656
rect 8941 6647 8999 6653
rect 8941 6644 8953 6647
rect 8904 6616 8953 6644
rect 8904 6604 8910 6616
rect 8941 6613 8953 6616
rect 8987 6613 8999 6647
rect 8941 6607 8999 6613
rect 9125 6647 9183 6653
rect 9125 6613 9137 6647
rect 9171 6644 9183 6647
rect 9306 6644 9312 6656
rect 9171 6616 9312 6644
rect 9171 6613 9183 6616
rect 9125 6607 9183 6613
rect 9306 6604 9312 6616
rect 9364 6604 9370 6656
rect 12802 6604 12808 6656
rect 12860 6644 12866 6656
rect 13188 6644 13216 6811
rect 13722 6808 13728 6820
rect 13780 6808 13786 6860
rect 14636 6851 14694 6857
rect 13832 6820 14044 6848
rect 13832 6780 13860 6820
rect 13372 6752 13860 6780
rect 13909 6783 13967 6789
rect 13372 6721 13400 6752
rect 13909 6749 13921 6783
rect 13955 6749 13967 6783
rect 13909 6743 13967 6749
rect 13357 6715 13415 6721
rect 13357 6681 13369 6715
rect 13403 6681 13415 6715
rect 13357 6675 13415 6681
rect 13722 6672 13728 6724
rect 13780 6712 13786 6724
rect 13924 6712 13952 6743
rect 13780 6684 13952 6712
rect 13780 6672 13786 6684
rect 12860 6616 13216 6644
rect 14016 6644 14044 6820
rect 14636 6817 14648 6851
rect 14682 6848 14694 6851
rect 14918 6848 14924 6860
rect 14682 6820 14924 6848
rect 14682 6817 14694 6820
rect 14636 6811 14694 6817
rect 14918 6808 14924 6820
rect 14976 6808 14982 6860
rect 17589 6851 17647 6857
rect 17589 6848 17601 6851
rect 15488 6820 17601 6848
rect 14093 6783 14151 6789
rect 14093 6749 14105 6783
rect 14139 6780 14151 6783
rect 14182 6780 14188 6792
rect 14139 6752 14188 6780
rect 14139 6749 14151 6752
rect 14093 6743 14151 6749
rect 14182 6740 14188 6752
rect 14240 6740 14246 6792
rect 14366 6780 14372 6792
rect 14327 6752 14372 6780
rect 14366 6740 14372 6752
rect 14424 6740 14430 6792
rect 15488 6644 15516 6820
rect 17589 6817 17601 6820
rect 17635 6817 17647 6851
rect 17589 6811 17647 6817
rect 17773 6851 17831 6857
rect 17773 6817 17785 6851
rect 17819 6848 17831 6851
rect 17862 6848 17868 6860
rect 17819 6820 17868 6848
rect 17819 6817 17831 6820
rect 17773 6811 17831 6817
rect 17862 6808 17868 6820
rect 17920 6808 17926 6860
rect 17957 6851 18015 6857
rect 17957 6817 17969 6851
rect 18003 6817 18015 6851
rect 17957 6811 18015 6817
rect 18141 6851 18199 6857
rect 18141 6817 18153 6851
rect 18187 6848 18199 6851
rect 18230 6848 18236 6860
rect 18187 6820 18236 6848
rect 18187 6817 18199 6820
rect 18141 6811 18199 6817
rect 15654 6740 15660 6792
rect 15712 6780 15718 6792
rect 15841 6783 15899 6789
rect 15841 6780 15853 6783
rect 15712 6752 15853 6780
rect 15712 6740 15718 6752
rect 15841 6749 15853 6752
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 17402 6740 17408 6792
rect 17460 6780 17466 6792
rect 17972 6780 18000 6811
rect 18230 6808 18236 6820
rect 18288 6808 18294 6860
rect 18322 6808 18328 6860
rect 18380 6848 18386 6860
rect 18380 6820 18425 6848
rect 18380 6808 18386 6820
rect 17460 6752 18000 6780
rect 17460 6740 17466 6752
rect 18506 6712 18512 6724
rect 18467 6684 18512 6712
rect 18506 6672 18512 6684
rect 18564 6672 18570 6724
rect 14016 6616 15516 6644
rect 12860 6604 12866 6616
rect 15562 6604 15568 6656
rect 15620 6644 15626 6656
rect 15749 6647 15807 6653
rect 15749 6644 15761 6647
rect 15620 6616 15761 6644
rect 15620 6604 15626 6616
rect 15749 6613 15761 6616
rect 15795 6613 15807 6647
rect 15749 6607 15807 6613
rect 17221 6647 17279 6653
rect 17221 6613 17233 6647
rect 17267 6644 17279 6647
rect 17678 6644 17684 6656
rect 17267 6616 17684 6644
rect 17267 6613 17279 6616
rect 17221 6607 17279 6613
rect 17678 6604 17684 6616
rect 17736 6604 17742 6656
rect 1104 6554 18860 6576
rect 1104 6502 3947 6554
rect 3999 6502 4011 6554
rect 4063 6502 4075 6554
rect 4127 6502 4139 6554
rect 4191 6502 9878 6554
rect 9930 6502 9942 6554
rect 9994 6502 10006 6554
rect 10058 6502 10070 6554
rect 10122 6502 15808 6554
rect 15860 6502 15872 6554
rect 15924 6502 15936 6554
rect 15988 6502 16000 6554
rect 16052 6502 18860 6554
rect 1104 6480 18860 6502
rect 1765 6443 1823 6449
rect 1765 6409 1777 6443
rect 1811 6440 1823 6443
rect 2314 6440 2320 6452
rect 1811 6412 2320 6440
rect 1811 6409 1823 6412
rect 1765 6403 1823 6409
rect 2314 6400 2320 6412
rect 2372 6440 2378 6452
rect 2372 6412 3004 6440
rect 2372 6400 2378 6412
rect 2774 6372 2780 6384
rect 2735 6344 2780 6372
rect 2774 6332 2780 6344
rect 2832 6332 2838 6384
rect 2976 6372 3004 6412
rect 3050 6400 3056 6452
rect 3108 6440 3114 6452
rect 6457 6443 6515 6449
rect 6457 6440 6469 6443
rect 3108 6412 6469 6440
rect 3108 6400 3114 6412
rect 6457 6409 6469 6412
rect 6503 6409 6515 6443
rect 6457 6403 6515 6409
rect 8202 6400 8208 6452
rect 8260 6440 8266 6452
rect 10686 6440 10692 6452
rect 8260 6412 10692 6440
rect 8260 6400 8266 6412
rect 10686 6400 10692 6412
rect 10744 6400 10750 6452
rect 11514 6440 11520 6452
rect 11475 6412 11520 6440
rect 11514 6400 11520 6412
rect 11572 6400 11578 6452
rect 11974 6400 11980 6452
rect 12032 6440 12038 6452
rect 13446 6440 13452 6452
rect 12032 6412 13452 6440
rect 12032 6400 12038 6412
rect 13446 6400 13452 6412
rect 13504 6400 13510 6452
rect 13722 6400 13728 6452
rect 13780 6440 13786 6452
rect 13909 6443 13967 6449
rect 13909 6440 13921 6443
rect 13780 6412 13921 6440
rect 13780 6400 13786 6412
rect 13909 6409 13921 6412
rect 13955 6409 13967 6443
rect 13909 6403 13967 6409
rect 13998 6400 14004 6452
rect 14056 6440 14062 6452
rect 14056 6412 14320 6440
rect 14056 6400 14062 6412
rect 3142 6372 3148 6384
rect 2976 6344 3148 6372
rect 3142 6332 3148 6344
rect 3200 6332 3206 6384
rect 5350 6332 5356 6384
rect 5408 6372 5414 6384
rect 6733 6375 6791 6381
rect 6733 6372 6745 6375
rect 5408 6344 6745 6372
rect 5408 6332 5414 6344
rect 6733 6341 6745 6344
rect 6779 6372 6791 6375
rect 7742 6372 7748 6384
rect 6779 6344 7748 6372
rect 6779 6341 6791 6344
rect 6733 6335 6791 6341
rect 7742 6332 7748 6344
rect 7800 6332 7806 6384
rect 10502 6332 10508 6384
rect 10560 6332 10566 6384
rect 11054 6332 11060 6384
rect 11112 6372 11118 6384
rect 12345 6375 12403 6381
rect 12345 6372 12357 6375
rect 11112 6344 12357 6372
rect 11112 6332 11118 6344
rect 12345 6341 12357 6344
rect 12391 6341 12403 6375
rect 12345 6335 12403 6341
rect 12710 6332 12716 6384
rect 12768 6372 12774 6384
rect 14292 6372 14320 6412
rect 14550 6400 14556 6452
rect 14608 6440 14614 6452
rect 14829 6443 14887 6449
rect 14829 6440 14841 6443
rect 14608 6412 14841 6440
rect 14608 6400 14614 6412
rect 14829 6409 14841 6412
rect 14875 6409 14887 6443
rect 14829 6403 14887 6409
rect 16574 6400 16580 6452
rect 16632 6440 16638 6452
rect 17862 6440 17868 6452
rect 16632 6412 17868 6440
rect 16632 6400 16638 6412
rect 14918 6372 14924 6384
rect 12768 6344 14228 6372
rect 14292 6344 14924 6372
rect 12768 6332 12774 6344
rect 2225 6307 2283 6313
rect 2225 6273 2237 6307
rect 2271 6304 2283 6307
rect 2271 6276 2728 6304
rect 2271 6273 2283 6276
rect 2225 6267 2283 6273
rect 1486 6236 1492 6248
rect 1447 6208 1492 6236
rect 1486 6196 1492 6208
rect 1544 6196 1550 6248
rect 2409 6239 2467 6245
rect 2409 6205 2421 6239
rect 2455 6236 2467 6239
rect 2590 6236 2596 6248
rect 2455 6208 2596 6236
rect 2455 6205 2467 6208
rect 2409 6199 2467 6205
rect 2590 6196 2596 6208
rect 2648 6196 2654 6248
rect 2700 6168 2728 6276
rect 4172 6276 4476 6304
rect 3602 6196 3608 6248
rect 3660 6236 3666 6248
rect 4172 6236 4200 6276
rect 3660 6208 4200 6236
rect 4249 6239 4307 6245
rect 3660 6196 3666 6208
rect 4249 6205 4261 6239
rect 4295 6236 4307 6239
rect 4338 6236 4344 6248
rect 4295 6208 4344 6236
rect 4295 6205 4307 6208
rect 4249 6199 4307 6205
rect 4338 6196 4344 6208
rect 4396 6196 4402 6248
rect 4448 6236 4476 6276
rect 6546 6264 6552 6316
rect 6604 6304 6610 6316
rect 7469 6307 7527 6313
rect 7469 6304 7481 6307
rect 6604 6276 7481 6304
rect 6604 6264 6610 6276
rect 7469 6273 7481 6276
rect 7515 6273 7527 6307
rect 7469 6267 7527 6273
rect 8846 6264 8852 6316
rect 8904 6264 8910 6316
rect 9306 6264 9312 6316
rect 9364 6264 9370 6316
rect 9398 6264 9404 6316
rect 9456 6264 9462 6316
rect 10137 6307 10195 6313
rect 10137 6273 10149 6307
rect 10183 6304 10195 6307
rect 10226 6304 10232 6316
rect 10183 6276 10232 6304
rect 10183 6273 10195 6276
rect 10137 6267 10195 6273
rect 10226 6264 10232 6276
rect 10284 6264 10290 6316
rect 10520 6304 10548 6332
rect 14200 6316 14228 6344
rect 14918 6332 14924 6344
rect 14976 6332 14982 6384
rect 17034 6372 17040 6384
rect 15672 6344 17040 6372
rect 10686 6304 10692 6316
rect 10336 6276 10692 6304
rect 5813 6239 5871 6245
rect 5813 6236 5825 6239
rect 4448 6208 5825 6236
rect 5813 6205 5825 6208
rect 5859 6205 5871 6239
rect 5994 6236 6000 6248
rect 5955 6208 6000 6236
rect 5813 6199 5871 6205
rect 5994 6196 6000 6208
rect 6052 6196 6058 6248
rect 6454 6196 6460 6248
rect 6512 6236 6518 6248
rect 6641 6239 6699 6245
rect 6641 6236 6653 6239
rect 6512 6208 6653 6236
rect 6512 6196 6518 6208
rect 6641 6205 6653 6208
rect 6687 6205 6699 6239
rect 6641 6199 6699 6205
rect 7837 6239 7895 6245
rect 7837 6205 7849 6239
rect 7883 6236 7895 6239
rect 7926 6236 7932 6248
rect 7883 6208 7932 6236
rect 7883 6205 7895 6208
rect 7837 6199 7895 6205
rect 7926 6196 7932 6208
rect 7984 6236 7990 6248
rect 8864 6236 8892 6264
rect 9122 6236 9128 6248
rect 7984 6208 9128 6236
rect 7984 6196 7990 6208
rect 9122 6196 9128 6208
rect 9180 6196 9186 6248
rect 2700 6140 2912 6168
rect 2317 6103 2375 6109
rect 2317 6069 2329 6103
rect 2363 6100 2375 6103
rect 2590 6100 2596 6112
rect 2363 6072 2596 6100
rect 2363 6069 2375 6072
rect 2317 6063 2375 6069
rect 2590 6060 2596 6072
rect 2648 6060 2654 6112
rect 2884 6109 2912 6140
rect 2958 6128 2964 6180
rect 3016 6168 3022 6180
rect 3970 6168 3976 6180
rect 4028 6177 4034 6180
rect 3016 6140 3976 6168
rect 3016 6128 3022 6140
rect 3970 6128 3976 6140
rect 4028 6131 4040 6177
rect 4586 6171 4644 6177
rect 4586 6168 4598 6171
rect 4080 6140 4598 6168
rect 4028 6128 4034 6131
rect 2869 6103 2927 6109
rect 2869 6069 2881 6103
rect 2915 6100 2927 6103
rect 4080 6100 4108 6140
rect 4586 6137 4598 6140
rect 4632 6137 4644 6171
rect 4586 6131 4644 6137
rect 4724 6140 5856 6168
rect 2915 6072 4108 6100
rect 2915 6069 2927 6072
rect 2869 6063 2927 6069
rect 4154 6060 4160 6112
rect 4212 6100 4218 6112
rect 4724 6100 4752 6140
rect 4212 6072 4752 6100
rect 4212 6060 4218 6072
rect 5534 6060 5540 6112
rect 5592 6100 5598 6112
rect 5721 6103 5779 6109
rect 5721 6100 5733 6103
rect 5592 6072 5733 6100
rect 5592 6060 5598 6072
rect 5721 6069 5733 6072
rect 5767 6069 5779 6103
rect 5828 6100 5856 6140
rect 6086 6128 6092 6180
rect 6144 6168 6150 6180
rect 7285 6171 7343 6177
rect 6144 6140 6960 6168
rect 6144 6128 6150 6140
rect 6932 6109 6960 6140
rect 7285 6137 7297 6171
rect 7331 6168 7343 6171
rect 8104 6171 8162 6177
rect 7331 6140 8064 6168
rect 7331 6137 7343 6140
rect 7285 6131 7343 6137
rect 6181 6103 6239 6109
rect 6181 6100 6193 6103
rect 5828 6072 6193 6100
rect 5721 6063 5779 6069
rect 6181 6069 6193 6072
rect 6227 6069 6239 6103
rect 6181 6063 6239 6069
rect 6917 6103 6975 6109
rect 6917 6069 6929 6103
rect 6963 6069 6975 6103
rect 6917 6063 6975 6069
rect 7374 6060 7380 6112
rect 7432 6100 7438 6112
rect 8036 6100 8064 6140
rect 8104 6137 8116 6171
rect 8150 6168 8162 6171
rect 8846 6168 8852 6180
rect 8150 6140 8852 6168
rect 8150 6137 8162 6140
rect 8104 6131 8162 6137
rect 8846 6128 8852 6140
rect 8904 6168 8910 6180
rect 9324 6168 9352 6264
rect 9416 6236 9444 6264
rect 10336 6245 10364 6276
rect 10686 6264 10692 6276
rect 10744 6264 10750 6316
rect 10965 6307 11023 6313
rect 10965 6273 10977 6307
rect 11011 6304 11023 6307
rect 12158 6304 12164 6316
rect 11011 6276 12164 6304
rect 11011 6273 11023 6276
rect 10965 6267 11023 6273
rect 12158 6264 12164 6276
rect 12216 6264 12222 6316
rect 12618 6264 12624 6316
rect 12676 6304 12682 6316
rect 12897 6307 12955 6313
rect 12897 6304 12909 6307
rect 12676 6276 12909 6304
rect 12676 6264 12682 6276
rect 12897 6273 12909 6276
rect 12943 6273 12955 6307
rect 12897 6267 12955 6273
rect 13357 6307 13415 6313
rect 13357 6273 13369 6307
rect 13403 6304 13415 6307
rect 13998 6304 14004 6316
rect 13403 6276 14004 6304
rect 13403 6273 13415 6276
rect 13357 6267 13415 6273
rect 13998 6264 14004 6276
rect 14056 6304 14062 6316
rect 14093 6307 14151 6313
rect 14093 6304 14105 6307
rect 14056 6276 14105 6304
rect 14056 6264 14062 6276
rect 14093 6273 14105 6276
rect 14139 6273 14151 6307
rect 14093 6267 14151 6273
rect 14182 6264 14188 6316
rect 14240 6304 14246 6316
rect 15473 6307 15531 6313
rect 15473 6304 15485 6307
rect 14240 6276 15485 6304
rect 14240 6264 14246 6276
rect 15473 6273 15485 6276
rect 15519 6304 15531 6307
rect 15562 6304 15568 6316
rect 15519 6276 15568 6304
rect 15519 6273 15531 6276
rect 15473 6267 15531 6273
rect 15562 6264 15568 6276
rect 15620 6264 15626 6316
rect 9585 6239 9643 6245
rect 9585 6236 9597 6239
rect 9416 6208 9597 6236
rect 9585 6205 9597 6208
rect 9631 6205 9643 6239
rect 9585 6199 9643 6205
rect 10321 6239 10379 6245
rect 10321 6205 10333 6239
rect 10367 6205 10379 6239
rect 10321 6199 10379 6205
rect 10502 6196 10508 6248
rect 10560 6236 10566 6248
rect 12069 6239 12127 6245
rect 12069 6236 12081 6239
rect 10560 6208 12081 6236
rect 10560 6196 10566 6208
rect 12069 6205 12081 6208
rect 12115 6205 12127 6239
rect 12069 6199 12127 6205
rect 12710 6196 12716 6248
rect 12768 6236 12774 6248
rect 12805 6239 12863 6245
rect 12805 6236 12817 6239
rect 12768 6208 12817 6236
rect 12768 6196 12774 6208
rect 12805 6205 12817 6208
rect 12851 6205 12863 6239
rect 13449 6239 13507 6245
rect 12805 6199 12863 6205
rect 12912 6208 13400 6236
rect 8904 6140 9352 6168
rect 9861 6171 9919 6177
rect 8904 6128 8910 6140
rect 9861 6137 9873 6171
rect 9907 6168 9919 6171
rect 11514 6168 11520 6180
rect 9907 6140 11520 6168
rect 9907 6137 9919 6140
rect 9861 6131 9919 6137
rect 11514 6128 11520 6140
rect 11572 6128 11578 6180
rect 12912 6168 12940 6208
rect 12268 6140 12940 6168
rect 13372 6168 13400 6208
rect 13449 6205 13461 6239
rect 13495 6236 13507 6239
rect 13538 6236 13544 6248
rect 13495 6208 13544 6236
rect 13495 6205 13507 6208
rect 13449 6199 13507 6205
rect 13538 6196 13544 6208
rect 13596 6196 13602 6248
rect 13630 6196 13636 6248
rect 13688 6236 13694 6248
rect 14369 6239 14427 6245
rect 14369 6236 14381 6239
rect 13688 6208 14381 6236
rect 13688 6196 13694 6208
rect 14369 6205 14381 6208
rect 14415 6236 14427 6239
rect 15672 6236 15700 6344
rect 17034 6332 17040 6344
rect 17092 6332 17098 6384
rect 16206 6304 16212 6316
rect 16167 6276 16212 6304
rect 16206 6264 16212 6276
rect 16264 6264 16270 6316
rect 16850 6304 16856 6316
rect 16316 6276 16856 6304
rect 14415 6208 15700 6236
rect 16117 6239 16175 6245
rect 14415 6205 14427 6208
rect 14369 6199 14427 6205
rect 16117 6205 16129 6239
rect 16163 6236 16175 6239
rect 16316 6236 16344 6276
rect 16850 6264 16856 6276
rect 16908 6264 16914 6316
rect 16942 6264 16948 6316
rect 17000 6264 17006 6316
rect 17512 6313 17540 6412
rect 17862 6400 17868 6412
rect 17920 6400 17926 6452
rect 17497 6307 17555 6313
rect 17497 6273 17509 6307
rect 17543 6273 17555 6307
rect 17678 6304 17684 6316
rect 17639 6276 17684 6304
rect 17497 6267 17555 6273
rect 17678 6264 17684 6276
rect 17736 6264 17742 6316
rect 16574 6236 16580 6248
rect 16163 6208 16344 6236
rect 16535 6208 16580 6236
rect 16163 6205 16175 6208
rect 16117 6199 16175 6205
rect 16574 6196 16580 6208
rect 16632 6196 16638 6248
rect 16960 6236 16988 6264
rect 16684 6208 16988 6236
rect 13722 6168 13728 6180
rect 13372 6140 13728 6168
rect 8386 6100 8392 6112
rect 7432 6072 7477 6100
rect 8036 6072 8392 6100
rect 7432 6060 7438 6072
rect 8386 6060 8392 6072
rect 8444 6060 8450 6112
rect 9214 6100 9220 6112
rect 9175 6072 9220 6100
rect 9214 6060 9220 6072
rect 9272 6060 9278 6112
rect 9306 6060 9312 6112
rect 9364 6100 9370 6112
rect 9401 6103 9459 6109
rect 9401 6100 9413 6103
rect 9364 6072 9413 6100
rect 9364 6060 9370 6072
rect 9401 6069 9413 6072
rect 9447 6069 9459 6103
rect 9401 6063 9459 6069
rect 9674 6060 9680 6112
rect 9732 6100 9738 6112
rect 10229 6103 10287 6109
rect 10229 6100 10241 6103
rect 9732 6072 10241 6100
rect 9732 6060 9738 6072
rect 10229 6069 10241 6072
rect 10275 6069 10287 6103
rect 10686 6100 10692 6112
rect 10647 6072 10692 6100
rect 10229 6063 10287 6069
rect 10686 6060 10692 6072
rect 10744 6060 10750 6112
rect 10962 6060 10968 6112
rect 11020 6100 11026 6112
rect 11057 6103 11115 6109
rect 11057 6100 11069 6103
rect 11020 6072 11069 6100
rect 11020 6060 11026 6072
rect 11057 6069 11069 6072
rect 11103 6069 11115 6103
rect 11057 6063 11115 6069
rect 11149 6103 11207 6109
rect 11149 6069 11161 6103
rect 11195 6100 11207 6103
rect 11330 6100 11336 6112
rect 11195 6072 11336 6100
rect 11195 6069 11207 6072
rect 11149 6063 11207 6069
rect 11330 6060 11336 6072
rect 11388 6100 11394 6112
rect 11606 6100 11612 6112
rect 11388 6072 11612 6100
rect 11388 6060 11394 6072
rect 11606 6060 11612 6072
rect 11664 6060 11670 6112
rect 11790 6100 11796 6112
rect 11751 6072 11796 6100
rect 11790 6060 11796 6072
rect 11848 6060 11854 6112
rect 12268 6109 12296 6140
rect 13722 6128 13728 6140
rect 13780 6128 13786 6180
rect 15289 6171 15347 6177
rect 15289 6168 15301 6171
rect 14752 6140 15301 6168
rect 12253 6103 12311 6109
rect 12253 6069 12265 6103
rect 12299 6069 12311 6103
rect 12253 6063 12311 6069
rect 12526 6060 12532 6112
rect 12584 6100 12590 6112
rect 12713 6103 12771 6109
rect 12713 6100 12725 6103
rect 12584 6072 12725 6100
rect 12584 6060 12590 6072
rect 12713 6069 12725 6072
rect 12759 6069 12771 6103
rect 12713 6063 12771 6069
rect 13446 6060 13452 6112
rect 13504 6100 13510 6112
rect 13541 6103 13599 6109
rect 13541 6100 13553 6103
rect 13504 6072 13553 6100
rect 13504 6060 13510 6072
rect 13541 6069 13553 6072
rect 13587 6069 13599 6103
rect 13541 6063 13599 6069
rect 13814 6060 13820 6112
rect 13872 6100 13878 6112
rect 14182 6100 14188 6112
rect 13872 6072 14188 6100
rect 13872 6060 13878 6072
rect 14182 6060 14188 6072
rect 14240 6100 14246 6112
rect 14752 6109 14780 6140
rect 15289 6137 15301 6140
rect 15335 6137 15347 6171
rect 15289 6131 15347 6137
rect 16025 6171 16083 6177
rect 16025 6137 16037 6171
rect 16071 6168 16083 6171
rect 16684 6168 16712 6208
rect 17126 6196 17132 6248
rect 17184 6236 17190 6248
rect 18325 6239 18383 6245
rect 18325 6236 18337 6239
rect 17184 6208 18337 6236
rect 17184 6196 17190 6208
rect 18325 6205 18337 6208
rect 18371 6205 18383 6239
rect 18325 6199 18383 6205
rect 17957 6171 18015 6177
rect 17957 6168 17969 6171
rect 16071 6140 16712 6168
rect 16776 6140 17969 6168
rect 16071 6137 16083 6140
rect 16025 6131 16083 6137
rect 14277 6103 14335 6109
rect 14277 6100 14289 6103
rect 14240 6072 14289 6100
rect 14240 6060 14246 6072
rect 14277 6069 14289 6072
rect 14323 6069 14335 6103
rect 14277 6063 14335 6069
rect 14737 6103 14795 6109
rect 14737 6069 14749 6103
rect 14783 6069 14795 6103
rect 14737 6063 14795 6069
rect 15102 6060 15108 6112
rect 15160 6100 15166 6112
rect 15197 6103 15255 6109
rect 15197 6100 15209 6103
rect 15160 6072 15209 6100
rect 15160 6060 15166 6072
rect 15197 6069 15209 6072
rect 15243 6069 15255 6103
rect 15197 6063 15255 6069
rect 15378 6060 15384 6112
rect 15436 6100 15442 6112
rect 16776 6109 16804 6140
rect 17957 6137 17969 6140
rect 18003 6137 18015 6171
rect 18506 6168 18512 6180
rect 18467 6140 18512 6168
rect 17957 6131 18015 6137
rect 18506 6128 18512 6140
rect 18564 6128 18570 6180
rect 15657 6103 15715 6109
rect 15657 6100 15669 6103
rect 15436 6072 15669 6100
rect 15436 6060 15442 6072
rect 15657 6069 15669 6072
rect 15703 6069 15715 6103
rect 15657 6063 15715 6069
rect 16761 6103 16819 6109
rect 16761 6069 16773 6103
rect 16807 6069 16819 6103
rect 17034 6100 17040 6112
rect 16995 6072 17040 6100
rect 16761 6063 16819 6069
rect 17034 6060 17040 6072
rect 17092 6060 17098 6112
rect 17218 6060 17224 6112
rect 17276 6100 17282 6112
rect 17405 6103 17463 6109
rect 17405 6100 17417 6103
rect 17276 6072 17417 6100
rect 17276 6060 17282 6072
rect 17405 6069 17417 6072
rect 17451 6069 17463 6103
rect 17405 6063 17463 6069
rect 17862 6060 17868 6112
rect 17920 6100 17926 6112
rect 18049 6103 18107 6109
rect 18049 6100 18061 6103
rect 17920 6072 18061 6100
rect 17920 6060 17926 6072
rect 18049 6069 18061 6072
rect 18095 6069 18107 6103
rect 18049 6063 18107 6069
rect 1104 6010 18860 6032
rect 1104 5958 6912 6010
rect 6964 5958 6976 6010
rect 7028 5958 7040 6010
rect 7092 5958 7104 6010
rect 7156 5958 12843 6010
rect 12895 5958 12907 6010
rect 12959 5958 12971 6010
rect 13023 5958 13035 6010
rect 13087 5958 18860 6010
rect 1104 5936 18860 5958
rect 2317 5899 2375 5905
rect 2317 5865 2329 5899
rect 2363 5896 2375 5899
rect 2869 5899 2927 5905
rect 2869 5896 2881 5899
rect 2363 5868 2881 5896
rect 2363 5865 2375 5868
rect 2317 5859 2375 5865
rect 2869 5865 2881 5868
rect 2915 5865 2927 5899
rect 2869 5859 2927 5865
rect 3237 5899 3295 5905
rect 3237 5865 3249 5899
rect 3283 5896 3295 5899
rect 3786 5896 3792 5908
rect 3283 5868 3792 5896
rect 3283 5865 3295 5868
rect 3237 5859 3295 5865
rect 3786 5856 3792 5868
rect 3844 5896 3850 5908
rect 4430 5896 4436 5908
rect 3844 5868 4436 5896
rect 3844 5856 3850 5868
rect 4430 5856 4436 5868
rect 4488 5856 4494 5908
rect 5997 5899 6055 5905
rect 5997 5865 6009 5899
rect 6043 5896 6055 5899
rect 6086 5896 6092 5908
rect 6043 5868 6092 5896
rect 6043 5865 6055 5868
rect 5997 5859 6055 5865
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 6365 5899 6423 5905
rect 6365 5865 6377 5899
rect 6411 5865 6423 5899
rect 6546 5896 6552 5908
rect 6507 5868 6552 5896
rect 6365 5859 6423 5865
rect 1489 5831 1547 5837
rect 1489 5797 1501 5831
rect 1535 5828 1547 5831
rect 1535 5800 2544 5828
rect 1535 5797 1547 5800
rect 1489 5791 1547 5797
rect 1578 5720 1584 5772
rect 1636 5760 1642 5772
rect 2406 5760 2412 5772
rect 1636 5732 2412 5760
rect 1636 5720 1642 5732
rect 2406 5720 2412 5732
rect 2464 5720 2470 5772
rect 2516 5760 2544 5800
rect 2590 5788 2596 5840
rect 2648 5828 2654 5840
rect 3697 5831 3755 5837
rect 3697 5828 3709 5831
rect 2648 5800 3709 5828
rect 2648 5788 2654 5800
rect 3697 5797 3709 5800
rect 3743 5797 3755 5831
rect 3697 5791 3755 5797
rect 3970 5788 3976 5840
rect 4028 5828 4034 5840
rect 6380 5828 6408 5859
rect 6546 5856 6552 5868
rect 6604 5856 6610 5908
rect 7374 5856 7380 5908
rect 7432 5896 7438 5908
rect 8021 5899 8079 5905
rect 8021 5896 8033 5899
rect 7432 5868 8033 5896
rect 7432 5856 7438 5868
rect 8021 5865 8033 5868
rect 8067 5865 8079 5899
rect 8021 5859 8079 5865
rect 8202 5856 8208 5908
rect 8260 5896 8266 5908
rect 8849 5899 8907 5905
rect 8849 5896 8861 5899
rect 8260 5868 8861 5896
rect 8260 5856 8266 5868
rect 8849 5865 8861 5868
rect 8895 5865 8907 5899
rect 8849 5859 8907 5865
rect 8938 5856 8944 5908
rect 8996 5896 9002 5908
rect 10965 5899 11023 5905
rect 10965 5896 10977 5899
rect 8996 5868 10977 5896
rect 8996 5856 9002 5868
rect 10965 5865 10977 5868
rect 11011 5896 11023 5899
rect 11011 5868 11100 5896
rect 11011 5865 11023 5868
rect 10965 5859 11023 5865
rect 11072 5828 11100 5868
rect 11146 5856 11152 5908
rect 11204 5896 11210 5908
rect 11425 5899 11483 5905
rect 11425 5896 11437 5899
rect 11204 5868 11437 5896
rect 11204 5856 11210 5868
rect 11425 5865 11437 5868
rect 11471 5865 11483 5899
rect 11790 5896 11796 5908
rect 11751 5868 11796 5896
rect 11425 5859 11483 5865
rect 11790 5856 11796 5868
rect 11848 5856 11854 5908
rect 12342 5856 12348 5908
rect 12400 5896 12406 5908
rect 14090 5896 14096 5908
rect 12400 5868 13768 5896
rect 14051 5868 14096 5896
rect 12400 5856 12406 5868
rect 13630 5828 13636 5840
rect 4028 5800 4476 5828
rect 6380 5800 11008 5828
rect 11072 5800 13636 5828
rect 4028 5788 4034 5800
rect 2866 5760 2872 5772
rect 2516 5732 2872 5760
rect 2866 5720 2872 5732
rect 2924 5760 2930 5772
rect 4062 5760 4068 5772
rect 2924 5732 4068 5760
rect 2924 5720 2930 5732
rect 4062 5720 4068 5732
rect 4120 5720 4126 5772
rect 4249 5763 4307 5769
rect 4249 5760 4261 5763
rect 4172 5732 4261 5760
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5692 2283 5695
rect 3234 5692 3240 5704
rect 2271 5664 3240 5692
rect 2271 5661 2283 5664
rect 2225 5655 2283 5661
rect 3234 5652 3240 5664
rect 3292 5652 3298 5704
rect 3329 5695 3387 5701
rect 3329 5661 3341 5695
rect 3375 5661 3387 5695
rect 3510 5692 3516 5704
rect 3471 5664 3516 5692
rect 3329 5655 3387 5661
rect 1765 5627 1823 5633
rect 1765 5593 1777 5627
rect 1811 5624 1823 5627
rect 2682 5624 2688 5636
rect 1811 5596 2688 5624
rect 1811 5593 1823 5596
rect 1765 5587 1823 5593
rect 2682 5584 2688 5596
rect 2740 5584 2746 5636
rect 2958 5584 2964 5636
rect 3016 5624 3022 5636
rect 3344 5624 3372 5655
rect 3510 5652 3516 5664
rect 3568 5652 3574 5704
rect 3016 5596 3372 5624
rect 3016 5584 3022 5596
rect 3418 5584 3424 5636
rect 3476 5624 3482 5636
rect 4172 5624 4200 5732
rect 4249 5729 4261 5732
rect 4295 5729 4307 5763
rect 4249 5723 4307 5729
rect 4338 5692 4344 5704
rect 4299 5664 4344 5692
rect 4338 5652 4344 5664
rect 4396 5652 4402 5704
rect 4448 5701 4476 5800
rect 5169 5763 5227 5769
rect 5169 5729 5181 5763
rect 5215 5760 5227 5763
rect 6178 5760 6184 5772
rect 5215 5732 6184 5760
rect 5215 5729 5227 5732
rect 5169 5723 5227 5729
rect 6178 5720 6184 5732
rect 6236 5760 6242 5772
rect 6638 5760 6644 5772
rect 6236 5732 6644 5760
rect 6236 5720 6242 5732
rect 6638 5720 6644 5732
rect 6696 5720 6702 5772
rect 7650 5720 7656 5772
rect 7708 5769 7714 5772
rect 7708 5760 7720 5769
rect 7708 5732 7753 5760
rect 7708 5723 7720 5732
rect 7708 5720 7714 5723
rect 8294 5720 8300 5772
rect 8352 5760 8358 5772
rect 8389 5763 8447 5769
rect 8389 5760 8401 5763
rect 8352 5732 8401 5760
rect 8352 5720 8358 5732
rect 8389 5729 8401 5732
rect 8435 5729 8447 5763
rect 8389 5723 8447 5729
rect 8478 5720 8484 5772
rect 8536 5760 8542 5772
rect 8754 5760 8760 5772
rect 8536 5732 8760 5760
rect 8536 5720 8542 5732
rect 8754 5720 8760 5732
rect 8812 5720 8818 5772
rect 9214 5760 9220 5772
rect 9048 5732 9220 5760
rect 4433 5695 4491 5701
rect 4433 5661 4445 5695
rect 4479 5661 4491 5695
rect 5261 5695 5319 5701
rect 5261 5692 5273 5695
rect 4433 5655 4491 5661
rect 4540 5664 5273 5692
rect 3476 5596 4200 5624
rect 3476 5584 3482 5596
rect 4246 5584 4252 5636
rect 4304 5624 4310 5636
rect 4540 5624 4568 5664
rect 5261 5661 5273 5664
rect 5307 5692 5319 5695
rect 5350 5692 5356 5704
rect 5307 5664 5356 5692
rect 5307 5661 5319 5664
rect 5261 5655 5319 5661
rect 5350 5652 5356 5664
rect 5408 5652 5414 5704
rect 5445 5695 5503 5701
rect 5445 5661 5457 5695
rect 5491 5692 5503 5695
rect 5534 5692 5540 5704
rect 5491 5664 5540 5692
rect 5491 5661 5503 5664
rect 5445 5655 5503 5661
rect 5534 5652 5540 5664
rect 5592 5652 5598 5704
rect 5626 5652 5632 5704
rect 5684 5692 5690 5704
rect 5721 5695 5779 5701
rect 5721 5692 5733 5695
rect 5684 5664 5733 5692
rect 5684 5652 5690 5664
rect 5721 5661 5733 5664
rect 5767 5661 5779 5695
rect 5902 5692 5908 5704
rect 5863 5664 5908 5692
rect 5721 5655 5779 5661
rect 5902 5652 5908 5664
rect 5960 5652 5966 5704
rect 7926 5692 7932 5704
rect 7839 5664 7932 5692
rect 7926 5652 7932 5664
rect 7984 5652 7990 5704
rect 8202 5652 8208 5704
rect 8260 5692 8266 5704
rect 8570 5692 8576 5704
rect 8260 5664 8576 5692
rect 8260 5652 8266 5664
rect 8570 5652 8576 5664
rect 8628 5652 8634 5704
rect 4304 5596 4568 5624
rect 4304 5584 4310 5596
rect 2777 5559 2835 5565
rect 2777 5525 2789 5559
rect 2823 5556 2835 5559
rect 2866 5556 2872 5568
rect 2823 5528 2872 5556
rect 2823 5525 2835 5528
rect 2777 5519 2835 5525
rect 2866 5516 2872 5528
rect 2924 5516 2930 5568
rect 3697 5559 3755 5565
rect 3697 5525 3709 5559
rect 3743 5556 3755 5559
rect 3881 5559 3939 5565
rect 3881 5556 3893 5559
rect 3743 5528 3893 5556
rect 3743 5525 3755 5528
rect 3697 5519 3755 5525
rect 3881 5525 3893 5528
rect 3927 5525 3939 5559
rect 4798 5556 4804 5568
rect 4759 5528 4804 5556
rect 3881 5519 3939 5525
rect 4798 5516 4804 5528
rect 4856 5516 4862 5568
rect 6086 5516 6092 5568
rect 6144 5556 6150 5568
rect 6730 5556 6736 5568
rect 6144 5528 6736 5556
rect 6144 5516 6150 5528
rect 6730 5516 6736 5528
rect 6788 5556 6794 5568
rect 7944 5556 7972 5652
rect 8294 5584 8300 5636
rect 8352 5624 8358 5636
rect 9048 5624 9076 5732
rect 9214 5720 9220 5732
rect 9272 5760 9278 5772
rect 9381 5763 9439 5769
rect 9381 5760 9393 5763
rect 9272 5732 9393 5760
rect 9272 5720 9278 5732
rect 9381 5729 9393 5732
rect 9427 5729 9439 5763
rect 9381 5723 9439 5729
rect 10778 5720 10784 5772
rect 10836 5760 10842 5772
rect 10873 5763 10931 5769
rect 10873 5760 10885 5763
rect 10836 5732 10885 5760
rect 10836 5720 10842 5732
rect 10873 5729 10885 5732
rect 10919 5729 10931 5763
rect 10873 5723 10931 5729
rect 9122 5652 9128 5704
rect 9180 5692 9186 5704
rect 9180 5664 9225 5692
rect 9180 5652 9186 5664
rect 10226 5652 10232 5704
rect 10284 5692 10290 5704
rect 10689 5695 10747 5701
rect 10689 5692 10701 5695
rect 10284 5664 10701 5692
rect 10284 5652 10290 5664
rect 10689 5661 10701 5664
rect 10735 5661 10747 5695
rect 10980 5692 11008 5800
rect 13630 5788 13636 5800
rect 13688 5788 13694 5840
rect 13740 5828 13768 5868
rect 14090 5856 14096 5868
rect 14148 5856 14154 5908
rect 14734 5896 14740 5908
rect 14695 5868 14740 5896
rect 14734 5856 14740 5868
rect 14792 5856 14798 5908
rect 15102 5896 15108 5908
rect 15063 5868 15108 5896
rect 15102 5856 15108 5868
rect 15160 5856 15166 5908
rect 15933 5899 15991 5905
rect 15933 5865 15945 5899
rect 15979 5896 15991 5899
rect 17034 5896 17040 5908
rect 15979 5868 17040 5896
rect 15979 5865 15991 5868
rect 15933 5859 15991 5865
rect 17034 5856 17040 5868
rect 17092 5856 17098 5908
rect 18138 5896 18144 5908
rect 18099 5868 18144 5896
rect 18138 5856 18144 5868
rect 18196 5856 18202 5908
rect 13740 5800 14136 5828
rect 14108 5772 14136 5800
rect 14366 5788 14372 5840
rect 14424 5828 14430 5840
rect 15010 5828 15016 5840
rect 14424 5800 15016 5828
rect 14424 5788 14430 5800
rect 15010 5788 15016 5800
rect 15068 5828 15074 5840
rect 15654 5828 15660 5840
rect 15068 5800 15660 5828
rect 15068 5788 15074 5800
rect 15654 5788 15660 5800
rect 15712 5828 15718 5840
rect 16752 5831 16810 5837
rect 15712 5800 16528 5828
rect 15712 5788 15718 5800
rect 11698 5720 11704 5772
rect 11756 5760 11762 5772
rect 12509 5763 12567 5769
rect 12509 5760 12521 5763
rect 11756 5732 12521 5760
rect 11756 5720 11762 5732
rect 12509 5729 12521 5732
rect 12555 5729 12567 5763
rect 12509 5723 12567 5729
rect 13262 5720 13268 5772
rect 13320 5760 13326 5772
rect 13725 5763 13783 5769
rect 13725 5760 13737 5763
rect 13320 5732 13737 5760
rect 13320 5720 13326 5732
rect 13725 5729 13737 5732
rect 13771 5729 13783 5763
rect 13725 5723 13783 5729
rect 14090 5720 14096 5772
rect 14148 5760 14154 5772
rect 14645 5763 14703 5769
rect 14645 5760 14657 5763
rect 14148 5732 14657 5760
rect 14148 5720 14154 5732
rect 14645 5729 14657 5732
rect 14691 5729 14703 5763
rect 14645 5723 14703 5729
rect 14918 5720 14924 5772
rect 14976 5760 14982 5772
rect 15102 5760 15108 5772
rect 14976 5732 15108 5760
rect 14976 5720 14982 5732
rect 15102 5720 15108 5732
rect 15160 5760 15166 5772
rect 16025 5763 16083 5769
rect 16025 5760 16037 5763
rect 15160 5732 16037 5760
rect 15160 5720 15166 5732
rect 16025 5729 16037 5732
rect 16071 5729 16083 5763
rect 16025 5723 16083 5729
rect 16114 5720 16120 5772
rect 16172 5760 16178 5772
rect 16390 5760 16396 5772
rect 16172 5732 16396 5760
rect 16172 5720 16178 5732
rect 16390 5720 16396 5732
rect 16448 5720 16454 5772
rect 16500 5704 16528 5800
rect 16752 5797 16764 5831
rect 16798 5828 16810 5831
rect 17678 5828 17684 5840
rect 16798 5800 17684 5828
rect 16798 5797 16810 5800
rect 16752 5791 16810 5797
rect 17678 5788 17684 5800
rect 17736 5788 17742 5840
rect 18506 5828 18512 5840
rect 18467 5800 18512 5828
rect 18506 5788 18512 5800
rect 18564 5788 18570 5840
rect 17034 5720 17040 5772
rect 17092 5760 17098 5772
rect 18325 5763 18383 5769
rect 18325 5760 18337 5763
rect 17092 5732 18337 5760
rect 17092 5720 17098 5732
rect 18325 5729 18337 5732
rect 18371 5729 18383 5763
rect 18325 5723 18383 5729
rect 11238 5692 11244 5704
rect 10980 5664 11244 5692
rect 10689 5655 10747 5661
rect 11238 5652 11244 5664
rect 11296 5652 11302 5704
rect 11885 5695 11943 5701
rect 11885 5661 11897 5695
rect 11931 5692 11943 5695
rect 11974 5692 11980 5704
rect 11931 5664 11980 5692
rect 11931 5661 11943 5664
rect 11885 5655 11943 5661
rect 11974 5652 11980 5664
rect 12032 5652 12038 5704
rect 12069 5695 12127 5701
rect 12069 5661 12081 5695
rect 12115 5692 12127 5695
rect 12158 5692 12164 5704
rect 12115 5664 12164 5692
rect 12115 5661 12127 5664
rect 12069 5655 12127 5661
rect 12158 5652 12164 5664
rect 12216 5652 12222 5704
rect 12253 5695 12311 5701
rect 12253 5661 12265 5695
rect 12299 5661 12311 5695
rect 13998 5692 14004 5704
rect 12253 5655 12311 5661
rect 13648 5664 14004 5692
rect 8352 5596 9076 5624
rect 8352 5584 8358 5596
rect 6788 5528 7972 5556
rect 6788 5516 6794 5528
rect 8754 5516 8760 5568
rect 8812 5556 8818 5568
rect 10318 5556 10324 5568
rect 8812 5528 10324 5556
rect 8812 5516 8818 5528
rect 10318 5516 10324 5528
rect 10376 5516 10382 5568
rect 10505 5559 10563 5565
rect 10505 5525 10517 5559
rect 10551 5556 10563 5559
rect 10778 5556 10784 5568
rect 10551 5528 10784 5556
rect 10551 5525 10563 5528
rect 10505 5519 10563 5525
rect 10778 5516 10784 5528
rect 10836 5516 10842 5568
rect 11330 5556 11336 5568
rect 11291 5528 11336 5556
rect 11330 5516 11336 5528
rect 11388 5516 11394 5568
rect 11422 5516 11428 5568
rect 11480 5556 11486 5568
rect 11790 5556 11796 5568
rect 11480 5528 11796 5556
rect 11480 5516 11486 5528
rect 11790 5516 11796 5528
rect 11848 5556 11854 5568
rect 12268 5556 12296 5655
rect 13648 5633 13676 5664
rect 13998 5652 14004 5664
rect 14056 5692 14062 5704
rect 14461 5695 14519 5701
rect 14461 5692 14473 5695
rect 14056 5664 14473 5692
rect 14056 5652 14062 5664
rect 14461 5661 14473 5664
rect 14507 5661 14519 5695
rect 15562 5692 15568 5704
rect 15523 5664 15568 5692
rect 14461 5655 14519 5661
rect 15562 5652 15568 5664
rect 15620 5652 15626 5704
rect 15841 5695 15899 5701
rect 15841 5661 15853 5695
rect 15887 5661 15899 5695
rect 16482 5692 16488 5704
rect 16443 5664 16488 5692
rect 15841 5655 15899 5661
rect 13633 5627 13691 5633
rect 13633 5593 13645 5627
rect 13679 5593 13691 5627
rect 13633 5587 13691 5593
rect 13814 5584 13820 5636
rect 13872 5624 13878 5636
rect 13909 5627 13967 5633
rect 13909 5624 13921 5627
rect 13872 5596 13921 5624
rect 13872 5584 13878 5596
rect 13909 5593 13921 5596
rect 13955 5624 13967 5627
rect 14918 5624 14924 5636
rect 13955 5596 14924 5624
rect 13955 5593 13967 5596
rect 13909 5587 13967 5593
rect 14918 5584 14924 5596
rect 14976 5584 14982 5636
rect 15856 5624 15884 5655
rect 16482 5652 16488 5664
rect 16540 5652 16546 5704
rect 16206 5624 16212 5636
rect 15856 5596 16212 5624
rect 16206 5584 16212 5596
rect 16264 5624 16270 5636
rect 16264 5596 16528 5624
rect 16264 5584 16270 5596
rect 13170 5556 13176 5568
rect 11848 5528 13176 5556
rect 11848 5516 11854 5528
rect 13170 5516 13176 5528
rect 13228 5516 13234 5568
rect 13998 5516 14004 5568
rect 14056 5556 14062 5568
rect 14182 5556 14188 5568
rect 14056 5528 14188 5556
rect 14056 5516 14062 5528
rect 14182 5516 14188 5528
rect 14240 5516 14246 5568
rect 15194 5556 15200 5568
rect 15155 5528 15200 5556
rect 15194 5516 15200 5528
rect 15252 5516 15258 5568
rect 16390 5556 16396 5568
rect 16351 5528 16396 5556
rect 16390 5516 16396 5528
rect 16448 5516 16454 5568
rect 16500 5556 16528 5596
rect 17770 5556 17776 5568
rect 16500 5528 17776 5556
rect 17770 5516 17776 5528
rect 17828 5556 17834 5568
rect 17865 5559 17923 5565
rect 17865 5556 17877 5559
rect 17828 5528 17877 5556
rect 17828 5516 17834 5528
rect 17865 5525 17877 5528
rect 17911 5525 17923 5559
rect 17865 5519 17923 5525
rect 1104 5466 18860 5488
rect 1104 5414 3947 5466
rect 3999 5414 4011 5466
rect 4063 5414 4075 5466
rect 4127 5414 4139 5466
rect 4191 5414 9878 5466
rect 9930 5414 9942 5466
rect 9994 5414 10006 5466
rect 10058 5414 10070 5466
rect 10122 5414 15808 5466
rect 15860 5414 15872 5466
rect 15924 5414 15936 5466
rect 15988 5414 16000 5466
rect 16052 5414 18860 5466
rect 1104 5392 18860 5414
rect 1486 5352 1492 5364
rect 1447 5324 1492 5352
rect 1486 5312 1492 5324
rect 1544 5312 1550 5364
rect 2317 5355 2375 5361
rect 2317 5321 2329 5355
rect 2363 5352 2375 5355
rect 4338 5352 4344 5364
rect 2363 5324 4344 5352
rect 2363 5321 2375 5324
rect 2317 5315 2375 5321
rect 4338 5312 4344 5324
rect 4396 5312 4402 5364
rect 7558 5352 7564 5364
rect 5000 5324 7564 5352
rect 3602 5244 3608 5296
rect 3660 5284 3666 5296
rect 5000 5284 5028 5324
rect 7558 5312 7564 5324
rect 7616 5312 7622 5364
rect 8386 5352 8392 5364
rect 8347 5324 8392 5352
rect 8386 5312 8392 5324
rect 8444 5312 8450 5364
rect 11698 5352 11704 5364
rect 11659 5324 11704 5352
rect 11698 5312 11704 5324
rect 11756 5312 11762 5364
rect 13170 5352 13176 5364
rect 13131 5324 13176 5352
rect 13170 5312 13176 5324
rect 13228 5312 13234 5364
rect 15010 5352 15016 5364
rect 13832 5324 15016 5352
rect 5994 5284 6000 5296
rect 3660 5256 5028 5284
rect 5955 5256 6000 5284
rect 3660 5244 3666 5256
rect 5994 5244 6000 5256
rect 6052 5244 6058 5296
rect 6454 5244 6460 5296
rect 6512 5284 6518 5296
rect 6512 5256 8248 5284
rect 6512 5244 6518 5256
rect 1765 5219 1823 5225
rect 1765 5185 1777 5219
rect 1811 5216 1823 5219
rect 7377 5219 7435 5225
rect 1811 5188 2544 5216
rect 1811 5185 1823 5188
rect 1765 5179 1823 5185
rect 2130 5108 2136 5160
rect 2188 5148 2194 5160
rect 2409 5151 2467 5157
rect 2409 5148 2421 5151
rect 2188 5120 2421 5148
rect 2188 5108 2194 5120
rect 2409 5117 2421 5120
rect 2455 5117 2467 5151
rect 2516 5148 2544 5188
rect 7377 5185 7389 5219
rect 7423 5216 7435 5219
rect 7650 5216 7656 5228
rect 7423 5188 7656 5216
rect 7423 5185 7435 5188
rect 7377 5179 7435 5185
rect 7650 5176 7656 5188
rect 7708 5216 7714 5228
rect 8110 5216 8116 5228
rect 7708 5188 8116 5216
rect 7708 5176 7714 5188
rect 8110 5176 8116 5188
rect 8168 5176 8174 5228
rect 3234 5148 3240 5160
rect 2516 5120 3240 5148
rect 2409 5111 2467 5117
rect 3234 5108 3240 5120
rect 3292 5108 3298 5160
rect 3878 5148 3884 5160
rect 3839 5120 3884 5148
rect 3878 5108 3884 5120
rect 3936 5108 3942 5160
rect 4433 5151 4491 5157
rect 4433 5117 4445 5151
rect 4479 5148 4491 5151
rect 4522 5148 4528 5160
rect 4479 5120 4528 5148
rect 4479 5117 4491 5120
rect 4433 5111 4491 5117
rect 4522 5108 4528 5120
rect 4580 5108 4586 5160
rect 5905 5151 5963 5157
rect 5905 5117 5917 5151
rect 5951 5148 5963 5151
rect 6086 5148 6092 5160
rect 5951 5120 6092 5148
rect 5951 5117 5963 5120
rect 5905 5111 5963 5117
rect 6086 5108 6092 5120
rect 6144 5108 6150 5160
rect 6181 5151 6239 5157
rect 6181 5117 6193 5151
rect 6227 5148 6239 5151
rect 6454 5148 6460 5160
rect 6227 5120 6460 5148
rect 6227 5117 6239 5120
rect 6181 5111 6239 5117
rect 6454 5108 6460 5120
rect 6512 5108 6518 5160
rect 6641 5151 6699 5157
rect 6641 5117 6653 5151
rect 6687 5117 6699 5151
rect 7098 5148 7104 5160
rect 7059 5120 7104 5148
rect 6641 5111 6699 5117
rect 2676 5083 2734 5089
rect 2676 5080 2688 5083
rect 2595 5052 2688 5080
rect 2676 5049 2688 5052
rect 2722 5080 2734 5083
rect 3510 5080 3516 5092
rect 2722 5052 3516 5080
rect 2722 5049 2734 5052
rect 2676 5043 2734 5049
rect 1762 4972 1768 5024
rect 1820 5012 1826 5024
rect 1857 5015 1915 5021
rect 1857 5012 1869 5015
rect 1820 4984 1869 5012
rect 1820 4972 1826 4984
rect 1857 4981 1869 4984
rect 1903 4981 1915 5015
rect 1857 4975 1915 4981
rect 1946 4972 1952 5024
rect 2004 5012 2010 5024
rect 2004 4984 2049 5012
rect 2004 4972 2010 4984
rect 2314 4972 2320 5024
rect 2372 5012 2378 5024
rect 2700 5012 2728 5043
rect 3510 5040 3516 5052
rect 3568 5040 3574 5092
rect 3694 5040 3700 5092
rect 3752 5080 3758 5092
rect 4065 5083 4123 5089
rect 4065 5080 4077 5083
rect 3752 5052 4077 5080
rect 3752 5040 3758 5052
rect 4065 5049 4077 5052
rect 4111 5049 4123 5083
rect 4065 5043 4123 5049
rect 4154 5040 4160 5092
rect 4212 5080 4218 5092
rect 4212 5052 5212 5080
rect 4212 5040 4218 5052
rect 2372 4984 2728 5012
rect 2372 4972 2378 4984
rect 3234 4972 3240 5024
rect 3292 5012 3298 5024
rect 3789 5015 3847 5021
rect 3789 5012 3801 5015
rect 3292 4984 3801 5012
rect 3292 4972 3298 4984
rect 3789 4981 3801 4984
rect 3835 4981 3847 5015
rect 4246 5012 4252 5024
rect 4207 4984 4252 5012
rect 3789 4975 3847 4981
rect 4246 4972 4252 4984
rect 4304 4972 4310 5024
rect 4525 5015 4583 5021
rect 4525 4981 4537 5015
rect 4571 5012 4583 5015
rect 5074 5012 5080 5024
rect 4571 4984 5080 5012
rect 4571 4981 4583 4984
rect 4525 4975 4583 4981
rect 5074 4972 5080 4984
rect 5132 4972 5138 5024
rect 5184 5012 5212 5052
rect 5534 5040 5540 5092
rect 5592 5080 5598 5092
rect 5638 5083 5696 5089
rect 5638 5080 5650 5083
rect 5592 5052 5650 5080
rect 5592 5040 5598 5052
rect 5638 5049 5650 5052
rect 5684 5049 5696 5083
rect 6656 5080 6684 5111
rect 7098 5108 7104 5120
rect 7156 5108 7162 5160
rect 7282 5108 7288 5160
rect 7340 5148 7346 5160
rect 7929 5151 7987 5157
rect 7929 5148 7941 5151
rect 7340 5120 7941 5148
rect 7340 5108 7346 5120
rect 7929 5117 7941 5120
rect 7975 5148 7987 5151
rect 8018 5148 8024 5160
rect 7975 5120 8024 5148
rect 7975 5117 7987 5120
rect 7929 5111 7987 5117
rect 8018 5108 8024 5120
rect 8076 5108 8082 5160
rect 8220 5148 8248 5256
rect 8754 5244 8760 5296
rect 8812 5284 8818 5296
rect 9217 5287 9275 5293
rect 9217 5284 9229 5287
rect 8812 5256 9229 5284
rect 8812 5244 8818 5256
rect 9217 5253 9229 5256
rect 9263 5253 9275 5287
rect 9217 5247 9275 5253
rect 9674 5244 9680 5296
rect 9732 5244 9738 5296
rect 8570 5176 8576 5228
rect 8628 5216 8634 5228
rect 8941 5219 8999 5225
rect 8941 5216 8953 5219
rect 8628 5188 8953 5216
rect 8628 5176 8634 5188
rect 8941 5185 8953 5188
rect 8987 5185 8999 5219
rect 8941 5179 8999 5185
rect 9122 5176 9128 5228
rect 9180 5216 9186 5228
rect 9692 5216 9720 5244
rect 10134 5216 10140 5228
rect 9180 5188 10140 5216
rect 9180 5176 9186 5188
rect 10134 5176 10140 5188
rect 10192 5176 10198 5228
rect 11146 5216 11152 5228
rect 11059 5188 11152 5216
rect 11146 5176 11152 5188
rect 11204 5216 11210 5228
rect 11790 5216 11796 5228
rect 11204 5188 11796 5216
rect 11204 5176 11210 5188
rect 11790 5176 11796 5188
rect 11848 5176 11854 5228
rect 13081 5219 13139 5225
rect 13081 5185 13093 5219
rect 13127 5216 13139 5219
rect 13832 5216 13860 5324
rect 15010 5312 15016 5324
rect 15068 5352 15074 5364
rect 15105 5355 15163 5361
rect 15105 5352 15117 5355
rect 15068 5324 15117 5352
rect 15068 5312 15074 5324
rect 15105 5321 15117 5324
rect 15151 5321 15163 5355
rect 15105 5315 15163 5321
rect 16485 5355 16543 5361
rect 16485 5321 16497 5355
rect 16531 5352 16543 5355
rect 17034 5352 17040 5364
rect 16531 5324 17040 5352
rect 16531 5321 16543 5324
rect 16485 5315 16543 5321
rect 17034 5312 17040 5324
rect 17092 5312 17098 5364
rect 15381 5287 15439 5293
rect 15381 5253 15393 5287
rect 15427 5284 15439 5287
rect 17402 5284 17408 5296
rect 15427 5256 17408 5284
rect 15427 5253 15439 5256
rect 15381 5247 15439 5253
rect 17402 5244 17408 5256
rect 17460 5244 17466 5296
rect 17678 5244 17684 5296
rect 17736 5284 17742 5296
rect 17736 5256 17816 5284
rect 17736 5244 17742 5256
rect 13127 5188 13860 5216
rect 14829 5219 14887 5225
rect 13127 5185 13139 5188
rect 13081 5179 13139 5185
rect 14829 5185 14841 5219
rect 14875 5216 14887 5219
rect 15010 5216 15016 5228
rect 14875 5188 15016 5216
rect 14875 5185 14887 5188
rect 14829 5179 14887 5185
rect 15010 5176 15016 5188
rect 15068 5176 15074 5228
rect 16117 5219 16175 5225
rect 16117 5185 16129 5219
rect 16163 5216 16175 5219
rect 16206 5216 16212 5228
rect 16163 5188 16212 5216
rect 16163 5185 16175 5188
rect 16117 5179 16175 5185
rect 16206 5176 16212 5188
rect 16264 5176 16270 5228
rect 16666 5216 16672 5228
rect 16592 5188 16672 5216
rect 8849 5151 8907 5157
rect 8849 5148 8861 5151
rect 8220 5120 8861 5148
rect 8849 5117 8861 5120
rect 8895 5117 8907 5151
rect 8849 5111 8907 5117
rect 9401 5151 9459 5157
rect 9401 5117 9413 5151
rect 9447 5148 9459 5151
rect 9490 5148 9496 5160
rect 9447 5120 9496 5148
rect 9447 5117 9459 5120
rect 9401 5111 9459 5117
rect 7742 5080 7748 5092
rect 6656 5052 7748 5080
rect 5638 5043 5696 5049
rect 7742 5040 7748 5052
rect 7800 5040 7806 5092
rect 8110 5040 8116 5092
rect 8168 5080 8174 5092
rect 8757 5083 8815 5089
rect 8757 5080 8769 5083
rect 8168 5052 8769 5080
rect 8168 5040 8174 5052
rect 8757 5049 8769 5052
rect 8803 5049 8815 5083
rect 8864 5080 8892 5111
rect 9490 5108 9496 5120
rect 9548 5108 9554 5160
rect 9582 5108 9588 5160
rect 9640 5148 9646 5160
rect 9677 5151 9735 5157
rect 9677 5148 9689 5151
rect 9640 5120 9689 5148
rect 9640 5108 9646 5120
rect 9677 5117 9689 5120
rect 9723 5117 9735 5151
rect 9677 5111 9735 5117
rect 10612 5120 11192 5148
rect 10612 5080 10640 5120
rect 8864 5052 10640 5080
rect 8757 5043 8815 5049
rect 10778 5040 10784 5092
rect 10836 5080 10842 5092
rect 10882 5083 10940 5089
rect 10882 5080 10894 5083
rect 10836 5052 10894 5080
rect 10836 5040 10842 5052
rect 10882 5049 10894 5052
rect 10928 5049 10940 5083
rect 11164 5080 11192 5120
rect 11238 5108 11244 5160
rect 11296 5148 11302 5160
rect 11425 5151 11483 5157
rect 11425 5148 11437 5151
rect 11296 5120 11437 5148
rect 11296 5108 11302 5120
rect 11425 5117 11437 5120
rect 11471 5117 11483 5151
rect 11425 5111 11483 5117
rect 11974 5108 11980 5160
rect 12032 5148 12038 5160
rect 13357 5151 13415 5157
rect 12032 5120 13032 5148
rect 12032 5108 12038 5120
rect 11790 5080 11796 5092
rect 11164 5052 11796 5080
rect 10882 5043 10940 5049
rect 11790 5040 11796 5052
rect 11848 5040 11854 5092
rect 12618 5040 12624 5092
rect 12676 5080 12682 5092
rect 12814 5083 12872 5089
rect 12814 5080 12826 5083
rect 12676 5052 12826 5080
rect 12676 5040 12682 5052
rect 12814 5049 12826 5052
rect 12860 5049 12872 5083
rect 13004 5080 13032 5120
rect 13357 5117 13369 5151
rect 13403 5148 13415 5151
rect 13814 5148 13820 5160
rect 13403 5120 13820 5148
rect 13403 5117 13415 5120
rect 13357 5111 13415 5117
rect 13814 5108 13820 5120
rect 13872 5108 13878 5160
rect 14182 5108 14188 5160
rect 14240 5148 14246 5160
rect 14562 5151 14620 5157
rect 14562 5148 14574 5151
rect 14240 5120 14574 5148
rect 14240 5108 14246 5120
rect 14562 5117 14574 5120
rect 14608 5117 14620 5151
rect 14562 5111 14620 5117
rect 14918 5108 14924 5160
rect 14976 5148 14982 5160
rect 15194 5148 15200 5160
rect 14976 5120 15021 5148
rect 15107 5120 15200 5148
rect 14976 5108 14982 5120
rect 15194 5108 15200 5120
rect 15252 5108 15258 5160
rect 15470 5148 15476 5160
rect 15396 5120 15476 5148
rect 15212 5080 15240 5108
rect 13004 5052 14504 5080
rect 12814 5043 12872 5049
rect 6457 5015 6515 5021
rect 6457 5012 6469 5015
rect 5184 4984 6469 5012
rect 6457 4981 6469 4984
rect 6503 4981 6515 5015
rect 6457 4975 6515 4981
rect 6638 4972 6644 5024
rect 6696 5012 6702 5024
rect 6733 5015 6791 5021
rect 6733 5012 6745 5015
rect 6696 4984 6745 5012
rect 6696 4972 6702 4984
rect 6733 4981 6745 4984
rect 6779 4981 6791 5015
rect 6733 4975 6791 4981
rect 7193 5015 7251 5021
rect 7193 4981 7205 5015
rect 7239 5012 7251 5015
rect 7282 5012 7288 5024
rect 7239 4984 7288 5012
rect 7239 4981 7251 4984
rect 7193 4975 7251 4981
rect 7282 4972 7288 4984
rect 7340 4972 7346 5024
rect 7374 4972 7380 5024
rect 7432 5012 7438 5024
rect 7561 5015 7619 5021
rect 7561 5012 7573 5015
rect 7432 4984 7573 5012
rect 7432 4972 7438 4984
rect 7561 4981 7573 4984
rect 7607 4981 7619 5015
rect 7561 4975 7619 4981
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 8021 5015 8079 5021
rect 8021 5012 8033 5015
rect 7708 4984 8033 5012
rect 7708 4972 7714 4984
rect 8021 4981 8033 4984
rect 8067 4981 8079 5015
rect 8021 4975 8079 4981
rect 8386 4972 8392 5024
rect 8444 5012 8450 5024
rect 9122 5012 9128 5024
rect 8444 4984 9128 5012
rect 8444 4972 8450 4984
rect 9122 4972 9128 4984
rect 9180 4972 9186 5024
rect 9490 5012 9496 5024
rect 9451 4984 9496 5012
rect 9490 4972 9496 4984
rect 9548 4972 9554 5024
rect 9674 4972 9680 5024
rect 9732 5012 9738 5024
rect 9769 5015 9827 5021
rect 9769 5012 9781 5015
rect 9732 4984 9781 5012
rect 9732 4972 9738 4984
rect 9769 4981 9781 4984
rect 9815 4981 9827 5015
rect 11238 5012 11244 5024
rect 11199 4984 11244 5012
rect 9769 4975 9827 4981
rect 11238 4972 11244 4984
rect 11296 4972 11302 5024
rect 12829 5012 12857 5043
rect 13449 5015 13507 5021
rect 13449 5012 13461 5015
rect 12829 4984 13461 5012
rect 13449 4981 13461 4984
rect 13495 4981 13507 5015
rect 14476 5012 14504 5052
rect 15028 5052 15240 5080
rect 15028 5012 15056 5052
rect 14476 4984 15056 5012
rect 13449 4975 13507 4981
rect 15194 4972 15200 5024
rect 15252 5012 15258 5024
rect 15396 5012 15424 5120
rect 15470 5108 15476 5120
rect 15528 5108 15534 5160
rect 15654 5108 15660 5160
rect 15712 5148 15718 5160
rect 15841 5151 15899 5157
rect 15841 5148 15853 5151
rect 15712 5120 15853 5148
rect 15712 5108 15718 5120
rect 15841 5117 15853 5120
rect 15887 5117 15899 5151
rect 16298 5148 16304 5160
rect 16259 5120 16304 5148
rect 15841 5111 15899 5117
rect 16298 5108 16304 5120
rect 16356 5108 16362 5160
rect 16592 5157 16620 5188
rect 16666 5176 16672 5188
rect 16724 5176 16730 5228
rect 17788 5225 17816 5256
rect 17773 5219 17831 5225
rect 17773 5185 17785 5219
rect 17819 5216 17831 5219
rect 17862 5216 17868 5228
rect 17819 5188 17868 5216
rect 17819 5185 17831 5188
rect 17773 5179 17831 5185
rect 17862 5176 17868 5188
rect 17920 5176 17926 5228
rect 16577 5151 16635 5157
rect 16577 5117 16589 5151
rect 16623 5117 16635 5151
rect 16945 5151 17003 5157
rect 16945 5148 16957 5151
rect 16577 5111 16635 5117
rect 16684 5120 16957 5148
rect 15930 5080 15936 5092
rect 15891 5052 15936 5080
rect 15930 5040 15936 5052
rect 15988 5040 15994 5092
rect 16316 5080 16344 5108
rect 16684 5080 16712 5120
rect 16945 5117 16957 5120
rect 16991 5117 17003 5151
rect 16945 5111 17003 5117
rect 18046 5108 18052 5160
rect 18104 5148 18110 5160
rect 18141 5151 18199 5157
rect 18141 5148 18153 5151
rect 18104 5120 18153 5148
rect 18104 5108 18110 5120
rect 18141 5117 18153 5120
rect 18187 5117 18199 5151
rect 18141 5111 18199 5117
rect 18325 5083 18383 5089
rect 18325 5080 18337 5083
rect 16316 5052 16712 5080
rect 16776 5052 18337 5080
rect 15252 4984 15424 5012
rect 15252 4972 15258 4984
rect 15470 4972 15476 5024
rect 15528 5012 15534 5024
rect 16776 5021 16804 5052
rect 18325 5049 18337 5052
rect 18371 5049 18383 5083
rect 18506 5080 18512 5092
rect 18467 5052 18512 5080
rect 18325 5043 18383 5049
rect 18506 5040 18512 5052
rect 18564 5040 18570 5092
rect 16761 5015 16819 5021
rect 15528 4984 15573 5012
rect 15528 4972 15534 4984
rect 16761 4981 16773 5015
rect 16807 4981 16819 5015
rect 16761 4975 16819 4981
rect 17129 5015 17187 5021
rect 17129 4981 17141 5015
rect 17175 5012 17187 5015
rect 17310 5012 17316 5024
rect 17175 4984 17316 5012
rect 17175 4981 17187 4984
rect 17129 4975 17187 4981
rect 17310 4972 17316 4984
rect 17368 4972 17374 5024
rect 17402 4972 17408 5024
rect 17460 5012 17466 5024
rect 17497 5015 17555 5021
rect 17497 5012 17509 5015
rect 17460 4984 17509 5012
rect 17460 4972 17466 4984
rect 17497 4981 17509 4984
rect 17543 4981 17555 5015
rect 17497 4975 17555 4981
rect 17589 5015 17647 5021
rect 17589 4981 17601 5015
rect 17635 5012 17647 5015
rect 17678 5012 17684 5024
rect 17635 4984 17684 5012
rect 17635 4981 17647 4984
rect 17589 4975 17647 4981
rect 17678 4972 17684 4984
rect 17736 4972 17742 5024
rect 17954 5012 17960 5024
rect 17915 4984 17960 5012
rect 17954 4972 17960 4984
rect 18012 4972 18018 5024
rect 1104 4922 18860 4944
rect 1104 4870 6912 4922
rect 6964 4870 6976 4922
rect 7028 4870 7040 4922
rect 7092 4870 7104 4922
rect 7156 4870 12843 4922
rect 12895 4870 12907 4922
rect 12959 4870 12971 4922
rect 13023 4870 13035 4922
rect 13087 4870 18860 4922
rect 1104 4848 18860 4870
rect 1765 4811 1823 4817
rect 1765 4777 1777 4811
rect 1811 4808 1823 4811
rect 1946 4808 1952 4820
rect 1811 4780 1952 4808
rect 1811 4777 1823 4780
rect 1765 4771 1823 4777
rect 1946 4768 1952 4780
rect 2004 4768 2010 4820
rect 2038 4768 2044 4820
rect 2096 4808 2102 4820
rect 2225 4811 2283 4817
rect 2225 4808 2237 4811
rect 2096 4780 2237 4808
rect 2096 4768 2102 4780
rect 2225 4777 2237 4780
rect 2271 4777 2283 4811
rect 2225 4771 2283 4777
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 2961 4811 3019 4817
rect 2961 4808 2973 4811
rect 2832 4780 2973 4808
rect 2832 4768 2838 4780
rect 2961 4777 2973 4780
rect 3007 4808 3019 4811
rect 3007 4780 5764 4808
rect 3007 4777 3019 4780
rect 2961 4771 3019 4777
rect 1581 4743 1639 4749
rect 1581 4709 1593 4743
rect 1627 4740 1639 4743
rect 4154 4740 4160 4752
rect 1627 4712 4160 4740
rect 1627 4709 1639 4712
rect 1581 4703 1639 4709
rect 4154 4700 4160 4712
rect 4212 4700 4218 4752
rect 4985 4743 5043 4749
rect 4985 4740 4997 4743
rect 4816 4712 4997 4740
rect 4816 4684 4844 4712
rect 4985 4709 4997 4712
rect 5031 4709 5043 4743
rect 4985 4703 5043 4709
rect 5166 4700 5172 4752
rect 5224 4740 5230 4752
rect 5736 4740 5764 4780
rect 5902 4768 5908 4820
rect 5960 4808 5966 4820
rect 6181 4811 6239 4817
rect 6181 4808 6193 4811
rect 5960 4780 6193 4808
rect 5960 4768 5966 4780
rect 6181 4777 6193 4780
rect 6227 4777 6239 4811
rect 6638 4808 6644 4820
rect 6599 4780 6644 4808
rect 6181 4771 6239 4777
rect 6638 4768 6644 4780
rect 6696 4768 6702 4820
rect 7009 4811 7067 4817
rect 7009 4777 7021 4811
rect 7055 4808 7067 4811
rect 7282 4808 7288 4820
rect 7055 4780 7288 4808
rect 7055 4777 7067 4780
rect 7009 4771 7067 4777
rect 7282 4768 7288 4780
rect 7340 4768 7346 4820
rect 8110 4808 8116 4820
rect 8071 4780 8116 4808
rect 8110 4768 8116 4780
rect 8168 4768 8174 4820
rect 8481 4811 8539 4817
rect 8481 4777 8493 4811
rect 8527 4808 8539 4811
rect 9585 4811 9643 4817
rect 9585 4808 9597 4811
rect 8527 4780 9597 4808
rect 8527 4777 8539 4780
rect 8481 4771 8539 4777
rect 9585 4777 9597 4780
rect 9631 4777 9643 4811
rect 9950 4808 9956 4820
rect 9911 4780 9956 4808
rect 9585 4771 9643 4777
rect 9950 4768 9956 4780
rect 10008 4768 10014 4820
rect 10045 4811 10103 4817
rect 10045 4777 10057 4811
rect 10091 4808 10103 4811
rect 10594 4808 10600 4820
rect 10091 4780 10600 4808
rect 10091 4777 10103 4780
rect 10045 4771 10103 4777
rect 10594 4768 10600 4780
rect 10652 4768 10658 4820
rect 10781 4811 10839 4817
rect 10781 4777 10793 4811
rect 10827 4808 10839 4811
rect 11054 4808 11060 4820
rect 10827 4780 11060 4808
rect 10827 4777 10839 4780
rect 10781 4771 10839 4777
rect 11054 4768 11060 4780
rect 11112 4768 11118 4820
rect 11517 4811 11575 4817
rect 11517 4777 11529 4811
rect 11563 4808 11575 4811
rect 11790 4808 11796 4820
rect 11563 4780 11796 4808
rect 11563 4777 11575 4780
rect 11517 4771 11575 4777
rect 11790 4768 11796 4780
rect 11848 4768 11854 4820
rect 11977 4811 12035 4817
rect 11977 4777 11989 4811
rect 12023 4808 12035 4811
rect 12526 4808 12532 4820
rect 12023 4780 12532 4808
rect 12023 4777 12035 4780
rect 11977 4771 12035 4777
rect 12526 4768 12532 4780
rect 12584 4768 12590 4820
rect 12710 4768 12716 4820
rect 12768 4808 12774 4820
rect 12805 4811 12863 4817
rect 12805 4808 12817 4811
rect 12768 4780 12817 4808
rect 12768 4768 12774 4780
rect 12805 4777 12817 4780
rect 12851 4777 12863 4811
rect 12805 4771 12863 4777
rect 13357 4811 13415 4817
rect 13357 4777 13369 4811
rect 13403 4808 13415 4811
rect 13630 4808 13636 4820
rect 13403 4780 13636 4808
rect 13403 4777 13415 4780
rect 13357 4771 13415 4777
rect 13630 4768 13636 4780
rect 13688 4768 13694 4820
rect 14185 4811 14243 4817
rect 14185 4777 14197 4811
rect 14231 4808 14243 4811
rect 14550 4808 14556 4820
rect 14231 4780 14556 4808
rect 14231 4777 14243 4780
rect 14185 4771 14243 4777
rect 14550 4768 14556 4780
rect 14608 4768 14614 4820
rect 14734 4768 14740 4820
rect 14792 4808 14798 4820
rect 17402 4808 17408 4820
rect 14792 4780 17408 4808
rect 14792 4768 14798 4780
rect 17402 4768 17408 4780
rect 17460 4768 17466 4820
rect 17494 4768 17500 4820
rect 17552 4768 17558 4820
rect 6549 4743 6607 4749
rect 5224 4712 5580 4740
rect 5736 4712 6500 4740
rect 5224 4700 5230 4712
rect 2133 4675 2191 4681
rect 2133 4641 2145 4675
rect 2179 4672 2191 4675
rect 3421 4675 3479 4681
rect 3421 4672 3433 4675
rect 2179 4644 3433 4672
rect 2179 4641 2191 4644
rect 2133 4635 2191 4641
rect 3421 4641 3433 4644
rect 3467 4672 3479 4675
rect 3602 4672 3608 4684
rect 3467 4644 3608 4672
rect 3467 4641 3479 4644
rect 3421 4635 3479 4641
rect 3602 4632 3608 4644
rect 3660 4632 3666 4684
rect 3786 4632 3792 4684
rect 3844 4672 3850 4684
rect 4065 4675 4123 4681
rect 4065 4672 4077 4675
rect 3844 4644 4077 4672
rect 3844 4632 3850 4644
rect 4065 4641 4077 4644
rect 4111 4641 4123 4675
rect 4065 4635 4123 4641
rect 4341 4675 4399 4681
rect 4341 4641 4353 4675
rect 4387 4641 4399 4675
rect 4341 4635 4399 4641
rect 2314 4604 2320 4616
rect 2275 4576 2320 4604
rect 2314 4564 2320 4576
rect 2372 4564 2378 4616
rect 3053 4607 3111 4613
rect 3053 4573 3065 4607
rect 3099 4604 3111 4607
rect 3142 4604 3148 4616
rect 3099 4576 3148 4604
rect 3099 4573 3111 4576
rect 3053 4567 3111 4573
rect 3142 4564 3148 4576
rect 3200 4564 3206 4616
rect 3237 4607 3295 4613
rect 3237 4573 3249 4607
rect 3283 4604 3295 4607
rect 3510 4604 3516 4616
rect 3283 4576 3516 4604
rect 3283 4573 3295 4576
rect 3237 4567 3295 4573
rect 3510 4564 3516 4576
rect 3568 4564 3574 4616
rect 4356 4604 4384 4635
rect 4798 4632 4804 4684
rect 4856 4632 4862 4684
rect 4893 4675 4951 4681
rect 4893 4641 4905 4675
rect 4939 4672 4951 4675
rect 5442 4672 5448 4684
rect 4939 4644 5448 4672
rect 4939 4641 4951 4644
rect 4893 4635 4951 4641
rect 5442 4632 5448 4644
rect 5500 4632 5506 4684
rect 5552 4681 5580 4712
rect 6472 4684 6500 4712
rect 6549 4709 6561 4743
rect 6595 4740 6607 4743
rect 7190 4740 7196 4752
rect 6595 4712 7196 4740
rect 6595 4709 6607 4712
rect 6549 4703 6607 4709
rect 7190 4700 7196 4712
rect 7248 4700 7254 4752
rect 7466 4740 7472 4752
rect 7392 4712 7472 4740
rect 5537 4675 5595 4681
rect 5537 4641 5549 4675
rect 5583 4672 5595 4675
rect 5813 4675 5871 4681
rect 5583 4644 5764 4672
rect 5583 4641 5595 4644
rect 5537 4635 5595 4641
rect 5166 4604 5172 4616
rect 4356 4576 5028 4604
rect 5127 4576 5172 4604
rect 1762 4496 1768 4548
rect 1820 4536 1826 4548
rect 2593 4539 2651 4545
rect 2593 4536 2605 4539
rect 1820 4508 2605 4536
rect 1820 4496 1826 4508
rect 2593 4505 2605 4508
rect 2639 4505 2651 4539
rect 2593 4499 2651 4505
rect 2866 4496 2872 4548
rect 2924 4536 2930 4548
rect 3881 4539 3939 4545
rect 3881 4536 3893 4539
rect 2924 4508 3893 4536
rect 2924 4496 2930 4508
rect 3881 4505 3893 4508
rect 3927 4505 3939 4539
rect 3881 4499 3939 4505
rect 4157 4539 4215 4545
rect 4157 4505 4169 4539
rect 4203 4536 4215 4539
rect 4798 4536 4804 4548
rect 4203 4508 4804 4536
rect 4203 4505 4215 4508
rect 4157 4499 4215 4505
rect 4798 4496 4804 4508
rect 4856 4496 4862 4548
rect 5000 4536 5028 4576
rect 5166 4564 5172 4576
rect 5224 4564 5230 4616
rect 5350 4564 5356 4616
rect 5408 4604 5414 4616
rect 5408 4576 5672 4604
rect 5408 4564 5414 4576
rect 5258 4536 5264 4548
rect 5000 4508 5264 4536
rect 5258 4496 5264 4508
rect 5316 4496 5322 4548
rect 5644 4545 5672 4576
rect 5629 4539 5687 4545
rect 5629 4505 5641 4539
rect 5675 4505 5687 4539
rect 5736 4536 5764 4644
rect 5813 4641 5825 4675
rect 5859 4641 5871 4675
rect 5813 4635 5871 4641
rect 6089 4675 6147 4681
rect 6089 4641 6101 4675
rect 6135 4672 6147 4675
rect 6135 4644 6408 4672
rect 6135 4641 6147 4644
rect 6089 4635 6147 4641
rect 5828 4604 5856 4635
rect 6270 4604 6276 4616
rect 5828 4576 6276 4604
rect 6270 4564 6276 4576
rect 6328 4564 6334 4616
rect 6380 4536 6408 4644
rect 6454 4632 6460 4684
rect 6512 4672 6518 4684
rect 7392 4681 7420 4712
rect 7466 4700 7472 4712
rect 7524 4700 7530 4752
rect 7837 4743 7895 4749
rect 7837 4709 7849 4743
rect 7883 4740 7895 4743
rect 10689 4743 10747 4749
rect 7883 4712 10548 4740
rect 7883 4709 7895 4712
rect 7837 4703 7895 4709
rect 7377 4675 7435 4681
rect 7377 4672 7389 4675
rect 6512 4644 7389 4672
rect 6512 4632 6518 4644
rect 7377 4641 7389 4644
rect 7423 4641 7435 4675
rect 8386 4672 8392 4684
rect 7377 4635 7435 4641
rect 7484 4644 8392 4672
rect 6546 4564 6552 4616
rect 6604 4604 6610 4616
rect 6733 4607 6791 4613
rect 6733 4604 6745 4607
rect 6604 4576 6745 4604
rect 6604 4564 6610 4576
rect 6733 4573 6745 4576
rect 6779 4573 6791 4607
rect 6733 4567 6791 4573
rect 6822 4564 6828 4616
rect 6880 4604 6886 4616
rect 7484 4613 7512 4644
rect 8386 4632 8392 4644
rect 8444 4632 8450 4684
rect 8570 4672 8576 4684
rect 8531 4644 8576 4672
rect 8570 4632 8576 4644
rect 8628 4632 8634 4684
rect 8662 4632 8668 4684
rect 8720 4672 8726 4684
rect 9309 4675 9367 4681
rect 9309 4672 9321 4675
rect 8720 4644 9321 4672
rect 8720 4632 8726 4644
rect 9309 4641 9321 4644
rect 9355 4641 9367 4675
rect 9309 4635 9367 4641
rect 9398 4632 9404 4684
rect 9456 4672 9462 4684
rect 10410 4672 10416 4684
rect 9456 4644 9501 4672
rect 9876 4644 10416 4672
rect 9456 4632 9462 4644
rect 7469 4607 7527 4613
rect 7469 4604 7481 4607
rect 6880 4576 7481 4604
rect 6880 4564 6886 4576
rect 7469 4573 7481 4576
rect 7515 4573 7527 4607
rect 7469 4567 7527 4573
rect 7558 4564 7564 4616
rect 7616 4604 7622 4616
rect 8297 4607 8355 4613
rect 7616 4576 7661 4604
rect 7616 4564 7622 4576
rect 8297 4573 8309 4607
rect 8343 4604 8355 4607
rect 9876 4604 9904 4644
rect 10410 4632 10416 4644
rect 10468 4632 10474 4684
rect 10226 4604 10232 4616
rect 8343 4576 9904 4604
rect 10187 4576 10232 4604
rect 8343 4573 8355 4576
rect 8297 4567 8355 4573
rect 10226 4564 10232 4576
rect 10284 4564 10290 4616
rect 7837 4539 7895 4545
rect 7837 4536 7849 4539
rect 5736 4508 6040 4536
rect 6380 4508 7849 4536
rect 5629 4499 5687 4505
rect 1486 4468 1492 4480
rect 1447 4440 1492 4468
rect 1486 4428 1492 4440
rect 1544 4428 1550 4480
rect 3602 4468 3608 4480
rect 3563 4440 3608 4468
rect 3602 4428 3608 4440
rect 3660 4428 3666 4480
rect 4522 4468 4528 4480
rect 4483 4440 4528 4468
rect 4522 4428 4528 4440
rect 4580 4428 4586 4480
rect 4706 4428 4712 4480
rect 4764 4468 4770 4480
rect 5353 4471 5411 4477
rect 5353 4468 5365 4471
rect 4764 4440 5365 4468
rect 4764 4428 4770 4440
rect 5353 4437 5365 4440
rect 5399 4437 5411 4471
rect 5353 4431 5411 4437
rect 5718 4428 5724 4480
rect 5776 4468 5782 4480
rect 5905 4471 5963 4477
rect 5905 4468 5917 4471
rect 5776 4440 5917 4468
rect 5776 4428 5782 4440
rect 5905 4437 5917 4440
rect 5951 4437 5963 4471
rect 6012 4468 6040 4508
rect 7837 4505 7849 4508
rect 7883 4505 7895 4539
rect 7837 4499 7895 4505
rect 8386 4496 8392 4548
rect 8444 4536 8450 4548
rect 9125 4539 9183 4545
rect 9125 4536 9137 4539
rect 8444 4508 9137 4536
rect 8444 4496 8450 4508
rect 9125 4505 9137 4508
rect 9171 4505 9183 4539
rect 9125 4499 9183 4505
rect 9950 4496 9956 4548
rect 10008 4496 10014 4548
rect 10520 4536 10548 4712
rect 10689 4709 10701 4743
rect 10735 4740 10747 4743
rect 11422 4740 11428 4752
rect 10735 4712 11428 4740
rect 10735 4709 10747 4712
rect 10689 4703 10747 4709
rect 11422 4700 11428 4712
rect 11480 4700 11486 4752
rect 11609 4743 11667 4749
rect 11609 4709 11621 4743
rect 11655 4740 11667 4743
rect 13725 4743 13783 4749
rect 13725 4740 13737 4743
rect 11655 4712 13737 4740
rect 11655 4709 11667 4712
rect 11609 4703 11667 4709
rect 13725 4709 13737 4712
rect 13771 4709 13783 4743
rect 13725 4703 13783 4709
rect 14921 4743 14979 4749
rect 14921 4709 14933 4743
rect 14967 4740 14979 4743
rect 15102 4740 15108 4752
rect 14967 4712 15108 4740
rect 14967 4709 14979 4712
rect 14921 4703 14979 4709
rect 15102 4700 15108 4712
rect 15160 4700 15166 4752
rect 15280 4743 15338 4749
rect 15280 4709 15292 4743
rect 15326 4740 15338 4743
rect 16206 4740 16212 4752
rect 15326 4712 16212 4740
rect 15326 4709 15338 4712
rect 15280 4703 15338 4709
rect 16206 4700 16212 4712
rect 16264 4740 16270 4752
rect 16666 4740 16672 4752
rect 16264 4712 16672 4740
rect 16264 4700 16270 4712
rect 16666 4700 16672 4712
rect 16724 4700 16730 4752
rect 17512 4740 17540 4768
rect 18325 4743 18383 4749
rect 18325 4740 18337 4743
rect 17512 4712 18337 4740
rect 18325 4709 18337 4712
rect 18371 4709 18383 4743
rect 18325 4703 18383 4709
rect 11698 4672 11704 4684
rect 10612 4644 11704 4672
rect 10612 4613 10640 4644
rect 11698 4632 11704 4644
rect 11756 4632 11762 4684
rect 12250 4632 12256 4684
rect 12308 4672 12314 4684
rect 12434 4672 12440 4684
rect 12308 4644 12440 4672
rect 12308 4632 12314 4644
rect 12434 4632 12440 4644
rect 12492 4632 12498 4684
rect 13170 4632 13176 4684
rect 13228 4672 13234 4684
rect 13265 4675 13323 4681
rect 13265 4672 13277 4675
rect 13228 4644 13277 4672
rect 13228 4632 13234 4644
rect 13265 4641 13277 4644
rect 13311 4672 13323 4675
rect 14553 4675 14611 4681
rect 13311 4644 14504 4672
rect 13311 4641 13323 4644
rect 13265 4635 13323 4641
rect 10597 4607 10655 4613
rect 10597 4573 10609 4607
rect 10643 4573 10655 4607
rect 10597 4567 10655 4573
rect 11425 4607 11483 4613
rect 11425 4573 11437 4607
rect 11471 4604 11483 4607
rect 12161 4607 12219 4613
rect 12161 4604 12173 4607
rect 11471 4576 12173 4604
rect 11471 4573 11483 4576
rect 11425 4567 11483 4573
rect 12161 4573 12173 4576
rect 12207 4573 12219 4607
rect 12161 4567 12219 4573
rect 12345 4607 12403 4613
rect 12345 4573 12357 4607
rect 12391 4604 12403 4607
rect 12526 4604 12532 4616
rect 12391 4576 12532 4604
rect 12391 4573 12403 4576
rect 12345 4567 12403 4573
rect 10962 4536 10968 4548
rect 10520 4508 10968 4536
rect 10962 4496 10968 4508
rect 11020 4496 11026 4548
rect 12176 4536 12204 4567
rect 12526 4564 12532 4576
rect 12584 4564 12590 4616
rect 13541 4607 13599 4613
rect 13541 4573 13553 4607
rect 13587 4573 13599 4607
rect 13541 4567 13599 4573
rect 12176 4508 13400 4536
rect 6546 4468 6552 4480
rect 6012 4440 6552 4468
rect 5905 4431 5963 4437
rect 6546 4428 6552 4440
rect 6604 4428 6610 4480
rect 8938 4468 8944 4480
rect 8899 4440 8944 4468
rect 8938 4428 8944 4440
rect 8996 4428 9002 4480
rect 9214 4428 9220 4480
rect 9272 4468 9278 4480
rect 9968 4468 9996 4496
rect 9272 4440 9996 4468
rect 9272 4428 9278 4440
rect 11054 4428 11060 4480
rect 11112 4468 11118 4480
rect 11149 4471 11207 4477
rect 11149 4468 11161 4471
rect 11112 4440 11161 4468
rect 11112 4428 11118 4440
rect 11149 4437 11161 4440
rect 11195 4437 11207 4471
rect 11149 4431 11207 4437
rect 11698 4428 11704 4480
rect 11756 4468 11762 4480
rect 11974 4468 11980 4480
rect 11756 4440 11980 4468
rect 11756 4428 11762 4440
rect 11974 4428 11980 4440
rect 12032 4428 12038 4480
rect 12250 4428 12256 4480
rect 12308 4468 12314 4480
rect 12897 4471 12955 4477
rect 12897 4468 12909 4471
rect 12308 4440 12909 4468
rect 12308 4428 12314 4440
rect 12897 4437 12909 4440
rect 12943 4437 12955 4471
rect 13372 4468 13400 4508
rect 13556 4468 13584 4567
rect 14366 4536 14372 4548
rect 14327 4508 14372 4536
rect 14366 4496 14372 4508
rect 14424 4496 14430 4548
rect 13814 4468 13820 4480
rect 13372 4440 13820 4468
rect 12897 4431 12955 4437
rect 13814 4428 13820 4440
rect 13872 4468 13878 4480
rect 14182 4468 14188 4480
rect 13872 4440 14188 4468
rect 13872 4428 13878 4440
rect 14182 4428 14188 4440
rect 14240 4428 14246 4480
rect 14476 4468 14504 4644
rect 14553 4641 14565 4675
rect 14599 4672 14611 4675
rect 14737 4675 14795 4681
rect 14737 4672 14749 4675
rect 14599 4644 14749 4672
rect 14599 4641 14611 4644
rect 14553 4635 14611 4641
rect 14737 4641 14749 4644
rect 14783 4672 14795 4675
rect 16298 4672 16304 4684
rect 14783 4644 16304 4672
rect 14783 4641 14795 4644
rect 14737 4635 14795 4641
rect 16298 4632 16304 4644
rect 16356 4632 16362 4684
rect 16574 4672 16580 4684
rect 16535 4644 16580 4672
rect 16574 4632 16580 4644
rect 16632 4632 16638 4684
rect 16853 4675 16911 4681
rect 16853 4641 16865 4675
rect 16899 4641 16911 4675
rect 16853 4635 16911 4641
rect 15010 4604 15016 4616
rect 14971 4576 15016 4604
rect 15010 4564 15016 4576
rect 15068 4564 15074 4616
rect 16868 4536 16896 4635
rect 16942 4632 16948 4684
rect 17000 4672 17006 4684
rect 17497 4675 17555 4681
rect 17497 4672 17509 4675
rect 17000 4644 17509 4672
rect 17000 4632 17006 4644
rect 17497 4641 17509 4644
rect 17543 4641 17555 4675
rect 17957 4675 18015 4681
rect 17957 4672 17969 4675
rect 17497 4635 17555 4641
rect 17604 4644 17969 4672
rect 17126 4604 17132 4616
rect 15948 4508 16896 4536
rect 16960 4576 17132 4604
rect 15948 4468 15976 4508
rect 14476 4440 15976 4468
rect 16206 4428 16212 4480
rect 16264 4468 16270 4480
rect 16393 4471 16451 4477
rect 16393 4468 16405 4471
rect 16264 4440 16405 4468
rect 16264 4428 16270 4440
rect 16393 4437 16405 4440
rect 16439 4437 16451 4471
rect 16393 4431 16451 4437
rect 16761 4471 16819 4477
rect 16761 4437 16773 4471
rect 16807 4468 16819 4471
rect 16960 4468 16988 4576
rect 17126 4564 17132 4576
rect 17184 4564 17190 4616
rect 17402 4564 17408 4616
rect 17460 4604 17466 4616
rect 17604 4613 17632 4644
rect 17957 4641 17969 4644
rect 18003 4641 18015 4675
rect 18506 4672 18512 4684
rect 18467 4644 18512 4672
rect 17957 4635 18015 4641
rect 18506 4632 18512 4644
rect 18564 4632 18570 4684
rect 17589 4607 17647 4613
rect 17589 4604 17601 4607
rect 17460 4576 17601 4604
rect 17460 4564 17466 4576
rect 17589 4573 17601 4576
rect 17635 4573 17647 4607
rect 17589 4567 17647 4573
rect 17773 4607 17831 4613
rect 17773 4573 17785 4607
rect 17819 4604 17831 4607
rect 17862 4604 17868 4616
rect 17819 4576 17868 4604
rect 17819 4573 17831 4576
rect 17773 4567 17831 4573
rect 17862 4564 17868 4576
rect 17920 4564 17926 4616
rect 17037 4539 17095 4545
rect 17037 4505 17049 4539
rect 17083 4536 17095 4539
rect 18046 4536 18052 4548
rect 17083 4508 18052 4536
rect 17083 4505 17095 4508
rect 17037 4499 17095 4505
rect 18046 4496 18052 4508
rect 18104 4496 18110 4548
rect 16807 4440 16988 4468
rect 16807 4437 16819 4440
rect 16761 4431 16819 4437
rect 17126 4428 17132 4480
rect 17184 4468 17190 4480
rect 18141 4471 18199 4477
rect 17184 4440 17229 4468
rect 17184 4428 17190 4440
rect 18141 4437 18153 4471
rect 18187 4468 18199 4471
rect 18322 4468 18328 4480
rect 18187 4440 18328 4468
rect 18187 4437 18199 4440
rect 18141 4431 18199 4437
rect 18322 4428 18328 4440
rect 18380 4428 18386 4480
rect 1104 4378 18860 4400
rect 1104 4326 3947 4378
rect 3999 4326 4011 4378
rect 4063 4326 4075 4378
rect 4127 4326 4139 4378
rect 4191 4326 9878 4378
rect 9930 4326 9942 4378
rect 9994 4326 10006 4378
rect 10058 4326 10070 4378
rect 10122 4326 15808 4378
rect 15860 4326 15872 4378
rect 15924 4326 15936 4378
rect 15988 4326 16000 4378
rect 16052 4326 18860 4378
rect 1104 4304 18860 4326
rect 382 4224 388 4276
rect 440 4264 446 4276
rect 3326 4264 3332 4276
rect 440 4236 3332 4264
rect 440 4224 446 4236
rect 3326 4224 3332 4236
rect 3384 4224 3390 4276
rect 5166 4264 5172 4276
rect 5079 4236 5172 4264
rect 5166 4224 5172 4236
rect 5224 4264 5230 4276
rect 6270 4264 6276 4276
rect 5224 4236 5948 4264
rect 6183 4236 6276 4264
rect 5224 4224 5230 4236
rect 2406 4156 2412 4208
rect 2464 4196 2470 4208
rect 2501 4199 2559 4205
rect 2501 4196 2513 4199
rect 2464 4168 2513 4196
rect 2464 4156 2470 4168
rect 2501 4165 2513 4168
rect 2547 4165 2559 4199
rect 2501 4159 2559 4165
rect 4154 4156 4160 4208
rect 4212 4196 4218 4208
rect 4430 4196 4436 4208
rect 4212 4168 4436 4196
rect 4212 4156 4218 4168
rect 4430 4156 4436 4168
rect 4488 4156 4494 4208
rect 2130 4128 2136 4140
rect 2091 4100 2136 4128
rect 2130 4088 2136 4100
rect 2188 4088 2194 4140
rect 2590 4128 2596 4140
rect 2516 4100 2596 4128
rect 1578 4060 1584 4072
rect 1539 4032 1584 4060
rect 1578 4020 1584 4032
rect 1636 4020 1642 4072
rect 2516 4060 2544 4100
rect 2590 4088 2596 4100
rect 2648 4088 2654 4140
rect 3970 4088 3976 4140
rect 4028 4128 4034 4140
rect 5184 4137 5212 4224
rect 5350 4196 5356 4208
rect 5311 4168 5356 4196
rect 5350 4156 5356 4168
rect 5408 4156 5414 4208
rect 5920 4140 5948 4236
rect 6270 4224 6276 4236
rect 6328 4264 6334 4276
rect 7650 4264 7656 4276
rect 6328 4236 7656 4264
rect 6328 4224 6334 4236
rect 7650 4224 7656 4236
rect 7708 4224 7714 4276
rect 7834 4224 7840 4276
rect 7892 4224 7898 4276
rect 8202 4224 8208 4276
rect 8260 4264 8266 4276
rect 8297 4267 8355 4273
rect 8297 4264 8309 4267
rect 8260 4236 8309 4264
rect 8260 4224 8266 4236
rect 8297 4233 8309 4236
rect 8343 4233 8355 4267
rect 10962 4264 10968 4276
rect 8297 4227 8355 4233
rect 8404 4236 10088 4264
rect 6730 4196 6736 4208
rect 6691 4168 6736 4196
rect 6730 4156 6736 4168
rect 6788 4156 6794 4208
rect 7852 4196 7880 4224
rect 8404 4196 8432 4236
rect 10060 4208 10088 4236
rect 10152 4236 10968 4264
rect 7852 4168 8432 4196
rect 9784 4168 9996 4196
rect 5169 4131 5227 4137
rect 5169 4128 5181 4131
rect 4028 4100 5181 4128
rect 4028 4088 4034 4100
rect 5169 4097 5181 4100
rect 5215 4097 5227 4131
rect 5810 4128 5816 4140
rect 5771 4100 5816 4128
rect 5169 4091 5227 4097
rect 5810 4088 5816 4100
rect 5868 4088 5874 4140
rect 5902 4088 5908 4140
rect 5960 4128 5966 4140
rect 5960 4100 6005 4128
rect 5960 4088 5966 4100
rect 6086 4088 6092 4140
rect 6144 4128 6150 4140
rect 9784 4137 9812 4168
rect 6917 4131 6975 4137
rect 6917 4128 6929 4131
rect 6144 4100 6929 4128
rect 6144 4088 6150 4100
rect 6917 4097 6929 4100
rect 6963 4097 6975 4131
rect 6917 4091 6975 4097
rect 9769 4131 9827 4137
rect 9769 4097 9781 4131
rect 9815 4097 9827 4131
rect 9968 4128 9996 4168
rect 10042 4156 10048 4208
rect 10100 4156 10106 4208
rect 10152 4128 10180 4236
rect 10962 4224 10968 4236
rect 11020 4224 11026 4276
rect 11054 4224 11060 4276
rect 11112 4264 11118 4276
rect 14734 4264 14740 4276
rect 11112 4236 14740 4264
rect 11112 4224 11118 4236
rect 14734 4224 14740 4236
rect 14792 4224 14798 4276
rect 16485 4267 16543 4273
rect 16485 4233 16497 4267
rect 16531 4264 16543 4267
rect 16574 4264 16580 4276
rect 16531 4236 16580 4264
rect 16531 4233 16543 4236
rect 16485 4227 16543 4233
rect 16574 4224 16580 4236
rect 16632 4224 16638 4276
rect 10410 4156 10416 4208
rect 10468 4196 10474 4208
rect 10594 4196 10600 4208
rect 10468 4168 10600 4196
rect 10468 4156 10474 4168
rect 10594 4156 10600 4168
rect 10652 4196 10658 4208
rect 10652 4168 11192 4196
rect 10652 4156 10658 4168
rect 9968 4100 10180 4128
rect 9769 4091 9827 4097
rect 10226 4088 10232 4140
rect 10284 4128 10290 4140
rect 10284 4100 10456 4128
rect 10284 4088 10290 4100
rect 2958 4060 2964 4072
rect 2424 4032 2544 4060
rect 2919 4032 2964 4060
rect 1949 3995 2007 4001
rect 1949 3961 1961 3995
rect 1995 3961 2007 3995
rect 1949 3955 2007 3961
rect 2317 3995 2375 4001
rect 2317 3961 2329 3995
rect 2363 3992 2375 3995
rect 2424 3992 2452 4032
rect 2958 4020 2964 4032
rect 3016 4020 3022 4072
rect 3228 4063 3286 4069
rect 3228 4029 3240 4063
rect 3274 4029 3286 4063
rect 3228 4023 3286 4029
rect 2363 3964 2452 3992
rect 2363 3961 2375 3964
rect 2317 3955 2375 3961
rect 1486 3924 1492 3936
rect 1447 3896 1492 3924
rect 1486 3884 1492 3896
rect 1544 3884 1550 3936
rect 1854 3924 1860 3936
rect 1815 3896 1860 3924
rect 1854 3884 1860 3896
rect 1912 3884 1918 3936
rect 1964 3924 1992 3955
rect 2498 3952 2504 4004
rect 2556 3992 2562 4004
rect 2685 3995 2743 4001
rect 2685 3992 2697 3995
rect 2556 3964 2697 3992
rect 2556 3952 2562 3964
rect 2685 3961 2697 3964
rect 2731 3961 2743 3995
rect 3243 3992 3271 4023
rect 3510 4020 3516 4072
rect 3568 4060 3574 4072
rect 5718 4060 5724 4072
rect 3568 4032 5724 4060
rect 3568 4020 3574 4032
rect 5718 4020 5724 4032
rect 5776 4020 5782 4072
rect 6178 4020 6184 4072
rect 6236 4060 6242 4072
rect 6638 4060 6644 4072
rect 6236 4032 6644 4060
rect 6236 4020 6242 4032
rect 6638 4020 6644 4032
rect 6696 4020 6702 4072
rect 7184 4063 7242 4069
rect 7184 4029 7196 4063
rect 7230 4060 7242 4063
rect 7558 4060 7564 4072
rect 7230 4032 7564 4060
rect 7230 4029 7242 4032
rect 7184 4023 7242 4029
rect 7558 4020 7564 4032
rect 7616 4020 7622 4072
rect 9513 4063 9571 4069
rect 9513 4029 9525 4063
rect 9559 4060 9571 4063
rect 9674 4060 9680 4072
rect 9559 4032 9680 4060
rect 9559 4029 9571 4032
rect 9513 4023 9571 4029
rect 9674 4020 9680 4032
rect 9732 4020 9738 4072
rect 9950 4020 9956 4072
rect 10008 4060 10014 4072
rect 10045 4063 10103 4069
rect 10045 4060 10057 4063
rect 10008 4032 10057 4060
rect 10008 4020 10014 4032
rect 10045 4029 10057 4032
rect 10091 4029 10103 4063
rect 10045 4023 10103 4029
rect 10321 4063 10379 4069
rect 10321 4029 10333 4063
rect 10367 4029 10379 4063
rect 10321 4023 10379 4029
rect 3970 3992 3976 4004
rect 3243 3964 3976 3992
rect 2685 3955 2743 3961
rect 3970 3952 3976 3964
rect 4028 3952 4034 4004
rect 4062 3952 4068 4004
rect 4120 3992 4126 4004
rect 4706 3992 4712 4004
rect 4120 3964 4712 3992
rect 4120 3952 4126 3964
rect 4706 3952 4712 3964
rect 4764 3952 4770 4004
rect 5258 3952 5264 4004
rect 5316 3992 5322 4004
rect 10336 3992 10364 4023
rect 5316 3964 9904 3992
rect 5316 3952 5322 3964
rect 3510 3924 3516 3936
rect 1964 3896 3516 3924
rect 3510 3884 3516 3896
rect 3568 3884 3574 3936
rect 4338 3924 4344 3936
rect 4299 3896 4344 3924
rect 4338 3884 4344 3896
rect 4396 3884 4402 3936
rect 4430 3884 4436 3936
rect 4488 3924 4494 3936
rect 4525 3927 4583 3933
rect 4525 3924 4537 3927
rect 4488 3896 4537 3924
rect 4488 3884 4494 3896
rect 4525 3893 4537 3896
rect 4571 3893 4583 3927
rect 4525 3887 4583 3893
rect 4614 3884 4620 3936
rect 4672 3924 4678 3936
rect 4893 3927 4951 3933
rect 4893 3924 4905 3927
rect 4672 3896 4905 3924
rect 4672 3884 4678 3896
rect 4893 3893 4905 3896
rect 4939 3893 4951 3927
rect 4893 3887 4951 3893
rect 4985 3927 5043 3933
rect 4985 3893 4997 3927
rect 5031 3924 5043 3927
rect 5074 3924 5080 3936
rect 5031 3896 5080 3924
rect 5031 3893 5043 3896
rect 4985 3887 5043 3893
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 5721 3927 5779 3933
rect 5721 3893 5733 3927
rect 5767 3924 5779 3927
rect 6270 3924 6276 3936
rect 5767 3896 6276 3924
rect 5767 3893 5779 3896
rect 5721 3887 5779 3893
rect 6270 3884 6276 3896
rect 6328 3884 6334 3936
rect 6454 3924 6460 3936
rect 6415 3896 6460 3924
rect 6454 3884 6460 3896
rect 6512 3884 6518 3936
rect 8110 3884 8116 3936
rect 8168 3924 8174 3936
rect 8389 3927 8447 3933
rect 8389 3924 8401 3927
rect 8168 3896 8401 3924
rect 8168 3884 8174 3896
rect 8389 3893 8401 3896
rect 8435 3893 8447 3927
rect 8389 3887 8447 3893
rect 8478 3884 8484 3936
rect 8536 3924 8542 3936
rect 9766 3924 9772 3936
rect 8536 3896 9772 3924
rect 8536 3884 8542 3896
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 9876 3933 9904 3964
rect 9968 3964 10364 3992
rect 10428 3992 10456 4100
rect 10686 4088 10692 4140
rect 10744 4128 10750 4140
rect 11164 4137 11192 4168
rect 11422 4156 11428 4208
rect 11480 4196 11486 4208
rect 11885 4199 11943 4205
rect 11885 4196 11897 4199
rect 11480 4168 11897 4196
rect 11480 4156 11486 4168
rect 11885 4165 11897 4168
rect 11931 4165 11943 4199
rect 13541 4199 13599 4205
rect 13541 4196 13553 4199
rect 11885 4159 11943 4165
rect 12360 4168 13553 4196
rect 11057 4131 11115 4137
rect 11057 4128 11069 4131
rect 10744 4100 11069 4128
rect 10744 4088 10750 4100
rect 11057 4097 11069 4100
rect 11103 4097 11115 4131
rect 11057 4091 11115 4097
rect 11149 4131 11207 4137
rect 11149 4097 11161 4131
rect 11195 4097 11207 4131
rect 11149 4091 11207 4097
rect 11517 4131 11575 4137
rect 11517 4097 11529 4131
rect 11563 4128 11575 4131
rect 12158 4128 12164 4140
rect 11563 4100 12164 4128
rect 11563 4097 11575 4100
rect 11517 4091 11575 4097
rect 12158 4088 12164 4100
rect 12216 4088 12222 4140
rect 12360 4137 12388 4168
rect 13541 4165 13553 4168
rect 13587 4165 13599 4199
rect 13541 4159 13599 4165
rect 12345 4131 12403 4137
rect 12345 4097 12357 4131
rect 12391 4097 12403 4131
rect 12345 4091 12403 4097
rect 12529 4131 12587 4137
rect 12529 4097 12541 4131
rect 12575 4128 12587 4131
rect 12618 4128 12624 4140
rect 12575 4100 12624 4128
rect 12575 4097 12587 4100
rect 12529 4091 12587 4097
rect 12618 4088 12624 4100
rect 12676 4088 12682 4140
rect 12710 4088 12716 4140
rect 12768 4128 12774 4140
rect 12805 4131 12863 4137
rect 12805 4128 12817 4131
rect 12768 4100 12817 4128
rect 12768 4088 12774 4100
rect 12805 4097 12817 4100
rect 12851 4097 12863 4131
rect 12805 4091 12863 4097
rect 13814 4088 13820 4140
rect 13872 4128 13878 4140
rect 14093 4131 14151 4137
rect 14093 4128 14105 4131
rect 13872 4100 14105 4128
rect 13872 4088 13878 4100
rect 14093 4097 14105 4100
rect 14139 4097 14151 4131
rect 15102 4128 15108 4140
rect 14093 4091 14151 4097
rect 14200 4100 15108 4128
rect 10505 4063 10563 4069
rect 10505 4029 10517 4063
rect 10551 4060 10563 4063
rect 10965 4063 11023 4069
rect 10551 4032 10925 4060
rect 10551 4029 10563 4032
rect 10505 4023 10563 4029
rect 10897 3992 10925 4032
rect 10965 4029 10977 4063
rect 11011 4060 11023 4063
rect 11330 4060 11336 4072
rect 11011 4032 11336 4060
rect 11011 4029 11023 4032
rect 10965 4023 11023 4029
rect 11330 4020 11336 4032
rect 11388 4020 11394 4072
rect 12250 4060 12256 4072
rect 12211 4032 12256 4060
rect 12250 4020 12256 4032
rect 12308 4020 12314 4072
rect 13078 4060 13084 4072
rect 13039 4032 13084 4060
rect 13078 4020 13084 4032
rect 13136 4020 13142 4072
rect 13630 4020 13636 4072
rect 13688 4060 13694 4072
rect 13909 4063 13967 4069
rect 13909 4060 13921 4063
rect 13688 4032 13921 4060
rect 13688 4020 13694 4032
rect 13909 4029 13921 4032
rect 13955 4060 13967 4063
rect 14200 4060 14228 4100
rect 15102 4088 15108 4100
rect 15160 4088 15166 4140
rect 16301 4131 16359 4137
rect 16301 4097 16313 4131
rect 16347 4128 16359 4131
rect 16482 4128 16488 4140
rect 16347 4100 16488 4128
rect 16347 4097 16359 4100
rect 16301 4091 16359 4097
rect 16482 4088 16488 4100
rect 16540 4088 16546 4140
rect 17126 4088 17132 4140
rect 17184 4128 17190 4140
rect 17405 4131 17463 4137
rect 17405 4128 17417 4131
rect 17184 4100 17417 4128
rect 17184 4088 17190 4100
rect 17405 4097 17417 4100
rect 17451 4097 17463 4131
rect 17405 4091 17463 4097
rect 17589 4131 17647 4137
rect 17589 4097 17601 4131
rect 17635 4128 17647 4131
rect 17770 4128 17776 4140
rect 17635 4100 17776 4128
rect 17635 4097 17647 4100
rect 17589 4091 17647 4097
rect 17770 4088 17776 4100
rect 17828 4088 17834 4140
rect 18138 4128 18144 4140
rect 18099 4100 18144 4128
rect 18138 4088 18144 4100
rect 18196 4088 18202 4140
rect 13955 4032 14228 4060
rect 13955 4029 13967 4032
rect 13909 4023 13967 4029
rect 14366 4020 14372 4072
rect 14424 4060 14430 4072
rect 14553 4063 14611 4069
rect 14553 4060 14565 4063
rect 14424 4032 14565 4060
rect 14424 4020 14430 4032
rect 14553 4029 14565 4032
rect 14599 4029 14611 4063
rect 14553 4023 14611 4029
rect 14642 4020 14648 4072
rect 14700 4060 14706 4072
rect 14829 4063 14887 4069
rect 14829 4060 14841 4063
rect 14700 4032 14841 4060
rect 14700 4020 14706 4032
rect 14829 4029 14841 4032
rect 14875 4029 14887 4063
rect 14829 4023 14887 4029
rect 16045 4063 16103 4069
rect 16045 4029 16057 4063
rect 16091 4060 16103 4063
rect 16206 4060 16212 4072
rect 16091 4032 16212 4060
rect 16091 4029 16103 4032
rect 16045 4023 16103 4029
rect 16206 4020 16212 4032
rect 16264 4020 16270 4072
rect 16577 4063 16635 4069
rect 16577 4029 16589 4063
rect 16623 4029 16635 4063
rect 17310 4060 17316 4072
rect 17271 4032 17316 4060
rect 16577 4023 16635 4029
rect 11606 3992 11612 4004
rect 10428 3964 10732 3992
rect 10897 3964 11612 3992
rect 9968 3936 9996 3964
rect 9861 3927 9919 3933
rect 9861 3893 9873 3927
rect 9907 3893 9919 3927
rect 9861 3887 9919 3893
rect 9950 3884 9956 3936
rect 10008 3884 10014 3936
rect 10137 3927 10195 3933
rect 10137 3893 10149 3927
rect 10183 3924 10195 3927
rect 10226 3924 10232 3936
rect 10183 3896 10232 3924
rect 10183 3893 10195 3896
rect 10137 3887 10195 3893
rect 10226 3884 10232 3896
rect 10284 3884 10290 3936
rect 10594 3924 10600 3936
rect 10555 3896 10600 3924
rect 10594 3884 10600 3896
rect 10652 3884 10658 3936
rect 10704 3924 10732 3964
rect 11606 3952 11612 3964
rect 11664 3952 11670 4004
rect 14001 3995 14059 4001
rect 14001 3992 14013 3995
rect 13464 3964 14013 3992
rect 11793 3927 11851 3933
rect 11793 3924 11805 3927
rect 10704 3896 11805 3924
rect 11793 3893 11805 3896
rect 11839 3924 11851 3927
rect 12989 3927 13047 3933
rect 12989 3924 13001 3927
rect 11839 3896 13001 3924
rect 11839 3893 11851 3896
rect 11793 3887 11851 3893
rect 12989 3893 13001 3896
rect 13035 3924 13047 3927
rect 13170 3924 13176 3936
rect 13035 3896 13176 3924
rect 13035 3893 13047 3896
rect 12989 3887 13047 3893
rect 13170 3884 13176 3896
rect 13228 3884 13234 3936
rect 13464 3933 13492 3964
rect 14001 3961 14013 3964
rect 14047 3961 14059 3995
rect 16592 3992 16620 4023
rect 17310 4020 17316 4032
rect 17368 4020 17374 4072
rect 17957 4063 18015 4069
rect 17957 4029 17969 4063
rect 18003 4060 18015 4063
rect 18046 4060 18052 4072
rect 18003 4032 18052 4060
rect 18003 4029 18015 4032
rect 17957 4023 18015 4029
rect 18046 4020 18052 4032
rect 18104 4020 18110 4072
rect 18325 3995 18383 4001
rect 18325 3992 18337 3995
rect 14001 3955 14059 3961
rect 14108 3964 16620 3992
rect 16776 3964 18337 3992
rect 13449 3927 13507 3933
rect 13449 3893 13461 3927
rect 13495 3893 13507 3927
rect 13449 3887 13507 3893
rect 13538 3884 13544 3936
rect 13596 3924 13602 3936
rect 14108 3924 14136 3964
rect 14366 3924 14372 3936
rect 13596 3896 14136 3924
rect 14327 3896 14372 3924
rect 13596 3884 13602 3896
rect 14366 3884 14372 3896
rect 14424 3884 14430 3936
rect 14642 3924 14648 3936
rect 14603 3896 14648 3924
rect 14642 3884 14648 3896
rect 14700 3884 14706 3936
rect 14918 3924 14924 3936
rect 14879 3896 14924 3924
rect 14918 3884 14924 3896
rect 14976 3884 14982 3936
rect 16776 3933 16804 3964
rect 18325 3961 18337 3964
rect 18371 3961 18383 3995
rect 18506 3992 18512 4004
rect 18467 3964 18512 3992
rect 18325 3955 18383 3961
rect 18506 3952 18512 3964
rect 18564 3952 18570 4004
rect 16761 3927 16819 3933
rect 16761 3893 16773 3927
rect 16807 3893 16819 3927
rect 16942 3924 16948 3936
rect 16903 3896 16948 3924
rect 16761 3887 16819 3893
rect 16942 3884 16948 3896
rect 17000 3884 17006 3936
rect 1104 3834 18860 3856
rect 1104 3782 6912 3834
rect 6964 3782 6976 3834
rect 7028 3782 7040 3834
rect 7092 3782 7104 3834
rect 7156 3782 12843 3834
rect 12895 3782 12907 3834
rect 12959 3782 12971 3834
rect 13023 3782 13035 3834
rect 13087 3782 18860 3834
rect 1104 3760 18860 3782
rect 1397 3723 1455 3729
rect 1397 3689 1409 3723
rect 1443 3720 1455 3723
rect 2314 3720 2320 3732
rect 1443 3692 2320 3720
rect 1443 3689 1455 3692
rect 1397 3683 1455 3689
rect 2314 3680 2320 3692
rect 2372 3680 2378 3732
rect 4982 3720 4988 3732
rect 3068 3692 4988 3720
rect 2590 3661 2596 3664
rect 2532 3655 2596 3661
rect 2532 3621 2544 3655
rect 2578 3621 2596 3655
rect 2532 3615 2596 3621
rect 2590 3612 2596 3615
rect 2648 3612 2654 3664
rect 2038 3544 2044 3596
rect 2096 3584 2102 3596
rect 2777 3587 2835 3593
rect 2777 3584 2789 3587
rect 2096 3556 2789 3584
rect 2096 3544 2102 3556
rect 2777 3553 2789 3556
rect 2823 3584 2835 3587
rect 2958 3584 2964 3596
rect 2823 3556 2964 3584
rect 2823 3553 2835 3556
rect 2777 3547 2835 3553
rect 2958 3544 2964 3556
rect 3016 3544 3022 3596
rect 3068 3525 3096 3692
rect 4982 3680 4988 3692
rect 5040 3680 5046 3732
rect 5074 3680 5080 3732
rect 5132 3720 5138 3732
rect 6730 3720 6736 3732
rect 5132 3692 6736 3720
rect 5132 3680 5138 3692
rect 6730 3680 6736 3692
rect 6788 3680 6794 3732
rect 7469 3723 7527 3729
rect 7469 3689 7481 3723
rect 7515 3720 7527 3723
rect 7558 3720 7564 3732
rect 7515 3692 7564 3720
rect 7515 3689 7527 3692
rect 7469 3683 7527 3689
rect 7558 3680 7564 3692
rect 7616 3680 7622 3732
rect 8573 3723 8631 3729
rect 8573 3689 8585 3723
rect 8619 3720 8631 3723
rect 8938 3720 8944 3732
rect 8619 3692 8944 3720
rect 8619 3689 8631 3692
rect 8573 3683 8631 3689
rect 8938 3680 8944 3692
rect 8996 3680 9002 3732
rect 9122 3720 9128 3732
rect 9083 3692 9128 3720
rect 9122 3680 9128 3692
rect 9180 3720 9186 3732
rect 10873 3723 10931 3729
rect 9180 3692 10732 3720
rect 9180 3680 9186 3692
rect 3970 3612 3976 3664
rect 4028 3652 4034 3664
rect 4065 3655 4123 3661
rect 4065 3652 4077 3655
rect 4028 3624 4077 3652
rect 4028 3612 4034 3624
rect 4065 3621 4077 3624
rect 4111 3621 4123 3655
rect 4065 3615 4123 3621
rect 4338 3612 4344 3664
rect 4396 3652 4402 3664
rect 4614 3652 4620 3664
rect 4396 3624 4620 3652
rect 4396 3612 4402 3624
rect 4614 3612 4620 3624
rect 4672 3652 4678 3664
rect 4862 3655 4920 3661
rect 4862 3652 4874 3655
rect 4672 3624 4874 3652
rect 4672 3612 4678 3624
rect 4862 3621 4874 3624
rect 4908 3621 4920 3655
rect 5258 3652 5264 3664
rect 4862 3615 4920 3621
rect 5092 3624 5264 3652
rect 3329 3587 3387 3593
rect 3329 3553 3341 3587
rect 3375 3553 3387 3587
rect 3329 3547 3387 3553
rect 3053 3519 3111 3525
rect 3053 3485 3065 3519
rect 3099 3485 3111 3519
rect 3234 3516 3240 3528
rect 3195 3488 3240 3516
rect 3053 3479 3111 3485
rect 3234 3476 3240 3488
rect 3292 3476 3298 3528
rect 3344 3448 3372 3547
rect 3418 3544 3424 3596
rect 3476 3584 3482 3596
rect 4249 3587 4307 3593
rect 4249 3584 4261 3587
rect 3476 3556 4261 3584
rect 3476 3544 3482 3556
rect 4249 3553 4261 3556
rect 4295 3553 4307 3587
rect 4249 3547 4307 3553
rect 4433 3587 4491 3593
rect 4433 3553 4445 3587
rect 4479 3584 4491 3587
rect 5092 3584 5120 3624
rect 5258 3612 5264 3624
rect 5316 3612 5322 3664
rect 8478 3652 8484 3664
rect 5920 3624 8484 3652
rect 4479 3556 5120 3584
rect 4479 3553 4491 3556
rect 4433 3547 4491 3553
rect 5166 3544 5172 3596
rect 5224 3584 5230 3596
rect 5920 3584 5948 3624
rect 8478 3612 8484 3624
rect 8536 3612 8542 3664
rect 8665 3655 8723 3661
rect 8665 3621 8677 3655
rect 8711 3652 8723 3655
rect 10594 3652 10600 3664
rect 8711 3624 10600 3652
rect 8711 3621 8723 3624
rect 8665 3615 8723 3621
rect 10594 3612 10600 3624
rect 10652 3612 10658 3664
rect 10704 3652 10732 3692
rect 10873 3689 10885 3723
rect 10919 3720 10931 3723
rect 11422 3720 11428 3732
rect 10919 3692 11428 3720
rect 10919 3689 10931 3692
rect 10873 3683 10931 3689
rect 11422 3680 11428 3692
rect 11480 3680 11486 3732
rect 13814 3720 13820 3732
rect 13775 3692 13820 3720
rect 13814 3680 13820 3692
rect 13872 3680 13878 3732
rect 15562 3680 15568 3732
rect 15620 3720 15626 3732
rect 15841 3723 15899 3729
rect 15841 3720 15853 3723
rect 15620 3692 15853 3720
rect 15620 3680 15626 3692
rect 15841 3689 15853 3692
rect 15887 3689 15899 3723
rect 16301 3723 16359 3729
rect 16301 3720 16313 3723
rect 15841 3683 15899 3689
rect 15948 3692 16313 3720
rect 12710 3661 12716 3664
rect 11210 3655 11268 3661
rect 11210 3652 11222 3655
rect 10704 3624 11222 3652
rect 11210 3621 11222 3624
rect 11256 3621 11268 3655
rect 12704 3652 12716 3661
rect 11210 3615 11268 3621
rect 12459 3624 12716 3652
rect 5224 3556 5948 3584
rect 5224 3544 5230 3556
rect 5994 3544 6000 3596
rect 6052 3584 6058 3596
rect 6345 3587 6403 3593
rect 6345 3584 6357 3587
rect 6052 3556 6357 3584
rect 6052 3544 6058 3556
rect 6345 3553 6357 3556
rect 6391 3553 6403 3587
rect 6345 3547 6403 3553
rect 6730 3544 6736 3596
rect 6788 3584 6794 3596
rect 7745 3587 7803 3593
rect 7745 3584 7757 3587
rect 6788 3556 7757 3584
rect 6788 3544 6794 3556
rect 7745 3553 7757 3556
rect 7791 3553 7803 3587
rect 7745 3547 7803 3553
rect 8021 3587 8079 3593
rect 8021 3553 8033 3587
rect 8067 3584 8079 3587
rect 8570 3584 8576 3596
rect 8067 3556 8576 3584
rect 8067 3553 8079 3556
rect 8021 3547 8079 3553
rect 4154 3476 4160 3528
rect 4212 3516 4218 3528
rect 4617 3519 4675 3525
rect 4617 3516 4629 3519
rect 4212 3488 4629 3516
rect 4212 3476 4218 3488
rect 4617 3485 4629 3488
rect 4663 3485 4675 3519
rect 6086 3516 6092 3528
rect 6047 3488 6092 3516
rect 4617 3479 4675 3485
rect 6086 3476 6092 3488
rect 6144 3476 6150 3528
rect 7760 3516 7788 3547
rect 8570 3544 8576 3556
rect 8628 3544 8634 3596
rect 9030 3584 9036 3596
rect 8680 3556 9036 3584
rect 8680 3516 8708 3556
rect 9030 3544 9036 3556
rect 9088 3544 9094 3596
rect 9214 3544 9220 3596
rect 9272 3584 9278 3596
rect 10249 3587 10307 3593
rect 10249 3584 10261 3587
rect 9272 3556 10261 3584
rect 9272 3544 9278 3556
rect 10249 3553 10261 3556
rect 10295 3584 10307 3587
rect 11974 3584 11980 3596
rect 10295 3556 11980 3584
rect 10295 3553 10307 3556
rect 10249 3547 10307 3553
rect 11974 3544 11980 3556
rect 12032 3544 12038 3596
rect 12459 3584 12487 3624
rect 12704 3615 12716 3624
rect 12710 3612 12716 3615
rect 12768 3612 12774 3664
rect 14921 3655 14979 3661
rect 14921 3621 14933 3655
rect 14967 3652 14979 3655
rect 15948 3652 15976 3692
rect 16301 3689 16313 3692
rect 16347 3689 16359 3723
rect 16301 3683 16359 3689
rect 16482 3680 16488 3732
rect 16540 3720 16546 3732
rect 16669 3723 16727 3729
rect 16669 3720 16681 3723
rect 16540 3692 16681 3720
rect 16540 3680 16546 3692
rect 16669 3689 16681 3692
rect 16715 3689 16727 3723
rect 16669 3683 16727 3689
rect 16761 3723 16819 3729
rect 16761 3689 16773 3723
rect 16807 3720 16819 3723
rect 16942 3720 16948 3732
rect 16807 3692 16948 3720
rect 16807 3689 16819 3692
rect 16761 3683 16819 3689
rect 16942 3680 16948 3692
rect 17000 3680 17006 3732
rect 17497 3723 17555 3729
rect 17497 3689 17509 3723
rect 17543 3720 17555 3723
rect 17543 3692 18368 3720
rect 17543 3689 17555 3692
rect 17497 3683 17555 3689
rect 17678 3652 17684 3664
rect 14967 3624 15976 3652
rect 16040 3624 17684 3652
rect 14967 3621 14979 3624
rect 14921 3615 14979 3621
rect 12360 3556 12487 3584
rect 8846 3516 8852 3528
rect 7760 3488 8708 3516
rect 8807 3488 8852 3516
rect 8846 3476 8852 3488
rect 8904 3476 8910 3528
rect 10505 3519 10563 3525
rect 10505 3485 10517 3519
rect 10551 3516 10563 3519
rect 10962 3516 10968 3528
rect 11020 3525 11026 3528
rect 10551 3488 10968 3516
rect 10551 3485 10563 3488
rect 10505 3479 10563 3485
rect 10962 3476 10968 3488
rect 11020 3516 11030 3525
rect 11020 3488 11113 3516
rect 11020 3479 11030 3488
rect 11020 3476 11026 3479
rect 3344 3420 4384 3448
rect 4356 3392 4384 3420
rect 7742 3408 7748 3460
rect 7800 3448 7806 3460
rect 9214 3448 9220 3460
rect 7800 3420 9220 3448
rect 7800 3408 7806 3420
rect 9214 3408 9220 3420
rect 9272 3408 9278 3460
rect 12360 3457 12388 3556
rect 13906 3544 13912 3596
rect 13964 3584 13970 3596
rect 14093 3587 14151 3593
rect 14093 3584 14105 3587
rect 13964 3556 14105 3584
rect 13964 3544 13970 3556
rect 14093 3553 14105 3556
rect 14139 3553 14151 3587
rect 14550 3584 14556 3596
rect 14511 3556 14556 3584
rect 14093 3547 14151 3553
rect 14550 3544 14556 3556
rect 14608 3544 14614 3596
rect 15013 3587 15071 3593
rect 15013 3553 15025 3587
rect 15059 3584 15071 3587
rect 15286 3584 15292 3596
rect 15059 3556 15292 3584
rect 15059 3553 15071 3556
rect 15013 3547 15071 3553
rect 15286 3544 15292 3556
rect 15344 3544 15350 3596
rect 15654 3544 15660 3596
rect 15712 3584 15718 3596
rect 15933 3587 15991 3593
rect 15933 3584 15945 3587
rect 15712 3556 15945 3584
rect 15712 3544 15718 3556
rect 15933 3553 15945 3556
rect 15979 3553 15991 3587
rect 15933 3547 15991 3553
rect 12434 3476 12440 3528
rect 12492 3516 12498 3528
rect 12492 3488 12537 3516
rect 12492 3476 12498 3488
rect 14182 3476 14188 3528
rect 14240 3516 14246 3528
rect 14737 3519 14795 3525
rect 14737 3516 14749 3519
rect 14240 3488 14749 3516
rect 14240 3476 14246 3488
rect 14737 3485 14749 3488
rect 14783 3516 14795 3519
rect 14918 3516 14924 3528
rect 14783 3488 14924 3516
rect 14783 3485 14795 3488
rect 14737 3479 14795 3485
rect 14918 3476 14924 3488
rect 14976 3476 14982 3528
rect 16040 3516 16068 3624
rect 16206 3544 16212 3596
rect 16264 3584 16270 3596
rect 16390 3584 16396 3596
rect 16264 3556 16396 3584
rect 16264 3544 16270 3556
rect 16390 3544 16396 3556
rect 16448 3584 16454 3596
rect 17328 3593 17356 3624
rect 17678 3612 17684 3624
rect 17736 3612 17742 3664
rect 17954 3652 17960 3664
rect 17915 3624 17960 3652
rect 17954 3612 17960 3624
rect 18012 3612 18018 3664
rect 18340 3661 18368 3692
rect 18325 3655 18383 3661
rect 18325 3621 18337 3655
rect 18371 3621 18383 3655
rect 18325 3615 18383 3621
rect 17313 3587 17371 3593
rect 16448 3556 16896 3584
rect 16448 3544 16454 3556
rect 15304 3488 16068 3516
rect 16117 3519 16175 3525
rect 12345 3451 12403 3457
rect 12345 3417 12357 3451
rect 12391 3417 12403 3451
rect 14369 3451 14427 3457
rect 14369 3448 14381 3451
rect 12345 3411 12403 3417
rect 13372 3420 14381 3448
rect 3694 3380 3700 3392
rect 3655 3352 3700 3380
rect 3694 3340 3700 3352
rect 3752 3340 3758 3392
rect 3786 3340 3792 3392
rect 3844 3380 3850 3392
rect 3973 3383 4031 3389
rect 3973 3380 3985 3383
rect 3844 3352 3985 3380
rect 3844 3340 3850 3352
rect 3973 3349 3985 3352
rect 4019 3349 4031 3383
rect 3973 3343 4031 3349
rect 4338 3340 4344 3392
rect 4396 3340 4402 3392
rect 4982 3340 4988 3392
rect 5040 3380 5046 3392
rect 5994 3380 6000 3392
rect 5040 3352 6000 3380
rect 5040 3340 5046 3352
rect 5994 3340 6000 3352
rect 6052 3340 6058 3392
rect 6086 3340 6092 3392
rect 6144 3380 6150 3392
rect 7561 3383 7619 3389
rect 7561 3380 7573 3383
rect 6144 3352 7573 3380
rect 6144 3340 6150 3352
rect 7561 3349 7573 3352
rect 7607 3349 7619 3383
rect 7834 3380 7840 3392
rect 7795 3352 7840 3380
rect 7561 3343 7619 3349
rect 7834 3340 7840 3352
rect 7892 3340 7898 3392
rect 8205 3383 8263 3389
rect 8205 3349 8217 3383
rect 8251 3380 8263 3383
rect 8478 3380 8484 3392
rect 8251 3352 8484 3380
rect 8251 3349 8263 3352
rect 8205 3343 8263 3349
rect 8478 3340 8484 3352
rect 8536 3340 8542 3392
rect 9766 3340 9772 3392
rect 9824 3380 9830 3392
rect 13372 3380 13400 3420
rect 14369 3417 14381 3420
rect 14415 3417 14427 3451
rect 14369 3411 14427 3417
rect 9824 3352 13400 3380
rect 9824 3340 9830 3352
rect 13906 3340 13912 3392
rect 13964 3380 13970 3392
rect 13964 3352 14009 3380
rect 13964 3340 13970 3352
rect 14090 3340 14096 3392
rect 14148 3380 14154 3392
rect 15304 3380 15332 3488
rect 16117 3485 16129 3519
rect 16163 3516 16175 3519
rect 16666 3516 16672 3528
rect 16163 3488 16672 3516
rect 16163 3485 16175 3488
rect 16117 3479 16175 3485
rect 16666 3476 16672 3488
rect 16724 3476 16730 3528
rect 16868 3525 16896 3556
rect 17313 3553 17325 3587
rect 17359 3553 17371 3587
rect 17313 3547 17371 3553
rect 17494 3544 17500 3596
rect 17552 3584 17558 3596
rect 17589 3587 17647 3593
rect 17589 3584 17601 3587
rect 17552 3556 17601 3584
rect 17552 3544 17558 3556
rect 17589 3553 17601 3556
rect 17635 3553 17647 3587
rect 18138 3584 18144 3596
rect 18099 3556 18144 3584
rect 17589 3547 17647 3553
rect 18138 3544 18144 3556
rect 18196 3544 18202 3596
rect 16853 3519 16911 3525
rect 16853 3485 16865 3519
rect 16899 3485 16911 3519
rect 16853 3479 16911 3485
rect 15381 3451 15439 3457
rect 15381 3417 15393 3451
rect 15427 3448 15439 3451
rect 16206 3448 16212 3460
rect 15427 3420 16212 3448
rect 15427 3417 15439 3420
rect 15381 3411 15439 3417
rect 16206 3408 16212 3420
rect 16264 3408 16270 3460
rect 16298 3408 16304 3460
rect 16356 3448 16362 3460
rect 16758 3448 16764 3460
rect 16356 3420 16764 3448
rect 16356 3408 16362 3420
rect 16758 3408 16764 3420
rect 16816 3408 16822 3460
rect 18506 3448 18512 3460
rect 18467 3420 18512 3448
rect 18506 3408 18512 3420
rect 18564 3408 18570 3460
rect 14148 3352 15332 3380
rect 15473 3383 15531 3389
rect 14148 3340 14154 3352
rect 15473 3349 15485 3383
rect 15519 3380 15531 3383
rect 15654 3380 15660 3392
rect 15519 3352 15660 3380
rect 15519 3349 15531 3352
rect 15473 3343 15531 3349
rect 15654 3340 15660 3352
rect 15712 3340 15718 3392
rect 16666 3340 16672 3392
rect 16724 3380 16730 3392
rect 17129 3383 17187 3389
rect 17129 3380 17141 3383
rect 16724 3352 17141 3380
rect 16724 3340 16730 3352
rect 17129 3349 17141 3352
rect 17175 3380 17187 3383
rect 17402 3380 17408 3392
rect 17175 3352 17408 3380
rect 17175 3349 17187 3352
rect 17129 3343 17187 3349
rect 17402 3340 17408 3352
rect 17460 3340 17466 3392
rect 17773 3383 17831 3389
rect 17773 3349 17785 3383
rect 17819 3380 17831 3383
rect 17954 3380 17960 3392
rect 17819 3352 17960 3380
rect 17819 3349 17831 3352
rect 17773 3343 17831 3349
rect 17954 3340 17960 3352
rect 18012 3340 18018 3392
rect 1104 3290 18860 3312
rect 1104 3238 3947 3290
rect 3999 3238 4011 3290
rect 4063 3238 4075 3290
rect 4127 3238 4139 3290
rect 4191 3238 9878 3290
rect 9930 3238 9942 3290
rect 9994 3238 10006 3290
rect 10058 3238 10070 3290
rect 10122 3238 15808 3290
rect 15860 3238 15872 3290
rect 15924 3238 15936 3290
rect 15988 3238 16000 3290
rect 16052 3238 18860 3290
rect 1104 3216 18860 3238
rect 1670 3136 1676 3188
rect 1728 3176 1734 3188
rect 1857 3179 1915 3185
rect 1857 3176 1869 3179
rect 1728 3148 1869 3176
rect 1728 3136 1734 3148
rect 1857 3145 1869 3148
rect 1903 3145 1915 3179
rect 1857 3139 1915 3145
rect 2225 3179 2283 3185
rect 2225 3145 2237 3179
rect 2271 3176 2283 3179
rect 2958 3176 2964 3188
rect 2271 3148 2964 3176
rect 2271 3145 2283 3148
rect 2225 3139 2283 3145
rect 2958 3136 2964 3148
rect 3016 3136 3022 3188
rect 3234 3136 3240 3188
rect 3292 3176 3298 3188
rect 4065 3179 4123 3185
rect 4065 3176 4077 3179
rect 3292 3148 4077 3176
rect 3292 3136 3298 3148
rect 4065 3145 4077 3148
rect 4111 3145 4123 3179
rect 7834 3176 7840 3188
rect 4065 3139 4123 3145
rect 4172 3148 7840 3176
rect 1394 3108 1400 3120
rect 1355 3080 1400 3108
rect 1394 3068 1400 3080
rect 1452 3068 1458 3120
rect 2501 3043 2559 3049
rect 2501 3009 2513 3043
rect 2547 3040 2559 3043
rect 3142 3040 3148 3052
rect 2547 3012 3148 3040
rect 2547 3009 2559 3012
rect 2501 3003 2559 3009
rect 3142 3000 3148 3012
rect 3200 3000 3206 3052
rect 4172 3040 4200 3148
rect 7834 3136 7840 3148
rect 7892 3136 7898 3188
rect 9122 3136 9128 3188
rect 9180 3136 9186 3188
rect 9214 3136 9220 3188
rect 9272 3176 9278 3188
rect 12529 3179 12587 3185
rect 12529 3176 12541 3179
rect 9272 3148 12541 3176
rect 9272 3136 9278 3148
rect 12529 3145 12541 3148
rect 12575 3145 12587 3179
rect 12529 3139 12587 3145
rect 13170 3136 13176 3188
rect 13228 3176 13234 3188
rect 15286 3176 15292 3188
rect 13228 3148 13584 3176
rect 15247 3148 15292 3176
rect 13228 3136 13234 3148
rect 9140 3108 9168 3136
rect 7576 3080 9168 3108
rect 4522 3040 4528 3052
rect 3436 3012 4200 3040
rect 4483 3012 4528 3040
rect 1946 2972 1952 2984
rect 1907 2944 1952 2972
rect 1946 2932 1952 2944
rect 2004 2932 2010 2984
rect 2314 2972 2320 2984
rect 2275 2944 2320 2972
rect 2314 2932 2320 2944
rect 2372 2932 2378 2984
rect 2685 2975 2743 2981
rect 2685 2941 2697 2975
rect 2731 2972 2743 2975
rect 2774 2972 2780 2984
rect 2731 2944 2780 2972
rect 2731 2941 2743 2944
rect 2685 2935 2743 2941
rect 2774 2932 2780 2944
rect 2832 2932 2838 2984
rect 2869 2975 2927 2981
rect 2869 2941 2881 2975
rect 2915 2972 2927 2975
rect 3234 2972 3240 2984
rect 2915 2944 3240 2972
rect 2915 2941 2927 2944
rect 2869 2935 2927 2941
rect 3234 2932 3240 2944
rect 3292 2932 3298 2984
rect 3436 2981 3464 3012
rect 4522 3000 4528 3012
rect 4580 3000 4586 3052
rect 4614 3000 4620 3052
rect 4672 3040 4678 3052
rect 4890 3040 4896 3052
rect 4672 3012 4717 3040
rect 4851 3012 4896 3040
rect 4672 3000 4678 3012
rect 4890 3000 4896 3012
rect 4948 3000 4954 3052
rect 5721 3043 5779 3049
rect 5721 3009 5733 3043
rect 5767 3040 5779 3043
rect 5902 3040 5908 3052
rect 5767 3012 5908 3040
rect 5767 3009 5779 3012
rect 5721 3003 5779 3009
rect 5902 3000 5908 3012
rect 5960 3000 5966 3052
rect 6546 3040 6552 3052
rect 6507 3012 6552 3040
rect 6546 3000 6552 3012
rect 6604 3000 6610 3052
rect 7576 3049 7604 3080
rect 10318 3068 10324 3120
rect 10376 3108 10382 3120
rect 13446 3108 13452 3120
rect 10376 3080 13452 3108
rect 10376 3068 10382 3080
rect 13446 3068 13452 3080
rect 13504 3068 13510 3120
rect 13556 3108 13584 3148
rect 15286 3136 15292 3148
rect 15344 3136 15350 3188
rect 15562 3136 15568 3188
rect 15620 3176 15626 3188
rect 16850 3176 16856 3188
rect 15620 3148 16856 3176
rect 15620 3136 15626 3148
rect 16850 3136 16856 3148
rect 16908 3136 16914 3188
rect 17037 3111 17095 3117
rect 17037 3108 17049 3111
rect 13556 3080 17049 3108
rect 17037 3077 17049 3080
rect 17083 3108 17095 3111
rect 17678 3108 17684 3120
rect 17083 3080 17684 3108
rect 17083 3077 17095 3080
rect 17037 3071 17095 3077
rect 17678 3068 17684 3080
rect 17736 3068 17742 3120
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3009 7619 3043
rect 8294 3040 8300 3052
rect 8255 3012 8300 3040
rect 7561 3003 7619 3009
rect 8294 3000 8300 3012
rect 8352 3000 8358 3052
rect 8478 3040 8484 3052
rect 8439 3012 8484 3040
rect 8478 3000 8484 3012
rect 8536 3000 8542 3052
rect 8846 3000 8852 3052
rect 8904 3040 8910 3052
rect 9585 3043 9643 3049
rect 9585 3040 9597 3043
rect 8904 3012 9597 3040
rect 8904 3000 8910 3012
rect 9585 3009 9597 3012
rect 9631 3009 9643 3043
rect 9585 3003 9643 3009
rect 9674 3000 9680 3052
rect 9732 3040 9738 3052
rect 10505 3043 10563 3049
rect 9732 3012 10456 3040
rect 9732 3000 9738 3012
rect 3421 2975 3479 2981
rect 3421 2941 3433 2975
rect 3467 2941 3479 2975
rect 3421 2935 3479 2941
rect 3789 2975 3847 2981
rect 3789 2941 3801 2975
rect 3835 2972 3847 2975
rect 4246 2972 4252 2984
rect 3835 2944 4252 2972
rect 3835 2941 3847 2944
rect 3789 2935 3847 2941
rect 4246 2932 4252 2944
rect 4304 2932 4310 2984
rect 4430 2972 4436 2984
rect 4391 2944 4436 2972
rect 4430 2932 4436 2944
rect 4488 2932 4494 2984
rect 4798 2972 4804 2984
rect 4540 2944 4804 2972
rect 1581 2907 1639 2913
rect 1581 2873 1593 2907
rect 1627 2904 1639 2907
rect 2222 2904 2228 2916
rect 1627 2876 2228 2904
rect 1627 2873 1639 2876
rect 1581 2867 1639 2873
rect 2222 2864 2228 2876
rect 2280 2864 2286 2916
rect 3053 2907 3111 2913
rect 3053 2873 3065 2907
rect 3099 2904 3111 2907
rect 4540 2904 4568 2944
rect 4798 2932 4804 2944
rect 4856 2932 4862 2984
rect 5534 2932 5540 2984
rect 5592 2972 5598 2984
rect 6181 2975 6239 2981
rect 6181 2972 6193 2975
rect 5592 2944 6193 2972
rect 5592 2932 5598 2944
rect 6181 2941 6193 2944
rect 6227 2941 6239 2975
rect 6730 2972 6736 2984
rect 6691 2944 6736 2972
rect 6181 2935 6239 2941
rect 6730 2932 6736 2944
rect 6788 2932 6794 2984
rect 7101 2975 7159 2981
rect 7101 2941 7113 2975
rect 7147 2972 7159 2975
rect 9766 2972 9772 2984
rect 7147 2944 9772 2972
rect 7147 2941 7159 2944
rect 7101 2935 7159 2941
rect 9766 2932 9772 2944
rect 9824 2932 9830 2984
rect 10428 2972 10456 3012
rect 10505 3009 10517 3043
rect 10551 3040 10563 3043
rect 10686 3040 10692 3052
rect 10551 3012 10692 3040
rect 10551 3009 10563 3012
rect 10505 3003 10563 3009
rect 10686 3000 10692 3012
rect 10744 3040 10750 3052
rect 11241 3043 11299 3049
rect 11241 3040 11253 3043
rect 10744 3012 11253 3040
rect 10744 3000 10750 3012
rect 11241 3009 11253 3012
rect 11287 3009 11299 3043
rect 11790 3040 11796 3052
rect 11241 3003 11299 3009
rect 11348 3012 11796 3040
rect 11348 2972 11376 3012
rect 11790 3000 11796 3012
rect 11848 3000 11854 3052
rect 11974 3000 11980 3052
rect 12032 3040 12038 3052
rect 13081 3043 13139 3049
rect 13081 3040 13093 3043
rect 12032 3012 13093 3040
rect 12032 3000 12038 3012
rect 13081 3009 13093 3012
rect 13127 3009 13139 3043
rect 14642 3040 14648 3052
rect 13081 3003 13139 3009
rect 13648 3012 14648 3040
rect 10428 2944 11376 2972
rect 11422 2932 11428 2984
rect 11480 2972 11486 2984
rect 12069 2975 12127 2981
rect 12069 2972 12081 2975
rect 11480 2944 12081 2972
rect 11480 2932 11486 2944
rect 12069 2941 12081 2944
rect 12115 2941 12127 2975
rect 12069 2935 12127 2941
rect 12158 2932 12164 2984
rect 12216 2972 12222 2984
rect 13354 2972 13360 2984
rect 12216 2944 13360 2972
rect 12216 2932 12222 2944
rect 13354 2932 13360 2944
rect 13412 2932 13418 2984
rect 13648 2981 13676 3012
rect 14642 3000 14648 3012
rect 14700 3000 14706 3052
rect 15470 3000 15476 3052
rect 15528 3040 15534 3052
rect 15749 3043 15807 3049
rect 15749 3040 15761 3043
rect 15528 3012 15761 3040
rect 15528 3000 15534 3012
rect 15749 3009 15761 3012
rect 15795 3009 15807 3043
rect 15749 3003 15807 3009
rect 15933 3043 15991 3049
rect 15933 3009 15945 3043
rect 15979 3040 15991 3043
rect 16390 3040 16396 3052
rect 15979 3012 16396 3040
rect 15979 3009 15991 3012
rect 15933 3003 15991 3009
rect 16390 3000 16396 3012
rect 16448 3000 16454 3052
rect 16482 3000 16488 3052
rect 16540 3040 16546 3052
rect 16540 3012 17264 3040
rect 16540 3000 16546 3012
rect 13633 2975 13691 2981
rect 13633 2941 13645 2975
rect 13679 2941 13691 2975
rect 13633 2935 13691 2941
rect 14093 2975 14151 2981
rect 14093 2941 14105 2975
rect 14139 2972 14151 2975
rect 14274 2972 14280 2984
rect 14139 2944 14280 2972
rect 14139 2941 14151 2944
rect 14093 2935 14151 2941
rect 14274 2932 14280 2944
rect 14332 2932 14338 2984
rect 14369 2975 14427 2981
rect 14369 2941 14381 2975
rect 14415 2972 14427 2975
rect 14458 2972 14464 2984
rect 14415 2944 14464 2972
rect 14415 2941 14427 2944
rect 14369 2935 14427 2941
rect 14458 2932 14464 2944
rect 14516 2932 14522 2984
rect 14737 2975 14795 2981
rect 14737 2941 14749 2975
rect 14783 2972 14795 2975
rect 14826 2972 14832 2984
rect 14783 2944 14832 2972
rect 14783 2941 14795 2944
rect 14737 2935 14795 2941
rect 14826 2932 14832 2944
rect 14884 2932 14890 2984
rect 15105 2975 15163 2981
rect 15105 2941 15117 2975
rect 15151 2972 15163 2975
rect 15378 2972 15384 2984
rect 15151 2944 15384 2972
rect 15151 2941 15163 2944
rect 15105 2935 15163 2941
rect 15378 2932 15384 2944
rect 15436 2932 15442 2984
rect 15654 2972 15660 2984
rect 15615 2944 15660 2972
rect 15654 2932 15660 2944
rect 15712 2932 15718 2984
rect 16206 2932 16212 2984
rect 16264 2972 16270 2984
rect 16301 2975 16359 2981
rect 16301 2972 16313 2975
rect 16264 2944 16313 2972
rect 16264 2932 16270 2944
rect 16301 2941 16313 2944
rect 16347 2941 16359 2975
rect 16666 2972 16672 2984
rect 16301 2935 16359 2941
rect 16408 2944 16672 2972
rect 3099 2876 4568 2904
rect 5445 2907 5503 2913
rect 3099 2873 3111 2876
rect 3053 2867 3111 2873
rect 5445 2873 5457 2907
rect 5491 2904 5503 2907
rect 5905 2907 5963 2913
rect 5905 2904 5917 2907
rect 5491 2876 5917 2904
rect 5491 2873 5503 2876
rect 5445 2867 5503 2873
rect 5905 2873 5917 2876
rect 5951 2873 5963 2907
rect 5905 2867 5963 2873
rect 7285 2907 7343 2913
rect 7285 2873 7297 2907
rect 7331 2904 7343 2907
rect 8478 2904 8484 2916
rect 7331 2876 8484 2904
rect 7331 2873 7343 2876
rect 7285 2867 7343 2873
rect 8478 2864 8484 2876
rect 8536 2864 8542 2916
rect 8573 2907 8631 2913
rect 8573 2873 8585 2907
rect 8619 2904 8631 2907
rect 9401 2907 9459 2913
rect 8619 2876 9076 2904
rect 8619 2873 8631 2876
rect 8573 2867 8631 2873
rect 3326 2836 3332 2848
rect 3287 2808 3332 2836
rect 3326 2796 3332 2808
rect 3384 2796 3390 2848
rect 3694 2836 3700 2848
rect 3655 2808 3700 2836
rect 3694 2796 3700 2808
rect 3752 2796 3758 2848
rect 5074 2836 5080 2848
rect 5035 2808 5080 2836
rect 5074 2796 5080 2808
rect 5132 2796 5138 2848
rect 5537 2839 5595 2845
rect 5537 2805 5549 2839
rect 5583 2836 5595 2839
rect 5626 2836 5632 2848
rect 5583 2808 5632 2836
rect 5583 2805 5595 2808
rect 5537 2799 5595 2805
rect 5626 2796 5632 2808
rect 5684 2796 5690 2848
rect 6825 2839 6883 2845
rect 6825 2805 6837 2839
rect 6871 2836 6883 2839
rect 7466 2836 7472 2848
rect 6871 2808 7472 2836
rect 6871 2805 6883 2808
rect 6825 2799 6883 2805
rect 7466 2796 7472 2808
rect 7524 2796 7530 2848
rect 7650 2836 7656 2848
rect 7611 2808 7656 2836
rect 7650 2796 7656 2808
rect 7708 2796 7714 2848
rect 7742 2796 7748 2848
rect 7800 2836 7806 2848
rect 8113 2839 8171 2845
rect 7800 2808 7845 2836
rect 7800 2796 7806 2808
rect 8113 2805 8125 2839
rect 8159 2836 8171 2839
rect 8662 2836 8668 2848
rect 8159 2808 8668 2836
rect 8159 2805 8171 2808
rect 8113 2799 8171 2805
rect 8662 2796 8668 2808
rect 8720 2796 8726 2848
rect 8846 2796 8852 2848
rect 8904 2836 8910 2848
rect 9048 2845 9076 2876
rect 9401 2873 9413 2907
rect 9447 2904 9459 2907
rect 11057 2907 11115 2913
rect 9447 2876 10732 2904
rect 9447 2873 9459 2876
rect 9401 2867 9459 2873
rect 8941 2839 8999 2845
rect 8941 2836 8953 2839
rect 8904 2808 8953 2836
rect 8904 2796 8910 2808
rect 8941 2805 8953 2808
rect 8987 2805 8999 2839
rect 8941 2799 8999 2805
rect 9033 2839 9091 2845
rect 9033 2805 9045 2839
rect 9079 2805 9091 2839
rect 9033 2799 9091 2805
rect 9493 2839 9551 2845
rect 9493 2805 9505 2839
rect 9539 2836 9551 2839
rect 9861 2839 9919 2845
rect 9861 2836 9873 2839
rect 9539 2808 9873 2836
rect 9539 2805 9551 2808
rect 9493 2799 9551 2805
rect 9861 2805 9873 2808
rect 9907 2805 9919 2839
rect 9861 2799 9919 2805
rect 9950 2796 9956 2848
rect 10008 2836 10014 2848
rect 10229 2839 10287 2845
rect 10229 2836 10241 2839
rect 10008 2808 10241 2836
rect 10008 2796 10014 2808
rect 10229 2805 10241 2808
rect 10275 2805 10287 2839
rect 10229 2799 10287 2805
rect 10321 2839 10379 2845
rect 10321 2805 10333 2839
rect 10367 2836 10379 2839
rect 10410 2836 10416 2848
rect 10367 2808 10416 2836
rect 10367 2805 10379 2808
rect 10321 2799 10379 2805
rect 10410 2796 10416 2808
rect 10468 2796 10474 2848
rect 10704 2845 10732 2876
rect 11057 2873 11069 2907
rect 11103 2904 11115 2907
rect 11514 2904 11520 2916
rect 11103 2876 11520 2904
rect 11103 2873 11115 2876
rect 11057 2867 11115 2873
rect 11514 2864 11520 2876
rect 11572 2864 11578 2916
rect 11882 2864 11888 2916
rect 11940 2904 11946 2916
rect 11977 2907 12035 2913
rect 11977 2904 11989 2907
rect 11940 2876 11989 2904
rect 11940 2864 11946 2876
rect 11977 2873 11989 2876
rect 12023 2873 12035 2907
rect 12897 2907 12955 2913
rect 12897 2904 12909 2907
rect 11977 2867 12035 2873
rect 12452 2876 12909 2904
rect 10689 2839 10747 2845
rect 10689 2805 10701 2839
rect 10735 2805 10747 2839
rect 10689 2799 10747 2805
rect 11149 2839 11207 2845
rect 11149 2805 11161 2839
rect 11195 2836 11207 2839
rect 12066 2836 12072 2848
rect 11195 2808 12072 2836
rect 11195 2805 11207 2808
rect 11149 2799 11207 2805
rect 12066 2796 12072 2808
rect 12124 2796 12130 2848
rect 12452 2845 12480 2876
rect 12897 2873 12909 2876
rect 12943 2873 12955 2907
rect 12897 2867 12955 2873
rect 13817 2907 13875 2913
rect 13817 2873 13829 2907
rect 13863 2904 13875 2907
rect 15470 2904 15476 2916
rect 13863 2876 15476 2904
rect 13863 2873 13875 2876
rect 13817 2867 13875 2873
rect 15470 2864 15476 2876
rect 15528 2864 15534 2916
rect 16022 2904 16028 2916
rect 15856 2876 16028 2904
rect 12437 2839 12495 2845
rect 12437 2805 12449 2839
rect 12483 2805 12495 2839
rect 12437 2799 12495 2805
rect 12618 2796 12624 2848
rect 12676 2836 12682 2848
rect 12989 2839 13047 2845
rect 12989 2836 13001 2839
rect 12676 2808 13001 2836
rect 12676 2796 12682 2808
rect 12989 2805 13001 2808
rect 13035 2805 13047 2839
rect 12989 2799 13047 2805
rect 13449 2839 13507 2845
rect 13449 2805 13461 2839
rect 13495 2836 13507 2839
rect 13630 2836 13636 2848
rect 13495 2808 13636 2836
rect 13495 2805 13507 2808
rect 13449 2799 13507 2805
rect 13630 2796 13636 2808
rect 13688 2796 13694 2848
rect 13906 2836 13912 2848
rect 13867 2808 13912 2836
rect 13906 2796 13912 2808
rect 13964 2796 13970 2848
rect 14185 2839 14243 2845
rect 14185 2805 14197 2839
rect 14231 2836 14243 2839
rect 14274 2836 14280 2848
rect 14231 2808 14280 2836
rect 14231 2805 14243 2808
rect 14185 2799 14243 2805
rect 14274 2796 14280 2808
rect 14332 2796 14338 2848
rect 14550 2836 14556 2848
rect 14511 2808 14556 2836
rect 14550 2796 14556 2808
rect 14608 2796 14614 2848
rect 14918 2836 14924 2848
rect 14879 2808 14924 2836
rect 14918 2796 14924 2808
rect 14976 2796 14982 2848
rect 15194 2796 15200 2848
rect 15252 2836 15258 2848
rect 15562 2836 15568 2848
rect 15252 2808 15568 2836
rect 15252 2796 15258 2808
rect 15562 2796 15568 2808
rect 15620 2836 15626 2848
rect 15856 2836 15884 2876
rect 16022 2864 16028 2876
rect 16080 2864 16086 2916
rect 15620 2808 15884 2836
rect 15620 2796 15626 2808
rect 15930 2796 15936 2848
rect 15988 2836 15994 2848
rect 16117 2839 16175 2845
rect 16117 2836 16129 2839
rect 15988 2808 16129 2836
rect 15988 2796 15994 2808
rect 16117 2805 16129 2808
rect 16163 2805 16175 2839
rect 16117 2799 16175 2805
rect 16206 2796 16212 2848
rect 16264 2836 16270 2848
rect 16408 2845 16436 2944
rect 16666 2932 16672 2944
rect 16724 2932 16730 2984
rect 16761 2975 16819 2981
rect 16761 2941 16773 2975
rect 16807 2972 16819 2975
rect 16850 2972 16856 2984
rect 16807 2944 16856 2972
rect 16807 2941 16819 2944
rect 16761 2935 16819 2941
rect 16850 2932 16856 2944
rect 16908 2932 16914 2984
rect 17236 2981 17264 3012
rect 17221 2975 17279 2981
rect 17221 2941 17233 2975
rect 17267 2941 17279 2975
rect 17586 2972 17592 2984
rect 17547 2944 17592 2972
rect 17221 2935 17279 2941
rect 17586 2932 17592 2944
rect 17644 2932 17650 2984
rect 17954 2972 17960 2984
rect 17915 2944 17960 2972
rect 17954 2932 17960 2944
rect 18012 2932 18018 2984
rect 18322 2972 18328 2984
rect 18283 2944 18328 2972
rect 18322 2932 18328 2944
rect 18380 2932 18386 2984
rect 16482 2864 16488 2916
rect 16540 2904 16546 2916
rect 17773 2907 17831 2913
rect 16540 2876 17080 2904
rect 16540 2864 16546 2876
rect 16393 2839 16451 2845
rect 16393 2836 16405 2839
rect 16264 2808 16405 2836
rect 16264 2796 16270 2808
rect 16393 2805 16405 2808
rect 16439 2805 16451 2839
rect 16574 2836 16580 2848
rect 16535 2808 16580 2836
rect 16393 2799 16451 2805
rect 16574 2796 16580 2808
rect 16632 2796 16638 2848
rect 17052 2836 17080 2876
rect 17773 2873 17785 2907
rect 17819 2904 17831 2907
rect 17862 2904 17868 2916
rect 17819 2876 17868 2904
rect 17819 2873 17831 2876
rect 17773 2867 17831 2873
rect 17862 2864 17868 2876
rect 17920 2864 17926 2916
rect 18138 2904 18144 2916
rect 18099 2876 18144 2904
rect 18138 2864 18144 2876
rect 18196 2864 18202 2916
rect 17313 2839 17371 2845
rect 17313 2836 17325 2839
rect 17052 2808 17325 2836
rect 17313 2805 17325 2808
rect 17359 2805 17371 2839
rect 18414 2836 18420 2848
rect 18375 2808 18420 2836
rect 17313 2799 17371 2805
rect 18414 2796 18420 2808
rect 18472 2796 18478 2848
rect 1104 2746 18860 2768
rect 1104 2694 6912 2746
rect 6964 2694 6976 2746
rect 7028 2694 7040 2746
rect 7092 2694 7104 2746
rect 7156 2694 12843 2746
rect 12895 2694 12907 2746
rect 12959 2694 12971 2746
rect 13023 2694 13035 2746
rect 13087 2694 18860 2746
rect 1104 2672 18860 2694
rect 2593 2635 2651 2641
rect 2593 2601 2605 2635
rect 2639 2632 2651 2635
rect 2866 2632 2872 2644
rect 2639 2604 2872 2632
rect 2639 2601 2651 2604
rect 2593 2595 2651 2601
rect 2866 2592 2872 2604
rect 2924 2592 2930 2644
rect 2961 2635 3019 2641
rect 2961 2601 2973 2635
rect 3007 2632 3019 2635
rect 3050 2632 3056 2644
rect 3007 2604 3056 2632
rect 3007 2601 3019 2604
rect 2961 2595 3019 2601
rect 3050 2592 3056 2604
rect 3108 2592 3114 2644
rect 3436 2604 3740 2632
rect 1949 2567 2007 2573
rect 1949 2533 1961 2567
rect 1995 2564 2007 2567
rect 3436 2564 3464 2604
rect 3602 2564 3608 2576
rect 1995 2536 3464 2564
rect 3563 2536 3608 2564
rect 1995 2533 2007 2536
rect 1949 2527 2007 2533
rect 3602 2524 3608 2536
rect 3660 2524 3666 2576
rect 3712 2564 3740 2604
rect 4338 2592 4344 2644
rect 4396 2632 4402 2644
rect 4433 2635 4491 2641
rect 4433 2632 4445 2635
rect 4396 2604 4445 2632
rect 4396 2592 4402 2604
rect 4433 2601 4445 2604
rect 4479 2601 4491 2635
rect 4433 2595 4491 2601
rect 4801 2635 4859 2641
rect 4801 2601 4813 2635
rect 4847 2632 4859 2635
rect 5074 2632 5080 2644
rect 4847 2604 5080 2632
rect 4847 2601 4859 2604
rect 4801 2595 4859 2601
rect 5074 2592 5080 2604
rect 5132 2592 5138 2644
rect 5721 2635 5779 2641
rect 5721 2601 5733 2635
rect 5767 2632 5779 2635
rect 6546 2632 6552 2644
rect 5767 2604 6552 2632
rect 5767 2601 5779 2604
rect 5721 2595 5779 2601
rect 6546 2592 6552 2604
rect 6604 2592 6610 2644
rect 7469 2635 7527 2641
rect 7469 2601 7481 2635
rect 7515 2632 7527 2635
rect 7650 2632 7656 2644
rect 7515 2604 7656 2632
rect 7515 2601 7527 2604
rect 7469 2595 7527 2601
rect 7650 2592 7656 2604
rect 7708 2592 7714 2644
rect 7837 2635 7895 2641
rect 7837 2601 7849 2635
rect 7883 2632 7895 2635
rect 8297 2635 8355 2641
rect 8297 2632 8309 2635
rect 7883 2604 8309 2632
rect 7883 2601 7895 2604
rect 7837 2595 7895 2601
rect 8297 2601 8309 2604
rect 8343 2601 8355 2635
rect 8297 2595 8355 2601
rect 8662 2592 8668 2644
rect 8720 2592 8726 2644
rect 8757 2635 8815 2641
rect 8757 2601 8769 2635
rect 8803 2632 8815 2635
rect 9030 2632 9036 2644
rect 8803 2604 9036 2632
rect 8803 2601 8815 2604
rect 8757 2595 8815 2601
rect 9030 2592 9036 2604
rect 9088 2592 9094 2644
rect 9309 2635 9367 2641
rect 9309 2601 9321 2635
rect 9355 2632 9367 2635
rect 9582 2632 9588 2644
rect 9355 2604 9588 2632
rect 9355 2601 9367 2604
rect 9309 2595 9367 2601
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 9683 2604 9996 2632
rect 4893 2567 4951 2573
rect 3712 2536 4476 2564
rect 1578 2496 1584 2508
rect 1539 2468 1584 2496
rect 1578 2456 1584 2468
rect 1636 2456 1642 2508
rect 2314 2496 2320 2508
rect 2275 2468 2320 2496
rect 2314 2456 2320 2468
rect 2372 2456 2378 2508
rect 2682 2496 2688 2508
rect 2643 2468 2688 2496
rect 2682 2456 2688 2468
rect 2740 2456 2746 2508
rect 3237 2499 3295 2505
rect 3237 2465 3249 2499
rect 3283 2496 3295 2499
rect 3510 2496 3516 2508
rect 3283 2468 3516 2496
rect 3283 2465 3295 2468
rect 3237 2459 3295 2465
rect 3510 2456 3516 2468
rect 3568 2456 3574 2508
rect 4157 2499 4215 2505
rect 4157 2465 4169 2499
rect 4203 2496 4215 2499
rect 4338 2496 4344 2508
rect 4203 2468 4344 2496
rect 4203 2465 4215 2468
rect 4157 2459 4215 2465
rect 4338 2456 4344 2468
rect 4396 2456 4402 2508
rect 4448 2496 4476 2536
rect 4893 2533 4905 2567
rect 4939 2564 4951 2567
rect 5350 2564 5356 2576
rect 4939 2536 5356 2564
rect 4939 2533 4951 2536
rect 4893 2527 4951 2533
rect 5350 2524 5356 2536
rect 5408 2524 5414 2576
rect 5445 2567 5503 2573
rect 5445 2533 5457 2567
rect 5491 2564 5503 2567
rect 8570 2564 8576 2576
rect 5491 2536 8576 2564
rect 5491 2533 5503 2536
rect 5445 2527 5503 2533
rect 8570 2524 8576 2536
rect 8628 2524 8634 2576
rect 8680 2564 8708 2592
rect 9683 2564 9711 2604
rect 8680 2536 9711 2564
rect 9766 2524 9772 2576
rect 9824 2564 9830 2576
rect 9968 2564 9996 2604
rect 11238 2592 11244 2644
rect 11296 2632 11302 2644
rect 11609 2635 11667 2641
rect 11609 2632 11621 2635
rect 11296 2604 11621 2632
rect 11296 2592 11302 2604
rect 11609 2601 11621 2604
rect 11655 2632 11667 2635
rect 12253 2635 12311 2641
rect 12253 2632 12265 2635
rect 11655 2604 12265 2632
rect 11655 2601 11667 2604
rect 11609 2595 11667 2601
rect 12253 2601 12265 2604
rect 12299 2601 12311 2635
rect 12618 2632 12624 2644
rect 12579 2604 12624 2632
rect 12253 2595 12311 2601
rect 12618 2592 12624 2604
rect 12676 2592 12682 2644
rect 13906 2632 13912 2644
rect 12912 2604 13912 2632
rect 10502 2564 10508 2576
rect 9824 2536 9869 2564
rect 9968 2536 10508 2564
rect 9824 2524 9830 2536
rect 10502 2524 10508 2536
rect 10560 2524 10566 2576
rect 12912 2573 12940 2604
rect 13906 2592 13912 2604
rect 13964 2592 13970 2644
rect 14274 2632 14280 2644
rect 14016 2604 14280 2632
rect 11425 2567 11483 2573
rect 11425 2533 11437 2567
rect 11471 2564 11483 2567
rect 12897 2567 12955 2573
rect 11471 2536 12480 2564
rect 11471 2533 11483 2536
rect 11425 2527 11483 2533
rect 5994 2496 6000 2508
rect 4448 2468 5120 2496
rect 5955 2468 6000 2496
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2428 1823 2431
rect 2774 2428 2780 2440
rect 1811 2400 2780 2428
rect 1811 2397 1823 2400
rect 1765 2391 1823 2397
rect 2774 2388 2780 2400
rect 2832 2388 2838 2440
rect 4706 2388 4712 2440
rect 4764 2428 4770 2440
rect 4985 2431 5043 2437
rect 4985 2428 4997 2431
rect 4764 2400 4997 2428
rect 4764 2388 4770 2400
rect 4985 2397 4997 2400
rect 5031 2397 5043 2431
rect 5092 2428 5120 2468
rect 5994 2456 6000 2468
rect 6052 2456 6058 2508
rect 6362 2496 6368 2508
rect 6323 2468 6368 2496
rect 6362 2456 6368 2468
rect 6420 2456 6426 2508
rect 6917 2499 6975 2505
rect 6917 2465 6929 2499
rect 6963 2465 6975 2499
rect 6917 2459 6975 2465
rect 7193 2499 7251 2505
rect 7193 2465 7205 2499
rect 7239 2496 7251 2499
rect 8202 2496 8208 2508
rect 7239 2468 8208 2496
rect 7239 2465 7251 2468
rect 7193 2459 7251 2465
rect 5092 2400 6224 2428
rect 4985 2391 5043 2397
rect 1210 2320 1216 2372
rect 1268 2360 1274 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 1268 2332 1409 2360
rect 1268 2320 1274 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 2130 2360 2136 2372
rect 2091 2332 2136 2360
rect 1397 2323 1455 2329
rect 2130 2320 2136 2332
rect 2188 2320 2194 2372
rect 3050 2360 3056 2372
rect 3011 2332 3056 2360
rect 3050 2320 3056 2332
rect 3108 2320 3114 2372
rect 3418 2360 3424 2372
rect 3379 2332 3424 2360
rect 3418 2320 3424 2332
rect 3476 2320 3482 2372
rect 3786 2320 3792 2372
rect 3844 2360 3850 2372
rect 3973 2363 4031 2369
rect 3973 2360 3985 2363
rect 3844 2332 3985 2360
rect 3844 2320 3850 2332
rect 3973 2329 3985 2332
rect 4019 2329 4031 2363
rect 5810 2360 5816 2372
rect 5771 2332 5816 2360
rect 3973 2323 4031 2329
rect 5810 2320 5816 2332
rect 5868 2320 5874 2372
rect 6196 2369 6224 2400
rect 6181 2363 6239 2369
rect 6181 2329 6193 2363
rect 6227 2329 6239 2363
rect 6730 2360 6736 2372
rect 6691 2332 6736 2360
rect 6181 2323 6239 2329
rect 6730 2320 6736 2332
rect 6788 2320 6794 2372
rect 4890 2252 4896 2304
rect 4948 2292 4954 2304
rect 5353 2295 5411 2301
rect 5353 2292 5365 2295
rect 4948 2264 5365 2292
rect 4948 2252 4954 2264
rect 5353 2261 5365 2264
rect 5399 2261 5411 2295
rect 5353 2255 5411 2261
rect 5534 2252 5540 2304
rect 5592 2292 5598 2304
rect 6641 2295 6699 2301
rect 6641 2292 6653 2295
rect 5592 2264 6653 2292
rect 5592 2252 5598 2264
rect 6641 2261 6653 2264
rect 6687 2292 6699 2295
rect 6822 2292 6828 2304
rect 6687 2264 6828 2292
rect 6687 2261 6699 2264
rect 6641 2255 6699 2261
rect 6822 2252 6828 2264
rect 6880 2252 6886 2304
rect 6932 2292 6960 2459
rect 8202 2456 8208 2468
rect 8260 2456 8266 2508
rect 8294 2456 8300 2508
rect 8352 2496 8358 2508
rect 8665 2499 8723 2505
rect 8665 2496 8677 2499
rect 8352 2468 8677 2496
rect 8352 2456 8358 2468
rect 8665 2465 8677 2468
rect 8711 2465 8723 2499
rect 9674 2496 9680 2508
rect 8665 2459 8723 2465
rect 9324 2468 9680 2496
rect 7929 2431 7987 2437
rect 7929 2397 7941 2431
rect 7975 2397 7987 2431
rect 8110 2428 8116 2440
rect 8071 2400 8116 2428
rect 7929 2391 7987 2397
rect 7377 2363 7435 2369
rect 7377 2329 7389 2363
rect 7423 2360 7435 2363
rect 7558 2360 7564 2372
rect 7423 2332 7564 2360
rect 7423 2329 7435 2332
rect 7377 2323 7435 2329
rect 7558 2320 7564 2332
rect 7616 2320 7622 2372
rect 7944 2360 7972 2391
rect 8110 2388 8116 2400
rect 8168 2388 8174 2440
rect 8941 2431 8999 2437
rect 8941 2397 8953 2431
rect 8987 2428 8999 2431
rect 9324 2428 9352 2468
rect 9674 2456 9680 2468
rect 9732 2456 9738 2508
rect 9861 2499 9919 2505
rect 9861 2465 9873 2499
rect 9907 2496 9919 2499
rect 10594 2496 10600 2508
rect 9907 2468 10272 2496
rect 10555 2468 10600 2496
rect 9907 2465 9919 2468
rect 9861 2459 9919 2465
rect 8987 2400 9352 2428
rect 8987 2397 8999 2400
rect 8941 2391 8999 2397
rect 9582 2388 9588 2440
rect 9640 2428 9646 2440
rect 9950 2428 9956 2440
rect 9640 2400 9956 2428
rect 9640 2388 9646 2400
rect 9950 2388 9956 2400
rect 10008 2388 10014 2440
rect 10045 2431 10103 2437
rect 10045 2397 10057 2431
rect 10091 2397 10103 2431
rect 10045 2391 10103 2397
rect 9401 2363 9459 2369
rect 9401 2360 9413 2363
rect 7944 2332 9413 2360
rect 9401 2329 9413 2332
rect 9447 2329 9459 2363
rect 9401 2323 9459 2329
rect 9674 2320 9680 2372
rect 9732 2360 9738 2372
rect 10060 2360 10088 2391
rect 10244 2369 10272 2468
rect 10594 2456 10600 2468
rect 10652 2456 10658 2508
rect 12158 2496 12164 2508
rect 12119 2468 12164 2496
rect 12158 2456 12164 2468
rect 12216 2456 12222 2508
rect 10689 2431 10747 2437
rect 10689 2397 10701 2431
rect 10735 2397 10747 2431
rect 10689 2391 10747 2397
rect 9732 2332 10088 2360
rect 10229 2363 10287 2369
rect 9732 2320 9738 2332
rect 10229 2329 10241 2363
rect 10275 2329 10287 2363
rect 10229 2323 10287 2329
rect 9306 2292 9312 2304
rect 6932 2264 9312 2292
rect 9306 2252 9312 2264
rect 9364 2252 9370 2304
rect 10704 2292 10732 2391
rect 10778 2388 10784 2440
rect 10836 2428 10842 2440
rect 10836 2400 10881 2428
rect 10836 2388 10842 2400
rect 11790 2388 11796 2440
rect 11848 2428 11854 2440
rect 11977 2431 12035 2437
rect 11977 2428 11989 2431
rect 11848 2400 11989 2428
rect 11848 2388 11854 2400
rect 11977 2397 11989 2400
rect 12023 2397 12035 2431
rect 12452 2428 12480 2536
rect 12897 2533 12909 2567
rect 12943 2533 12955 2567
rect 12897 2527 12955 2533
rect 13265 2567 13323 2573
rect 13265 2533 13277 2567
rect 13311 2564 13323 2567
rect 14016 2564 14044 2604
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 15102 2592 15108 2644
rect 15160 2632 15166 2644
rect 15289 2635 15347 2641
rect 15289 2632 15301 2635
rect 15160 2604 15301 2632
rect 15160 2592 15166 2604
rect 15289 2601 15301 2604
rect 15335 2632 15347 2635
rect 16301 2635 16359 2641
rect 15335 2604 16252 2632
rect 15335 2601 15347 2604
rect 15289 2595 15347 2601
rect 13311 2536 14044 2564
rect 14093 2567 14151 2573
rect 13311 2533 13323 2536
rect 13265 2527 13323 2533
rect 14093 2533 14105 2567
rect 14139 2564 14151 2567
rect 14550 2564 14556 2576
rect 14139 2536 14556 2564
rect 14139 2533 14151 2536
rect 14093 2527 14151 2533
rect 14550 2524 14556 2536
rect 14608 2524 14614 2576
rect 14918 2524 14924 2576
rect 14976 2564 14982 2576
rect 15013 2567 15071 2573
rect 15013 2564 15025 2567
rect 14976 2536 15025 2564
rect 14976 2524 14982 2536
rect 15013 2533 15025 2536
rect 15059 2533 15071 2567
rect 15930 2564 15936 2576
rect 15891 2536 15936 2564
rect 15013 2527 15071 2533
rect 15930 2524 15936 2536
rect 15988 2524 15994 2576
rect 13446 2496 13452 2508
rect 13407 2468 13452 2496
rect 13446 2456 13452 2468
rect 13504 2456 13510 2508
rect 13633 2499 13691 2505
rect 13633 2465 13645 2499
rect 13679 2496 13691 2499
rect 13722 2496 13728 2508
rect 13679 2468 13728 2496
rect 13679 2465 13691 2468
rect 13633 2459 13691 2465
rect 13722 2456 13728 2468
rect 13780 2456 13786 2508
rect 14734 2496 14740 2508
rect 14695 2468 14740 2496
rect 14734 2456 14740 2468
rect 14792 2456 14798 2508
rect 15473 2499 15531 2505
rect 15473 2465 15485 2499
rect 15519 2465 15531 2499
rect 15473 2459 15531 2465
rect 15488 2428 15516 2459
rect 16022 2456 16028 2508
rect 16080 2496 16086 2508
rect 16117 2499 16175 2505
rect 16117 2496 16129 2499
rect 16080 2468 16129 2496
rect 16080 2456 16086 2468
rect 16117 2465 16129 2468
rect 16163 2465 16175 2499
rect 16224 2496 16252 2604
rect 16301 2601 16313 2635
rect 16347 2632 16359 2635
rect 18141 2635 18199 2641
rect 16347 2604 16528 2632
rect 16347 2601 16359 2604
rect 16301 2595 16359 2601
rect 16500 2573 16528 2604
rect 18141 2601 18153 2635
rect 18187 2601 18199 2635
rect 18141 2595 18199 2601
rect 16485 2567 16543 2573
rect 16485 2533 16497 2567
rect 16531 2533 16543 2567
rect 16850 2564 16856 2576
rect 16811 2536 16856 2564
rect 16485 2527 16543 2533
rect 16850 2524 16856 2536
rect 16908 2524 16914 2576
rect 16942 2524 16948 2576
rect 17000 2564 17006 2576
rect 17313 2567 17371 2573
rect 17313 2564 17325 2567
rect 17000 2536 17325 2564
rect 17000 2524 17006 2536
rect 17313 2533 17325 2536
rect 17359 2533 17371 2567
rect 17770 2564 17776 2576
rect 17731 2536 17776 2564
rect 17313 2527 17371 2533
rect 17770 2524 17776 2536
rect 17828 2524 17834 2576
rect 18156 2564 18184 2595
rect 18325 2567 18383 2573
rect 18325 2564 18337 2567
rect 18156 2536 18337 2564
rect 18325 2533 18337 2536
rect 18371 2533 18383 2567
rect 18325 2527 18383 2533
rect 17494 2496 17500 2508
rect 16224 2468 17500 2496
rect 16117 2459 16175 2465
rect 17494 2456 17500 2468
rect 17552 2456 17558 2508
rect 17678 2456 17684 2508
rect 17736 2496 17742 2508
rect 17957 2499 18015 2505
rect 17957 2496 17969 2499
rect 17736 2468 17969 2496
rect 17736 2456 17742 2468
rect 17957 2465 17969 2468
rect 18003 2465 18015 2499
rect 17957 2459 18015 2465
rect 16574 2428 16580 2440
rect 12452 2400 14596 2428
rect 15488 2400 16580 2428
rect 11977 2391 12035 2397
rect 11238 2360 11244 2372
rect 11199 2332 11244 2360
rect 11238 2320 11244 2332
rect 11296 2320 11302 2372
rect 12250 2320 12256 2372
rect 12308 2360 12314 2372
rect 12713 2363 12771 2369
rect 12713 2360 12725 2363
rect 12308 2332 12725 2360
rect 12308 2320 12314 2332
rect 12713 2329 12725 2332
rect 12759 2329 12771 2363
rect 13078 2360 13084 2372
rect 13039 2332 13084 2360
rect 12713 2323 12771 2329
rect 13078 2320 13084 2332
rect 13136 2320 13142 2372
rect 13906 2360 13912 2372
rect 13867 2332 13912 2360
rect 13906 2320 13912 2332
rect 13964 2320 13970 2372
rect 14568 2369 14596 2400
rect 16574 2388 16580 2400
rect 16632 2388 16638 2440
rect 19426 2428 19432 2440
rect 17328 2400 19432 2428
rect 14553 2363 14611 2369
rect 14553 2329 14565 2363
rect 14599 2329 14611 2363
rect 14826 2360 14832 2372
rect 14787 2332 14832 2360
rect 14553 2323 14611 2329
rect 14826 2320 14832 2332
rect 14884 2320 14890 2372
rect 15654 2320 15660 2372
rect 15712 2360 15718 2372
rect 15749 2363 15807 2369
rect 15749 2360 15761 2363
rect 15712 2332 15761 2360
rect 15712 2320 15718 2332
rect 15749 2329 15761 2332
rect 15795 2329 15807 2363
rect 15749 2323 15807 2329
rect 16669 2363 16727 2369
rect 16669 2329 16681 2363
rect 16715 2360 16727 2363
rect 16850 2360 16856 2372
rect 16715 2332 16856 2360
rect 16715 2329 16727 2332
rect 16669 2323 16727 2329
rect 16850 2320 16856 2332
rect 16908 2320 16914 2372
rect 17034 2360 17040 2372
rect 16995 2332 17040 2360
rect 17034 2320 17040 2332
rect 17092 2320 17098 2372
rect 11146 2292 11152 2304
rect 10704 2264 11152 2292
rect 11146 2252 11152 2264
rect 11204 2252 11210 2304
rect 11330 2252 11336 2304
rect 11388 2292 11394 2304
rect 13814 2292 13820 2304
rect 11388 2264 13820 2292
rect 11388 2252 11394 2264
rect 13814 2252 13820 2264
rect 13872 2252 13878 2304
rect 14090 2252 14096 2304
rect 14148 2292 14154 2304
rect 14274 2292 14280 2304
rect 14148 2264 14280 2292
rect 14148 2252 14154 2264
rect 14274 2252 14280 2264
rect 14332 2252 14338 2304
rect 15565 2295 15623 2301
rect 15565 2261 15577 2295
rect 15611 2292 15623 2295
rect 17328 2292 17356 2400
rect 19426 2388 19432 2400
rect 19484 2388 19490 2440
rect 17586 2360 17592 2372
rect 17547 2332 17592 2360
rect 17586 2320 17592 2332
rect 17644 2320 17650 2372
rect 18506 2360 18512 2372
rect 18467 2332 18512 2360
rect 18506 2320 18512 2332
rect 18564 2320 18570 2372
rect 15611 2264 17356 2292
rect 17405 2295 17463 2301
rect 15611 2261 15623 2264
rect 15565 2255 15623 2261
rect 17405 2261 17417 2295
rect 17451 2292 17463 2295
rect 18414 2292 18420 2304
rect 17451 2264 18420 2292
rect 17451 2261 17463 2264
rect 17405 2255 17463 2261
rect 18414 2252 18420 2264
rect 18472 2252 18478 2304
rect 1104 2202 18860 2224
rect 1104 2150 3947 2202
rect 3999 2150 4011 2202
rect 4063 2150 4075 2202
rect 4127 2150 4139 2202
rect 4191 2150 9878 2202
rect 9930 2150 9942 2202
rect 9994 2150 10006 2202
rect 10058 2150 10070 2202
rect 10122 2150 15808 2202
rect 15860 2150 15872 2202
rect 15924 2150 15936 2202
rect 15988 2150 16000 2202
rect 16052 2150 18860 2202
rect 1104 2128 18860 2150
rect 5994 2048 6000 2100
rect 6052 2088 6058 2100
rect 9490 2088 9496 2100
rect 6052 2060 9496 2088
rect 6052 2048 6058 2060
rect 9490 2048 9496 2060
rect 9548 2048 9554 2100
rect 11146 2048 11152 2100
rect 11204 2088 11210 2100
rect 14458 2088 14464 2100
rect 11204 2060 14464 2088
rect 11204 2048 11210 2060
rect 14458 2048 14464 2060
rect 14516 2088 14522 2100
rect 16206 2088 16212 2100
rect 14516 2060 16212 2088
rect 14516 2048 14522 2060
rect 16206 2048 16212 2060
rect 16264 2048 16270 2100
rect 1578 1980 1584 2032
rect 1636 2020 1642 2032
rect 1636 1992 7604 2020
rect 1636 1980 1642 1992
rect 2314 1912 2320 1964
rect 2372 1952 2378 1964
rect 7576 1952 7604 1992
rect 8202 1980 8208 2032
rect 8260 2020 8266 2032
rect 11330 2020 11336 2032
rect 8260 1992 11336 2020
rect 8260 1980 8266 1992
rect 11330 1980 11336 1992
rect 11388 1980 11394 2032
rect 2372 1924 2774 1952
rect 7576 1924 12434 1952
rect 2372 1912 2378 1924
rect 2746 1680 2774 1924
rect 6638 1844 6644 1896
rect 6696 1884 6702 1896
rect 10594 1884 10600 1896
rect 6696 1856 10600 1884
rect 6696 1844 6702 1856
rect 10594 1844 10600 1856
rect 10652 1844 10658 1896
rect 4338 1776 4344 1828
rect 4396 1816 4402 1828
rect 11054 1816 11060 1828
rect 4396 1788 11060 1816
rect 4396 1776 4402 1788
rect 11054 1776 11060 1788
rect 11112 1776 11118 1828
rect 3510 1708 3516 1760
rect 3568 1748 3574 1760
rect 10226 1748 10232 1760
rect 3568 1720 10232 1748
rect 3568 1708 3574 1720
rect 10226 1708 10232 1720
rect 10284 1708 10290 1760
rect 12406 1748 12434 1924
rect 14182 1748 14188 1760
rect 12406 1720 14188 1748
rect 14182 1708 14188 1720
rect 14240 1708 14246 1760
rect 8386 1680 8392 1692
rect 2746 1652 8392 1680
rect 8386 1640 8392 1652
rect 8444 1640 8450 1692
rect 6822 1572 6828 1624
rect 6880 1612 6886 1624
rect 9766 1612 9772 1624
rect 6880 1584 9772 1612
rect 6880 1572 6886 1584
rect 9766 1572 9772 1584
rect 9824 1612 9830 1624
rect 14274 1612 14280 1624
rect 9824 1584 14280 1612
rect 9824 1572 9830 1584
rect 14274 1572 14280 1584
rect 14332 1572 14338 1624
rect 5902 1504 5908 1556
rect 5960 1544 5966 1556
rect 12158 1544 12164 1556
rect 5960 1516 12164 1544
rect 5960 1504 5966 1516
rect 12158 1504 12164 1516
rect 12216 1504 12222 1556
rect 7466 1368 7472 1420
rect 7524 1408 7530 1420
rect 9398 1408 9404 1420
rect 7524 1380 9404 1408
rect 7524 1368 7530 1380
rect 9398 1368 9404 1380
rect 9456 1368 9462 1420
<< via1 >>
rect 1492 14764 1544 14816
rect 2964 14764 3016 14816
rect 11888 14764 11940 14816
rect 17500 14764 17552 14816
rect 6912 14662 6964 14714
rect 6976 14662 7028 14714
rect 7040 14662 7092 14714
rect 7104 14662 7156 14714
rect 12843 14662 12895 14714
rect 12907 14662 12959 14714
rect 12971 14662 13023 14714
rect 13035 14662 13087 14714
rect 1860 14603 1912 14612
rect 1860 14569 1869 14603
rect 1869 14569 1903 14603
rect 1903 14569 1912 14603
rect 1860 14560 1912 14569
rect 2228 14603 2280 14612
rect 2228 14569 2237 14603
rect 2237 14569 2271 14603
rect 2271 14569 2280 14603
rect 2228 14560 2280 14569
rect 2780 14560 2832 14612
rect 4436 14603 4488 14612
rect 4436 14569 4445 14603
rect 4445 14569 4479 14603
rect 4479 14569 4488 14603
rect 4436 14560 4488 14569
rect 14464 14560 14516 14612
rect 17868 14560 17920 14612
rect 1492 14535 1544 14544
rect 1492 14501 1501 14535
rect 1501 14501 1535 14535
rect 1535 14501 1544 14535
rect 1492 14492 1544 14501
rect 2044 14492 2096 14544
rect 2320 14467 2372 14476
rect 2320 14433 2329 14467
rect 2329 14433 2363 14467
rect 2363 14433 2372 14467
rect 2320 14424 2372 14433
rect 2688 14467 2740 14476
rect 2688 14433 2697 14467
rect 2697 14433 2731 14467
rect 2731 14433 2740 14467
rect 2688 14424 2740 14433
rect 3332 14492 3384 14544
rect 4160 14492 4212 14544
rect 3056 14467 3108 14476
rect 3056 14433 3065 14467
rect 3065 14433 3099 14467
rect 3099 14433 3108 14467
rect 3056 14424 3108 14433
rect 3516 14467 3568 14476
rect 3516 14433 3525 14467
rect 3525 14433 3559 14467
rect 3559 14433 3568 14467
rect 3516 14424 3568 14433
rect 3884 14467 3936 14476
rect 3884 14433 3893 14467
rect 3893 14433 3927 14467
rect 3927 14433 3936 14467
rect 3884 14424 3936 14433
rect 4252 14424 4304 14476
rect 5908 14535 5960 14544
rect 5908 14501 5917 14535
rect 5917 14501 5951 14535
rect 5951 14501 5960 14535
rect 5908 14492 5960 14501
rect 9864 14535 9916 14544
rect 9864 14501 9873 14535
rect 9873 14501 9907 14535
rect 9907 14501 9916 14535
rect 9864 14492 9916 14501
rect 17500 14535 17552 14544
rect 6092 14467 6144 14476
rect 6092 14433 6101 14467
rect 6101 14433 6135 14467
rect 6135 14433 6144 14467
rect 6092 14424 6144 14433
rect 9772 14424 9824 14476
rect 16120 14467 16172 14476
rect 16120 14433 16129 14467
rect 16129 14433 16163 14467
rect 16163 14433 16172 14467
rect 16120 14424 16172 14433
rect 16488 14424 16540 14476
rect 16948 14467 17000 14476
rect 16948 14433 16957 14467
rect 16957 14433 16991 14467
rect 16991 14433 17000 14467
rect 16948 14424 17000 14433
rect 17500 14501 17509 14535
rect 17509 14501 17543 14535
rect 17543 14501 17552 14535
rect 17500 14492 17552 14501
rect 17684 14535 17736 14544
rect 17684 14501 17693 14535
rect 17693 14501 17727 14535
rect 17727 14501 17736 14535
rect 17684 14492 17736 14501
rect 18144 14467 18196 14476
rect 2504 14356 2556 14408
rect 18144 14433 18153 14467
rect 18153 14433 18187 14467
rect 18187 14433 18196 14467
rect 18144 14424 18196 14433
rect 18420 14467 18472 14476
rect 18420 14433 18429 14467
rect 18429 14433 18463 14467
rect 18463 14433 18472 14467
rect 18420 14424 18472 14433
rect 2872 14288 2924 14340
rect 9588 14288 9640 14340
rect 2044 14220 2096 14272
rect 3424 14220 3476 14272
rect 3792 14220 3844 14272
rect 4252 14220 4304 14272
rect 4344 14220 4396 14272
rect 15384 14288 15436 14340
rect 16580 14288 16632 14340
rect 17500 14288 17552 14340
rect 18512 14288 18564 14340
rect 17408 14263 17460 14272
rect 17408 14229 17417 14263
rect 17417 14229 17451 14263
rect 17451 14229 17460 14263
rect 17408 14220 17460 14229
rect 18328 14263 18380 14272
rect 18328 14229 18337 14263
rect 18337 14229 18371 14263
rect 18371 14229 18380 14263
rect 18328 14220 18380 14229
rect 3947 14118 3999 14170
rect 4011 14118 4063 14170
rect 4075 14118 4127 14170
rect 4139 14118 4191 14170
rect 9878 14118 9930 14170
rect 9942 14118 9994 14170
rect 10006 14118 10058 14170
rect 10070 14118 10122 14170
rect 15808 14118 15860 14170
rect 15872 14118 15924 14170
rect 15936 14118 15988 14170
rect 16000 14118 16052 14170
rect 1860 14059 1912 14068
rect 1860 14025 1869 14059
rect 1869 14025 1903 14059
rect 1903 14025 1912 14059
rect 1860 14016 1912 14025
rect 2320 14016 2372 14068
rect 2872 14016 2924 14068
rect 9772 14059 9824 14068
rect 2136 13991 2188 14000
rect 2136 13957 2145 13991
rect 2145 13957 2179 13991
rect 2179 13957 2188 13991
rect 2136 13948 2188 13957
rect 2504 13991 2556 14000
rect 2504 13957 2513 13991
rect 2513 13957 2547 13991
rect 2547 13957 2556 13991
rect 2504 13948 2556 13957
rect 3332 13991 3384 14000
rect 3332 13957 3341 13991
rect 3341 13957 3375 13991
rect 3375 13957 3384 13991
rect 3332 13948 3384 13957
rect 3700 13948 3752 14000
rect 1400 13855 1452 13864
rect 1400 13821 1409 13855
rect 1409 13821 1443 13855
rect 1443 13821 1452 13855
rect 1400 13812 1452 13821
rect 3148 13880 3200 13932
rect 3608 13880 3660 13932
rect 1584 13787 1636 13796
rect 1584 13753 1593 13787
rect 1593 13753 1627 13787
rect 1627 13753 1636 13787
rect 1584 13744 1636 13753
rect 1952 13787 2004 13796
rect 1952 13753 1961 13787
rect 1961 13753 1995 13787
rect 1995 13753 2004 13787
rect 1952 13744 2004 13753
rect 4436 13948 4488 14000
rect 9772 14025 9781 14059
rect 9781 14025 9815 14059
rect 9815 14025 9824 14059
rect 9772 14016 9824 14025
rect 13912 14016 13964 14068
rect 15016 14016 15068 14068
rect 15292 13948 15344 14000
rect 9588 13855 9640 13864
rect 9588 13821 9597 13855
rect 9597 13821 9631 13855
rect 9631 13821 9640 13855
rect 9588 13812 9640 13821
rect 16488 14016 16540 14068
rect 18144 14016 18196 14068
rect 16948 13948 17000 14000
rect 17224 13948 17276 14000
rect 17776 13948 17828 14000
rect 16120 13880 16172 13932
rect 16212 13855 16264 13864
rect 16212 13821 16221 13855
rect 16221 13821 16255 13855
rect 16255 13821 16264 13855
rect 17132 13855 17184 13864
rect 16212 13812 16264 13821
rect 3792 13744 3844 13796
rect 17132 13821 17141 13855
rect 17141 13821 17175 13855
rect 17175 13821 17184 13855
rect 17132 13812 17184 13821
rect 17684 13880 17736 13932
rect 17960 13880 18012 13932
rect 18420 13855 18472 13864
rect 17316 13787 17368 13796
rect 17316 13753 17325 13787
rect 17325 13753 17359 13787
rect 17359 13753 17368 13787
rect 18420 13821 18429 13855
rect 18429 13821 18463 13855
rect 18463 13821 18472 13855
rect 18420 13812 18472 13821
rect 17316 13744 17368 13753
rect 17776 13744 17828 13796
rect 3424 13676 3476 13728
rect 16304 13676 16356 13728
rect 6912 13574 6964 13626
rect 6976 13574 7028 13626
rect 7040 13574 7092 13626
rect 7104 13574 7156 13626
rect 12843 13574 12895 13626
rect 12907 13574 12959 13626
rect 12971 13574 13023 13626
rect 13035 13574 13087 13626
rect 1584 13472 1636 13524
rect 1952 13472 2004 13524
rect 2964 13515 3016 13524
rect 2964 13481 2973 13515
rect 2973 13481 3007 13515
rect 3007 13481 3016 13515
rect 2964 13472 3016 13481
rect 6092 13515 6144 13524
rect 6092 13481 6101 13515
rect 6101 13481 6135 13515
rect 6135 13481 6144 13515
rect 6092 13472 6144 13481
rect 14280 13472 14332 13524
rect 16396 13515 16448 13524
rect 16396 13481 16405 13515
rect 16405 13481 16439 13515
rect 16439 13481 16448 13515
rect 16396 13472 16448 13481
rect 17224 13472 17276 13524
rect 17592 13472 17644 13524
rect 17776 13472 17828 13524
rect 18236 13472 18288 13524
rect 3792 13404 3844 13456
rect 1492 13379 1544 13388
rect 1492 13345 1501 13379
rect 1501 13345 1535 13379
rect 1535 13345 1544 13379
rect 1492 13336 1544 13345
rect 2044 13336 2096 13388
rect 4252 13336 4304 13388
rect 6184 13336 6236 13388
rect 18420 13447 18472 13456
rect 18420 13413 18429 13447
rect 18429 13413 18463 13447
rect 18463 13413 18472 13447
rect 18420 13404 18472 13413
rect 18052 13379 18104 13388
rect 18052 13345 18061 13379
rect 18061 13345 18095 13379
rect 18095 13345 18104 13379
rect 18052 13336 18104 13345
rect 16396 13268 16448 13320
rect 16672 13268 16724 13320
rect 16948 13200 17000 13252
rect 7840 13132 7892 13184
rect 17316 13132 17368 13184
rect 17592 13175 17644 13184
rect 17592 13141 17601 13175
rect 17601 13141 17635 13175
rect 17635 13141 17644 13175
rect 17592 13132 17644 13141
rect 3947 13030 3999 13082
rect 4011 13030 4063 13082
rect 4075 13030 4127 13082
rect 4139 13030 4191 13082
rect 9878 13030 9930 13082
rect 9942 13030 9994 13082
rect 10006 13030 10058 13082
rect 10070 13030 10122 13082
rect 15808 13030 15860 13082
rect 15872 13030 15924 13082
rect 15936 13030 15988 13082
rect 16000 13030 16052 13082
rect 8484 12928 8536 12980
rect 15292 12928 15344 12980
rect 15568 12928 15620 12980
rect 16304 12971 16356 12980
rect 16304 12937 16313 12971
rect 16313 12937 16347 12971
rect 16347 12937 16356 12971
rect 16304 12928 16356 12937
rect 16856 12928 16908 12980
rect 18328 12928 18380 12980
rect 5080 12860 5132 12912
rect 9772 12860 9824 12912
rect 10232 12860 10284 12912
rect 11520 12860 11572 12912
rect 12440 12860 12492 12912
rect 17316 12860 17368 12912
rect 1400 12656 1452 12708
rect 15292 12792 15344 12844
rect 3424 12724 3476 12776
rect 17500 12724 17552 12776
rect 18420 12767 18472 12776
rect 1860 12699 1912 12708
rect 1860 12665 1869 12699
rect 1869 12665 1903 12699
rect 1903 12665 1912 12699
rect 1860 12656 1912 12665
rect 2228 12699 2280 12708
rect 2228 12665 2237 12699
rect 2237 12665 2271 12699
rect 2271 12665 2280 12699
rect 2228 12656 2280 12665
rect 2964 12656 3016 12708
rect 8116 12656 8168 12708
rect 10324 12656 10376 12708
rect 14556 12656 14608 12708
rect 17868 12699 17920 12708
rect 2136 12588 2188 12640
rect 3608 12631 3660 12640
rect 3608 12597 3617 12631
rect 3617 12597 3651 12631
rect 3651 12597 3660 12631
rect 3608 12588 3660 12597
rect 4804 12588 4856 12640
rect 9036 12588 9088 12640
rect 10784 12588 10836 12640
rect 14832 12588 14884 12640
rect 16488 12588 16540 12640
rect 16764 12631 16816 12640
rect 16764 12597 16773 12631
rect 16773 12597 16807 12631
rect 16807 12597 16816 12631
rect 16764 12588 16816 12597
rect 17500 12631 17552 12640
rect 17500 12597 17509 12631
rect 17509 12597 17543 12631
rect 17543 12597 17552 12631
rect 17500 12588 17552 12597
rect 17868 12665 17877 12699
rect 17877 12665 17911 12699
rect 17911 12665 17920 12699
rect 17868 12656 17920 12665
rect 18052 12699 18104 12708
rect 18052 12665 18061 12699
rect 18061 12665 18095 12699
rect 18095 12665 18104 12699
rect 18052 12656 18104 12665
rect 18144 12656 18196 12708
rect 18420 12733 18429 12767
rect 18429 12733 18463 12767
rect 18463 12733 18472 12767
rect 18420 12724 18472 12733
rect 6912 12486 6964 12538
rect 6976 12486 7028 12538
rect 7040 12486 7092 12538
rect 7104 12486 7156 12538
rect 12843 12486 12895 12538
rect 12907 12486 12959 12538
rect 12971 12486 13023 12538
rect 13035 12486 13087 12538
rect 5264 12384 5316 12436
rect 5908 12384 5960 12436
rect 9772 12384 9824 12436
rect 10692 12384 10744 12436
rect 12164 12384 12216 12436
rect 1676 12316 1728 12368
rect 3608 12316 3660 12368
rect 12256 12316 12308 12368
rect 1492 12291 1544 12300
rect 1492 12257 1501 12291
rect 1501 12257 1535 12291
rect 1535 12257 1544 12291
rect 1492 12248 1544 12257
rect 1768 12248 1820 12300
rect 6184 12248 6236 12300
rect 7748 12248 7800 12300
rect 11796 12248 11848 12300
rect 11888 12248 11940 12300
rect 16948 12384 17000 12436
rect 17040 12384 17092 12436
rect 15384 12359 15436 12368
rect 15384 12325 15393 12359
rect 15393 12325 15427 12359
rect 15427 12325 15436 12359
rect 15384 12316 15436 12325
rect 13912 12248 13964 12300
rect 14832 12291 14884 12300
rect 14832 12257 14841 12291
rect 14841 12257 14875 12291
rect 14875 12257 14884 12291
rect 14832 12248 14884 12257
rect 15292 12291 15344 12300
rect 15292 12257 15301 12291
rect 15301 12257 15335 12291
rect 15335 12257 15344 12291
rect 15292 12248 15344 12257
rect 4528 12180 4580 12232
rect 4620 12180 4672 12232
rect 5356 12223 5408 12232
rect 5356 12189 5365 12223
rect 5365 12189 5399 12223
rect 5399 12189 5408 12223
rect 5356 12180 5408 12189
rect 5632 12180 5684 12232
rect 7840 12180 7892 12232
rect 9036 12180 9088 12232
rect 9404 12223 9456 12232
rect 1860 12112 1912 12164
rect 2780 12112 2832 12164
rect 2872 12112 2924 12164
rect 2044 12044 2096 12096
rect 3056 12087 3108 12096
rect 3056 12053 3065 12087
rect 3065 12053 3099 12087
rect 3099 12053 3108 12087
rect 3056 12044 3108 12053
rect 3608 12044 3660 12096
rect 4252 12044 4304 12096
rect 4804 12087 4856 12096
rect 4804 12053 4813 12087
rect 4813 12053 4847 12087
rect 4847 12053 4856 12087
rect 4804 12044 4856 12053
rect 9404 12189 9413 12223
rect 9413 12189 9447 12223
rect 9447 12189 9456 12223
rect 9404 12180 9456 12189
rect 9680 12180 9732 12232
rect 10416 12180 10468 12232
rect 10600 12223 10652 12232
rect 10600 12189 10609 12223
rect 10609 12189 10643 12223
rect 10643 12189 10652 12223
rect 10600 12180 10652 12189
rect 11152 12180 11204 12232
rect 13820 12180 13872 12232
rect 16672 12316 16724 12368
rect 15660 12248 15712 12300
rect 17224 12248 17276 12300
rect 5724 12044 5776 12096
rect 6184 12087 6236 12096
rect 6184 12053 6193 12087
rect 6193 12053 6227 12087
rect 6227 12053 6236 12087
rect 6184 12044 6236 12053
rect 6460 12044 6512 12096
rect 6552 12087 6604 12096
rect 6552 12053 6561 12087
rect 6561 12053 6595 12087
rect 6595 12053 6604 12087
rect 6552 12044 6604 12053
rect 7840 12044 7892 12096
rect 8024 12087 8076 12096
rect 8024 12053 8033 12087
rect 8033 12053 8067 12087
rect 8067 12053 8076 12087
rect 8024 12044 8076 12053
rect 9588 12112 9640 12164
rect 9772 12044 9824 12096
rect 10232 12087 10284 12096
rect 10232 12053 10241 12087
rect 10241 12053 10275 12087
rect 10275 12053 10284 12087
rect 10232 12044 10284 12053
rect 10784 12087 10836 12096
rect 10784 12053 10793 12087
rect 10793 12053 10827 12087
rect 10827 12053 10836 12087
rect 10784 12044 10836 12053
rect 11152 12044 11204 12096
rect 11336 12044 11388 12096
rect 11980 12044 12032 12096
rect 13176 12112 13228 12164
rect 16580 12180 16632 12232
rect 16948 12112 17000 12164
rect 17500 12180 17552 12232
rect 13268 12044 13320 12096
rect 14464 12044 14516 12096
rect 14740 12044 14792 12096
rect 16120 12044 16172 12096
rect 16396 12087 16448 12096
rect 16396 12053 16405 12087
rect 16405 12053 16439 12087
rect 16439 12053 16448 12087
rect 16396 12044 16448 12053
rect 17040 12044 17092 12096
rect 17408 12044 17460 12096
rect 18420 12112 18472 12164
rect 17868 12044 17920 12096
rect 18052 12087 18104 12096
rect 18052 12053 18061 12087
rect 18061 12053 18095 12087
rect 18095 12053 18104 12087
rect 18052 12044 18104 12053
rect 3947 11942 3999 11994
rect 4011 11942 4063 11994
rect 4075 11942 4127 11994
rect 4139 11942 4191 11994
rect 9878 11942 9930 11994
rect 9942 11942 9994 11994
rect 10006 11942 10058 11994
rect 10070 11942 10122 11994
rect 15808 11942 15860 11994
rect 15872 11942 15924 11994
rect 15936 11942 15988 11994
rect 16000 11942 16052 11994
rect 3516 11840 3568 11892
rect 5540 11840 5592 11892
rect 6552 11840 6604 11892
rect 8116 11840 8168 11892
rect 8668 11840 8720 11892
rect 10324 11840 10376 11892
rect 10784 11840 10836 11892
rect 14280 11883 14332 11892
rect 14280 11849 14289 11883
rect 14289 11849 14323 11883
rect 14323 11849 14332 11883
rect 14280 11840 14332 11849
rect 14372 11840 14424 11892
rect 15016 11883 15068 11892
rect 9588 11772 9640 11824
rect 9956 11772 10008 11824
rect 12072 11815 12124 11824
rect 12072 11781 12081 11815
rect 12081 11781 12115 11815
rect 12115 11781 12124 11815
rect 15016 11849 15025 11883
rect 15025 11849 15059 11883
rect 15059 11849 15068 11883
rect 15016 11840 15068 11849
rect 15108 11840 15160 11892
rect 16396 11840 16448 11892
rect 12072 11772 12124 11781
rect 2228 11747 2280 11756
rect 2228 11713 2237 11747
rect 2237 11713 2271 11747
rect 2271 11713 2280 11747
rect 2228 11704 2280 11713
rect 1676 11636 1728 11688
rect 2136 11636 2188 11688
rect 2596 11704 2648 11756
rect 2780 11636 2832 11688
rect 3056 11636 3108 11688
rect 3516 11636 3568 11688
rect 3976 11679 4028 11688
rect 3976 11645 3985 11679
rect 3985 11645 4019 11679
rect 4019 11645 4028 11679
rect 3976 11636 4028 11645
rect 4252 11636 4304 11688
rect 4988 11679 5040 11688
rect 4988 11645 4997 11679
rect 4997 11645 5031 11679
rect 5031 11645 5040 11679
rect 4988 11636 5040 11645
rect 5448 11636 5500 11688
rect 5632 11679 5684 11688
rect 5632 11645 5641 11679
rect 5641 11645 5675 11679
rect 5675 11645 5684 11679
rect 5632 11636 5684 11645
rect 6092 11704 6144 11756
rect 6552 11704 6604 11756
rect 7748 11704 7800 11756
rect 6644 11679 6696 11688
rect 6644 11645 6653 11679
rect 6653 11645 6687 11679
rect 6687 11645 6696 11679
rect 6644 11636 6696 11645
rect 1400 11568 1452 11620
rect 5356 11568 5408 11620
rect 1952 11543 2004 11552
rect 1952 11509 1961 11543
rect 1961 11509 1995 11543
rect 1995 11509 2004 11543
rect 1952 11500 2004 11509
rect 2320 11543 2372 11552
rect 2320 11509 2329 11543
rect 2329 11509 2363 11543
rect 2363 11509 2372 11543
rect 2320 11500 2372 11509
rect 2412 11543 2464 11552
rect 2412 11509 2421 11543
rect 2421 11509 2455 11543
rect 2455 11509 2464 11543
rect 2412 11500 2464 11509
rect 2780 11543 2832 11552
rect 2780 11509 2789 11543
rect 2789 11509 2823 11543
rect 2823 11509 2832 11543
rect 3240 11543 3292 11552
rect 2780 11500 2832 11509
rect 3240 11509 3249 11543
rect 3249 11509 3283 11543
rect 3283 11509 3292 11543
rect 3240 11500 3292 11509
rect 3424 11500 3476 11552
rect 3608 11500 3660 11552
rect 4252 11543 4304 11552
rect 4252 11509 4261 11543
rect 4261 11509 4295 11543
rect 4295 11509 4304 11543
rect 4252 11500 4304 11509
rect 5724 11568 5776 11620
rect 6460 11568 6512 11620
rect 7380 11636 7432 11688
rect 7288 11568 7340 11620
rect 6276 11543 6328 11552
rect 6276 11509 6285 11543
rect 6285 11509 6319 11543
rect 6319 11509 6328 11543
rect 6276 11500 6328 11509
rect 6736 11543 6788 11552
rect 6736 11509 6745 11543
rect 6745 11509 6779 11543
rect 6779 11509 6788 11543
rect 6736 11500 6788 11509
rect 7472 11500 7524 11552
rect 7564 11500 7616 11552
rect 9312 11704 9364 11756
rect 9496 11704 9548 11756
rect 10600 11704 10652 11756
rect 12440 11704 12492 11756
rect 16856 11840 16908 11892
rect 17224 11883 17276 11892
rect 17224 11849 17233 11883
rect 17233 11849 17267 11883
rect 17267 11849 17276 11883
rect 17224 11840 17276 11849
rect 16672 11772 16724 11824
rect 17132 11772 17184 11824
rect 8300 11679 8352 11688
rect 8300 11645 8309 11679
rect 8309 11645 8343 11679
rect 8343 11645 8352 11679
rect 8300 11636 8352 11645
rect 15476 11704 15528 11756
rect 16580 11704 16632 11756
rect 8024 11568 8076 11620
rect 14924 11636 14976 11688
rect 15016 11636 15068 11688
rect 16212 11636 16264 11688
rect 17040 11679 17092 11688
rect 17040 11645 17049 11679
rect 17049 11645 17083 11679
rect 17083 11645 17092 11679
rect 17040 11636 17092 11645
rect 17500 11679 17552 11688
rect 17500 11645 17509 11679
rect 17509 11645 17543 11679
rect 17543 11645 17552 11679
rect 17500 11636 17552 11645
rect 8760 11568 8812 11620
rect 9496 11568 9548 11620
rect 8116 11500 8168 11552
rect 9312 11500 9364 11552
rect 9772 11543 9824 11552
rect 9772 11509 9781 11543
rect 9781 11509 9815 11543
rect 9815 11509 9824 11543
rect 9772 11500 9824 11509
rect 9864 11500 9916 11552
rect 10140 11543 10192 11552
rect 10140 11509 10149 11543
rect 10149 11509 10183 11543
rect 10183 11509 10192 11543
rect 10140 11500 10192 11509
rect 10232 11543 10284 11552
rect 10232 11509 10241 11543
rect 10241 11509 10275 11543
rect 10275 11509 10284 11543
rect 12164 11568 12216 11620
rect 15292 11568 15344 11620
rect 18144 11568 18196 11620
rect 18420 11611 18472 11620
rect 18420 11577 18429 11611
rect 18429 11577 18463 11611
rect 18463 11577 18472 11611
rect 18420 11568 18472 11577
rect 10232 11500 10284 11509
rect 11244 11500 11296 11552
rect 11428 11543 11480 11552
rect 11428 11509 11437 11543
rect 11437 11509 11471 11543
rect 11471 11509 11480 11543
rect 11428 11500 11480 11509
rect 12072 11500 12124 11552
rect 13268 11500 13320 11552
rect 16396 11500 16448 11552
rect 16764 11500 16816 11552
rect 16856 11500 16908 11552
rect 17500 11500 17552 11552
rect 6912 11398 6964 11450
rect 6976 11398 7028 11450
rect 7040 11398 7092 11450
rect 7104 11398 7156 11450
rect 12843 11398 12895 11450
rect 12907 11398 12959 11450
rect 12971 11398 13023 11450
rect 13035 11398 13087 11450
rect 4528 11296 4580 11348
rect 6092 11296 6144 11348
rect 7288 11296 7340 11348
rect 7564 11339 7616 11348
rect 7564 11305 7573 11339
rect 7573 11305 7607 11339
rect 7607 11305 7616 11339
rect 7564 11296 7616 11305
rect 8024 11296 8076 11348
rect 9772 11296 9824 11348
rect 10140 11296 10192 11348
rect 10968 11296 11020 11348
rect 11060 11296 11112 11348
rect 13176 11296 13228 11348
rect 13360 11296 13412 11348
rect 13820 11296 13872 11348
rect 14924 11296 14976 11348
rect 17684 11296 17736 11348
rect 3332 11228 3384 11280
rect 1492 11203 1544 11212
rect 1492 11169 1501 11203
rect 1501 11169 1535 11203
rect 1535 11169 1544 11203
rect 1492 11160 1544 11169
rect 1860 11203 1912 11212
rect 1860 11169 1869 11203
rect 1869 11169 1903 11203
rect 1903 11169 1912 11203
rect 1860 11160 1912 11169
rect 3148 11160 3200 11212
rect 3792 11092 3844 11144
rect 4528 11092 4580 11144
rect 4712 11092 4764 11144
rect 6828 11135 6880 11144
rect 6828 11101 6837 11135
rect 6837 11101 6871 11135
rect 6871 11101 6880 11135
rect 6828 11092 6880 11101
rect 1584 11024 1636 11076
rect 4344 11067 4396 11076
rect 4344 11033 4353 11067
rect 4353 11033 4387 11067
rect 4387 11033 4396 11067
rect 4344 11024 4396 11033
rect 4436 11067 4488 11076
rect 4436 11033 4445 11067
rect 4445 11033 4479 11067
rect 4479 11033 4488 11067
rect 4436 11024 4488 11033
rect 5724 11024 5776 11076
rect 7564 11092 7616 11144
rect 8208 11228 8260 11280
rect 8760 11228 8812 11280
rect 9312 11203 9364 11212
rect 8208 11092 8260 11144
rect 9312 11169 9321 11203
rect 9321 11169 9355 11203
rect 9355 11169 9364 11203
rect 9312 11160 9364 11169
rect 8484 11135 8536 11144
rect 8484 11101 8493 11135
rect 8493 11101 8527 11135
rect 8527 11101 8536 11135
rect 8484 11092 8536 11101
rect 9128 11135 9180 11144
rect 9128 11101 9137 11135
rect 9137 11101 9171 11135
rect 9171 11101 9180 11135
rect 9128 11092 9180 11101
rect 9220 11092 9272 11144
rect 9772 11092 9824 11144
rect 8760 11024 8812 11076
rect 9404 11024 9456 11076
rect 10600 11203 10652 11212
rect 10600 11169 10618 11203
rect 10618 11169 10652 11203
rect 10600 11160 10652 11169
rect 11428 11228 11480 11280
rect 12624 11228 12676 11280
rect 14556 11228 14608 11280
rect 17776 11228 17828 11280
rect 18972 11271 19024 11280
rect 18972 11237 18981 11271
rect 18981 11237 19015 11271
rect 19015 11237 19024 11271
rect 18972 11228 19024 11237
rect 11336 11203 11388 11212
rect 11336 11169 11345 11203
rect 11345 11169 11379 11203
rect 11379 11169 11388 11203
rect 11336 11160 11388 11169
rect 12072 11160 12124 11212
rect 15200 11160 15252 11212
rect 16488 11160 16540 11212
rect 16764 11203 16816 11212
rect 16764 11169 16773 11203
rect 16773 11169 16807 11203
rect 16807 11169 16816 11203
rect 16764 11160 16816 11169
rect 17040 11203 17092 11212
rect 17040 11169 17049 11203
rect 17049 11169 17083 11203
rect 17083 11169 17092 11203
rect 17040 11160 17092 11169
rect 17408 11203 17460 11212
rect 17408 11169 17417 11203
rect 17417 11169 17451 11203
rect 17451 11169 17460 11203
rect 17408 11160 17460 11169
rect 12532 11092 12584 11144
rect 13912 11092 13964 11144
rect 14188 11092 14240 11144
rect 18144 11135 18196 11144
rect 11612 11024 11664 11076
rect 11796 11067 11848 11076
rect 11796 11033 11805 11067
rect 11805 11033 11839 11067
rect 11839 11033 11848 11067
rect 11796 11024 11848 11033
rect 1952 10999 2004 11008
rect 1952 10965 1961 10999
rect 1961 10965 1995 10999
rect 1995 10965 2004 10999
rect 1952 10956 2004 10965
rect 2228 10956 2280 11008
rect 2688 10956 2740 11008
rect 4804 10956 4856 11008
rect 5080 10999 5132 11008
rect 5080 10965 5089 10999
rect 5089 10965 5123 10999
rect 5123 10965 5132 10999
rect 5080 10956 5132 10965
rect 6460 10956 6512 11008
rect 6828 10956 6880 11008
rect 7288 10956 7340 11008
rect 7840 10956 7892 11008
rect 11428 10956 11480 11008
rect 11704 10956 11756 11008
rect 12348 10956 12400 11008
rect 13268 11067 13320 11076
rect 13268 11033 13277 11067
rect 13277 11033 13311 11067
rect 13311 11033 13320 11067
rect 13268 11024 13320 11033
rect 13452 11024 13504 11076
rect 15016 11067 15068 11076
rect 14096 10956 14148 11008
rect 15016 11033 15025 11067
rect 15025 11033 15059 11067
rect 15059 11033 15068 11067
rect 15016 11024 15068 11033
rect 16396 11024 16448 11076
rect 16672 11024 16724 11076
rect 18144 11101 18153 11135
rect 18153 11101 18187 11135
rect 18187 11101 18196 11135
rect 18144 11092 18196 11101
rect 17684 11024 17736 11076
rect 16488 10999 16540 11008
rect 16488 10965 16497 10999
rect 16497 10965 16531 10999
rect 16531 10965 16540 10999
rect 16488 10956 16540 10965
rect 16856 10999 16908 11008
rect 16856 10965 16865 10999
rect 16865 10965 16899 10999
rect 16899 10965 16908 10999
rect 16856 10956 16908 10965
rect 3947 10854 3999 10906
rect 4011 10854 4063 10906
rect 4075 10854 4127 10906
rect 4139 10854 4191 10906
rect 9878 10854 9930 10906
rect 9942 10854 9994 10906
rect 10006 10854 10058 10906
rect 10070 10854 10122 10906
rect 15808 10854 15860 10906
rect 15872 10854 15924 10906
rect 15936 10854 15988 10906
rect 16000 10854 16052 10906
rect 2320 10795 2372 10804
rect 2320 10761 2329 10795
rect 2329 10761 2363 10795
rect 2363 10761 2372 10795
rect 2320 10752 2372 10761
rect 2504 10752 2556 10804
rect 6000 10752 6052 10804
rect 6184 10752 6236 10804
rect 2412 10684 2464 10736
rect 3148 10616 3200 10668
rect 5448 10684 5500 10736
rect 7472 10752 7524 10804
rect 8484 10752 8536 10804
rect 9680 10752 9732 10804
rect 10324 10752 10376 10804
rect 11980 10795 12032 10804
rect 11980 10761 11989 10795
rect 11989 10761 12023 10795
rect 12023 10761 12032 10795
rect 11980 10752 12032 10761
rect 5724 10659 5776 10668
rect 5724 10625 5733 10659
rect 5733 10625 5767 10659
rect 5767 10625 5776 10659
rect 5724 10616 5776 10625
rect 7564 10616 7616 10668
rect 8668 10684 8720 10736
rect 9128 10727 9180 10736
rect 9128 10693 9137 10727
rect 9137 10693 9171 10727
rect 9171 10693 9180 10727
rect 9128 10684 9180 10693
rect 9220 10616 9272 10668
rect 3240 10548 3292 10600
rect 3792 10548 3844 10600
rect 5448 10591 5500 10600
rect 5448 10557 5457 10591
rect 5457 10557 5491 10591
rect 5491 10557 5500 10591
rect 5448 10548 5500 10557
rect 2504 10480 2556 10532
rect 2596 10480 2648 10532
rect 2872 10480 2924 10532
rect 4252 10480 4304 10532
rect 4896 10480 4948 10532
rect 6184 10548 6236 10600
rect 6460 10591 6512 10600
rect 6460 10557 6469 10591
rect 6469 10557 6503 10591
rect 6503 10557 6512 10591
rect 6460 10548 6512 10557
rect 6552 10548 6604 10600
rect 8208 10548 8260 10600
rect 8392 10548 8444 10600
rect 11336 10684 11388 10736
rect 11428 10727 11480 10736
rect 11428 10693 11437 10727
rect 11437 10693 11471 10727
rect 11471 10693 11480 10727
rect 14372 10752 14424 10804
rect 15200 10752 15252 10804
rect 16948 10752 17000 10804
rect 17224 10752 17276 10804
rect 11428 10684 11480 10693
rect 10140 10659 10192 10668
rect 10140 10625 10149 10659
rect 10149 10625 10183 10659
rect 10183 10625 10192 10659
rect 10140 10616 10192 10625
rect 10600 10616 10652 10668
rect 10784 10616 10836 10668
rect 11060 10616 11112 10668
rect 11704 10659 11756 10668
rect 11704 10625 11713 10659
rect 11713 10625 11747 10659
rect 11747 10625 11756 10659
rect 11704 10616 11756 10625
rect 10324 10548 10376 10600
rect 11152 10548 11204 10600
rect 11612 10548 11664 10600
rect 15016 10548 15068 10600
rect 16948 10591 17000 10600
rect 16948 10557 16957 10591
rect 16957 10557 16991 10591
rect 16991 10557 17000 10591
rect 16948 10548 17000 10557
rect 3240 10455 3292 10464
rect 3240 10421 3249 10455
rect 3249 10421 3283 10455
rect 3283 10421 3292 10455
rect 3240 10412 3292 10421
rect 3516 10412 3568 10464
rect 5816 10455 5868 10464
rect 5816 10421 5825 10455
rect 5825 10421 5859 10455
rect 5859 10421 5868 10455
rect 5816 10412 5868 10421
rect 6276 10455 6328 10464
rect 6276 10421 6285 10455
rect 6285 10421 6319 10455
rect 6319 10421 6328 10455
rect 6276 10412 6328 10421
rect 7748 10412 7800 10464
rect 7840 10455 7892 10464
rect 7840 10421 7849 10455
rect 7849 10421 7883 10455
rect 7883 10421 7892 10455
rect 9680 10480 9732 10532
rect 9864 10523 9916 10532
rect 9864 10489 9873 10523
rect 9873 10489 9907 10523
rect 9907 10489 9916 10523
rect 9864 10480 9916 10489
rect 12532 10523 12584 10532
rect 12532 10489 12566 10523
rect 12566 10489 12584 10523
rect 12532 10480 12584 10489
rect 7840 10412 7892 10421
rect 8760 10455 8812 10464
rect 8760 10421 8769 10455
rect 8769 10421 8803 10455
rect 8803 10421 8812 10455
rect 8760 10412 8812 10421
rect 9312 10455 9364 10464
rect 9312 10421 9321 10455
rect 9321 10421 9355 10455
rect 9355 10421 9364 10455
rect 9312 10412 9364 10421
rect 10048 10412 10100 10464
rect 10416 10412 10468 10464
rect 10508 10412 10560 10464
rect 11336 10412 11388 10464
rect 11796 10412 11848 10464
rect 11980 10412 12032 10464
rect 12256 10412 12308 10464
rect 14924 10480 14976 10532
rect 15476 10480 15528 10532
rect 15660 10412 15712 10464
rect 16396 10480 16448 10532
rect 16488 10480 16540 10532
rect 17040 10412 17092 10464
rect 17868 10412 17920 10464
rect 18512 10455 18564 10464
rect 18512 10421 18521 10455
rect 18521 10421 18555 10455
rect 18555 10421 18564 10455
rect 18512 10412 18564 10421
rect 6912 10310 6964 10362
rect 6976 10310 7028 10362
rect 7040 10310 7092 10362
rect 7104 10310 7156 10362
rect 12843 10310 12895 10362
rect 12907 10310 12959 10362
rect 12971 10310 13023 10362
rect 13035 10310 13087 10362
rect 4804 10251 4856 10260
rect 4804 10217 4813 10251
rect 4813 10217 4847 10251
rect 4847 10217 4856 10251
rect 4804 10208 4856 10217
rect 5080 10208 5132 10260
rect 5908 10208 5960 10260
rect 6368 10208 6420 10260
rect 6552 10208 6604 10260
rect 7748 10208 7800 10260
rect 8668 10208 8720 10260
rect 9772 10251 9824 10260
rect 9772 10217 9781 10251
rect 9781 10217 9815 10251
rect 9815 10217 9824 10251
rect 9772 10208 9824 10217
rect 10232 10208 10284 10260
rect 10416 10208 10468 10260
rect 11704 10251 11756 10260
rect 11704 10217 11713 10251
rect 11713 10217 11747 10251
rect 11747 10217 11756 10251
rect 11704 10208 11756 10217
rect 5540 10183 5592 10192
rect 5540 10149 5549 10183
rect 5549 10149 5583 10183
rect 5583 10149 5592 10183
rect 5540 10140 5592 10149
rect 6092 10140 6144 10192
rect 13544 10208 13596 10260
rect 15292 10208 15344 10260
rect 17040 10208 17092 10260
rect 2688 10072 2740 10124
rect 3700 10072 3752 10124
rect 3792 10072 3844 10124
rect 4436 10072 4488 10124
rect 5632 10072 5684 10124
rect 6644 10115 6696 10124
rect 6644 10081 6653 10115
rect 6653 10081 6687 10115
rect 6687 10081 6696 10115
rect 6644 10072 6696 10081
rect 3148 10047 3200 10056
rect 3148 10013 3157 10047
rect 3157 10013 3191 10047
rect 3191 10013 3200 10047
rect 3148 10004 3200 10013
rect 4160 10047 4212 10056
rect 4160 10013 4169 10047
rect 4169 10013 4203 10047
rect 4203 10013 4212 10047
rect 4896 10047 4948 10056
rect 4160 10004 4212 10013
rect 4896 10013 4905 10047
rect 4905 10013 4939 10047
rect 4939 10013 4948 10047
rect 4896 10004 4948 10013
rect 5540 10004 5592 10056
rect 6368 10047 6420 10056
rect 6368 10013 6377 10047
rect 6377 10013 6411 10047
rect 6411 10013 6420 10047
rect 6368 10004 6420 10013
rect 6920 10004 6972 10056
rect 4712 9936 4764 9988
rect 1400 9911 1452 9920
rect 1400 9877 1409 9911
rect 1409 9877 1443 9911
rect 1443 9877 1452 9911
rect 1400 9868 1452 9877
rect 2136 9868 2188 9920
rect 2964 9868 3016 9920
rect 3516 9868 3568 9920
rect 5816 9936 5868 9988
rect 5080 9868 5132 9920
rect 7564 10004 7616 10056
rect 8024 10004 8076 10056
rect 8760 10115 8812 10124
rect 8760 10081 8769 10115
rect 8769 10081 8803 10115
rect 8803 10081 8812 10115
rect 8760 10072 8812 10081
rect 9496 10072 9548 10124
rect 10416 10072 10468 10124
rect 17132 10140 17184 10192
rect 17500 10140 17552 10192
rect 18236 10183 18288 10192
rect 18236 10149 18245 10183
rect 18245 10149 18279 10183
rect 18279 10149 18288 10183
rect 18236 10140 18288 10149
rect 10784 10072 10836 10124
rect 11612 10115 11664 10124
rect 11612 10081 11621 10115
rect 11621 10081 11655 10115
rect 11655 10081 11664 10115
rect 11612 10072 11664 10081
rect 12624 10072 12676 10124
rect 14556 10072 14608 10124
rect 14648 10072 14700 10124
rect 16120 10072 16172 10124
rect 16580 10072 16632 10124
rect 17040 10072 17092 10124
rect 17776 10072 17828 10124
rect 9312 10004 9364 10056
rect 10508 10004 10560 10056
rect 9772 9936 9824 9988
rect 10140 9936 10192 9988
rect 8300 9868 8352 9920
rect 9128 9868 9180 9920
rect 9220 9868 9272 9920
rect 12256 9868 12308 9920
rect 12532 9868 12584 9920
rect 13636 10047 13688 10056
rect 13636 10013 13645 10047
rect 13645 10013 13679 10047
rect 13679 10013 13688 10047
rect 13636 10004 13688 10013
rect 13820 10004 13872 10056
rect 14924 10047 14976 10056
rect 14924 10013 14933 10047
rect 14933 10013 14967 10047
rect 14967 10013 14976 10047
rect 14924 10004 14976 10013
rect 15200 10004 15252 10056
rect 14188 9936 14240 9988
rect 16488 9936 16540 9988
rect 18144 10004 18196 10056
rect 17408 9936 17460 9988
rect 18236 9936 18288 9988
rect 14464 9868 14516 9920
rect 16120 9911 16172 9920
rect 16120 9877 16129 9911
rect 16129 9877 16163 9911
rect 16163 9877 16172 9911
rect 16120 9868 16172 9877
rect 16580 9868 16632 9920
rect 17776 9911 17828 9920
rect 17776 9877 17785 9911
rect 17785 9877 17819 9911
rect 17819 9877 17828 9911
rect 17776 9868 17828 9877
rect 3947 9766 3999 9818
rect 4011 9766 4063 9818
rect 4075 9766 4127 9818
rect 4139 9766 4191 9818
rect 9878 9766 9930 9818
rect 9942 9766 9994 9818
rect 10006 9766 10058 9818
rect 10070 9766 10122 9818
rect 15808 9766 15860 9818
rect 15872 9766 15924 9818
rect 15936 9766 15988 9818
rect 16000 9766 16052 9818
rect 1400 9664 1452 9716
rect 2228 9596 2280 9648
rect 2872 9664 2924 9716
rect 2136 9503 2188 9512
rect 2136 9469 2145 9503
rect 2145 9469 2179 9503
rect 2179 9469 2188 9503
rect 2136 9460 2188 9469
rect 2780 9460 2832 9512
rect 3516 9571 3568 9580
rect 3516 9537 3525 9571
rect 3525 9537 3559 9571
rect 3559 9537 3568 9571
rect 3516 9528 3568 9537
rect 4252 9596 4304 9648
rect 1400 9392 1452 9444
rect 2688 9392 2740 9444
rect 3240 9460 3292 9512
rect 3148 9392 3200 9444
rect 4436 9528 4488 9580
rect 4896 9664 4948 9716
rect 5448 9664 5500 9716
rect 6460 9664 6512 9716
rect 7564 9664 7616 9716
rect 8300 9664 8352 9716
rect 9772 9664 9824 9716
rect 10784 9707 10836 9716
rect 10784 9673 10793 9707
rect 10793 9673 10827 9707
rect 10827 9673 10836 9707
rect 10784 9664 10836 9673
rect 11612 9664 11664 9716
rect 11796 9664 11848 9716
rect 12348 9664 12400 9716
rect 5080 9571 5132 9580
rect 3884 9503 3936 9512
rect 3884 9469 3893 9503
rect 3893 9469 3927 9503
rect 3927 9469 3936 9503
rect 3884 9460 3936 9469
rect 4344 9460 4396 9512
rect 5080 9537 5089 9571
rect 5089 9537 5123 9571
rect 5123 9537 5132 9571
rect 5080 9528 5132 9537
rect 5264 9528 5316 9580
rect 5632 9528 5684 9580
rect 1860 9324 1912 9376
rect 3700 9324 3752 9376
rect 4620 9324 4672 9376
rect 4804 9392 4856 9444
rect 5540 9460 5592 9512
rect 5816 9460 5868 9512
rect 6092 9460 6144 9512
rect 6460 9503 6512 9512
rect 6460 9469 6469 9503
rect 6469 9469 6503 9503
rect 6503 9469 6512 9503
rect 6460 9460 6512 9469
rect 7472 9528 7524 9580
rect 7748 9460 7800 9512
rect 9128 9528 9180 9580
rect 6184 9392 6236 9444
rect 6368 9392 6420 9444
rect 7288 9392 7340 9444
rect 7840 9392 7892 9444
rect 8576 9460 8628 9512
rect 9220 9460 9272 9512
rect 10692 9528 10744 9580
rect 11796 9571 11848 9580
rect 11796 9537 11805 9571
rect 11805 9537 11839 9571
rect 11839 9537 11848 9571
rect 11796 9528 11848 9537
rect 11888 9571 11940 9580
rect 11888 9537 11897 9571
rect 11897 9537 11931 9571
rect 11931 9537 11940 9571
rect 11888 9528 11940 9537
rect 12072 9460 12124 9512
rect 12256 9596 12308 9648
rect 13360 9596 13412 9648
rect 13636 9664 13688 9716
rect 14096 9664 14148 9716
rect 15292 9664 15344 9716
rect 16396 9664 16448 9716
rect 14280 9596 14332 9648
rect 14556 9639 14608 9648
rect 14556 9605 14565 9639
rect 14565 9605 14599 9639
rect 14599 9605 14608 9639
rect 14556 9596 14608 9605
rect 14924 9596 14976 9648
rect 15476 9639 15528 9648
rect 12348 9528 12400 9580
rect 12624 9528 12676 9580
rect 15200 9571 15252 9580
rect 15200 9537 15209 9571
rect 15209 9537 15243 9571
rect 15243 9537 15252 9571
rect 15200 9528 15252 9537
rect 15476 9605 15485 9639
rect 15485 9605 15519 9639
rect 15519 9605 15528 9639
rect 15476 9596 15528 9605
rect 16120 9528 16172 9580
rect 17868 9664 17920 9716
rect 18512 9639 18564 9648
rect 18512 9605 18521 9639
rect 18521 9605 18555 9639
rect 18555 9605 18564 9639
rect 18512 9596 18564 9605
rect 14096 9460 14148 9512
rect 14280 9460 14332 9512
rect 15108 9460 15160 9512
rect 15384 9460 15436 9512
rect 16212 9460 16264 9512
rect 16580 9460 16632 9512
rect 16948 9503 17000 9512
rect 16948 9469 16957 9503
rect 16957 9469 16991 9503
rect 16991 9469 17000 9503
rect 16948 9460 17000 9469
rect 5264 9367 5316 9376
rect 5264 9333 5273 9367
rect 5273 9333 5307 9367
rect 5307 9333 5316 9367
rect 5264 9324 5316 9333
rect 5816 9324 5868 9376
rect 8668 9324 8720 9376
rect 8852 9324 8904 9376
rect 10416 9392 10468 9444
rect 11152 9367 11204 9376
rect 11152 9333 11161 9367
rect 11161 9333 11195 9367
rect 11195 9333 11204 9367
rect 11152 9324 11204 9333
rect 16672 9392 16724 9444
rect 17224 9435 17276 9444
rect 17224 9401 17258 9435
rect 17258 9401 17276 9435
rect 17224 9392 17276 9401
rect 12348 9324 12400 9376
rect 12716 9324 12768 9376
rect 13176 9324 13228 9376
rect 13360 9324 13412 9376
rect 14004 9324 14056 9376
rect 14372 9324 14424 9376
rect 15752 9367 15804 9376
rect 15752 9333 15761 9367
rect 15761 9333 15795 9367
rect 15795 9333 15804 9367
rect 15752 9324 15804 9333
rect 18328 9367 18380 9376
rect 18328 9333 18337 9367
rect 18337 9333 18371 9367
rect 18371 9333 18380 9367
rect 18328 9324 18380 9333
rect 6912 9222 6964 9274
rect 6976 9222 7028 9274
rect 7040 9222 7092 9274
rect 7104 9222 7156 9274
rect 12843 9222 12895 9274
rect 12907 9222 12959 9274
rect 12971 9222 13023 9274
rect 13035 9222 13087 9274
rect 1400 9120 1452 9172
rect 3332 9120 3384 9172
rect 2872 9095 2924 9104
rect 2872 9061 2890 9095
rect 2890 9061 2924 9095
rect 2872 9052 2924 9061
rect 1492 9027 1544 9036
rect 1492 8993 1501 9027
rect 1501 8993 1535 9027
rect 1535 8993 1544 9027
rect 3424 9052 3476 9104
rect 3332 9027 3384 9036
rect 1492 8984 1544 8993
rect 3332 8993 3341 9027
rect 3341 8993 3375 9027
rect 3375 8993 3384 9027
rect 4528 9120 4580 9172
rect 4160 9052 4212 9104
rect 5448 9120 5500 9172
rect 6368 9163 6420 9172
rect 6368 9129 6377 9163
rect 6377 9129 6411 9163
rect 6411 9129 6420 9163
rect 6368 9120 6420 9129
rect 6736 9120 6788 9172
rect 9404 9120 9456 9172
rect 10324 9120 10376 9172
rect 12072 9163 12124 9172
rect 12072 9129 12081 9163
rect 12081 9129 12115 9163
rect 12115 9129 12124 9163
rect 12072 9120 12124 9129
rect 12348 9120 12400 9172
rect 4252 9027 4304 9036
rect 3332 8984 3384 8993
rect 4252 8993 4261 9027
rect 4261 8993 4295 9027
rect 4295 8993 4304 9027
rect 4252 8984 4304 8993
rect 3424 8916 3476 8968
rect 4068 8959 4120 8968
rect 4068 8925 4077 8959
rect 4077 8925 4111 8959
rect 4111 8925 4120 8959
rect 4068 8916 4120 8925
rect 4344 8916 4396 8968
rect 4436 8916 4488 8968
rect 5908 9052 5960 9104
rect 6092 9052 6144 9104
rect 8392 9052 8444 9104
rect 8484 9052 8536 9104
rect 9588 9052 9640 9104
rect 11244 9052 11296 9104
rect 12164 9052 12216 9104
rect 6276 8984 6328 9036
rect 7288 8984 7340 9036
rect 8208 8984 8260 9036
rect 8944 8984 8996 9036
rect 9128 8984 9180 9036
rect 9312 8984 9364 9036
rect 10692 8984 10744 9036
rect 7380 8959 7432 8968
rect 7380 8925 7389 8959
rect 7389 8925 7423 8959
rect 7423 8925 7432 8959
rect 7380 8916 7432 8925
rect 7472 8916 7524 8968
rect 8852 8959 8904 8968
rect 8852 8925 8861 8959
rect 8861 8925 8895 8959
rect 8895 8925 8904 8959
rect 8852 8916 8904 8925
rect 1768 8823 1820 8832
rect 1768 8789 1777 8823
rect 1777 8789 1811 8823
rect 1811 8789 1820 8823
rect 1768 8780 1820 8789
rect 3148 8780 3200 8832
rect 3240 8780 3292 8832
rect 3516 8780 3568 8832
rect 9128 8848 9180 8900
rect 4620 8780 4672 8832
rect 6368 8780 6420 8832
rect 6552 8780 6604 8832
rect 8208 8823 8260 8832
rect 8208 8789 8217 8823
rect 8217 8789 8251 8823
rect 8251 8789 8260 8823
rect 8208 8780 8260 8789
rect 8944 8780 8996 8832
rect 10232 8780 10284 8832
rect 10784 8848 10836 8900
rect 11704 8916 11756 8968
rect 12256 8984 12308 9036
rect 12624 9052 12676 9104
rect 13176 9120 13228 9172
rect 14648 9120 14700 9172
rect 15200 9120 15252 9172
rect 16948 9120 17000 9172
rect 17776 9163 17828 9172
rect 17776 9129 17785 9163
rect 17785 9129 17819 9163
rect 17819 9129 17828 9163
rect 17776 9120 17828 9129
rect 14372 9052 14424 9104
rect 15016 9052 15068 9104
rect 15844 9052 15896 9104
rect 15936 9052 15988 9104
rect 17684 9095 17736 9104
rect 17684 9061 17693 9095
rect 17693 9061 17727 9095
rect 17727 9061 17736 9095
rect 17684 9052 17736 9061
rect 13360 9027 13412 9036
rect 13360 8993 13369 9027
rect 13369 8993 13403 9027
rect 13403 8993 13412 9027
rect 13360 8984 13412 8993
rect 13728 8984 13780 9036
rect 14004 9027 14056 9036
rect 14004 8993 14013 9027
rect 14013 8993 14047 9027
rect 14047 8993 14056 9027
rect 14004 8984 14056 8993
rect 14648 9027 14700 9036
rect 12164 8848 12216 8900
rect 13176 8916 13228 8968
rect 13268 8916 13320 8968
rect 14648 8993 14682 9027
rect 14682 8993 14700 9027
rect 14648 8984 14700 8993
rect 15108 8984 15160 9036
rect 16856 8984 16908 9036
rect 18512 9027 18564 9036
rect 18512 8993 18521 9027
rect 18521 8993 18555 9027
rect 18555 8993 18564 9027
rect 18512 8984 18564 8993
rect 11796 8823 11848 8832
rect 11796 8789 11805 8823
rect 11805 8789 11839 8823
rect 11839 8789 11848 8823
rect 11796 8780 11848 8789
rect 12624 8780 12676 8832
rect 13360 8848 13412 8900
rect 14188 8916 14240 8968
rect 14372 8959 14424 8968
rect 14372 8925 14381 8959
rect 14381 8925 14415 8959
rect 14415 8925 14424 8959
rect 14372 8916 14424 8925
rect 15844 8959 15896 8968
rect 15844 8925 15853 8959
rect 15853 8925 15887 8959
rect 15887 8925 15896 8959
rect 15844 8916 15896 8925
rect 17040 8916 17092 8968
rect 17868 8959 17920 8968
rect 13636 8780 13688 8832
rect 13912 8823 13964 8832
rect 13912 8789 13921 8823
rect 13921 8789 13955 8823
rect 13955 8789 13964 8823
rect 13912 8780 13964 8789
rect 15660 8780 15712 8832
rect 16212 8780 16264 8832
rect 17868 8925 17877 8959
rect 17877 8925 17911 8959
rect 17911 8925 17920 8959
rect 17868 8916 17920 8925
rect 17224 8823 17276 8832
rect 17224 8789 17233 8823
rect 17233 8789 17267 8823
rect 17267 8789 17276 8823
rect 17224 8780 17276 8789
rect 17500 8780 17552 8832
rect 17868 8780 17920 8832
rect 3947 8678 3999 8730
rect 4011 8678 4063 8730
rect 4075 8678 4127 8730
rect 4139 8678 4191 8730
rect 9878 8678 9930 8730
rect 9942 8678 9994 8730
rect 10006 8678 10058 8730
rect 10070 8678 10122 8730
rect 15808 8678 15860 8730
rect 15872 8678 15924 8730
rect 15936 8678 15988 8730
rect 16000 8678 16052 8730
rect 2688 8576 2740 8628
rect 3700 8576 3752 8628
rect 5908 8508 5960 8560
rect 10416 8576 10468 8628
rect 10508 8576 10560 8628
rect 1768 8372 1820 8424
rect 2596 8415 2648 8424
rect 2596 8381 2614 8415
rect 2614 8381 2648 8415
rect 2596 8372 2648 8381
rect 4436 8415 4488 8424
rect 4436 8381 4445 8415
rect 4445 8381 4479 8415
rect 4479 8381 4488 8415
rect 4436 8372 4488 8381
rect 5080 8372 5132 8424
rect 2688 8304 2740 8356
rect 2780 8304 2832 8356
rect 3608 8304 3660 8356
rect 3792 8304 3844 8356
rect 8300 8508 8352 8560
rect 9496 8508 9548 8560
rect 10324 8508 10376 8560
rect 12164 8551 12216 8560
rect 12164 8517 12173 8551
rect 12173 8517 12207 8551
rect 12207 8517 12216 8551
rect 12164 8508 12216 8517
rect 10508 8440 10560 8492
rect 11612 8440 11664 8492
rect 11704 8440 11756 8492
rect 12532 8508 12584 8560
rect 13176 8551 13228 8560
rect 13176 8517 13185 8551
rect 13185 8517 13219 8551
rect 13219 8517 13228 8551
rect 13176 8508 13228 8517
rect 13268 8508 13320 8560
rect 14832 8508 14884 8560
rect 12624 8483 12676 8492
rect 12624 8449 12633 8483
rect 12633 8449 12667 8483
rect 12667 8449 12676 8483
rect 12624 8440 12676 8449
rect 13728 8440 13780 8492
rect 14648 8483 14700 8492
rect 14648 8449 14657 8483
rect 14657 8449 14691 8483
rect 14691 8449 14700 8483
rect 14648 8440 14700 8449
rect 15292 8483 15344 8492
rect 15292 8449 15301 8483
rect 15301 8449 15335 8483
rect 15335 8449 15344 8483
rect 15292 8440 15344 8449
rect 8760 8372 8812 8424
rect 8852 8372 8904 8424
rect 9312 8372 9364 8424
rect 9496 8372 9548 8424
rect 10692 8372 10744 8424
rect 11796 8372 11848 8424
rect 12348 8372 12400 8424
rect 12716 8415 12768 8424
rect 12716 8381 12725 8415
rect 12725 8381 12759 8415
rect 12759 8381 12768 8415
rect 12716 8372 12768 8381
rect 13452 8372 13504 8424
rect 6552 8304 6604 8356
rect 2044 8236 2096 8288
rect 4068 8236 4120 8288
rect 4160 8236 4212 8288
rect 5356 8236 5408 8288
rect 5724 8236 5776 8288
rect 6092 8236 6144 8288
rect 7380 8304 7432 8356
rect 7840 8236 7892 8288
rect 8300 8304 8352 8356
rect 10232 8304 10284 8356
rect 11888 8347 11940 8356
rect 11888 8313 11897 8347
rect 11897 8313 11931 8347
rect 11931 8313 11940 8347
rect 11888 8304 11940 8313
rect 12164 8304 12216 8356
rect 15108 8415 15160 8424
rect 9312 8236 9364 8288
rect 9680 8236 9732 8288
rect 10784 8236 10836 8288
rect 13820 8304 13872 8356
rect 14004 8304 14056 8356
rect 14280 8304 14332 8356
rect 14556 8236 14608 8288
rect 15108 8381 15117 8415
rect 15117 8381 15151 8415
rect 15151 8381 15160 8415
rect 15108 8372 15160 8381
rect 14924 8304 14976 8356
rect 16028 8483 16080 8492
rect 16028 8449 16037 8483
rect 16037 8449 16071 8483
rect 16071 8449 16080 8483
rect 16028 8440 16080 8449
rect 15936 8372 15988 8424
rect 17500 8576 17552 8628
rect 16672 8508 16724 8560
rect 17040 8508 17092 8560
rect 17224 8440 17276 8492
rect 16488 8372 16540 8424
rect 15660 8304 15712 8356
rect 18604 8372 18656 8424
rect 16948 8304 17000 8356
rect 17960 8347 18012 8356
rect 17960 8313 17969 8347
rect 17969 8313 18003 8347
rect 18003 8313 18012 8347
rect 17960 8304 18012 8313
rect 18144 8347 18196 8356
rect 18144 8313 18153 8347
rect 18153 8313 18187 8347
rect 18187 8313 18196 8347
rect 18144 8304 18196 8313
rect 17224 8236 17276 8288
rect 17408 8236 17460 8288
rect 6912 8134 6964 8186
rect 6976 8134 7028 8186
rect 7040 8134 7092 8186
rect 7104 8134 7156 8186
rect 12843 8134 12895 8186
rect 12907 8134 12959 8186
rect 12971 8134 13023 8186
rect 13035 8134 13087 8186
rect 3516 8032 3568 8084
rect 4068 8032 4120 8084
rect 5172 8032 5224 8084
rect 5264 8032 5316 8084
rect 5816 8032 5868 8084
rect 6092 8075 6144 8084
rect 6092 8041 6101 8075
rect 6101 8041 6135 8075
rect 6135 8041 6144 8075
rect 6092 8032 6144 8041
rect 7564 8032 7616 8084
rect 8392 8075 8444 8084
rect 8392 8041 8401 8075
rect 8401 8041 8435 8075
rect 8435 8041 8444 8075
rect 8392 8032 8444 8041
rect 8944 8075 8996 8084
rect 8944 8041 8953 8075
rect 8953 8041 8987 8075
rect 8987 8041 8996 8075
rect 8944 8032 8996 8041
rect 1492 8007 1544 8016
rect 1492 7973 1501 8007
rect 1501 7973 1535 8007
rect 1535 7973 1544 8007
rect 1492 7964 1544 7973
rect 3700 7964 3752 8016
rect 2688 7896 2740 7948
rect 2320 7871 2372 7880
rect 2320 7837 2329 7871
rect 2329 7837 2363 7871
rect 2363 7837 2372 7871
rect 2320 7828 2372 7837
rect 3148 7871 3200 7880
rect 1676 7803 1728 7812
rect 1676 7769 1685 7803
rect 1685 7769 1719 7803
rect 1719 7769 1728 7803
rect 1676 7760 1728 7769
rect 3148 7837 3157 7871
rect 3157 7837 3191 7871
rect 3191 7837 3200 7871
rect 3148 7828 3200 7837
rect 3608 7896 3660 7948
rect 3976 7896 4028 7948
rect 2596 7760 2648 7812
rect 4160 7828 4212 7880
rect 2044 7692 2096 7744
rect 2136 7692 2188 7744
rect 3700 7735 3752 7744
rect 3700 7701 3709 7735
rect 3709 7701 3743 7735
rect 3743 7701 3752 7735
rect 3700 7692 3752 7701
rect 3792 7692 3844 7744
rect 5908 7964 5960 8016
rect 6000 7896 6052 7948
rect 5080 7828 5132 7880
rect 5632 7828 5684 7880
rect 6460 7828 6512 7880
rect 6276 7760 6328 7812
rect 4896 7692 4948 7744
rect 6000 7735 6052 7744
rect 6000 7701 6009 7735
rect 6009 7701 6043 7735
rect 6043 7701 6052 7735
rect 6000 7692 6052 7701
rect 6552 7692 6604 7744
rect 7748 7964 7800 8016
rect 8852 7964 8904 8016
rect 12532 8032 12584 8084
rect 13728 8075 13780 8084
rect 13728 8041 13737 8075
rect 13737 8041 13771 8075
rect 13771 8041 13780 8075
rect 13728 8032 13780 8041
rect 14372 8032 14424 8084
rect 16212 8032 16264 8084
rect 8116 7896 8168 7948
rect 7748 7828 7800 7880
rect 7932 7828 7984 7880
rect 9864 7828 9916 7880
rect 7840 7760 7892 7812
rect 7564 7692 7616 7744
rect 9588 7760 9640 7812
rect 8024 7692 8076 7744
rect 9680 7692 9732 7744
rect 11520 7896 11572 7948
rect 11796 7871 11848 7880
rect 10600 7760 10652 7812
rect 11152 7760 11204 7812
rect 11796 7837 11805 7871
rect 11805 7837 11839 7871
rect 11839 7837 11848 7871
rect 11796 7828 11848 7837
rect 12900 7896 12952 7948
rect 17960 7964 18012 8016
rect 13820 7939 13872 7948
rect 12072 7828 12124 7880
rect 13820 7905 13829 7939
rect 13829 7905 13863 7939
rect 13863 7905 13872 7939
rect 13820 7896 13872 7905
rect 13912 7896 13964 7948
rect 15292 7896 15344 7948
rect 16304 7939 16356 7948
rect 16304 7905 16313 7939
rect 16313 7905 16347 7939
rect 16347 7905 16356 7939
rect 16304 7896 16356 7905
rect 16672 7896 16724 7948
rect 17776 7896 17828 7948
rect 16212 7871 16264 7880
rect 16212 7837 16221 7871
rect 16221 7837 16255 7871
rect 16255 7837 16264 7871
rect 16212 7828 16264 7837
rect 17684 7828 17736 7880
rect 11336 7692 11388 7744
rect 14280 7692 14332 7744
rect 14740 7692 14792 7744
rect 16856 7735 16908 7744
rect 16856 7701 16865 7735
rect 16865 7701 16899 7735
rect 16899 7701 16908 7735
rect 16856 7692 16908 7701
rect 16948 7692 17000 7744
rect 3947 7590 3999 7642
rect 4011 7590 4063 7642
rect 4075 7590 4127 7642
rect 4139 7590 4191 7642
rect 9878 7590 9930 7642
rect 9942 7590 9994 7642
rect 10006 7590 10058 7642
rect 10070 7590 10122 7642
rect 15808 7590 15860 7642
rect 15872 7590 15924 7642
rect 15936 7590 15988 7642
rect 16000 7590 16052 7642
rect 1952 7488 2004 7540
rect 3148 7488 3200 7540
rect 4252 7488 4304 7540
rect 4804 7531 4856 7540
rect 4804 7497 4813 7531
rect 4813 7497 4847 7531
rect 4847 7497 4856 7531
rect 4804 7488 4856 7497
rect 5816 7488 5868 7540
rect 8484 7488 8536 7540
rect 11888 7488 11940 7540
rect 16672 7531 16724 7540
rect 16672 7497 16681 7531
rect 16681 7497 16715 7531
rect 16715 7497 16724 7531
rect 16672 7488 16724 7497
rect 17776 7531 17828 7540
rect 17776 7497 17785 7531
rect 17785 7497 17819 7531
rect 17819 7497 17828 7531
rect 17776 7488 17828 7497
rect 2504 7420 2556 7472
rect 6184 7420 6236 7472
rect 2780 7352 2832 7404
rect 3148 7395 3200 7404
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 3608 7395 3660 7404
rect 3608 7361 3617 7395
rect 3617 7361 3651 7395
rect 3651 7361 3660 7395
rect 3608 7352 3660 7361
rect 3792 7352 3844 7404
rect 3976 7352 4028 7404
rect 6276 7352 6328 7404
rect 7840 7352 7892 7404
rect 8208 7352 8260 7404
rect 1400 7327 1452 7336
rect 1400 7293 1409 7327
rect 1409 7293 1443 7327
rect 1443 7293 1452 7327
rect 1400 7284 1452 7293
rect 2044 7327 2096 7336
rect 2044 7293 2053 7327
rect 2053 7293 2087 7327
rect 2087 7293 2096 7327
rect 2044 7284 2096 7293
rect 2136 7327 2188 7336
rect 2136 7293 2145 7327
rect 2145 7293 2179 7327
rect 2179 7293 2188 7327
rect 2136 7284 2188 7293
rect 4068 7284 4120 7336
rect 4160 7284 4212 7336
rect 4988 7284 5040 7336
rect 4344 7216 4396 7268
rect 4896 7216 4948 7268
rect 5448 7216 5500 7268
rect 5540 7216 5592 7268
rect 6460 7284 6512 7336
rect 7380 7284 7432 7336
rect 7564 7284 7616 7336
rect 8668 7352 8720 7404
rect 9680 7420 9732 7472
rect 11428 7420 11480 7472
rect 12900 7420 12952 7472
rect 13544 7420 13596 7472
rect 17684 7463 17736 7472
rect 17684 7429 17693 7463
rect 17693 7429 17727 7463
rect 17727 7429 17736 7463
rect 17684 7420 17736 7429
rect 9312 7352 9364 7404
rect 10416 7395 10468 7404
rect 10416 7361 10425 7395
rect 10425 7361 10459 7395
rect 10459 7361 10468 7395
rect 10416 7352 10468 7361
rect 11612 7352 11664 7404
rect 6736 7216 6788 7268
rect 9128 7284 9180 7336
rect 11336 7327 11388 7336
rect 11336 7293 11345 7327
rect 11345 7293 11379 7327
rect 11379 7293 11388 7327
rect 11336 7284 11388 7293
rect 13728 7395 13780 7404
rect 13728 7361 13737 7395
rect 13737 7361 13771 7395
rect 13771 7361 13780 7395
rect 13728 7352 13780 7361
rect 14372 7352 14424 7404
rect 16212 7352 16264 7404
rect 18328 7395 18380 7404
rect 18328 7361 18337 7395
rect 18337 7361 18371 7395
rect 18371 7361 18380 7395
rect 18328 7352 18380 7361
rect 2596 7191 2648 7200
rect 2596 7157 2605 7191
rect 2605 7157 2639 7191
rect 2639 7157 2648 7191
rect 2964 7191 3016 7200
rect 2596 7148 2648 7157
rect 2964 7157 2973 7191
rect 2973 7157 3007 7191
rect 3007 7157 3016 7191
rect 2964 7148 3016 7157
rect 3056 7191 3108 7200
rect 3056 7157 3065 7191
rect 3065 7157 3099 7191
rect 3099 7157 3108 7191
rect 3056 7148 3108 7157
rect 4712 7148 4764 7200
rect 6460 7148 6512 7200
rect 7748 7148 7800 7200
rect 8024 7148 8076 7200
rect 8668 7148 8720 7200
rect 9680 7148 9732 7200
rect 9864 7191 9916 7200
rect 9864 7157 9873 7191
rect 9873 7157 9907 7191
rect 9907 7157 9916 7191
rect 9864 7148 9916 7157
rect 11888 7216 11940 7268
rect 14096 7284 14148 7336
rect 14740 7327 14792 7336
rect 14740 7293 14774 7327
rect 14774 7293 14792 7327
rect 14740 7284 14792 7293
rect 15660 7284 15712 7336
rect 11336 7148 11388 7200
rect 12256 7148 12308 7200
rect 13268 7148 13320 7200
rect 14556 7216 14608 7268
rect 15292 7216 15344 7268
rect 15568 7216 15620 7268
rect 13820 7148 13872 7200
rect 14004 7191 14056 7200
rect 14004 7157 14013 7191
rect 14013 7157 14047 7191
rect 14047 7157 14056 7191
rect 14004 7148 14056 7157
rect 18328 7216 18380 7268
rect 15844 7191 15896 7200
rect 15844 7157 15853 7191
rect 15853 7157 15887 7191
rect 15887 7157 15896 7191
rect 15844 7148 15896 7157
rect 16028 7148 16080 7200
rect 16304 7191 16356 7200
rect 16304 7157 16313 7191
rect 16313 7157 16347 7191
rect 16347 7157 16356 7191
rect 16304 7148 16356 7157
rect 17132 7148 17184 7200
rect 17408 7148 17460 7200
rect 18144 7191 18196 7200
rect 18144 7157 18153 7191
rect 18153 7157 18187 7191
rect 18187 7157 18196 7191
rect 18144 7148 18196 7157
rect 6912 7046 6964 7098
rect 6976 7046 7028 7098
rect 7040 7046 7092 7098
rect 7104 7046 7156 7098
rect 12843 7046 12895 7098
rect 12907 7046 12959 7098
rect 12971 7046 13023 7098
rect 13035 7046 13087 7098
rect 2964 6987 3016 6996
rect 2964 6953 2973 6987
rect 2973 6953 3007 6987
rect 3007 6953 3016 6987
rect 2964 6944 3016 6953
rect 3976 6944 4028 6996
rect 4896 6944 4948 6996
rect 5172 6944 5224 6996
rect 11336 6944 11388 6996
rect 11520 6987 11572 6996
rect 11520 6953 11529 6987
rect 11529 6953 11563 6987
rect 11563 6953 11572 6987
rect 11520 6944 11572 6953
rect 4068 6876 4120 6928
rect 7380 6876 7432 6928
rect 7748 6876 7800 6928
rect 8208 6876 8260 6928
rect 8944 6876 8996 6928
rect 9680 6876 9732 6928
rect 12072 6944 12124 6996
rect 4160 6808 4212 6860
rect 3240 6740 3292 6792
rect 3056 6672 3108 6724
rect 5816 6808 5868 6860
rect 6552 6808 6604 6860
rect 6736 6740 6788 6792
rect 2136 6604 2188 6656
rect 2964 6604 3016 6656
rect 3148 6604 3200 6656
rect 3792 6604 3844 6656
rect 5448 6604 5500 6656
rect 6276 6604 6328 6656
rect 7196 6808 7248 6860
rect 7564 6808 7616 6860
rect 7840 6740 7892 6792
rect 8392 6808 8444 6860
rect 8760 6851 8812 6860
rect 8760 6817 8769 6851
rect 8769 6817 8803 6851
rect 8803 6817 8812 6851
rect 8760 6808 8812 6817
rect 8944 6740 8996 6792
rect 7472 6715 7524 6724
rect 7472 6681 7481 6715
rect 7481 6681 7515 6715
rect 7515 6681 7524 6715
rect 7472 6672 7524 6681
rect 9864 6808 9916 6860
rect 10416 6808 10468 6860
rect 11796 6876 11848 6928
rect 13544 6944 13596 6996
rect 13912 6944 13964 6996
rect 16488 6944 16540 6996
rect 16764 6944 16816 6996
rect 17408 6944 17460 6996
rect 11152 6851 11204 6860
rect 11152 6817 11161 6851
rect 11161 6817 11195 6851
rect 11195 6817 11204 6851
rect 11152 6808 11204 6817
rect 12164 6808 12216 6860
rect 12716 6851 12768 6860
rect 12716 6817 12734 6851
rect 12734 6817 12768 6851
rect 12716 6808 12768 6817
rect 15660 6876 15712 6928
rect 15844 6876 15896 6928
rect 16212 6876 16264 6928
rect 11520 6740 11572 6792
rect 11612 6740 11664 6792
rect 11980 6740 12032 6792
rect 13084 6740 13136 6792
rect 11428 6672 11480 6724
rect 8760 6604 8812 6656
rect 8852 6604 8904 6656
rect 9312 6604 9364 6656
rect 12808 6604 12860 6656
rect 13728 6808 13780 6860
rect 13728 6672 13780 6724
rect 14924 6808 14976 6860
rect 14188 6740 14240 6792
rect 14372 6783 14424 6792
rect 14372 6749 14381 6783
rect 14381 6749 14415 6783
rect 14415 6749 14424 6783
rect 14372 6740 14424 6749
rect 17868 6808 17920 6860
rect 15660 6740 15712 6792
rect 17408 6740 17460 6792
rect 18236 6808 18288 6860
rect 18328 6851 18380 6860
rect 18328 6817 18337 6851
rect 18337 6817 18371 6851
rect 18371 6817 18380 6851
rect 18328 6808 18380 6817
rect 18512 6715 18564 6724
rect 18512 6681 18521 6715
rect 18521 6681 18555 6715
rect 18555 6681 18564 6715
rect 18512 6672 18564 6681
rect 15568 6604 15620 6656
rect 17684 6604 17736 6656
rect 3947 6502 3999 6554
rect 4011 6502 4063 6554
rect 4075 6502 4127 6554
rect 4139 6502 4191 6554
rect 9878 6502 9930 6554
rect 9942 6502 9994 6554
rect 10006 6502 10058 6554
rect 10070 6502 10122 6554
rect 15808 6502 15860 6554
rect 15872 6502 15924 6554
rect 15936 6502 15988 6554
rect 16000 6502 16052 6554
rect 2320 6400 2372 6452
rect 2780 6375 2832 6384
rect 2780 6341 2789 6375
rect 2789 6341 2823 6375
rect 2823 6341 2832 6375
rect 2780 6332 2832 6341
rect 3056 6400 3108 6452
rect 8208 6400 8260 6452
rect 10692 6400 10744 6452
rect 11520 6443 11572 6452
rect 11520 6409 11529 6443
rect 11529 6409 11563 6443
rect 11563 6409 11572 6443
rect 11520 6400 11572 6409
rect 11980 6400 12032 6452
rect 13452 6400 13504 6452
rect 13728 6400 13780 6452
rect 14004 6400 14056 6452
rect 3148 6332 3200 6384
rect 5356 6332 5408 6384
rect 7748 6332 7800 6384
rect 10508 6332 10560 6384
rect 11060 6332 11112 6384
rect 12716 6332 12768 6384
rect 14556 6400 14608 6452
rect 16580 6400 16632 6452
rect 1492 6239 1544 6248
rect 1492 6205 1501 6239
rect 1501 6205 1535 6239
rect 1535 6205 1544 6239
rect 1492 6196 1544 6205
rect 2596 6196 2648 6248
rect 3608 6196 3660 6248
rect 4344 6239 4396 6248
rect 4344 6205 4353 6239
rect 4353 6205 4387 6239
rect 4387 6205 4396 6239
rect 4344 6196 4396 6205
rect 6552 6264 6604 6316
rect 8852 6264 8904 6316
rect 9312 6264 9364 6316
rect 9404 6264 9456 6316
rect 10232 6264 10284 6316
rect 14924 6332 14976 6384
rect 6000 6239 6052 6248
rect 6000 6205 6009 6239
rect 6009 6205 6043 6239
rect 6043 6205 6052 6239
rect 6000 6196 6052 6205
rect 6460 6196 6512 6248
rect 7932 6196 7984 6248
rect 9128 6196 9180 6248
rect 2596 6060 2648 6112
rect 2964 6128 3016 6180
rect 3976 6171 4028 6180
rect 3976 6137 3994 6171
rect 3994 6137 4028 6171
rect 3976 6128 4028 6137
rect 4160 6060 4212 6112
rect 5540 6060 5592 6112
rect 6092 6128 6144 6180
rect 7380 6103 7432 6112
rect 7380 6069 7389 6103
rect 7389 6069 7423 6103
rect 7423 6069 7432 6103
rect 8852 6128 8904 6180
rect 10692 6264 10744 6316
rect 12164 6264 12216 6316
rect 12624 6264 12676 6316
rect 14004 6264 14056 6316
rect 14188 6264 14240 6316
rect 15568 6264 15620 6316
rect 10508 6196 10560 6248
rect 12716 6196 12768 6248
rect 11520 6128 11572 6180
rect 13544 6196 13596 6248
rect 13636 6196 13688 6248
rect 17040 6332 17092 6384
rect 16212 6307 16264 6316
rect 16212 6273 16221 6307
rect 16221 6273 16255 6307
rect 16255 6273 16264 6307
rect 16212 6264 16264 6273
rect 16856 6264 16908 6316
rect 16948 6264 17000 6316
rect 17868 6400 17920 6452
rect 17684 6307 17736 6316
rect 17684 6273 17693 6307
rect 17693 6273 17727 6307
rect 17727 6273 17736 6307
rect 17684 6264 17736 6273
rect 16580 6239 16632 6248
rect 16580 6205 16589 6239
rect 16589 6205 16623 6239
rect 16623 6205 16632 6239
rect 16580 6196 16632 6205
rect 7380 6060 7432 6069
rect 8392 6060 8444 6112
rect 9220 6103 9272 6112
rect 9220 6069 9229 6103
rect 9229 6069 9263 6103
rect 9263 6069 9272 6103
rect 9220 6060 9272 6069
rect 9312 6060 9364 6112
rect 9680 6060 9732 6112
rect 10692 6103 10744 6112
rect 10692 6069 10701 6103
rect 10701 6069 10735 6103
rect 10735 6069 10744 6103
rect 10692 6060 10744 6069
rect 10968 6060 11020 6112
rect 11336 6060 11388 6112
rect 11612 6060 11664 6112
rect 11796 6103 11848 6112
rect 11796 6069 11805 6103
rect 11805 6069 11839 6103
rect 11839 6069 11848 6103
rect 11796 6060 11848 6069
rect 13728 6128 13780 6180
rect 12532 6060 12584 6112
rect 13452 6060 13504 6112
rect 13820 6060 13872 6112
rect 14188 6060 14240 6112
rect 17132 6196 17184 6248
rect 15108 6060 15160 6112
rect 15384 6060 15436 6112
rect 18512 6171 18564 6180
rect 18512 6137 18521 6171
rect 18521 6137 18555 6171
rect 18555 6137 18564 6171
rect 18512 6128 18564 6137
rect 17040 6103 17092 6112
rect 17040 6069 17049 6103
rect 17049 6069 17083 6103
rect 17083 6069 17092 6103
rect 17040 6060 17092 6069
rect 17224 6060 17276 6112
rect 17868 6060 17920 6112
rect 6912 5958 6964 6010
rect 6976 5958 7028 6010
rect 7040 5958 7092 6010
rect 7104 5958 7156 6010
rect 12843 5958 12895 6010
rect 12907 5958 12959 6010
rect 12971 5958 13023 6010
rect 13035 5958 13087 6010
rect 3792 5856 3844 5908
rect 4436 5856 4488 5908
rect 6092 5856 6144 5908
rect 6552 5899 6604 5908
rect 1584 5720 1636 5772
rect 2412 5763 2464 5772
rect 2412 5729 2421 5763
rect 2421 5729 2455 5763
rect 2455 5729 2464 5763
rect 2412 5720 2464 5729
rect 2596 5788 2648 5840
rect 3976 5788 4028 5840
rect 6552 5865 6561 5899
rect 6561 5865 6595 5899
rect 6595 5865 6604 5899
rect 6552 5856 6604 5865
rect 7380 5856 7432 5908
rect 8208 5856 8260 5908
rect 8944 5856 8996 5908
rect 11152 5856 11204 5908
rect 11796 5899 11848 5908
rect 11796 5865 11805 5899
rect 11805 5865 11839 5899
rect 11839 5865 11848 5899
rect 11796 5856 11848 5865
rect 12348 5856 12400 5908
rect 14096 5899 14148 5908
rect 2872 5720 2924 5772
rect 4068 5720 4120 5772
rect 3240 5652 3292 5704
rect 3516 5695 3568 5704
rect 2688 5584 2740 5636
rect 2964 5584 3016 5636
rect 3516 5661 3525 5695
rect 3525 5661 3559 5695
rect 3559 5661 3568 5695
rect 3516 5652 3568 5661
rect 3424 5584 3476 5636
rect 4344 5695 4396 5704
rect 4344 5661 4353 5695
rect 4353 5661 4387 5695
rect 4387 5661 4396 5695
rect 4344 5652 4396 5661
rect 6184 5720 6236 5772
rect 6644 5720 6696 5772
rect 7656 5763 7708 5772
rect 7656 5729 7674 5763
rect 7674 5729 7708 5763
rect 7656 5720 7708 5729
rect 8300 5720 8352 5772
rect 8484 5763 8536 5772
rect 8484 5729 8493 5763
rect 8493 5729 8527 5763
rect 8527 5729 8536 5763
rect 8484 5720 8536 5729
rect 8760 5720 8812 5772
rect 4252 5584 4304 5636
rect 5356 5652 5408 5704
rect 5540 5652 5592 5704
rect 5632 5652 5684 5704
rect 5908 5695 5960 5704
rect 5908 5661 5917 5695
rect 5917 5661 5951 5695
rect 5951 5661 5960 5695
rect 5908 5652 5960 5661
rect 7932 5695 7984 5704
rect 7932 5661 7941 5695
rect 7941 5661 7975 5695
rect 7975 5661 7984 5695
rect 7932 5652 7984 5661
rect 8208 5652 8260 5704
rect 8576 5695 8628 5704
rect 8576 5661 8585 5695
rect 8585 5661 8619 5695
rect 8619 5661 8628 5695
rect 8576 5652 8628 5661
rect 2872 5516 2924 5568
rect 4804 5559 4856 5568
rect 4804 5525 4813 5559
rect 4813 5525 4847 5559
rect 4847 5525 4856 5559
rect 4804 5516 4856 5525
rect 6092 5516 6144 5568
rect 6736 5516 6788 5568
rect 8300 5584 8352 5636
rect 9220 5720 9272 5772
rect 10784 5720 10836 5772
rect 9128 5695 9180 5704
rect 9128 5661 9137 5695
rect 9137 5661 9171 5695
rect 9171 5661 9180 5695
rect 9128 5652 9180 5661
rect 10232 5652 10284 5704
rect 13636 5788 13688 5840
rect 14096 5865 14105 5899
rect 14105 5865 14139 5899
rect 14139 5865 14148 5899
rect 14096 5856 14148 5865
rect 14740 5899 14792 5908
rect 14740 5865 14749 5899
rect 14749 5865 14783 5899
rect 14783 5865 14792 5899
rect 14740 5856 14792 5865
rect 15108 5899 15160 5908
rect 15108 5865 15117 5899
rect 15117 5865 15151 5899
rect 15151 5865 15160 5899
rect 15108 5856 15160 5865
rect 17040 5856 17092 5908
rect 18144 5899 18196 5908
rect 18144 5865 18153 5899
rect 18153 5865 18187 5899
rect 18187 5865 18196 5899
rect 18144 5856 18196 5865
rect 14372 5788 14424 5840
rect 15016 5788 15068 5840
rect 15660 5788 15712 5840
rect 11704 5720 11756 5772
rect 13268 5720 13320 5772
rect 14096 5720 14148 5772
rect 14924 5720 14976 5772
rect 15108 5720 15160 5772
rect 16120 5720 16172 5772
rect 16396 5720 16448 5772
rect 17684 5788 17736 5840
rect 18512 5831 18564 5840
rect 18512 5797 18521 5831
rect 18521 5797 18555 5831
rect 18555 5797 18564 5831
rect 18512 5788 18564 5797
rect 17040 5720 17092 5772
rect 11244 5652 11296 5704
rect 11980 5652 12032 5704
rect 12164 5652 12216 5704
rect 8760 5516 8812 5568
rect 10324 5516 10376 5568
rect 10784 5516 10836 5568
rect 11336 5559 11388 5568
rect 11336 5525 11345 5559
rect 11345 5525 11379 5559
rect 11379 5525 11388 5559
rect 11336 5516 11388 5525
rect 11428 5516 11480 5568
rect 11796 5516 11848 5568
rect 14004 5652 14056 5704
rect 15568 5695 15620 5704
rect 15568 5661 15577 5695
rect 15577 5661 15611 5695
rect 15611 5661 15620 5695
rect 15568 5652 15620 5661
rect 16488 5695 16540 5704
rect 13820 5584 13872 5636
rect 14924 5584 14976 5636
rect 16488 5661 16497 5695
rect 16497 5661 16531 5695
rect 16531 5661 16540 5695
rect 16488 5652 16540 5661
rect 16212 5584 16264 5636
rect 13176 5516 13228 5568
rect 14004 5516 14056 5568
rect 14188 5516 14240 5568
rect 15200 5559 15252 5568
rect 15200 5525 15209 5559
rect 15209 5525 15243 5559
rect 15243 5525 15252 5559
rect 15200 5516 15252 5525
rect 16396 5559 16448 5568
rect 16396 5525 16405 5559
rect 16405 5525 16439 5559
rect 16439 5525 16448 5559
rect 16396 5516 16448 5525
rect 17776 5516 17828 5568
rect 3947 5414 3999 5466
rect 4011 5414 4063 5466
rect 4075 5414 4127 5466
rect 4139 5414 4191 5466
rect 9878 5414 9930 5466
rect 9942 5414 9994 5466
rect 10006 5414 10058 5466
rect 10070 5414 10122 5466
rect 15808 5414 15860 5466
rect 15872 5414 15924 5466
rect 15936 5414 15988 5466
rect 16000 5414 16052 5466
rect 1492 5355 1544 5364
rect 1492 5321 1501 5355
rect 1501 5321 1535 5355
rect 1535 5321 1544 5355
rect 1492 5312 1544 5321
rect 4344 5312 4396 5364
rect 3608 5244 3660 5296
rect 7564 5312 7616 5364
rect 8392 5355 8444 5364
rect 8392 5321 8401 5355
rect 8401 5321 8435 5355
rect 8435 5321 8444 5355
rect 8392 5312 8444 5321
rect 11704 5355 11756 5364
rect 11704 5321 11713 5355
rect 11713 5321 11747 5355
rect 11747 5321 11756 5355
rect 11704 5312 11756 5321
rect 13176 5355 13228 5364
rect 13176 5321 13185 5355
rect 13185 5321 13219 5355
rect 13219 5321 13228 5355
rect 13176 5312 13228 5321
rect 6000 5287 6052 5296
rect 6000 5253 6009 5287
rect 6009 5253 6043 5287
rect 6043 5253 6052 5287
rect 6000 5244 6052 5253
rect 6460 5244 6512 5296
rect 2136 5108 2188 5160
rect 7656 5176 7708 5228
rect 8116 5219 8168 5228
rect 8116 5185 8125 5219
rect 8125 5185 8159 5219
rect 8159 5185 8168 5219
rect 8116 5176 8168 5185
rect 3240 5108 3292 5160
rect 3884 5151 3936 5160
rect 3884 5117 3893 5151
rect 3893 5117 3927 5151
rect 3927 5117 3936 5151
rect 3884 5108 3936 5117
rect 4528 5108 4580 5160
rect 6092 5108 6144 5160
rect 6460 5108 6512 5160
rect 7104 5151 7156 5160
rect 1768 4972 1820 5024
rect 1952 5015 2004 5024
rect 1952 4981 1961 5015
rect 1961 4981 1995 5015
rect 1995 4981 2004 5015
rect 1952 4972 2004 4981
rect 2320 4972 2372 5024
rect 3516 5040 3568 5092
rect 3700 5040 3752 5092
rect 4160 5040 4212 5092
rect 3240 4972 3292 5024
rect 4252 5015 4304 5024
rect 4252 4981 4261 5015
rect 4261 4981 4295 5015
rect 4295 4981 4304 5015
rect 4252 4972 4304 4981
rect 5080 4972 5132 5024
rect 5540 5040 5592 5092
rect 7104 5117 7113 5151
rect 7113 5117 7147 5151
rect 7147 5117 7156 5151
rect 7104 5108 7156 5117
rect 7288 5108 7340 5160
rect 8024 5108 8076 5160
rect 8760 5244 8812 5296
rect 9680 5244 9732 5296
rect 8576 5176 8628 5228
rect 9128 5176 9180 5228
rect 10140 5176 10192 5228
rect 11152 5219 11204 5228
rect 11152 5185 11161 5219
rect 11161 5185 11195 5219
rect 11195 5185 11204 5219
rect 11152 5176 11204 5185
rect 11796 5176 11848 5228
rect 15016 5312 15068 5364
rect 17040 5312 17092 5364
rect 17408 5244 17460 5296
rect 17684 5244 17736 5296
rect 15016 5176 15068 5228
rect 16212 5176 16264 5228
rect 7748 5040 7800 5092
rect 8116 5040 8168 5092
rect 9496 5108 9548 5160
rect 9588 5108 9640 5160
rect 10784 5040 10836 5092
rect 11244 5108 11296 5160
rect 11980 5108 12032 5160
rect 11796 5040 11848 5092
rect 12624 5040 12676 5092
rect 13820 5108 13872 5160
rect 14188 5108 14240 5160
rect 14924 5151 14976 5160
rect 14924 5117 14933 5151
rect 14933 5117 14967 5151
rect 14967 5117 14976 5151
rect 15200 5151 15252 5160
rect 14924 5108 14976 5117
rect 15200 5117 15209 5151
rect 15209 5117 15243 5151
rect 15243 5117 15252 5151
rect 15200 5108 15252 5117
rect 6644 4972 6696 5024
rect 7288 4972 7340 5024
rect 7380 4972 7432 5024
rect 7656 4972 7708 5024
rect 8392 4972 8444 5024
rect 9128 4972 9180 5024
rect 9496 5015 9548 5024
rect 9496 4981 9505 5015
rect 9505 4981 9539 5015
rect 9539 4981 9548 5015
rect 9496 4972 9548 4981
rect 9680 4972 9732 5024
rect 11244 5015 11296 5024
rect 11244 4981 11253 5015
rect 11253 4981 11287 5015
rect 11287 4981 11296 5015
rect 11244 4972 11296 4981
rect 15200 4972 15252 5024
rect 15476 5108 15528 5160
rect 15660 5108 15712 5160
rect 16304 5151 16356 5160
rect 16304 5117 16313 5151
rect 16313 5117 16347 5151
rect 16347 5117 16356 5151
rect 16304 5108 16356 5117
rect 16672 5176 16724 5228
rect 17868 5176 17920 5228
rect 15936 5083 15988 5092
rect 15936 5049 15945 5083
rect 15945 5049 15979 5083
rect 15979 5049 15988 5083
rect 15936 5040 15988 5049
rect 18052 5108 18104 5160
rect 15476 5015 15528 5024
rect 15476 4981 15485 5015
rect 15485 4981 15519 5015
rect 15519 4981 15528 5015
rect 18512 5083 18564 5092
rect 18512 5049 18521 5083
rect 18521 5049 18555 5083
rect 18555 5049 18564 5083
rect 18512 5040 18564 5049
rect 15476 4972 15528 4981
rect 17316 4972 17368 5024
rect 17408 4972 17460 5024
rect 17684 4972 17736 5024
rect 17960 5015 18012 5024
rect 17960 4981 17969 5015
rect 17969 4981 18003 5015
rect 18003 4981 18012 5015
rect 17960 4972 18012 4981
rect 6912 4870 6964 4922
rect 6976 4870 7028 4922
rect 7040 4870 7092 4922
rect 7104 4870 7156 4922
rect 12843 4870 12895 4922
rect 12907 4870 12959 4922
rect 12971 4870 13023 4922
rect 13035 4870 13087 4922
rect 1952 4768 2004 4820
rect 2044 4768 2096 4820
rect 2780 4768 2832 4820
rect 4160 4700 4212 4752
rect 5172 4700 5224 4752
rect 5908 4768 5960 4820
rect 6644 4811 6696 4820
rect 6644 4777 6653 4811
rect 6653 4777 6687 4811
rect 6687 4777 6696 4811
rect 6644 4768 6696 4777
rect 7288 4768 7340 4820
rect 8116 4811 8168 4820
rect 8116 4777 8125 4811
rect 8125 4777 8159 4811
rect 8159 4777 8168 4811
rect 8116 4768 8168 4777
rect 9956 4811 10008 4820
rect 9956 4777 9965 4811
rect 9965 4777 9999 4811
rect 9999 4777 10008 4811
rect 9956 4768 10008 4777
rect 10600 4768 10652 4820
rect 11060 4768 11112 4820
rect 11796 4768 11848 4820
rect 12532 4768 12584 4820
rect 12716 4768 12768 4820
rect 13636 4768 13688 4820
rect 14556 4768 14608 4820
rect 14740 4768 14792 4820
rect 17408 4768 17460 4820
rect 17500 4768 17552 4820
rect 3608 4632 3660 4684
rect 3792 4632 3844 4684
rect 2320 4607 2372 4616
rect 2320 4573 2329 4607
rect 2329 4573 2363 4607
rect 2363 4573 2372 4607
rect 2320 4564 2372 4573
rect 3148 4564 3200 4616
rect 3516 4564 3568 4616
rect 4804 4632 4856 4684
rect 5448 4632 5500 4684
rect 7196 4700 7248 4752
rect 5172 4607 5224 4616
rect 1768 4496 1820 4548
rect 2872 4496 2924 4548
rect 4804 4496 4856 4548
rect 5172 4573 5181 4607
rect 5181 4573 5215 4607
rect 5215 4573 5224 4607
rect 5172 4564 5224 4573
rect 5356 4564 5408 4616
rect 5264 4496 5316 4548
rect 6276 4564 6328 4616
rect 6460 4632 6512 4684
rect 7472 4700 7524 4752
rect 6552 4564 6604 4616
rect 6828 4564 6880 4616
rect 8392 4632 8444 4684
rect 8576 4675 8628 4684
rect 8576 4641 8585 4675
rect 8585 4641 8619 4675
rect 8619 4641 8628 4675
rect 8576 4632 8628 4641
rect 8668 4632 8720 4684
rect 9404 4675 9456 4684
rect 9404 4641 9413 4675
rect 9413 4641 9447 4675
rect 9447 4641 9456 4675
rect 9404 4632 9456 4641
rect 7564 4607 7616 4616
rect 7564 4573 7573 4607
rect 7573 4573 7607 4607
rect 7607 4573 7616 4607
rect 7564 4564 7616 4573
rect 10416 4632 10468 4684
rect 10232 4607 10284 4616
rect 10232 4573 10241 4607
rect 10241 4573 10275 4607
rect 10275 4573 10284 4607
rect 10232 4564 10284 4573
rect 1492 4471 1544 4480
rect 1492 4437 1501 4471
rect 1501 4437 1535 4471
rect 1535 4437 1544 4471
rect 1492 4428 1544 4437
rect 3608 4471 3660 4480
rect 3608 4437 3617 4471
rect 3617 4437 3651 4471
rect 3651 4437 3660 4471
rect 3608 4428 3660 4437
rect 4528 4471 4580 4480
rect 4528 4437 4537 4471
rect 4537 4437 4571 4471
rect 4571 4437 4580 4471
rect 4528 4428 4580 4437
rect 4712 4428 4764 4480
rect 5724 4428 5776 4480
rect 8392 4496 8444 4548
rect 9956 4496 10008 4548
rect 11428 4700 11480 4752
rect 15108 4700 15160 4752
rect 16212 4700 16264 4752
rect 16672 4700 16724 4752
rect 11704 4632 11756 4684
rect 12256 4632 12308 4684
rect 12440 4675 12492 4684
rect 12440 4641 12449 4675
rect 12449 4641 12483 4675
rect 12483 4641 12492 4675
rect 12440 4632 12492 4641
rect 13176 4632 13228 4684
rect 10968 4496 11020 4548
rect 12532 4564 12584 4616
rect 6552 4428 6604 4480
rect 8944 4471 8996 4480
rect 8944 4437 8953 4471
rect 8953 4437 8987 4471
rect 8987 4437 8996 4471
rect 8944 4428 8996 4437
rect 9220 4428 9272 4480
rect 11060 4428 11112 4480
rect 11704 4428 11756 4480
rect 11980 4428 12032 4480
rect 12256 4428 12308 4480
rect 14372 4539 14424 4548
rect 14372 4505 14381 4539
rect 14381 4505 14415 4539
rect 14415 4505 14424 4539
rect 14372 4496 14424 4505
rect 13820 4428 13872 4480
rect 14188 4428 14240 4480
rect 16304 4632 16356 4684
rect 16580 4675 16632 4684
rect 16580 4641 16589 4675
rect 16589 4641 16623 4675
rect 16623 4641 16632 4675
rect 16580 4632 16632 4641
rect 15016 4607 15068 4616
rect 15016 4573 15025 4607
rect 15025 4573 15059 4607
rect 15059 4573 15068 4607
rect 15016 4564 15068 4573
rect 16948 4632 17000 4684
rect 16212 4428 16264 4480
rect 17132 4564 17184 4616
rect 17408 4564 17460 4616
rect 18512 4675 18564 4684
rect 18512 4641 18521 4675
rect 18521 4641 18555 4675
rect 18555 4641 18564 4675
rect 18512 4632 18564 4641
rect 17868 4564 17920 4616
rect 18052 4496 18104 4548
rect 17132 4471 17184 4480
rect 17132 4437 17141 4471
rect 17141 4437 17175 4471
rect 17175 4437 17184 4471
rect 17132 4428 17184 4437
rect 18328 4428 18380 4480
rect 3947 4326 3999 4378
rect 4011 4326 4063 4378
rect 4075 4326 4127 4378
rect 4139 4326 4191 4378
rect 9878 4326 9930 4378
rect 9942 4326 9994 4378
rect 10006 4326 10058 4378
rect 10070 4326 10122 4378
rect 15808 4326 15860 4378
rect 15872 4326 15924 4378
rect 15936 4326 15988 4378
rect 16000 4326 16052 4378
rect 388 4224 440 4276
rect 3332 4224 3384 4276
rect 5172 4224 5224 4276
rect 6276 4267 6328 4276
rect 2412 4156 2464 4208
rect 4160 4156 4212 4208
rect 4436 4156 4488 4208
rect 2136 4131 2188 4140
rect 2136 4097 2145 4131
rect 2145 4097 2179 4131
rect 2179 4097 2188 4131
rect 2136 4088 2188 4097
rect 1584 4063 1636 4072
rect 1584 4029 1593 4063
rect 1593 4029 1627 4063
rect 1627 4029 1636 4063
rect 1584 4020 1636 4029
rect 2596 4088 2648 4140
rect 3976 4088 4028 4140
rect 5356 4199 5408 4208
rect 5356 4165 5365 4199
rect 5365 4165 5399 4199
rect 5399 4165 5408 4199
rect 5356 4156 5408 4165
rect 6276 4233 6285 4267
rect 6285 4233 6319 4267
rect 6319 4233 6328 4267
rect 6276 4224 6328 4233
rect 7656 4224 7708 4276
rect 7840 4224 7892 4276
rect 8208 4224 8260 4276
rect 6736 4199 6788 4208
rect 6736 4165 6745 4199
rect 6745 4165 6779 4199
rect 6779 4165 6788 4199
rect 6736 4156 6788 4165
rect 5816 4131 5868 4140
rect 5816 4097 5825 4131
rect 5825 4097 5859 4131
rect 5859 4097 5868 4131
rect 5816 4088 5868 4097
rect 5908 4131 5960 4140
rect 5908 4097 5917 4131
rect 5917 4097 5951 4131
rect 5951 4097 5960 4131
rect 5908 4088 5960 4097
rect 6092 4088 6144 4140
rect 10048 4156 10100 4208
rect 10968 4224 11020 4276
rect 11060 4224 11112 4276
rect 14740 4224 14792 4276
rect 16580 4224 16632 4276
rect 10416 4156 10468 4208
rect 10600 4156 10652 4208
rect 10232 4088 10284 4140
rect 2964 4063 3016 4072
rect 2964 4029 2973 4063
rect 2973 4029 3007 4063
rect 3007 4029 3016 4063
rect 2964 4020 3016 4029
rect 1492 3927 1544 3936
rect 1492 3893 1501 3927
rect 1501 3893 1535 3927
rect 1535 3893 1544 3927
rect 1492 3884 1544 3893
rect 1860 3927 1912 3936
rect 1860 3893 1869 3927
rect 1869 3893 1903 3927
rect 1903 3893 1912 3927
rect 1860 3884 1912 3893
rect 2504 3952 2556 4004
rect 3516 4020 3568 4072
rect 5724 4020 5776 4072
rect 6184 4020 6236 4072
rect 6644 4063 6696 4072
rect 6644 4029 6653 4063
rect 6653 4029 6687 4063
rect 6687 4029 6696 4063
rect 6644 4020 6696 4029
rect 7564 4020 7616 4072
rect 9680 4020 9732 4072
rect 9956 4020 10008 4072
rect 3976 3952 4028 4004
rect 4068 3952 4120 4004
rect 4712 3952 4764 4004
rect 5264 3952 5316 4004
rect 3516 3884 3568 3936
rect 4344 3927 4396 3936
rect 4344 3893 4353 3927
rect 4353 3893 4387 3927
rect 4387 3893 4396 3927
rect 4344 3884 4396 3893
rect 4436 3884 4488 3936
rect 4620 3884 4672 3936
rect 5080 3884 5132 3936
rect 6276 3884 6328 3936
rect 6460 3927 6512 3936
rect 6460 3893 6469 3927
rect 6469 3893 6503 3927
rect 6503 3893 6512 3927
rect 6460 3884 6512 3893
rect 8116 3884 8168 3936
rect 8484 3884 8536 3936
rect 9772 3884 9824 3936
rect 10692 4088 10744 4140
rect 11428 4156 11480 4208
rect 12164 4088 12216 4140
rect 12624 4088 12676 4140
rect 12716 4088 12768 4140
rect 13820 4088 13872 4140
rect 11336 4020 11388 4072
rect 12256 4063 12308 4072
rect 12256 4029 12265 4063
rect 12265 4029 12299 4063
rect 12299 4029 12308 4063
rect 12256 4020 12308 4029
rect 13084 4063 13136 4072
rect 13084 4029 13093 4063
rect 13093 4029 13127 4063
rect 13127 4029 13136 4063
rect 13084 4020 13136 4029
rect 13636 4020 13688 4072
rect 15108 4088 15160 4140
rect 16488 4088 16540 4140
rect 17132 4088 17184 4140
rect 17776 4088 17828 4140
rect 18144 4131 18196 4140
rect 18144 4097 18153 4131
rect 18153 4097 18187 4131
rect 18187 4097 18196 4131
rect 18144 4088 18196 4097
rect 14372 4020 14424 4072
rect 14648 4020 14700 4072
rect 16212 4020 16264 4072
rect 17316 4063 17368 4072
rect 9956 3884 10008 3936
rect 10232 3884 10284 3936
rect 10600 3927 10652 3936
rect 10600 3893 10609 3927
rect 10609 3893 10643 3927
rect 10643 3893 10652 3927
rect 10600 3884 10652 3893
rect 11612 3952 11664 4004
rect 13176 3884 13228 3936
rect 17316 4029 17325 4063
rect 17325 4029 17359 4063
rect 17359 4029 17368 4063
rect 17316 4020 17368 4029
rect 18052 4020 18104 4072
rect 13544 3884 13596 3936
rect 14372 3927 14424 3936
rect 14372 3893 14381 3927
rect 14381 3893 14415 3927
rect 14415 3893 14424 3927
rect 14372 3884 14424 3893
rect 14648 3927 14700 3936
rect 14648 3893 14657 3927
rect 14657 3893 14691 3927
rect 14691 3893 14700 3927
rect 14648 3884 14700 3893
rect 14924 3927 14976 3936
rect 14924 3893 14933 3927
rect 14933 3893 14967 3927
rect 14967 3893 14976 3927
rect 14924 3884 14976 3893
rect 18512 3995 18564 4004
rect 18512 3961 18521 3995
rect 18521 3961 18555 3995
rect 18555 3961 18564 3995
rect 18512 3952 18564 3961
rect 16948 3927 17000 3936
rect 16948 3893 16957 3927
rect 16957 3893 16991 3927
rect 16991 3893 17000 3927
rect 16948 3884 17000 3893
rect 6912 3782 6964 3834
rect 6976 3782 7028 3834
rect 7040 3782 7092 3834
rect 7104 3782 7156 3834
rect 12843 3782 12895 3834
rect 12907 3782 12959 3834
rect 12971 3782 13023 3834
rect 13035 3782 13087 3834
rect 2320 3680 2372 3732
rect 2596 3612 2648 3664
rect 2044 3544 2096 3596
rect 2964 3544 3016 3596
rect 4988 3680 5040 3732
rect 5080 3680 5132 3732
rect 6736 3680 6788 3732
rect 7564 3680 7616 3732
rect 8944 3680 8996 3732
rect 9128 3723 9180 3732
rect 9128 3689 9137 3723
rect 9137 3689 9171 3723
rect 9171 3689 9180 3723
rect 9128 3680 9180 3689
rect 3976 3612 4028 3664
rect 4344 3612 4396 3664
rect 4620 3612 4672 3664
rect 3240 3519 3292 3528
rect 3240 3485 3249 3519
rect 3249 3485 3283 3519
rect 3283 3485 3292 3519
rect 3240 3476 3292 3485
rect 3424 3544 3476 3596
rect 5264 3612 5316 3664
rect 5172 3544 5224 3596
rect 8484 3612 8536 3664
rect 10600 3612 10652 3664
rect 11428 3680 11480 3732
rect 13820 3723 13872 3732
rect 13820 3689 13829 3723
rect 13829 3689 13863 3723
rect 13863 3689 13872 3723
rect 13820 3680 13872 3689
rect 15568 3680 15620 3732
rect 12716 3655 12768 3664
rect 6000 3544 6052 3596
rect 6736 3544 6788 3596
rect 4160 3476 4212 3528
rect 6092 3519 6144 3528
rect 6092 3485 6101 3519
rect 6101 3485 6135 3519
rect 6135 3485 6144 3519
rect 6092 3476 6144 3485
rect 8576 3544 8628 3596
rect 9036 3544 9088 3596
rect 9220 3544 9272 3596
rect 11980 3544 12032 3596
rect 12716 3621 12750 3655
rect 12750 3621 12768 3655
rect 12716 3612 12768 3621
rect 16488 3680 16540 3732
rect 16948 3680 17000 3732
rect 8852 3519 8904 3528
rect 8852 3485 8861 3519
rect 8861 3485 8895 3519
rect 8895 3485 8904 3519
rect 8852 3476 8904 3485
rect 10968 3519 11020 3528
rect 10968 3485 10984 3519
rect 10984 3485 11018 3519
rect 11018 3485 11020 3519
rect 10968 3476 11020 3485
rect 7748 3408 7800 3460
rect 9220 3408 9272 3460
rect 13912 3544 13964 3596
rect 14556 3587 14608 3596
rect 14556 3553 14565 3587
rect 14565 3553 14599 3587
rect 14599 3553 14608 3587
rect 14556 3544 14608 3553
rect 15292 3544 15344 3596
rect 15660 3544 15712 3596
rect 12440 3519 12492 3528
rect 12440 3485 12449 3519
rect 12449 3485 12483 3519
rect 12483 3485 12492 3519
rect 12440 3476 12492 3485
rect 14188 3476 14240 3528
rect 14924 3476 14976 3528
rect 16212 3544 16264 3596
rect 16396 3544 16448 3596
rect 17684 3612 17736 3664
rect 17960 3655 18012 3664
rect 17960 3621 17969 3655
rect 17969 3621 18003 3655
rect 18003 3621 18012 3655
rect 17960 3612 18012 3621
rect 3700 3383 3752 3392
rect 3700 3349 3709 3383
rect 3709 3349 3743 3383
rect 3743 3349 3752 3383
rect 3700 3340 3752 3349
rect 3792 3340 3844 3392
rect 4344 3340 4396 3392
rect 4988 3340 5040 3392
rect 6000 3383 6052 3392
rect 6000 3349 6009 3383
rect 6009 3349 6043 3383
rect 6043 3349 6052 3383
rect 6000 3340 6052 3349
rect 6092 3340 6144 3392
rect 7840 3383 7892 3392
rect 7840 3349 7849 3383
rect 7849 3349 7883 3383
rect 7883 3349 7892 3383
rect 7840 3340 7892 3349
rect 8484 3340 8536 3392
rect 9772 3340 9824 3392
rect 13912 3383 13964 3392
rect 13912 3349 13921 3383
rect 13921 3349 13955 3383
rect 13955 3349 13964 3383
rect 13912 3340 13964 3349
rect 14096 3340 14148 3392
rect 16672 3476 16724 3528
rect 17500 3544 17552 3596
rect 18144 3587 18196 3596
rect 18144 3553 18153 3587
rect 18153 3553 18187 3587
rect 18187 3553 18196 3587
rect 18144 3544 18196 3553
rect 16212 3408 16264 3460
rect 16304 3408 16356 3460
rect 16764 3408 16816 3460
rect 18512 3451 18564 3460
rect 18512 3417 18521 3451
rect 18521 3417 18555 3451
rect 18555 3417 18564 3451
rect 18512 3408 18564 3417
rect 15660 3340 15712 3392
rect 16672 3340 16724 3392
rect 17408 3340 17460 3392
rect 17960 3340 18012 3392
rect 3947 3238 3999 3290
rect 4011 3238 4063 3290
rect 4075 3238 4127 3290
rect 4139 3238 4191 3290
rect 9878 3238 9930 3290
rect 9942 3238 9994 3290
rect 10006 3238 10058 3290
rect 10070 3238 10122 3290
rect 15808 3238 15860 3290
rect 15872 3238 15924 3290
rect 15936 3238 15988 3290
rect 16000 3238 16052 3290
rect 1676 3136 1728 3188
rect 2964 3136 3016 3188
rect 3240 3136 3292 3188
rect 1400 3111 1452 3120
rect 1400 3077 1409 3111
rect 1409 3077 1443 3111
rect 1443 3077 1452 3111
rect 1400 3068 1452 3077
rect 3148 3000 3200 3052
rect 7840 3136 7892 3188
rect 9128 3136 9180 3188
rect 9220 3136 9272 3188
rect 13176 3136 13228 3188
rect 15292 3179 15344 3188
rect 4528 3043 4580 3052
rect 1952 2975 2004 2984
rect 1952 2941 1961 2975
rect 1961 2941 1995 2975
rect 1995 2941 2004 2975
rect 1952 2932 2004 2941
rect 2320 2975 2372 2984
rect 2320 2941 2329 2975
rect 2329 2941 2363 2975
rect 2363 2941 2372 2975
rect 2320 2932 2372 2941
rect 2780 2932 2832 2984
rect 3240 2932 3292 2984
rect 4528 3009 4537 3043
rect 4537 3009 4571 3043
rect 4571 3009 4580 3043
rect 4528 3000 4580 3009
rect 4620 3043 4672 3052
rect 4620 3009 4629 3043
rect 4629 3009 4663 3043
rect 4663 3009 4672 3043
rect 4896 3043 4948 3052
rect 4620 3000 4672 3009
rect 4896 3009 4905 3043
rect 4905 3009 4939 3043
rect 4939 3009 4948 3043
rect 4896 3000 4948 3009
rect 5908 3000 5960 3052
rect 6552 3043 6604 3052
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 10324 3068 10376 3120
rect 13452 3068 13504 3120
rect 15292 3145 15301 3179
rect 15301 3145 15335 3179
rect 15335 3145 15344 3179
rect 15292 3136 15344 3145
rect 15568 3136 15620 3188
rect 16856 3136 16908 3188
rect 17684 3068 17736 3120
rect 8300 3043 8352 3052
rect 8300 3009 8309 3043
rect 8309 3009 8343 3043
rect 8343 3009 8352 3043
rect 8300 3000 8352 3009
rect 8484 3043 8536 3052
rect 8484 3009 8493 3043
rect 8493 3009 8527 3043
rect 8527 3009 8536 3043
rect 8484 3000 8536 3009
rect 8852 3000 8904 3052
rect 9680 3000 9732 3052
rect 4252 2932 4304 2984
rect 4436 2975 4488 2984
rect 4436 2941 4445 2975
rect 4445 2941 4479 2975
rect 4479 2941 4488 2975
rect 4436 2932 4488 2941
rect 2228 2864 2280 2916
rect 4804 2932 4856 2984
rect 5540 2932 5592 2984
rect 6736 2975 6788 2984
rect 6736 2941 6745 2975
rect 6745 2941 6779 2975
rect 6779 2941 6788 2975
rect 6736 2932 6788 2941
rect 9772 2932 9824 2984
rect 10692 3000 10744 3052
rect 11796 3043 11848 3052
rect 11796 3009 11805 3043
rect 11805 3009 11839 3043
rect 11839 3009 11848 3043
rect 11796 3000 11848 3009
rect 11980 3000 12032 3052
rect 11428 2932 11480 2984
rect 12164 2932 12216 2984
rect 13360 2932 13412 2984
rect 14648 3000 14700 3052
rect 15476 3000 15528 3052
rect 16396 3000 16448 3052
rect 16488 3000 16540 3052
rect 14280 2932 14332 2984
rect 14464 2932 14516 2984
rect 14832 2932 14884 2984
rect 15384 2932 15436 2984
rect 15660 2975 15712 2984
rect 15660 2941 15669 2975
rect 15669 2941 15703 2975
rect 15703 2941 15712 2975
rect 15660 2932 15712 2941
rect 16212 2932 16264 2984
rect 8484 2864 8536 2916
rect 3332 2839 3384 2848
rect 3332 2805 3341 2839
rect 3341 2805 3375 2839
rect 3375 2805 3384 2839
rect 3332 2796 3384 2805
rect 3700 2839 3752 2848
rect 3700 2805 3709 2839
rect 3709 2805 3743 2839
rect 3743 2805 3752 2839
rect 3700 2796 3752 2805
rect 5080 2839 5132 2848
rect 5080 2805 5089 2839
rect 5089 2805 5123 2839
rect 5123 2805 5132 2839
rect 5080 2796 5132 2805
rect 5632 2796 5684 2848
rect 7472 2796 7524 2848
rect 7656 2839 7708 2848
rect 7656 2805 7665 2839
rect 7665 2805 7699 2839
rect 7699 2805 7708 2839
rect 7656 2796 7708 2805
rect 7748 2839 7800 2848
rect 7748 2805 7757 2839
rect 7757 2805 7791 2839
rect 7791 2805 7800 2839
rect 7748 2796 7800 2805
rect 8668 2796 8720 2848
rect 8852 2796 8904 2848
rect 9956 2796 10008 2848
rect 10416 2796 10468 2848
rect 11520 2864 11572 2916
rect 11888 2864 11940 2916
rect 12072 2796 12124 2848
rect 15476 2864 15528 2916
rect 12624 2796 12676 2848
rect 13636 2796 13688 2848
rect 13912 2839 13964 2848
rect 13912 2805 13921 2839
rect 13921 2805 13955 2839
rect 13955 2805 13964 2839
rect 13912 2796 13964 2805
rect 14280 2796 14332 2848
rect 14556 2839 14608 2848
rect 14556 2805 14565 2839
rect 14565 2805 14599 2839
rect 14599 2805 14608 2839
rect 14556 2796 14608 2805
rect 14924 2839 14976 2848
rect 14924 2805 14933 2839
rect 14933 2805 14967 2839
rect 14967 2805 14976 2839
rect 14924 2796 14976 2805
rect 15200 2796 15252 2848
rect 15568 2796 15620 2848
rect 16028 2864 16080 2916
rect 15936 2796 15988 2848
rect 16212 2796 16264 2848
rect 16672 2932 16724 2984
rect 16856 2932 16908 2984
rect 17592 2975 17644 2984
rect 17592 2941 17601 2975
rect 17601 2941 17635 2975
rect 17635 2941 17644 2975
rect 17592 2932 17644 2941
rect 17960 2975 18012 2984
rect 17960 2941 17969 2975
rect 17969 2941 18003 2975
rect 18003 2941 18012 2975
rect 17960 2932 18012 2941
rect 18328 2975 18380 2984
rect 18328 2941 18337 2975
rect 18337 2941 18371 2975
rect 18371 2941 18380 2975
rect 18328 2932 18380 2941
rect 16488 2864 16540 2916
rect 16580 2839 16632 2848
rect 16580 2805 16589 2839
rect 16589 2805 16623 2839
rect 16623 2805 16632 2839
rect 16580 2796 16632 2805
rect 17868 2864 17920 2916
rect 18144 2907 18196 2916
rect 18144 2873 18153 2907
rect 18153 2873 18187 2907
rect 18187 2873 18196 2907
rect 18144 2864 18196 2873
rect 18420 2839 18472 2848
rect 18420 2805 18429 2839
rect 18429 2805 18463 2839
rect 18463 2805 18472 2839
rect 18420 2796 18472 2805
rect 6912 2694 6964 2746
rect 6976 2694 7028 2746
rect 7040 2694 7092 2746
rect 7104 2694 7156 2746
rect 12843 2694 12895 2746
rect 12907 2694 12959 2746
rect 12971 2694 13023 2746
rect 13035 2694 13087 2746
rect 2872 2592 2924 2644
rect 3056 2592 3108 2644
rect 3608 2567 3660 2576
rect 3608 2533 3617 2567
rect 3617 2533 3651 2567
rect 3651 2533 3660 2567
rect 3608 2524 3660 2533
rect 4344 2592 4396 2644
rect 5080 2592 5132 2644
rect 6552 2592 6604 2644
rect 7656 2592 7708 2644
rect 8668 2592 8720 2644
rect 9036 2592 9088 2644
rect 9588 2592 9640 2644
rect 1584 2499 1636 2508
rect 1584 2465 1593 2499
rect 1593 2465 1627 2499
rect 1627 2465 1636 2499
rect 1584 2456 1636 2465
rect 2320 2499 2372 2508
rect 2320 2465 2329 2499
rect 2329 2465 2363 2499
rect 2363 2465 2372 2499
rect 2320 2456 2372 2465
rect 2688 2499 2740 2508
rect 2688 2465 2697 2499
rect 2697 2465 2731 2499
rect 2731 2465 2740 2499
rect 2688 2456 2740 2465
rect 3516 2456 3568 2508
rect 4344 2456 4396 2508
rect 5356 2524 5408 2576
rect 8576 2524 8628 2576
rect 9772 2567 9824 2576
rect 9772 2533 9781 2567
rect 9781 2533 9815 2567
rect 9815 2533 9824 2567
rect 11244 2592 11296 2644
rect 12624 2635 12676 2644
rect 12624 2601 12633 2635
rect 12633 2601 12667 2635
rect 12667 2601 12676 2635
rect 12624 2592 12676 2601
rect 9772 2524 9824 2533
rect 10508 2524 10560 2576
rect 13912 2592 13964 2644
rect 6000 2499 6052 2508
rect 2780 2388 2832 2440
rect 4712 2388 4764 2440
rect 6000 2465 6009 2499
rect 6009 2465 6043 2499
rect 6043 2465 6052 2499
rect 6000 2456 6052 2465
rect 6368 2499 6420 2508
rect 6368 2465 6377 2499
rect 6377 2465 6411 2499
rect 6411 2465 6420 2499
rect 6368 2456 6420 2465
rect 1216 2320 1268 2372
rect 2136 2363 2188 2372
rect 2136 2329 2145 2363
rect 2145 2329 2179 2363
rect 2179 2329 2188 2363
rect 2136 2320 2188 2329
rect 3056 2363 3108 2372
rect 3056 2329 3065 2363
rect 3065 2329 3099 2363
rect 3099 2329 3108 2363
rect 3056 2320 3108 2329
rect 3424 2363 3476 2372
rect 3424 2329 3433 2363
rect 3433 2329 3467 2363
rect 3467 2329 3476 2363
rect 3424 2320 3476 2329
rect 3792 2320 3844 2372
rect 5816 2363 5868 2372
rect 5816 2329 5825 2363
rect 5825 2329 5859 2363
rect 5859 2329 5868 2363
rect 5816 2320 5868 2329
rect 6736 2363 6788 2372
rect 6736 2329 6745 2363
rect 6745 2329 6779 2363
rect 6779 2329 6788 2363
rect 6736 2320 6788 2329
rect 4896 2252 4948 2304
rect 5540 2252 5592 2304
rect 6828 2252 6880 2304
rect 8208 2456 8260 2508
rect 8300 2456 8352 2508
rect 8116 2431 8168 2440
rect 7564 2320 7616 2372
rect 8116 2397 8125 2431
rect 8125 2397 8159 2431
rect 8159 2397 8168 2431
rect 8116 2388 8168 2397
rect 9680 2456 9732 2508
rect 10600 2499 10652 2508
rect 9588 2388 9640 2440
rect 9956 2388 10008 2440
rect 9680 2320 9732 2372
rect 10600 2465 10609 2499
rect 10609 2465 10643 2499
rect 10643 2465 10652 2499
rect 10600 2456 10652 2465
rect 12164 2499 12216 2508
rect 12164 2465 12173 2499
rect 12173 2465 12207 2499
rect 12207 2465 12216 2499
rect 12164 2456 12216 2465
rect 9312 2252 9364 2304
rect 10784 2431 10836 2440
rect 10784 2397 10793 2431
rect 10793 2397 10827 2431
rect 10827 2397 10836 2431
rect 10784 2388 10836 2397
rect 11796 2388 11848 2440
rect 14280 2592 14332 2644
rect 15108 2592 15160 2644
rect 14556 2524 14608 2576
rect 14924 2524 14976 2576
rect 15936 2567 15988 2576
rect 15936 2533 15945 2567
rect 15945 2533 15979 2567
rect 15979 2533 15988 2567
rect 15936 2524 15988 2533
rect 13452 2499 13504 2508
rect 13452 2465 13461 2499
rect 13461 2465 13495 2499
rect 13495 2465 13504 2499
rect 13452 2456 13504 2465
rect 13728 2456 13780 2508
rect 14740 2499 14792 2508
rect 14740 2465 14749 2499
rect 14749 2465 14783 2499
rect 14783 2465 14792 2499
rect 14740 2456 14792 2465
rect 16028 2456 16080 2508
rect 16856 2567 16908 2576
rect 16856 2533 16865 2567
rect 16865 2533 16899 2567
rect 16899 2533 16908 2567
rect 16856 2524 16908 2533
rect 16948 2524 17000 2576
rect 17776 2567 17828 2576
rect 17776 2533 17785 2567
rect 17785 2533 17819 2567
rect 17819 2533 17828 2567
rect 17776 2524 17828 2533
rect 17500 2456 17552 2508
rect 17684 2456 17736 2508
rect 11244 2363 11296 2372
rect 11244 2329 11253 2363
rect 11253 2329 11287 2363
rect 11287 2329 11296 2363
rect 11244 2320 11296 2329
rect 12256 2320 12308 2372
rect 13084 2363 13136 2372
rect 13084 2329 13093 2363
rect 13093 2329 13127 2363
rect 13127 2329 13136 2363
rect 13084 2320 13136 2329
rect 13912 2363 13964 2372
rect 13912 2329 13921 2363
rect 13921 2329 13955 2363
rect 13955 2329 13964 2363
rect 13912 2320 13964 2329
rect 16580 2388 16632 2440
rect 14832 2363 14884 2372
rect 14832 2329 14841 2363
rect 14841 2329 14875 2363
rect 14875 2329 14884 2363
rect 14832 2320 14884 2329
rect 15660 2320 15712 2372
rect 16856 2320 16908 2372
rect 17040 2363 17092 2372
rect 17040 2329 17049 2363
rect 17049 2329 17083 2363
rect 17083 2329 17092 2363
rect 17040 2320 17092 2329
rect 11152 2295 11204 2304
rect 11152 2261 11161 2295
rect 11161 2261 11195 2295
rect 11195 2261 11204 2295
rect 11152 2252 11204 2261
rect 11336 2252 11388 2304
rect 13820 2252 13872 2304
rect 14096 2252 14148 2304
rect 14280 2295 14332 2304
rect 14280 2261 14289 2295
rect 14289 2261 14323 2295
rect 14323 2261 14332 2295
rect 14280 2252 14332 2261
rect 19432 2388 19484 2440
rect 17592 2363 17644 2372
rect 17592 2329 17601 2363
rect 17601 2329 17635 2363
rect 17635 2329 17644 2363
rect 17592 2320 17644 2329
rect 18512 2363 18564 2372
rect 18512 2329 18521 2363
rect 18521 2329 18555 2363
rect 18555 2329 18564 2363
rect 18512 2320 18564 2329
rect 18420 2252 18472 2304
rect 3947 2150 3999 2202
rect 4011 2150 4063 2202
rect 4075 2150 4127 2202
rect 4139 2150 4191 2202
rect 9878 2150 9930 2202
rect 9942 2150 9994 2202
rect 10006 2150 10058 2202
rect 10070 2150 10122 2202
rect 15808 2150 15860 2202
rect 15872 2150 15924 2202
rect 15936 2150 15988 2202
rect 16000 2150 16052 2202
rect 6000 2048 6052 2100
rect 9496 2048 9548 2100
rect 11152 2048 11204 2100
rect 14464 2048 14516 2100
rect 16212 2048 16264 2100
rect 1584 1980 1636 2032
rect 2320 1912 2372 1964
rect 8208 1980 8260 2032
rect 11336 1980 11388 2032
rect 6644 1844 6696 1896
rect 10600 1844 10652 1896
rect 4344 1776 4396 1828
rect 11060 1776 11112 1828
rect 3516 1708 3568 1760
rect 10232 1708 10284 1760
rect 14188 1708 14240 1760
rect 8392 1640 8444 1692
rect 6828 1572 6880 1624
rect 9772 1572 9824 1624
rect 14280 1572 14332 1624
rect 5908 1504 5960 1556
rect 12164 1504 12216 1556
rect 7472 1368 7524 1420
rect 9404 1368 9456 1420
<< metal2 >>
rect 1950 16400 2006 17200
rect 3054 16960 3110 16969
rect 3054 16895 3110 16904
rect 1490 16008 1546 16017
rect 1490 15943 1546 15952
rect 1504 14822 1532 15943
rect 1858 15056 1914 15065
rect 1858 14991 1914 15000
rect 1492 14816 1544 14822
rect 1492 14758 1544 14764
rect 1504 14550 1532 14758
rect 1872 14618 1900 14991
rect 1964 14634 1992 16400
rect 2964 14816 3016 14822
rect 2964 14758 3016 14764
rect 2226 14648 2282 14657
rect 1860 14612 1912 14618
rect 1964 14606 2084 14634
rect 1860 14554 1912 14560
rect 2056 14550 2084 14606
rect 2226 14583 2228 14592
rect 2280 14583 2282 14592
rect 2780 14612 2832 14618
rect 2228 14554 2280 14560
rect 2780 14554 2832 14560
rect 1492 14544 1544 14550
rect 1492 14486 1544 14492
rect 2044 14544 2096 14550
rect 2044 14486 2096 14492
rect 2320 14476 2372 14482
rect 2320 14418 2372 14424
rect 2688 14476 2740 14482
rect 2688 14418 2740 14424
rect 1858 14376 1914 14385
rect 1858 14311 1914 14320
rect 1872 14074 1900 14311
rect 2044 14272 2096 14278
rect 2044 14214 2096 14220
rect 1860 14068 1912 14074
rect 1860 14010 1912 14016
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 1412 13297 1440 13806
rect 1584 13796 1636 13802
rect 1584 13738 1636 13744
rect 1952 13796 2004 13802
rect 1952 13738 2004 13744
rect 1596 13530 1624 13738
rect 1964 13530 1992 13738
rect 1584 13524 1636 13530
rect 1584 13466 1636 13472
rect 1952 13524 2004 13530
rect 1952 13466 2004 13472
rect 2056 13394 2084 14214
rect 2332 14074 2360 14418
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 2700 14362 2728 14418
rect 2792 14362 2820 14554
rect 2320 14068 2372 14074
rect 2320 14010 2372 14016
rect 2516 14006 2544 14350
rect 2700 14334 2820 14362
rect 2136 14000 2188 14006
rect 2134 13968 2136 13977
rect 2504 14000 2556 14006
rect 2188 13968 2190 13977
rect 2504 13942 2556 13948
rect 2134 13903 2190 13912
rect 2792 13705 2820 14334
rect 2872 14340 2924 14346
rect 2872 14282 2924 14288
rect 2884 14074 2912 14282
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 2778 13696 2834 13705
rect 2778 13631 2834 13640
rect 2976 13530 3004 14758
rect 3068 14482 3096 16895
rect 3514 16688 3570 16697
rect 3514 16623 3570 16632
rect 3332 14544 3384 14550
rect 3332 14486 3384 14492
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 3068 14090 3096 14418
rect 3068 14062 3188 14090
rect 3160 13938 3188 14062
rect 3344 14006 3372 14486
rect 3528 14482 3556 16623
rect 5906 16400 5962 17200
rect 9862 16400 9918 17200
rect 13910 16400 13966 17200
rect 17314 16960 17370 16969
rect 17314 16895 17370 16904
rect 16210 16552 16266 16561
rect 16210 16487 16266 16496
rect 3882 16280 3938 16289
rect 3882 16215 3938 16224
rect 3896 14482 3924 16215
rect 4250 15600 4306 15609
rect 4250 15535 4306 15544
rect 4158 15328 4214 15337
rect 4158 15263 4214 15272
rect 4172 14550 4200 15263
rect 4160 14544 4212 14550
rect 4160 14486 4212 14492
rect 4264 14482 4292 15535
rect 4436 14612 4488 14618
rect 4436 14554 4488 14560
rect 3516 14476 3568 14482
rect 3516 14418 3568 14424
rect 3884 14476 3936 14482
rect 3884 14418 3936 14424
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 3424 14272 3476 14278
rect 3424 14214 3476 14220
rect 3332 14000 3384 14006
rect 3332 13942 3384 13948
rect 3148 13932 3200 13938
rect 3148 13874 3200 13880
rect 3436 13734 3464 14214
rect 3528 13954 3556 14418
rect 3896 14362 3924 14418
rect 3712 14334 3924 14362
rect 4264 14362 4292 14418
rect 4264 14334 4384 14362
rect 3712 14006 3740 14334
rect 4356 14278 4384 14334
rect 3792 14272 3844 14278
rect 3792 14214 3844 14220
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4344 14272 4396 14278
rect 4344 14214 4396 14220
rect 3700 14000 3752 14006
rect 3528 13938 3648 13954
rect 3700 13942 3752 13948
rect 3528 13932 3660 13938
rect 3528 13926 3608 13932
rect 3608 13874 3660 13880
rect 3804 13802 3832 14214
rect 3921 14172 4217 14192
rect 3977 14170 4001 14172
rect 4057 14170 4081 14172
rect 4137 14170 4161 14172
rect 3999 14118 4001 14170
rect 4063 14118 4075 14170
rect 4137 14118 4139 14170
rect 3977 14116 4001 14118
rect 4057 14116 4081 14118
rect 4137 14116 4161 14118
rect 3921 14096 4217 14116
rect 3792 13796 3844 13802
rect 3792 13738 3844 13744
rect 3424 13728 3476 13734
rect 3424 13670 3476 13676
rect 2964 13524 3016 13530
rect 2964 13466 3016 13472
rect 1492 13388 1544 13394
rect 1492 13330 1544 13336
rect 2044 13388 2096 13394
rect 2044 13330 2096 13336
rect 1398 13288 1454 13297
rect 1398 13223 1454 13232
rect 1504 12753 1532 13330
rect 2226 13016 2282 13025
rect 2226 12951 2282 12960
rect 1490 12744 1546 12753
rect 1400 12708 1452 12714
rect 2240 12714 2268 12951
rect 3436 12782 3464 13670
rect 3804 13462 3832 13738
rect 3792 13456 3844 13462
rect 3792 13398 3844 13404
rect 4264 13394 4292 14214
rect 4448 14006 4476 14554
rect 5920 14550 5948 16400
rect 6886 14716 7182 14736
rect 6942 14714 6966 14716
rect 7022 14714 7046 14716
rect 7102 14714 7126 14716
rect 6964 14662 6966 14714
rect 7028 14662 7040 14714
rect 7102 14662 7104 14714
rect 6942 14660 6966 14662
rect 7022 14660 7046 14662
rect 7102 14660 7126 14662
rect 6886 14640 7182 14660
rect 9876 14550 9904 16400
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 5908 14544 5960 14550
rect 5908 14486 5960 14492
rect 9864 14544 9916 14550
rect 9864 14486 9916 14492
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 4436 14000 4488 14006
rect 4436 13942 4488 13948
rect 6104 13530 6132 14418
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 9600 13870 9628 14282
rect 9784 14074 9812 14418
rect 9852 14172 10148 14192
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 9930 14118 9932 14170
rect 9994 14118 10006 14170
rect 10068 14118 10070 14170
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 9852 14096 10148 14116
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 6886 13628 7182 13648
rect 6942 13626 6966 13628
rect 7022 13626 7046 13628
rect 7102 13626 7126 13628
rect 6964 13574 6966 13626
rect 7028 13574 7040 13626
rect 7102 13574 7104 13626
rect 6942 13572 6966 13574
rect 7022 13572 7046 13574
rect 7102 13572 7126 13574
rect 6886 13552 7182 13572
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 4252 13388 4304 13394
rect 4252 13330 4304 13336
rect 6184 13388 6236 13394
rect 6184 13330 6236 13336
rect 3921 13084 4217 13104
rect 3977 13082 4001 13084
rect 4057 13082 4081 13084
rect 4137 13082 4161 13084
rect 3999 13030 4001 13082
rect 4063 13030 4075 13082
rect 4137 13030 4139 13082
rect 3977 13028 4001 13030
rect 4057 13028 4081 13030
rect 4137 13028 4161 13030
rect 3921 13008 4217 13028
rect 5080 12912 5132 12918
rect 5080 12854 5132 12860
rect 3424 12776 3476 12782
rect 3424 12718 3476 12724
rect 1490 12679 1546 12688
rect 1860 12708 1912 12714
rect 1400 12650 1452 12656
rect 1860 12650 1912 12656
rect 2228 12708 2280 12714
rect 2228 12650 2280 12656
rect 2964 12708 3016 12714
rect 2964 12650 3016 12656
rect 1412 12073 1440 12650
rect 1676 12368 1728 12374
rect 1872 12345 1900 12650
rect 2136 12640 2188 12646
rect 2136 12582 2188 12588
rect 1676 12310 1728 12316
rect 1858 12336 1914 12345
rect 1492 12300 1544 12306
rect 1492 12242 1544 12248
rect 1398 12064 1454 12073
rect 1398 11999 1454 12008
rect 1400 11620 1452 11626
rect 1400 11562 1452 11568
rect 1412 10985 1440 11562
rect 1504 11393 1532 12242
rect 1688 11694 1716 12310
rect 1768 12300 1820 12306
rect 1858 12271 1914 12280
rect 1768 12242 1820 12248
rect 1676 11688 1728 11694
rect 1780 11665 1808 12242
rect 1860 12164 1912 12170
rect 1860 12106 1912 12112
rect 1676 11630 1728 11636
rect 1766 11656 1822 11665
rect 1490 11384 1546 11393
rect 1490 11319 1546 11328
rect 1492 11212 1544 11218
rect 1492 11154 1544 11160
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 1504 10033 1532 11154
rect 1584 11076 1636 11082
rect 1584 11018 1636 11024
rect 1490 10024 1546 10033
rect 1490 9959 1546 9968
rect 1400 9920 1452 9926
rect 1400 9862 1452 9868
rect 1412 9722 1440 9862
rect 1400 9716 1452 9722
rect 1400 9658 1452 9664
rect 1400 9444 1452 9450
rect 1400 9386 1452 9392
rect 1412 9178 1440 9386
rect 1400 9172 1452 9178
rect 1400 9114 1452 9120
rect 1412 7721 1440 9114
rect 1492 9036 1544 9042
rect 1492 8978 1544 8984
rect 1504 8401 1532 8978
rect 1490 8392 1546 8401
rect 1490 8327 1546 8336
rect 1490 8120 1546 8129
rect 1490 8055 1546 8064
rect 1504 8022 1532 8055
rect 1492 8016 1544 8022
rect 1492 7958 1544 7964
rect 1398 7712 1454 7721
rect 1398 7647 1454 7656
rect 1398 7440 1454 7449
rect 1398 7375 1454 7384
rect 1412 7342 1440 7375
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 1490 6760 1546 6769
rect 1490 6695 1546 6704
rect 1504 6254 1532 6695
rect 1492 6248 1544 6254
rect 1492 6190 1544 6196
rect 1504 5370 1532 6190
rect 1596 5778 1624 11018
rect 1688 10441 1716 11630
rect 1766 11591 1822 11600
rect 1872 11218 1900 12106
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 1952 11552 2004 11558
rect 1952 11494 2004 11500
rect 1964 11257 1992 11494
rect 1950 11248 2006 11257
rect 1860 11212 1912 11218
rect 1950 11183 2006 11192
rect 1860 11154 1912 11160
rect 1872 10713 1900 11154
rect 1952 11008 2004 11014
rect 1952 10950 2004 10956
rect 1858 10704 1914 10713
rect 1858 10639 1914 10648
rect 1674 10432 1730 10441
rect 1674 10367 1730 10376
rect 1964 10033 1992 10950
rect 1950 10024 2006 10033
rect 1950 9959 2006 9968
rect 1860 9376 1912 9382
rect 1860 9318 1912 9324
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1780 8430 1808 8774
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 1676 7812 1728 7818
rect 1676 7754 1728 7760
rect 1688 7449 1716 7754
rect 1674 7440 1730 7449
rect 1674 7375 1730 7384
rect 1674 5808 1730 5817
rect 1584 5772 1636 5778
rect 1674 5743 1730 5752
rect 1584 5714 1636 5720
rect 1492 5364 1544 5370
rect 1492 5306 1544 5312
rect 1398 4720 1454 4729
rect 1398 4655 1454 4664
rect 1582 4720 1638 4729
rect 1582 4655 1638 4664
rect 388 4276 440 4282
rect 388 4218 440 4224
rect 400 800 428 4218
rect 1412 3126 1440 4655
rect 1492 4480 1544 4486
rect 1492 4422 1544 4428
rect 1504 4185 1532 4422
rect 1490 4176 1546 4185
rect 1490 4111 1546 4120
rect 1596 4078 1624 4655
rect 1584 4072 1636 4078
rect 1584 4014 1636 4020
rect 1492 3936 1544 3942
rect 1492 3878 1544 3884
rect 1504 3505 1532 3878
rect 1490 3496 1546 3505
rect 1490 3431 1546 3440
rect 1688 3194 1716 5743
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 1780 4554 1808 4966
rect 1872 4706 1900 9318
rect 2056 8294 2084 12038
rect 2148 11694 2176 12582
rect 2780 12164 2832 12170
rect 2780 12106 2832 12112
rect 2872 12164 2924 12170
rect 2872 12106 2924 12112
rect 2228 11756 2280 11762
rect 2228 11698 2280 11704
rect 2596 11756 2648 11762
rect 2596 11698 2648 11704
rect 2136 11688 2188 11694
rect 2136 11630 2188 11636
rect 2240 11014 2268 11698
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2412 11552 2464 11558
rect 2412 11494 2464 11500
rect 2228 11008 2280 11014
rect 2228 10950 2280 10956
rect 2332 10810 2360 11494
rect 2320 10804 2372 10810
rect 2320 10746 2372 10752
rect 2424 10742 2452 11494
rect 2504 10804 2556 10810
rect 2504 10746 2556 10752
rect 2412 10736 2464 10742
rect 2412 10678 2464 10684
rect 2516 10538 2544 10746
rect 2608 10538 2636 11698
rect 2792 11694 2820 12106
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2688 11008 2740 11014
rect 2688 10950 2740 10956
rect 2504 10532 2556 10538
rect 2504 10474 2556 10480
rect 2596 10532 2648 10538
rect 2596 10474 2648 10480
rect 2226 10296 2282 10305
rect 2226 10231 2282 10240
rect 2136 9920 2188 9926
rect 2136 9862 2188 9868
rect 2148 9518 2176 9862
rect 2240 9654 2268 10231
rect 2700 10130 2728 10950
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 2228 9648 2280 9654
rect 2228 9590 2280 9596
rect 2136 9512 2188 9518
rect 2136 9454 2188 9460
rect 2700 9450 2728 10066
rect 2792 9518 2820 11494
rect 2884 10538 2912 12106
rect 2872 10532 2924 10538
rect 2872 10474 2924 10480
rect 2976 9926 3004 12650
rect 3608 12640 3660 12646
rect 3608 12582 3660 12588
rect 4804 12640 4856 12646
rect 4804 12582 4856 12588
rect 3620 12374 3648 12582
rect 3608 12368 3660 12374
rect 3608 12310 3660 12316
rect 4528 12232 4580 12238
rect 4528 12174 4580 12180
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 3056 12096 3108 12102
rect 3056 12038 3108 12044
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 4252 12096 4304 12102
rect 4252 12038 4304 12044
rect 3068 11694 3096 12038
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3528 11694 3556 11834
rect 3056 11688 3108 11694
rect 3056 11630 3108 11636
rect 3516 11688 3568 11694
rect 3516 11630 3568 11636
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 3068 9761 3096 11630
rect 3240 11552 3292 11558
rect 3240 11494 3292 11500
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3148 11212 3200 11218
rect 3148 11154 3200 11160
rect 3160 10674 3188 11154
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3160 10062 3188 10610
rect 3252 10606 3280 11494
rect 3332 11280 3384 11286
rect 3332 11222 3384 11228
rect 3240 10600 3292 10606
rect 3240 10542 3292 10548
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3054 9752 3110 9761
rect 2872 9716 2924 9722
rect 3054 9687 3110 9696
rect 2872 9658 2924 9664
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2688 9444 2740 9450
rect 2688 9386 2740 9392
rect 2884 9110 2912 9658
rect 3252 9518 3280 10406
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 3148 9444 3200 9450
rect 3148 9386 3200 9392
rect 2872 9104 2924 9110
rect 2872 9046 2924 9052
rect 3160 8838 3188 9386
rect 3344 9178 3372 11222
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3436 9110 3464 11494
rect 3528 10470 3556 11630
rect 3620 11558 3648 12038
rect 3921 11996 4217 12016
rect 3977 11994 4001 11996
rect 4057 11994 4081 11996
rect 4137 11994 4161 11996
rect 3999 11942 4001 11994
rect 4063 11942 4075 11994
rect 4137 11942 4139 11994
rect 3977 11940 4001 11942
rect 4057 11940 4081 11942
rect 4137 11940 4161 11942
rect 3921 11920 4217 11940
rect 4264 11694 4292 12038
rect 3976 11688 4028 11694
rect 3974 11656 3976 11665
rect 4252 11688 4304 11694
rect 4028 11656 4030 11665
rect 4252 11630 4304 11636
rect 3974 11591 4030 11600
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3516 9920 3568 9926
rect 3516 9862 3568 9868
rect 3528 9586 3556 9862
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3424 9104 3476 9110
rect 3424 9046 3476 9052
rect 3332 9036 3384 9042
rect 3332 8978 3384 8984
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 3240 8832 3292 8838
rect 3344 8809 3372 8978
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3436 8820 3464 8910
rect 3516 8832 3568 8838
rect 3240 8774 3292 8780
rect 3330 8800 3386 8809
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2596 8424 2648 8430
rect 2596 8366 2648 8372
rect 2044 8288 2096 8294
rect 2044 8230 2096 8236
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 2044 7744 2096 7750
rect 2044 7686 2096 7692
rect 2136 7744 2188 7750
rect 2136 7686 2188 7692
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 1964 5556 1992 7482
rect 2056 7342 2084 7686
rect 2148 7342 2176 7686
rect 2044 7336 2096 7342
rect 2044 7278 2096 7284
rect 2136 7336 2188 7342
rect 2136 7278 2188 7284
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 1964 5528 2084 5556
rect 2056 5273 2084 5528
rect 2042 5264 2098 5273
rect 2042 5199 2098 5208
rect 1952 5024 2004 5030
rect 1952 4966 2004 4972
rect 1964 4826 1992 4966
rect 2056 4826 2084 5199
rect 2148 5166 2176 6598
rect 2332 6458 2360 7822
rect 2608 7818 2636 8366
rect 2700 8362 2728 8570
rect 3252 8537 3280 8774
rect 3330 8735 3386 8744
rect 3436 8792 3516 8820
rect 3436 8650 3464 8792
rect 3516 8774 3568 8780
rect 3344 8622 3464 8650
rect 3238 8528 3294 8537
rect 3238 8463 3294 8472
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2780 8356 2832 8362
rect 2780 8298 2832 8304
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 2596 7812 2648 7818
rect 2596 7754 2648 7760
rect 2504 7472 2556 7478
rect 2504 7414 2556 7420
rect 2320 6452 2372 6458
rect 2320 6394 2372 6400
rect 2410 6216 2466 6225
rect 2410 6151 2466 6160
rect 2318 5808 2374 5817
rect 2424 5778 2452 6151
rect 2318 5743 2374 5752
rect 2412 5772 2464 5778
rect 2136 5160 2188 5166
rect 2332 5114 2360 5743
rect 2412 5714 2464 5720
rect 2410 5400 2466 5409
rect 2410 5335 2466 5344
rect 2136 5102 2188 5108
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 2044 4820 2096 4826
rect 2044 4762 2096 4768
rect 2148 4706 2176 5102
rect 1872 4678 1992 4706
rect 1768 4548 1820 4554
rect 1768 4490 1820 4496
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 1872 3777 1900 3878
rect 1858 3768 1914 3777
rect 1858 3703 1914 3712
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 1400 3120 1452 3126
rect 1400 3062 1452 3068
rect 1964 2990 1992 4678
rect 2056 4678 2176 4706
rect 2240 5086 2360 5114
rect 2056 3602 2084 4678
rect 2134 4448 2190 4457
rect 2134 4383 2190 4392
rect 2148 4146 2176 4383
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2044 3596 2096 3602
rect 2044 3538 2096 3544
rect 1952 2984 2004 2990
rect 1952 2926 2004 2932
rect 2240 2922 2268 5086
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 2332 4622 2360 4966
rect 2320 4616 2372 4622
rect 2320 4558 2372 4564
rect 2332 3738 2360 4558
rect 2424 4214 2452 5335
rect 2412 4208 2464 4214
rect 2412 4150 2464 4156
rect 2516 4010 2544 7414
rect 2596 7200 2648 7206
rect 2596 7142 2648 7148
rect 2608 6254 2636 7142
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 2596 6112 2648 6118
rect 2596 6054 2648 6060
rect 2608 5846 2636 6054
rect 2596 5840 2648 5846
rect 2596 5782 2648 5788
rect 2700 5760 2728 7890
rect 2792 7410 2820 8298
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 3160 7546 3188 7822
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 3056 7200 3108 7206
rect 3056 7142 3108 7148
rect 2870 7032 2926 7041
rect 2976 7002 3004 7142
rect 2870 6967 2926 6976
rect 2964 6996 3016 7002
rect 2780 6384 2832 6390
rect 2778 6352 2780 6361
rect 2832 6352 2834 6361
rect 2778 6287 2834 6296
rect 2884 5778 2912 6967
rect 2964 6938 3016 6944
rect 3068 6730 3096 7142
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 3160 6662 3188 7346
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 2976 6186 3004 6598
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 2964 6180 3016 6186
rect 2964 6122 3016 6128
rect 2962 5944 3018 5953
rect 2962 5879 3018 5888
rect 2872 5772 2924 5778
rect 2700 5732 2820 5760
rect 2686 5672 2742 5681
rect 2686 5607 2688 5616
rect 2740 5607 2742 5616
rect 2688 5578 2740 5584
rect 2792 4826 2820 5732
rect 2872 5714 2924 5720
rect 2976 5642 3004 5879
rect 3068 5817 3096 6394
rect 3148 6384 3200 6390
rect 3148 6326 3200 6332
rect 3054 5808 3110 5817
rect 3054 5743 3110 5752
rect 2964 5636 3016 5642
rect 2964 5578 3016 5584
rect 2872 5568 2924 5574
rect 2870 5536 2872 5545
rect 2924 5536 2926 5545
rect 2870 5471 2926 5480
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 3160 4622 3188 6326
rect 3252 5710 3280 6734
rect 3240 5704 3292 5710
rect 3240 5646 3292 5652
rect 3252 5166 3280 5646
rect 3240 5160 3292 5166
rect 3240 5102 3292 5108
rect 3252 5030 3280 5102
rect 3240 5024 3292 5030
rect 3240 4966 3292 4972
rect 3148 4616 3200 4622
rect 2594 4584 2650 4593
rect 3068 4576 3148 4604
rect 2594 4519 2650 4528
rect 2872 4548 2924 4554
rect 2608 4146 2636 4519
rect 2872 4490 2924 4496
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 2594 4040 2650 4049
rect 2504 4004 2556 4010
rect 2594 3975 2650 3984
rect 2504 3946 2556 3952
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2608 3670 2636 3975
rect 2596 3664 2648 3670
rect 2596 3606 2648 3612
rect 2884 3074 2912 4490
rect 3068 4185 3096 4576
rect 3148 4558 3200 4564
rect 3344 4282 3372 8622
rect 3620 8514 3648 11494
rect 3792 11144 3844 11150
rect 3792 11086 3844 11092
rect 3804 10606 3832 11086
rect 3921 10908 4217 10928
rect 3977 10906 4001 10908
rect 4057 10906 4081 10908
rect 4137 10906 4161 10908
rect 3999 10854 4001 10906
rect 4063 10854 4075 10906
rect 4137 10854 4139 10906
rect 3977 10852 4001 10854
rect 4057 10852 4081 10854
rect 4137 10852 4161 10854
rect 3921 10832 4217 10852
rect 4264 10690 4292 11494
rect 4540 11354 4568 12174
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4528 11144 4580 11150
rect 4528 11086 4580 11092
rect 4344 11076 4396 11082
rect 4344 11018 4396 11024
rect 4436 11076 4488 11082
rect 4436 11018 4488 11024
rect 4172 10662 4292 10690
rect 3792 10600 3844 10606
rect 3792 10542 3844 10548
rect 3804 10282 3832 10542
rect 3712 10254 3832 10282
rect 3712 10130 3740 10254
rect 3700 10124 3752 10130
rect 3700 10066 3752 10072
rect 3792 10124 3844 10130
rect 3792 10066 3844 10072
rect 3700 9376 3752 9382
rect 3804 9353 3832 10066
rect 4172 10062 4200 10662
rect 4252 10532 4304 10538
rect 4252 10474 4304 10480
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 3921 9820 4217 9840
rect 3977 9818 4001 9820
rect 4057 9818 4081 9820
rect 4137 9818 4161 9820
rect 3999 9766 4001 9818
rect 4063 9766 4075 9818
rect 4137 9766 4139 9818
rect 3977 9764 4001 9766
rect 4057 9764 4081 9766
rect 4137 9764 4161 9766
rect 3921 9744 4217 9764
rect 4264 9654 4292 10474
rect 4252 9648 4304 9654
rect 4252 9590 4304 9596
rect 4356 9518 4384 11018
rect 4448 10130 4476 11018
rect 4436 10124 4488 10130
rect 4436 10066 4488 10072
rect 4434 10024 4490 10033
rect 4434 9959 4490 9968
rect 4448 9586 4476 9959
rect 4436 9580 4488 9586
rect 4436 9522 4488 9528
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 4344 9512 4396 9518
rect 4344 9454 4396 9460
rect 3700 9318 3752 9324
rect 3790 9344 3846 9353
rect 3712 8786 3740 9318
rect 3790 9279 3846 9288
rect 3896 9081 3924 9454
rect 4066 9344 4122 9353
rect 4066 9279 4122 9288
rect 3882 9072 3938 9081
rect 3882 9007 3938 9016
rect 4080 8974 4108 9279
rect 4160 9104 4212 9110
rect 4448 9081 4476 9522
rect 4540 9178 4568 11086
rect 4632 9382 4660 12174
rect 4816 12102 4844 12582
rect 4804 12096 4856 12102
rect 4802 12064 4804 12073
rect 4856 12064 4858 12073
rect 5092 12050 5120 12854
rect 5264 12436 5316 12442
rect 5368 12434 5856 12458
rect 5316 12430 5856 12434
rect 5316 12406 5396 12430
rect 5264 12378 5316 12384
rect 5356 12232 5408 12238
rect 5356 12174 5408 12180
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5092 12022 5304 12050
rect 4802 11999 4858 12008
rect 4816 11973 4844 11999
rect 5170 11928 5226 11937
rect 5170 11863 5226 11872
rect 4988 11688 5040 11694
rect 4988 11630 5040 11636
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4724 10169 4752 11086
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4816 10266 4844 10950
rect 4896 10532 4948 10538
rect 4896 10474 4948 10480
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4710 10160 4766 10169
rect 4710 10095 4766 10104
rect 4816 10033 4844 10202
rect 4908 10062 4936 10474
rect 4896 10056 4948 10062
rect 4802 10024 4858 10033
rect 4712 9988 4764 9994
rect 4896 9998 4948 10004
rect 4802 9959 4858 9968
rect 4712 9930 4764 9936
rect 4724 9489 4752 9930
rect 4816 9568 4844 9959
rect 4908 9761 4936 9998
rect 4894 9752 4950 9761
rect 4894 9687 4896 9696
rect 4948 9687 4950 9696
rect 4896 9658 4948 9664
rect 4816 9540 4936 9568
rect 4710 9480 4766 9489
rect 4710 9415 4766 9424
rect 4804 9444 4856 9450
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 4160 9046 4212 9052
rect 4434 9072 4490 9081
rect 4068 8968 4120 8974
rect 4172 8945 4200 9046
rect 4252 9036 4304 9042
rect 4632 9058 4660 9318
rect 4434 9007 4490 9016
rect 4540 9030 4660 9058
rect 4252 8978 4304 8984
rect 4068 8910 4120 8916
rect 4158 8936 4214 8945
rect 4158 8871 4214 8880
rect 3712 8758 3832 8786
rect 3700 8628 3752 8634
rect 3700 8570 3752 8576
rect 3436 8486 3648 8514
rect 3436 7449 3464 8486
rect 3608 8356 3660 8362
rect 3608 8298 3660 8304
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3422 7440 3478 7449
rect 3422 7375 3478 7384
rect 3436 5953 3464 7375
rect 3422 5944 3478 5953
rect 3422 5879 3478 5888
rect 3528 5794 3556 8026
rect 3620 7954 3648 8298
rect 3712 8022 3740 8570
rect 3804 8362 3832 8758
rect 3921 8732 4217 8752
rect 3977 8730 4001 8732
rect 4057 8730 4081 8732
rect 4137 8730 4161 8732
rect 3999 8678 4001 8730
rect 4063 8678 4075 8730
rect 4137 8678 4139 8730
rect 3977 8676 4001 8678
rect 4057 8676 4081 8678
rect 4137 8676 4161 8678
rect 3921 8656 4217 8676
rect 3792 8356 3844 8362
rect 3792 8298 3844 8304
rect 4068 8288 4120 8294
rect 3974 8256 4030 8265
rect 4068 8230 4120 8236
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 3974 8191 4030 8200
rect 3700 8016 3752 8022
rect 3700 7958 3752 7964
rect 3988 7954 4016 8191
rect 4080 8090 4108 8230
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 3608 7948 3660 7954
rect 3608 7890 3660 7896
rect 3976 7948 4028 7954
rect 3976 7890 4028 7896
rect 3620 7410 3648 7890
rect 4172 7886 4200 8230
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 3700 7744 3752 7750
rect 3700 7686 3752 7692
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3606 6488 3662 6497
rect 3606 6423 3662 6432
rect 3620 6254 3648 6423
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3528 5766 3648 5794
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 3424 5636 3476 5642
rect 3424 5578 3476 5584
rect 3436 5545 3464 5578
rect 3422 5536 3478 5545
rect 3422 5471 3478 5480
rect 3528 5098 3556 5646
rect 3620 5302 3648 5766
rect 3608 5296 3660 5302
rect 3608 5238 3660 5244
rect 3516 5092 3568 5098
rect 3516 5034 3568 5040
rect 3528 4622 3556 5034
rect 3620 4690 3648 5238
rect 3712 5098 3740 7686
rect 3804 7410 3832 7686
rect 3921 7644 4217 7664
rect 3977 7642 4001 7644
rect 4057 7642 4081 7644
rect 4137 7642 4161 7644
rect 3999 7590 4001 7642
rect 4063 7590 4075 7642
rect 4137 7590 4139 7642
rect 3977 7588 4001 7590
rect 4057 7588 4081 7590
rect 4137 7588 4161 7590
rect 3921 7568 4217 7588
rect 4264 7546 4292 8978
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3988 7002 4016 7346
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 4080 6934 4108 7278
rect 4068 6928 4120 6934
rect 4068 6870 4120 6876
rect 4172 6866 4200 7278
rect 4356 7274 4384 8910
rect 4448 8430 4476 8910
rect 4436 8424 4488 8430
rect 4436 8366 4488 8372
rect 4434 8256 4490 8265
rect 4434 8191 4490 8200
rect 4344 7268 4396 7274
rect 4344 7210 4396 7216
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3804 6089 3832 6598
rect 3921 6556 4217 6576
rect 3977 6554 4001 6556
rect 4057 6554 4081 6556
rect 4137 6554 4161 6556
rect 3999 6502 4001 6554
rect 4063 6502 4075 6554
rect 4137 6502 4139 6554
rect 3977 6500 4001 6502
rect 4057 6500 4081 6502
rect 4137 6500 4161 6502
rect 3921 6480 4217 6500
rect 4342 6488 4398 6497
rect 4342 6423 4398 6432
rect 4356 6254 4384 6423
rect 4344 6248 4396 6254
rect 4344 6190 4396 6196
rect 3976 6180 4028 6186
rect 3976 6122 4028 6128
rect 3790 6080 3846 6089
rect 3790 6015 3846 6024
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3700 5092 3752 5098
rect 3700 5034 3752 5040
rect 3804 4690 3832 5850
rect 3988 5846 4016 6122
rect 4160 6112 4212 6118
rect 4080 6072 4160 6100
rect 3976 5840 4028 5846
rect 3976 5782 4028 5788
rect 4080 5778 4108 6072
rect 4160 6054 4212 6060
rect 4356 5794 4384 6190
rect 4448 5914 4476 8191
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4068 5772 4120 5778
rect 4356 5766 4476 5794
rect 4068 5714 4120 5720
rect 4344 5704 4396 5710
rect 4250 5672 4306 5681
rect 4344 5646 4396 5652
rect 4250 5607 4252 5616
rect 4304 5607 4306 5616
rect 4252 5578 4304 5584
rect 3921 5468 4217 5488
rect 3977 5466 4001 5468
rect 4057 5466 4081 5468
rect 4137 5466 4161 5468
rect 3999 5414 4001 5466
rect 4063 5414 4075 5466
rect 4137 5414 4139 5466
rect 3977 5412 4001 5414
rect 4057 5412 4081 5414
rect 4137 5412 4161 5414
rect 3921 5392 4217 5412
rect 4356 5370 4384 5646
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 3884 5160 3936 5166
rect 3882 5128 3884 5137
rect 3936 5128 3938 5137
rect 3882 5063 3938 5072
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 4172 4758 4200 5034
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 4160 4752 4212 4758
rect 4160 4694 4212 4700
rect 3608 4684 3660 4690
rect 3608 4626 3660 4632
rect 3792 4684 3844 4690
rect 3792 4626 3844 4632
rect 3516 4616 3568 4622
rect 3516 4558 3568 4564
rect 3608 4480 3660 4486
rect 3608 4422 3660 4428
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 3054 4176 3110 4185
rect 3054 4111 3110 4120
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 2976 3913 3004 4014
rect 2962 3904 3018 3913
rect 2962 3839 3018 3848
rect 2976 3602 3004 3839
rect 2964 3596 3016 3602
rect 2964 3538 3016 3544
rect 2964 3188 3016 3194
rect 2964 3130 3016 3136
rect 2792 3046 2912 3074
rect 2792 2990 2820 3046
rect 2320 2984 2372 2990
rect 2318 2952 2320 2961
rect 2780 2984 2832 2990
rect 2372 2952 2374 2961
rect 2228 2916 2280 2922
rect 2780 2926 2832 2932
rect 2318 2887 2374 2896
rect 2228 2858 2280 2864
rect 2686 2680 2742 2689
rect 2686 2615 2742 2624
rect 2872 2644 2924 2650
rect 2700 2514 2728 2615
rect 2872 2586 2924 2592
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 2320 2508 2372 2514
rect 2320 2450 2372 2456
rect 2688 2508 2740 2514
rect 2688 2450 2740 2456
rect 1216 2372 1268 2378
rect 1216 2314 1268 2320
rect 1228 800 1256 2314
rect 1596 2038 1624 2450
rect 2136 2372 2188 2378
rect 2136 2314 2188 2320
rect 1584 2032 1636 2038
rect 1584 1974 1636 1980
rect 2148 800 2176 2314
rect 2332 1970 2360 2450
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 2320 1964 2372 1970
rect 2320 1906 2372 1912
rect 386 0 442 800
rect 1214 0 1270 800
rect 2134 0 2190 800
rect 2792 241 2820 2382
rect 2884 513 2912 2586
rect 2976 1193 3004 3130
rect 3068 2650 3096 4111
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 3528 3942 3556 4014
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 3424 3596 3476 3602
rect 3424 3538 3476 3544
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 3252 3194 3280 3470
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3436 3097 3464 3538
rect 3422 3088 3478 3097
rect 3148 3052 3200 3058
rect 3422 3023 3478 3032
rect 3148 2994 3200 3000
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 3056 2372 3108 2378
rect 3056 2314 3108 2320
rect 2962 1184 3018 1193
rect 2962 1119 3018 1128
rect 3068 800 3096 2314
rect 3160 1465 3188 2994
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 3252 1873 3280 2926
rect 3332 2848 3384 2854
rect 3332 2790 3384 2796
rect 3344 2145 3372 2790
rect 3620 2582 3648 4422
rect 3921 4380 4217 4400
rect 3977 4378 4001 4380
rect 4057 4378 4081 4380
rect 4137 4378 4161 4380
rect 3999 4326 4001 4378
rect 4063 4326 4075 4378
rect 4137 4326 4139 4378
rect 3977 4324 4001 4326
rect 4057 4324 4081 4326
rect 4137 4324 4161 4326
rect 3921 4304 4217 4324
rect 4160 4208 4212 4214
rect 4160 4150 4212 4156
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3988 4010 4016 4082
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 4068 4004 4120 4010
rect 4068 3946 4120 3952
rect 3976 3664 4028 3670
rect 4080 3652 4108 3946
rect 4172 3913 4200 4150
rect 4158 3904 4214 3913
rect 4158 3839 4214 3848
rect 4028 3624 4108 3652
rect 3976 3606 4028 3612
rect 4172 3534 4200 3839
rect 4160 3528 4212 3534
rect 3698 3496 3754 3505
rect 4160 3470 4212 3476
rect 3698 3431 3754 3440
rect 3712 3398 3740 3431
rect 3700 3392 3752 3398
rect 3700 3334 3752 3340
rect 3792 3392 3844 3398
rect 3792 3334 3844 3340
rect 3700 2848 3752 2854
rect 3804 2825 3832 3334
rect 3921 3292 4217 3312
rect 3977 3290 4001 3292
rect 4057 3290 4081 3292
rect 4137 3290 4161 3292
rect 3999 3238 4001 3290
rect 4063 3238 4075 3290
rect 4137 3238 4139 3290
rect 3977 3236 4001 3238
rect 4057 3236 4081 3238
rect 4137 3236 4161 3238
rect 3921 3216 4217 3236
rect 4264 2990 4292 4966
rect 4448 4214 4476 5766
rect 4540 5166 4568 9030
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 4528 4480 4580 4486
rect 4528 4422 4580 4428
rect 4436 4208 4488 4214
rect 4436 4150 4488 4156
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4436 3936 4488 3942
rect 4436 3878 4488 3884
rect 4356 3670 4384 3878
rect 4344 3664 4396 3670
rect 4344 3606 4396 3612
rect 4344 3392 4396 3398
rect 4344 3334 4396 3340
rect 4252 2984 4304 2990
rect 4252 2926 4304 2932
rect 3700 2790 3752 2796
rect 3790 2816 3846 2825
rect 3608 2576 3660 2582
rect 3608 2518 3660 2524
rect 3516 2508 3568 2514
rect 3516 2450 3568 2456
rect 3424 2372 3476 2378
rect 3424 2314 3476 2320
rect 3330 2136 3386 2145
rect 3330 2071 3386 2080
rect 3238 1864 3294 1873
rect 3238 1799 3294 1808
rect 3146 1456 3202 1465
rect 3146 1391 3202 1400
rect 2870 504 2926 513
rect 2870 439 2926 448
rect 2778 232 2834 241
rect 2778 167 2834 176
rect 3054 0 3110 800
rect 3436 785 3464 2314
rect 3528 1766 3556 2450
rect 3712 2417 3740 2790
rect 3790 2751 3846 2760
rect 4356 2650 4384 3334
rect 4448 2990 4476 3878
rect 4540 3058 4568 4422
rect 4632 4049 4660 8774
rect 4724 7206 4752 9415
rect 4804 9386 4856 9392
rect 4816 7546 4844 9386
rect 4908 7993 4936 9540
rect 4894 7984 4950 7993
rect 4894 7919 4950 7928
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 4908 7449 4936 7686
rect 4894 7440 4950 7449
rect 4894 7375 4950 7384
rect 5000 7342 5028 11630
rect 5080 11008 5132 11014
rect 5080 10950 5132 10956
rect 5092 10305 5120 10950
rect 5078 10296 5134 10305
rect 5078 10231 5080 10240
rect 5132 10231 5134 10240
rect 5080 10202 5132 10208
rect 5092 9926 5120 10202
rect 5080 9920 5132 9926
rect 5080 9862 5132 9868
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 5092 9353 5120 9522
rect 5078 9344 5134 9353
rect 5078 9279 5134 9288
rect 5092 8430 5120 9279
rect 5080 8424 5132 8430
rect 5080 8366 5132 8372
rect 5184 8265 5212 11863
rect 5276 9586 5304 12022
rect 5368 11937 5396 12174
rect 5354 11928 5410 11937
rect 5354 11863 5410 11872
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5448 11688 5500 11694
rect 5448 11630 5500 11636
rect 5356 11620 5408 11626
rect 5356 11562 5408 11568
rect 5368 10169 5396 11562
rect 5460 10742 5488 11630
rect 5448 10736 5500 10742
rect 5448 10678 5500 10684
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 5354 10160 5410 10169
rect 5354 10095 5410 10104
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5170 8256 5226 8265
rect 5170 8191 5226 8200
rect 5276 8090 5304 9318
rect 5368 8294 5396 10095
rect 5460 9722 5488 10542
rect 5552 10198 5580 11834
rect 5644 11694 5672 12174
rect 5724 12096 5776 12102
rect 5724 12038 5776 12044
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5644 10130 5672 11630
rect 5736 11626 5764 12038
rect 5724 11620 5776 11626
rect 5724 11562 5776 11568
rect 5724 11076 5776 11082
rect 5724 11018 5776 11024
rect 5736 10674 5764 11018
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 5722 10568 5778 10577
rect 5828 10554 5856 12430
rect 5908 12436 5960 12442
rect 6196 12434 6224 13330
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 6886 12540 7182 12560
rect 6942 12538 6966 12540
rect 7022 12538 7046 12540
rect 7102 12538 7126 12540
rect 6964 12486 6966 12538
rect 7028 12486 7040 12538
rect 7102 12486 7104 12538
rect 6942 12484 6966 12486
rect 7022 12484 7046 12486
rect 7102 12484 7126 12486
rect 6886 12464 7182 12484
rect 7852 12434 7880 13126
rect 9852 13084 10148 13104
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 9930 13030 9932 13082
rect 9994 13030 10006 13082
rect 10068 13030 10070 13082
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 9852 13008 10148 13028
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 8116 12708 8168 12714
rect 8116 12650 8168 12656
rect 8128 12434 8156 12650
rect 8496 12434 8524 12922
rect 9772 12912 9824 12918
rect 9772 12854 9824 12860
rect 10232 12912 10284 12918
rect 10232 12854 10284 12860
rect 11520 12912 11572 12918
rect 11520 12854 11572 12860
rect 9036 12640 9088 12646
rect 9036 12582 9088 12588
rect 6196 12406 6408 12434
rect 7852 12406 7972 12434
rect 5908 12378 5960 12384
rect 5920 12345 5948 12378
rect 5906 12336 5962 12345
rect 5906 12271 5962 12280
rect 6184 12300 6236 12306
rect 5920 10713 5948 12271
rect 6184 12242 6236 12248
rect 6196 12102 6224 12242
rect 6184 12096 6236 12102
rect 6184 12038 6236 12044
rect 6196 11801 6224 12038
rect 6182 11792 6238 11801
rect 6092 11756 6144 11762
rect 6182 11727 6238 11736
rect 6092 11698 6144 11704
rect 6104 11354 6132 11698
rect 6092 11348 6144 11354
rect 6092 11290 6144 11296
rect 6104 10985 6132 11290
rect 6090 10976 6146 10985
rect 6090 10911 6146 10920
rect 6196 10810 6224 11727
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 6288 11121 6316 11494
rect 6274 11112 6330 11121
rect 6274 11047 6330 11056
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 5906 10704 5962 10713
rect 5906 10639 5962 10648
rect 5828 10526 5948 10554
rect 5722 10503 5778 10512
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5552 9761 5580 9998
rect 5538 9752 5594 9761
rect 5448 9716 5500 9722
rect 5538 9687 5594 9696
rect 5448 9658 5500 9664
rect 5460 9178 5488 9658
rect 5630 9616 5686 9625
rect 5630 9551 5632 9560
rect 5684 9551 5686 9560
rect 5632 9522 5684 9528
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5552 9081 5580 9454
rect 5538 9072 5594 9081
rect 5538 9007 5594 9016
rect 5644 8922 5672 9522
rect 5460 8894 5672 8922
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 4896 7268 4948 7274
rect 4896 7210 4948 7216
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4908 7002 4936 7210
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 4816 4690 4844 5510
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4804 4548 4856 4554
rect 4804 4490 4856 4496
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 4618 4040 4674 4049
rect 4724 4010 4752 4422
rect 4618 3975 4674 3984
rect 4712 4004 4764 4010
rect 4712 3946 4764 3952
rect 4620 3936 4672 3942
rect 4618 3904 4620 3913
rect 4672 3904 4674 3913
rect 4618 3839 4674 3848
rect 4620 3664 4672 3670
rect 4620 3606 4672 3612
rect 4632 3058 4660 3606
rect 4528 3052 4580 3058
rect 4528 2994 4580 3000
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4436 2984 4488 2990
rect 4436 2926 4488 2932
rect 4632 2774 4660 2994
rect 4816 2990 4844 4490
rect 4908 3058 4936 6938
rect 5092 6882 5120 7822
rect 5184 7002 5212 8026
rect 5262 7984 5318 7993
rect 5262 7919 5318 7928
rect 5172 6996 5224 7002
rect 5172 6938 5224 6944
rect 5092 6854 5212 6882
rect 5080 5024 5132 5030
rect 5080 4966 5132 4972
rect 5092 4604 5120 4966
rect 5184 4758 5212 6854
rect 5276 6100 5304 7919
rect 5460 7274 5488 8894
rect 5736 8378 5764 10503
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5828 9994 5856 10406
rect 5920 10266 5948 10526
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 5816 9988 5868 9994
rect 5816 9930 5868 9936
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 5828 9382 5856 9454
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5920 9194 5948 10202
rect 5644 8350 5764 8378
rect 5828 9166 5948 9194
rect 5644 7886 5672 8350
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5448 7268 5500 7274
rect 5448 7210 5500 7216
rect 5540 7268 5592 7274
rect 5540 7210 5592 7216
rect 5448 6656 5500 6662
rect 5552 6610 5580 7210
rect 5500 6604 5580 6610
rect 5448 6598 5580 6604
rect 5460 6582 5580 6598
rect 5356 6384 5408 6390
rect 5356 6326 5408 6332
rect 5368 6225 5396 6326
rect 5354 6216 5410 6225
rect 5552 6202 5580 6582
rect 5736 6497 5764 8230
rect 5828 8090 5856 9166
rect 5908 9104 5960 9110
rect 5908 9046 5960 9052
rect 5920 8566 5948 9046
rect 5908 8560 5960 8566
rect 5908 8502 5960 8508
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 5828 7993 5856 8026
rect 5920 8022 5948 8502
rect 5908 8016 5960 8022
rect 5814 7984 5870 7993
rect 5908 7958 5960 7964
rect 6012 7954 6040 10746
rect 6184 10600 6236 10606
rect 6184 10542 6236 10548
rect 6092 10192 6144 10198
rect 6090 10160 6092 10169
rect 6144 10160 6146 10169
rect 6090 10095 6146 10104
rect 6196 9761 6224 10542
rect 6276 10464 6328 10470
rect 6276 10406 6328 10412
rect 6182 9752 6238 9761
rect 6182 9687 6238 9696
rect 6092 9512 6144 9518
rect 6092 9454 6144 9460
rect 6104 9110 6132 9454
rect 6184 9444 6236 9450
rect 6184 9386 6236 9392
rect 6092 9104 6144 9110
rect 6092 9046 6144 9052
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 6104 8090 6132 8230
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 5814 7919 5870 7928
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5828 6866 5856 7482
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 5722 6488 5778 6497
rect 5722 6423 5778 6432
rect 6012 6254 6040 7686
rect 6196 7478 6224 9386
rect 6288 9042 6316 10406
rect 6380 10266 6408 12406
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 6550 12200 6606 12209
rect 6550 12135 6606 12144
rect 6564 12102 6592 12135
rect 6460 12096 6512 12102
rect 6460 12038 6512 12044
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6472 11626 6500 12038
rect 6564 11898 6592 12038
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 7760 11762 7788 12242
rect 7840 12232 7892 12238
rect 7838 12200 7840 12209
rect 7892 12200 7894 12209
rect 7838 12135 7894 12144
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 6460 11620 6512 11626
rect 6460 11562 6512 11568
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6472 10606 6500 10950
rect 6564 10606 6592 11698
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 6460 10600 6512 10606
rect 6460 10542 6512 10548
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6380 9450 6408 9998
rect 6472 9722 6500 10542
rect 6656 10305 6684 11630
rect 7288 11620 7340 11626
rect 7288 11562 7340 11568
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6642 10296 6698 10305
rect 6552 10260 6604 10266
rect 6642 10231 6698 10240
rect 6552 10202 6604 10208
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6472 9518 6500 9658
rect 6460 9512 6512 9518
rect 6460 9454 6512 9460
rect 6368 9444 6420 9450
rect 6368 9386 6420 9392
rect 6380 9178 6408 9386
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 6276 7812 6328 7818
rect 6276 7754 6328 7760
rect 6184 7472 6236 7478
rect 6184 7414 6236 7420
rect 6288 7410 6316 7754
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6000 6248 6052 6254
rect 5552 6174 5672 6202
rect 6000 6190 6052 6196
rect 5354 6151 5410 6160
rect 5540 6112 5592 6118
rect 5276 6072 5396 6100
rect 5368 5710 5396 6072
rect 5540 6054 5592 6060
rect 5552 5710 5580 6054
rect 5644 5710 5672 6174
rect 6092 6180 6144 6186
rect 6092 6122 6144 6128
rect 6104 5914 6132 6122
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 5368 4808 5396 5646
rect 5552 5098 5580 5646
rect 5540 5092 5592 5098
rect 5540 5034 5592 5040
rect 5920 4826 5948 5646
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 6000 5296 6052 5302
rect 6000 5238 6052 5244
rect 5908 4820 5960 4826
rect 5368 4780 5580 4808
rect 5172 4752 5224 4758
rect 5172 4694 5224 4700
rect 5354 4720 5410 4729
rect 5354 4655 5410 4664
rect 5448 4684 5500 4690
rect 5368 4622 5396 4655
rect 5448 4626 5500 4632
rect 5172 4616 5224 4622
rect 5092 4576 5172 4604
rect 5172 4558 5224 4564
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5184 4282 5212 4558
rect 5264 4548 5316 4554
rect 5264 4490 5316 4496
rect 5276 4457 5304 4490
rect 5262 4448 5318 4457
rect 5262 4383 5318 4392
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 5356 4208 5408 4214
rect 5356 4150 5408 4156
rect 5264 4004 5316 4010
rect 5264 3946 5316 3952
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 5092 3738 5120 3878
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5000 3398 5028 3674
rect 5276 3670 5304 3946
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5184 3505 5212 3538
rect 5170 3496 5226 3505
rect 5170 3431 5226 3440
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 4632 2746 4752 2774
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 4344 2508 4396 2514
rect 4344 2450 4396 2456
rect 3698 2408 3754 2417
rect 3698 2343 3754 2352
rect 3792 2372 3844 2378
rect 3792 2314 3844 2320
rect 3516 1760 3568 1766
rect 3516 1702 3568 1708
rect 3804 1170 3832 2314
rect 3921 2204 4217 2224
rect 3977 2202 4001 2204
rect 4057 2202 4081 2204
rect 4137 2202 4161 2204
rect 3999 2150 4001 2202
rect 4063 2150 4075 2202
rect 4137 2150 4139 2202
rect 3977 2148 4001 2150
rect 4057 2148 4081 2150
rect 4137 2148 4161 2150
rect 3921 2128 4217 2148
rect 4356 1834 4384 2450
rect 4724 2446 4752 2746
rect 5092 2650 5120 2790
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 5368 2582 5396 4150
rect 5460 2774 5488 4626
rect 5552 2990 5580 4780
rect 5908 4762 5960 4768
rect 6012 4593 6040 5238
rect 6104 5166 6132 5510
rect 6092 5160 6144 5166
rect 6092 5102 6144 5108
rect 5998 4584 6054 4593
rect 5998 4519 6054 4528
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 5814 4448 5870 4457
rect 5736 4078 5764 4422
rect 5814 4383 5870 4392
rect 5828 4146 5856 4383
rect 6104 4146 6132 5102
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 6092 4140 6144 4146
rect 6092 4082 6144 4088
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5630 3088 5686 3097
rect 5630 3023 5686 3032
rect 5540 2984 5592 2990
rect 5540 2926 5592 2932
rect 5644 2854 5672 3023
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5828 2774 5856 4082
rect 5920 3058 5948 4082
rect 6000 3596 6052 3602
rect 6000 3538 6052 3544
rect 6012 3398 6040 3538
rect 6104 3534 6132 4082
rect 6196 4078 6224 5714
rect 6288 4622 6316 6598
rect 6276 4616 6328 4622
rect 6380 4593 6408 8774
rect 6472 8650 6500 9454
rect 6564 8838 6592 10202
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6472 8622 6592 8650
rect 6564 8362 6592 8622
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6472 7342 6500 7822
rect 6564 7750 6592 8298
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6460 7336 6512 7342
rect 6460 7278 6512 7284
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6472 6254 6500 7142
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 6564 6322 6592 6802
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6460 6248 6512 6254
rect 6460 6190 6512 6196
rect 6472 5302 6500 6190
rect 6564 5914 6592 6258
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 6460 5160 6512 5166
rect 6458 5128 6460 5137
rect 6512 5128 6514 5137
rect 6458 5063 6514 5072
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6276 4558 6328 4564
rect 6366 4584 6422 4593
rect 6366 4519 6422 4528
rect 6472 4468 6500 4626
rect 6564 4622 6592 5850
rect 6656 5778 6684 10066
rect 6748 9178 6776 11494
rect 6886 11452 7182 11472
rect 6942 11450 6966 11452
rect 7022 11450 7046 11452
rect 7102 11450 7126 11452
rect 6964 11398 6966 11450
rect 7028 11398 7040 11450
rect 7102 11398 7104 11450
rect 6942 11396 6966 11398
rect 7022 11396 7046 11398
rect 7102 11396 7126 11398
rect 6886 11376 7182 11396
rect 7300 11354 7328 11562
rect 7392 11393 7420 11630
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7378 11384 7434 11393
rect 7288 11348 7340 11354
rect 7378 11319 7434 11328
rect 7288 11290 7340 11296
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6840 11014 6868 11086
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 6886 10364 7182 10384
rect 6942 10362 6966 10364
rect 7022 10362 7046 10364
rect 7102 10362 7126 10364
rect 6964 10310 6966 10362
rect 7028 10310 7040 10362
rect 7102 10310 7104 10362
rect 6942 10308 6966 10310
rect 7022 10308 7046 10310
rect 7102 10308 7126 10310
rect 6886 10288 7182 10308
rect 6826 10160 6882 10169
rect 6826 10095 6882 10104
rect 6840 9364 6868 10095
rect 6920 10056 6972 10062
rect 6918 10024 6920 10033
rect 7300 10033 7328 10950
rect 7484 10810 7512 11494
rect 7576 11354 7604 11494
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7564 11144 7616 11150
rect 7564 11086 7616 11092
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7576 10674 7604 11086
rect 7852 11014 7880 12038
rect 7840 11008 7892 11014
rect 7668 10968 7840 10996
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7576 10062 7604 10610
rect 7564 10056 7616 10062
rect 6972 10024 6974 10033
rect 6918 9959 6974 9968
rect 7286 10024 7342 10033
rect 7564 9998 7616 10004
rect 7286 9959 7342 9968
rect 7576 9722 7604 9998
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7470 9616 7526 9625
rect 7470 9551 7472 9560
rect 7524 9551 7526 9560
rect 7472 9522 7524 9528
rect 7288 9444 7340 9450
rect 7288 9386 7340 9392
rect 6840 9336 7256 9364
rect 6886 9276 7182 9296
rect 6942 9274 6966 9276
rect 7022 9274 7046 9276
rect 7102 9274 7126 9276
rect 6964 9222 6966 9274
rect 7028 9222 7040 9274
rect 7102 9222 7104 9274
rect 6942 9220 6966 9222
rect 7022 9220 7046 9222
rect 7102 9220 7126 9222
rect 6886 9200 7182 9220
rect 6736 9172 6788 9178
rect 7228 9160 7256 9336
rect 6736 9114 6788 9120
rect 7208 9132 7256 9160
rect 7208 8276 7236 9132
rect 7300 9042 7328 9386
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7562 8936 7618 8945
rect 7286 8528 7342 8537
rect 7286 8463 7342 8472
rect 7208 8248 7256 8276
rect 6886 8188 7182 8208
rect 6942 8186 6966 8188
rect 7022 8186 7046 8188
rect 7102 8186 7126 8188
rect 6964 8134 6966 8186
rect 7028 8134 7040 8186
rect 7102 8134 7104 8186
rect 6942 8132 6966 8134
rect 7022 8132 7046 8134
rect 7102 8132 7126 8134
rect 6886 8112 7182 8132
rect 7228 8072 7256 8248
rect 7208 8044 7256 8072
rect 6736 7268 6788 7274
rect 6736 7210 6788 7216
rect 6748 6798 6776 7210
rect 7208 7188 7236 8044
rect 7208 7160 7256 7188
rect 6886 7100 7182 7120
rect 6942 7098 6966 7100
rect 7022 7098 7046 7100
rect 7102 7098 7126 7100
rect 6964 7046 6966 7098
rect 7028 7046 7040 7098
rect 7102 7046 7104 7098
rect 6942 7044 6966 7046
rect 7022 7044 7046 7046
rect 7102 7044 7126 7046
rect 6886 7024 7182 7044
rect 7228 6984 7256 7160
rect 7208 6956 7256 6984
rect 7208 6866 7236 6956
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 6644 5772 6696 5778
rect 6644 5714 6696 5720
rect 6748 5574 6776 6734
rect 6886 6012 7182 6032
rect 6942 6010 6966 6012
rect 7022 6010 7046 6012
rect 7102 6010 7126 6012
rect 6964 5958 6966 6010
rect 7028 5958 7040 6010
rect 7102 5958 7104 6010
rect 6942 5956 6966 5958
rect 7022 5956 7046 5958
rect 7102 5956 7126 5958
rect 6886 5936 7182 5956
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 7102 5264 7158 5273
rect 7102 5199 7158 5208
rect 7116 5166 7144 5199
rect 7300 5166 7328 8463
rect 7392 8362 7420 8910
rect 7380 8356 7432 8362
rect 7380 8298 7432 8304
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7392 6934 7420 7278
rect 7380 6928 7432 6934
rect 7380 6870 7432 6876
rect 7484 6730 7512 8910
rect 7562 8871 7618 8880
rect 7576 8090 7604 8871
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7576 7342 7604 7686
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 7472 6724 7524 6730
rect 7472 6666 7524 6672
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7392 5914 7420 6054
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7470 5672 7526 5681
rect 7470 5607 7526 5616
rect 7104 5160 7156 5166
rect 6734 5128 6790 5137
rect 7104 5102 7156 5108
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 6734 5063 6790 5072
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 6656 4826 6684 4966
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6274 4448 6330 4457
rect 6274 4383 6330 4392
rect 6380 4440 6500 4468
rect 6552 4480 6604 4486
rect 6550 4448 6552 4457
rect 6604 4448 6606 4457
rect 6288 4282 6316 4383
rect 6276 4276 6328 4282
rect 6276 4218 6328 4224
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 6288 3942 6316 4218
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 6000 3392 6052 3398
rect 6000 3334 6052 3340
rect 6092 3392 6144 3398
rect 6092 3334 6144 3340
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 6104 2961 6132 3334
rect 6090 2952 6146 2961
rect 6090 2887 6146 2896
rect 5460 2746 5580 2774
rect 5828 2746 5948 2774
rect 5356 2576 5408 2582
rect 5356 2518 5408 2524
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 5552 2310 5580 2746
rect 5816 2372 5868 2378
rect 5816 2314 5868 2320
rect 4896 2304 4948 2310
rect 4896 2246 4948 2252
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 4344 1828 4396 1834
rect 4344 1770 4396 1776
rect 3804 1142 4016 1170
rect 3988 800 4016 1142
rect 4908 800 4936 2246
rect 5828 800 5856 2314
rect 5920 1562 5948 2746
rect 6380 2514 6408 4440
rect 6550 4383 6606 4392
rect 6748 4298 6776 5063
rect 7288 5024 7340 5030
rect 7288 4966 7340 4972
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 6886 4924 7182 4944
rect 6942 4922 6966 4924
rect 7022 4922 7046 4924
rect 7102 4922 7126 4924
rect 6964 4870 6966 4922
rect 7028 4870 7040 4922
rect 7102 4870 7104 4922
rect 6942 4868 6966 4870
rect 7022 4868 7046 4870
rect 7102 4868 7126 4870
rect 6886 4848 7182 4868
rect 7300 4826 7328 4966
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7196 4752 7248 4758
rect 7392 4706 7420 4966
rect 7484 4758 7512 5607
rect 7576 5370 7604 6802
rect 7668 5896 7696 10968
rect 7840 10950 7892 10956
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 7760 10266 7788 10406
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7748 9512 7800 9518
rect 7748 9454 7800 9460
rect 7760 8022 7788 9454
rect 7852 9450 7880 10406
rect 7840 9444 7892 9450
rect 7840 9386 7892 9392
rect 7840 8288 7892 8294
rect 7840 8230 7892 8236
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 7760 7206 7788 7822
rect 7852 7818 7880 8230
rect 7944 7886 7972 12406
rect 8036 12406 8156 12434
rect 8404 12406 8524 12434
rect 8036 12102 8064 12406
rect 8114 12200 8170 12209
rect 8114 12135 8170 12144
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8036 11626 8064 12038
rect 8128 11898 8156 12135
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 8024 11620 8076 11626
rect 8024 11562 8076 11568
rect 8036 11354 8064 11562
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 8206 11520 8262 11529
rect 8024 11348 8076 11354
rect 8024 11290 8076 11296
rect 8022 10160 8078 10169
rect 8022 10095 8078 10104
rect 8036 10062 8064 10095
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 8128 7954 8156 11494
rect 8206 11455 8262 11464
rect 8220 11286 8248 11455
rect 8208 11280 8260 11286
rect 8208 11222 8260 11228
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 8220 10606 8248 11086
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 8206 10024 8262 10033
rect 8206 9959 8262 9968
rect 8220 9625 8248 9959
rect 8312 9926 8340 11630
rect 8404 10606 8432 12406
rect 9048 12238 9076 12582
rect 9784 12442 9812 12854
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 9036 12232 9088 12238
rect 9036 12174 9088 12180
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8496 10810 8524 11086
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8680 10742 8708 11834
rect 8760 11620 8812 11626
rect 8760 11562 8812 11568
rect 8772 11529 8800 11562
rect 8758 11520 8814 11529
rect 8758 11455 8814 11464
rect 8772 11286 8800 11455
rect 8760 11280 8812 11286
rect 8760 11222 8812 11228
rect 8760 11076 8812 11082
rect 8760 11018 8812 11024
rect 8668 10736 8720 10742
rect 8668 10678 8720 10684
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8680 10266 8708 10678
rect 8772 10470 8800 11018
rect 8760 10464 8812 10470
rect 8758 10432 8760 10441
rect 8812 10432 8814 10441
rect 8758 10367 8814 10376
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 9048 10169 9076 12174
rect 9218 11928 9274 11937
rect 9218 11863 9274 11872
rect 9232 11150 9260 11863
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9324 11558 9352 11698
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 9324 11218 9352 11494
rect 9312 11212 9364 11218
rect 9312 11154 9364 11160
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9140 10985 9168 11086
rect 9416 11082 9444 12174
rect 9588 12164 9640 12170
rect 9588 12106 9640 12112
rect 9600 11830 9628 12106
rect 9588 11824 9640 11830
rect 9588 11766 9640 11772
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9508 11626 9536 11698
rect 9496 11620 9548 11626
rect 9496 11562 9548 11568
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9126 10976 9182 10985
rect 9126 10911 9182 10920
rect 9140 10742 9168 10911
rect 9128 10736 9180 10742
rect 9128 10678 9180 10684
rect 9034 10160 9090 10169
rect 8760 10124 8812 10130
rect 9034 10095 9090 10104
rect 8760 10066 8812 10072
rect 8482 10024 8538 10033
rect 8482 9959 8538 9968
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 8312 9722 8340 9862
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8206 9616 8262 9625
rect 8206 9551 8262 9560
rect 8496 9110 8524 9959
rect 8574 9888 8630 9897
rect 8574 9823 8630 9832
rect 8588 9518 8616 9823
rect 8772 9674 8800 10066
rect 8680 9646 8800 9674
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8680 9382 8708 9646
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8852 9376 8904 9382
rect 8852 9318 8904 9324
rect 8392 9104 8444 9110
rect 8392 9046 8444 9052
rect 8484 9104 8536 9110
rect 8484 9046 8536 9052
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8220 8945 8248 8978
rect 8206 8936 8262 8945
rect 8206 8871 8262 8880
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 7840 7812 7892 7818
rect 7840 7754 7892 7760
rect 7852 7410 7880 7754
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7748 6928 7800 6934
rect 7748 6870 7800 6876
rect 7760 6390 7788 6870
rect 7852 6798 7880 7346
rect 8036 7206 8064 7686
rect 8220 7410 8248 8774
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8312 8362 8340 8502
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 8404 8090 8432 9046
rect 8864 8974 8892 9318
rect 8944 9036 8996 9042
rect 8944 8978 8996 8984
rect 8852 8968 8904 8974
rect 8482 8936 8538 8945
rect 8852 8910 8904 8916
rect 8482 8871 8538 8880
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8298 7984 8354 7993
rect 8298 7919 8354 7928
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8024 7200 8076 7206
rect 8024 7142 8076 7148
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7748 6384 7800 6390
rect 7748 6326 7800 6332
rect 7932 6248 7984 6254
rect 7932 6190 7984 6196
rect 7668 5868 7788 5896
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 7576 5012 7604 5306
rect 7668 5234 7696 5714
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7760 5098 7788 5868
rect 7944 5710 7972 6190
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 8036 5273 8064 7142
rect 8208 6928 8260 6934
rect 8208 6870 8260 6876
rect 8220 6458 8248 6870
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8220 5914 8248 6394
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8312 5778 8340 7919
rect 8404 6866 8432 8026
rect 8496 7546 8524 8871
rect 8864 8430 8892 8910
rect 8956 8838 8984 8978
rect 8944 8832 8996 8838
rect 8944 8774 8996 8780
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8680 7206 8708 7346
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8772 6866 8800 8366
rect 8956 8090 8984 8774
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8852 8016 8904 8022
rect 8850 7984 8852 7993
rect 8904 7984 8906 7993
rect 8850 7919 8906 7928
rect 8956 6934 8984 8026
rect 9048 7313 9076 10095
rect 9140 10033 9168 10678
rect 9220 10668 9272 10674
rect 9220 10610 9272 10616
rect 9126 10024 9182 10033
rect 9126 9959 9182 9968
rect 9232 9926 9260 10610
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9324 10062 9352 10406
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9312 10056 9364 10062
rect 9508 10033 9536 10066
rect 9312 9998 9364 10004
rect 9494 10024 9550 10033
rect 9494 9959 9550 9968
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 9220 9920 9272 9926
rect 9220 9862 9272 9868
rect 9140 9586 9168 9862
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 9140 9042 9168 9522
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 9128 9036 9180 9042
rect 9128 8978 9180 8984
rect 9128 8900 9180 8906
rect 9128 8842 9180 8848
rect 9140 7342 9168 8842
rect 9128 7336 9180 7342
rect 9034 7304 9090 7313
rect 9128 7278 9180 7284
rect 9034 7239 9090 7248
rect 8944 6928 8996 6934
rect 8944 6870 8996 6876
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 8772 6662 8800 6802
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8666 6352 8722 6361
rect 8864 6322 8892 6598
rect 8666 6287 8722 6296
rect 8852 6316 8904 6322
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8022 5264 8078 5273
rect 8220 5250 8248 5646
rect 8300 5636 8352 5642
rect 8300 5578 8352 5584
rect 8128 5234 8248 5250
rect 8022 5199 8078 5208
rect 8116 5228 8248 5234
rect 8168 5222 8248 5228
rect 8116 5170 8168 5176
rect 8024 5160 8076 5166
rect 8022 5128 8024 5137
rect 8076 5128 8078 5137
rect 7748 5092 7800 5098
rect 8022 5063 8078 5072
rect 8116 5092 8168 5098
rect 7748 5034 7800 5040
rect 8116 5034 8168 5040
rect 7656 5024 7708 5030
rect 7576 4984 7656 5012
rect 7656 4966 7708 4972
rect 7248 4700 7420 4706
rect 7196 4694 7420 4700
rect 7472 4752 7524 4758
rect 7472 4694 7524 4700
rect 7208 4678 7420 4694
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 7564 4616 7616 4622
rect 7564 4558 7616 4564
rect 6564 4270 6776 4298
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6472 2689 6500 3878
rect 6564 3058 6592 4270
rect 6736 4208 6788 4214
rect 6734 4176 6736 4185
rect 6840 4196 6868 4558
rect 6788 4176 6868 4196
rect 6790 4168 6868 4176
rect 6734 4111 6790 4120
rect 7576 4078 7604 4558
rect 7656 4276 7708 4282
rect 7760 4264 7788 5034
rect 8128 4826 8156 5034
rect 8116 4820 8168 4826
rect 8116 4762 8168 4768
rect 8220 4282 8248 5222
rect 7840 4276 7892 4282
rect 7760 4236 7840 4264
rect 7656 4218 7708 4224
rect 7840 4218 7892 4224
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 7668 4185 7696 4218
rect 7654 4176 7710 4185
rect 7654 4111 7710 4120
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6458 2680 6514 2689
rect 6564 2650 6592 2994
rect 6458 2615 6514 2624
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 6368 2508 6420 2514
rect 6368 2450 6420 2456
rect 6012 2106 6040 2450
rect 6000 2100 6052 2106
rect 6000 2042 6052 2048
rect 6656 1902 6684 4014
rect 6886 3836 7182 3856
rect 6942 3834 6966 3836
rect 7022 3834 7046 3836
rect 7102 3834 7126 3836
rect 6964 3782 6966 3834
rect 7028 3782 7040 3834
rect 7102 3782 7104 3834
rect 6942 3780 6966 3782
rect 7022 3780 7046 3782
rect 7102 3780 7126 3782
rect 6886 3760 7182 3780
rect 7576 3738 7604 4014
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 6748 3602 6776 3674
rect 8128 3641 8156 3878
rect 8114 3632 8170 3641
rect 6736 3596 6788 3602
rect 8114 3567 8170 3576
rect 6736 3538 6788 3544
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 6736 2984 6788 2990
rect 6734 2952 6736 2961
rect 6788 2952 6790 2961
rect 6734 2887 6790 2896
rect 7760 2854 7788 3402
rect 7840 3392 7892 3398
rect 7840 3334 7892 3340
rect 7852 3194 7880 3334
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7656 2848 7708 2854
rect 7656 2790 7708 2796
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 6886 2748 7182 2768
rect 6942 2746 6966 2748
rect 7022 2746 7046 2748
rect 7102 2746 7126 2748
rect 6964 2694 6966 2746
rect 7028 2694 7040 2746
rect 7102 2694 7104 2746
rect 6942 2692 6966 2694
rect 7022 2692 7046 2694
rect 7102 2692 7126 2694
rect 6886 2672 7182 2692
rect 6736 2372 6788 2378
rect 6736 2314 6788 2320
rect 6644 1896 6696 1902
rect 6644 1838 6696 1844
rect 5908 1556 5960 1562
rect 5908 1498 5960 1504
rect 6748 800 6776 2314
rect 6828 2304 6880 2310
rect 6828 2246 6880 2252
rect 6840 1630 6868 2246
rect 6828 1624 6880 1630
rect 6828 1566 6880 1572
rect 7484 1426 7512 2790
rect 7668 2650 7696 2790
rect 7656 2644 7708 2650
rect 7656 2586 7708 2592
rect 8128 2446 8156 3567
rect 8312 3058 8340 5578
rect 8404 5370 8432 6054
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 8392 5364 8444 5370
rect 8392 5306 8444 5312
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 8404 4690 8432 4966
rect 8392 4684 8444 4690
rect 8392 4626 8444 4632
rect 8392 4548 8444 4554
rect 8392 4490 8444 4496
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 8298 2544 8354 2553
rect 8208 2508 8260 2514
rect 8298 2479 8300 2488
rect 8208 2450 8260 2456
rect 8352 2479 8354 2488
rect 8300 2450 8352 2456
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 7564 2372 7616 2378
rect 7564 2314 7616 2320
rect 7472 1420 7524 1426
rect 7472 1362 7524 1368
rect 7576 800 7604 2314
rect 8220 2038 8248 2450
rect 8208 2032 8260 2038
rect 8208 1974 8260 1980
rect 8404 1698 8432 4490
rect 8496 4026 8524 5714
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8588 5234 8616 5646
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 8574 4720 8630 4729
rect 8680 4690 8708 6287
rect 8852 6258 8904 6264
rect 8852 6180 8904 6186
rect 8852 6122 8904 6128
rect 8760 5772 8812 5778
rect 8760 5714 8812 5720
rect 8772 5574 8800 5714
rect 8760 5568 8812 5574
rect 8760 5510 8812 5516
rect 8760 5296 8812 5302
rect 8760 5238 8812 5244
rect 8574 4655 8576 4664
rect 8628 4655 8630 4664
rect 8668 4684 8720 4690
rect 8576 4626 8628 4632
rect 8668 4626 8720 4632
rect 8496 3998 8616 4026
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8496 3670 8524 3878
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 8588 3602 8616 3998
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 8484 3392 8536 3398
rect 8484 3334 8536 3340
rect 8496 3058 8524 3334
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 8484 2916 8536 2922
rect 8484 2858 8536 2864
rect 8392 1692 8444 1698
rect 8392 1634 8444 1640
rect 8496 800 8524 2858
rect 8668 2848 8720 2854
rect 8668 2790 8720 2796
rect 8680 2650 8708 2790
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 8576 2576 8628 2582
rect 8772 2530 8800 5238
rect 8864 3534 8892 6122
rect 8956 5914 8984 6734
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 8956 3738 8984 4422
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 9048 3602 9076 7239
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 9232 6202 9260 9454
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9312 9036 9364 9042
rect 9312 8978 9364 8984
rect 9324 8430 9352 8978
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9312 8288 9364 8294
rect 9312 8230 9364 8236
rect 9324 7410 9352 8230
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9324 6322 9352 6598
rect 9416 6322 9444 9114
rect 9508 8566 9536 9959
rect 9600 9110 9628 11766
rect 9692 11132 9720 12174
rect 10244 12102 10272 12854
rect 10324 12708 10376 12714
rect 10324 12650 10376 12656
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 9784 11880 9812 12038
rect 9852 11996 10148 12016
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 9930 11942 9932 11994
rect 9994 11942 10006 11994
rect 10068 11942 10070 11994
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 9852 11920 10148 11940
rect 10336 11898 10364 12650
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 10692 12436 10744 12442
rect 10796 12434 10824 12582
rect 10796 12406 11192 12434
rect 10692 12378 10744 12384
rect 10598 12336 10654 12345
rect 10598 12271 10654 12280
rect 10612 12238 10640 12271
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10324 11892 10376 11898
rect 9784 11852 9904 11880
rect 9876 11558 9904 11852
rect 10324 11834 10376 11840
rect 9956 11824 10008 11830
rect 9956 11766 10008 11772
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9864 11552 9916 11558
rect 9968 11529 9996 11766
rect 10140 11552 10192 11558
rect 9864 11494 9916 11500
rect 9954 11520 10010 11529
rect 9784 11354 9812 11494
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9876 11257 9904 11494
rect 10140 11494 10192 11500
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 9954 11455 10010 11464
rect 10152 11354 10180 11494
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 9862 11248 9918 11257
rect 9862 11183 9918 11192
rect 9772 11144 9824 11150
rect 9692 11104 9772 11132
rect 9772 11086 9824 11092
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9692 10538 9720 10746
rect 9680 10532 9732 10538
rect 9680 10474 9732 10480
rect 9692 9602 9720 10474
rect 9784 10266 9812 11086
rect 9852 10908 10148 10928
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 9930 10854 9932 10906
rect 9994 10854 10006 10906
rect 10068 10854 10070 10906
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 9852 10832 10148 10852
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 9862 10568 9918 10577
rect 9862 10503 9864 10512
rect 9916 10503 9918 10512
rect 9864 10474 9916 10480
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 10060 10305 10088 10406
rect 10046 10296 10102 10305
rect 9772 10260 9824 10266
rect 10046 10231 10102 10240
rect 9772 10202 9824 10208
rect 10152 9994 10180 10610
rect 10244 10266 10272 11494
rect 10336 10810 10364 11834
rect 10428 11778 10456 12174
rect 10506 11792 10562 11801
rect 10428 11750 10506 11778
rect 10506 11727 10562 11736
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 10612 11218 10640 11698
rect 10600 11212 10652 11218
rect 10600 11154 10652 11160
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10612 10674 10640 11154
rect 10704 10792 10732 12378
rect 11164 12238 11192 12406
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 11164 12102 11192 12174
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 10796 11898 10824 12038
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 10704 10764 10916 10792
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10414 10568 10470 10577
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 10140 9988 10192 9994
rect 10140 9930 10192 9936
rect 9784 9722 9812 9930
rect 9852 9820 10148 9840
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 9930 9766 9932 9818
rect 9994 9766 10006 9818
rect 10068 9766 10070 9818
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 9852 9744 10148 9764
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9692 9574 9812 9602
rect 9588 9104 9640 9110
rect 9588 9046 9640 9052
rect 9496 8560 9548 8566
rect 9496 8502 9548 8508
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 9404 6316 9456 6322
rect 9404 6258 9456 6264
rect 9140 5710 9168 6190
rect 9232 6174 9444 6202
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 9232 5778 9260 6054
rect 9220 5772 9272 5778
rect 9220 5714 9272 5720
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9140 5030 9168 5170
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9220 4480 9272 4486
rect 9218 4448 9220 4457
rect 9272 4448 9274 4457
rect 9218 4383 9274 4392
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9036 3596 9088 3602
rect 9036 3538 9088 3544
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 8864 3058 8892 3470
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 8852 2848 8904 2854
rect 8850 2816 8852 2825
rect 8904 2816 8906 2825
rect 8850 2751 8906 2760
rect 9048 2650 9076 3538
rect 9140 3194 9168 3674
rect 9218 3632 9274 3641
rect 9218 3567 9220 3576
rect 9272 3567 9274 3576
rect 9220 3538 9272 3544
rect 9220 3460 9272 3466
rect 9220 3402 9272 3408
rect 9232 3194 9260 3402
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 8628 2524 8800 2530
rect 8576 2518 8800 2524
rect 8588 2502 8800 2518
rect 9324 2310 9352 6054
rect 9416 4729 9444 6174
rect 9508 5166 9536 8366
rect 9680 8288 9732 8294
rect 9680 8230 9732 8236
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9600 5166 9628 7754
rect 9692 7750 9720 8230
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9680 7472 9732 7478
rect 9680 7414 9732 7420
rect 9692 7206 9720 7414
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9680 6928 9732 6934
rect 9680 6870 9732 6876
rect 9692 6118 9720 6870
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9692 5302 9720 6054
rect 9680 5296 9732 5302
rect 9680 5238 9732 5244
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9402 4720 9458 4729
rect 9402 4655 9404 4664
rect 9456 4655 9458 4664
rect 9404 4626 9456 4632
rect 9416 4595 9444 4626
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 9508 2106 9536 4966
rect 9692 4078 9720 4966
rect 9784 4264 9812 9574
rect 10336 9178 10364 10542
rect 10414 10503 10470 10512
rect 10428 10470 10456 10503
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10520 10305 10548 10406
rect 10506 10296 10562 10305
rect 10416 10260 10468 10266
rect 10562 10254 10640 10282
rect 10506 10231 10562 10240
rect 10416 10202 10468 10208
rect 10428 10130 10456 10202
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10416 9444 10468 9450
rect 10416 9386 10468 9392
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 9852 8732 10148 8752
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 9930 8678 9932 8730
rect 9994 8678 10006 8730
rect 10068 8678 10070 8730
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 9852 8656 10148 8676
rect 10244 8362 10272 8774
rect 10428 8634 10456 9386
rect 10520 9081 10548 9998
rect 10506 9072 10562 9081
rect 10506 9007 10562 9016
rect 10520 8634 10548 9007
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10324 8560 10376 8566
rect 10324 8502 10376 8508
rect 10232 8356 10284 8362
rect 10232 8298 10284 8304
rect 9864 7880 9916 7886
rect 9862 7848 9864 7857
rect 9916 7848 9918 7857
rect 9862 7783 9918 7792
rect 9852 7644 10148 7664
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 9930 7590 9932 7642
rect 9994 7590 10006 7642
rect 10068 7590 10070 7642
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 9852 7568 10148 7588
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9876 6866 9904 7142
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9852 6556 10148 6576
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 9930 6502 9932 6554
rect 9994 6502 10006 6554
rect 10068 6502 10070 6554
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 9852 6480 10148 6500
rect 10244 6322 10272 8298
rect 10336 6848 10364 8502
rect 10428 7410 10456 8570
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10416 6860 10468 6866
rect 10336 6820 10416 6848
rect 10416 6802 10468 6808
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 10244 5710 10272 6258
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 9852 5468 10148 5488
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 9930 5414 9932 5466
rect 9994 5414 10006 5466
rect 10068 5414 10070 5466
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 9852 5392 10148 5412
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 9968 4554 9996 4762
rect 9956 4548 10008 4554
rect 9956 4490 10008 4496
rect 10152 4468 10180 5170
rect 10244 4622 10272 5646
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 10152 4440 10272 4468
rect 10336 4457 10364 5510
rect 10428 4690 10456 6802
rect 10520 6390 10548 8434
rect 10612 8412 10640 10254
rect 10796 10130 10824 10610
rect 10784 10124 10836 10130
rect 10784 10066 10836 10072
rect 10796 9722 10824 10066
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10690 9616 10746 9625
rect 10690 9551 10692 9560
rect 10744 9551 10746 9560
rect 10692 9522 10744 9528
rect 10704 9042 10732 9522
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10796 8906 10824 9658
rect 10784 8900 10836 8906
rect 10784 8842 10836 8848
rect 10692 8424 10744 8430
rect 10612 8384 10692 8412
rect 10692 8366 10744 8372
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10600 7812 10652 7818
rect 10600 7754 10652 7760
rect 10508 6384 10560 6390
rect 10508 6326 10560 6332
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 9852 4380 10148 4400
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 9930 4326 9932 4378
rect 9994 4326 10006 4378
rect 10068 4326 10070 4378
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 9852 4304 10148 4324
rect 9784 4236 9996 4264
rect 9968 4078 9996 4236
rect 10048 4208 10100 4214
rect 10100 4168 10180 4196
rect 10048 4150 10100 4156
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 10152 4026 10180 4168
rect 10244 4146 10272 4440
rect 10322 4448 10378 4457
rect 10322 4383 10378 4392
rect 10428 4214 10456 4626
rect 10416 4208 10468 4214
rect 10416 4150 10468 4156
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 9692 3058 9720 4014
rect 10152 3998 10456 4026
rect 9772 3936 9824 3942
rect 9956 3936 10008 3942
rect 9824 3896 9956 3924
rect 9772 3878 9824 3884
rect 9956 3878 10008 3884
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 9772 3392 9824 3398
rect 9772 3334 9824 3340
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9600 2446 9628 2586
rect 9692 2514 9720 2994
rect 9784 2990 9812 3334
rect 9852 3292 10148 3312
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 9930 3238 9932 3290
rect 9994 3238 10006 3290
rect 10068 3238 10070 3290
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 9852 3216 10148 3236
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 9968 2689 9996 2790
rect 9954 2680 10010 2689
rect 9954 2615 10010 2624
rect 9772 2576 9824 2582
rect 9772 2518 9824 2524
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 9692 2378 9720 2450
rect 9680 2372 9732 2378
rect 9680 2314 9732 2320
rect 9496 2100 9548 2106
rect 9496 2042 9548 2048
rect 9784 1630 9812 2518
rect 9968 2446 9996 2615
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 9852 2204 10148 2224
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 9930 2150 9932 2202
rect 9994 2150 10006 2202
rect 10068 2150 10070 2202
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 9852 2128 10148 2148
rect 10244 1766 10272 3878
rect 10324 3120 10376 3126
rect 10324 3062 10376 3068
rect 10232 1760 10284 1766
rect 10232 1702 10284 1708
rect 9772 1624 9824 1630
rect 9772 1566 9824 1572
rect 9404 1420 9456 1426
rect 9404 1362 9456 1368
rect 9416 800 9444 1362
rect 10336 800 10364 3062
rect 10428 2854 10456 3998
rect 10416 2848 10468 2854
rect 10416 2790 10468 2796
rect 10520 2582 10548 6190
rect 10612 4826 10640 7754
rect 10690 6624 10746 6633
rect 10690 6559 10746 6568
rect 10704 6458 10732 6559
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10690 6352 10746 6361
rect 10690 6287 10692 6296
rect 10744 6287 10746 6296
rect 10692 6258 10744 6264
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10600 4208 10652 4214
rect 10600 4150 10652 4156
rect 10612 4026 10640 4150
rect 10704 4146 10732 6054
rect 10796 5778 10824 8230
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10796 5098 10824 5510
rect 10784 5092 10836 5098
rect 10784 5034 10836 5040
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 10612 3998 10732 4026
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10612 3670 10640 3878
rect 10600 3664 10652 3670
rect 10600 3606 10652 3612
rect 10704 3058 10732 3998
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10508 2576 10560 2582
rect 10508 2518 10560 2524
rect 10598 2544 10654 2553
rect 10598 2479 10600 2488
rect 10652 2479 10654 2488
rect 10600 2450 10652 2456
rect 10612 1902 10640 2450
rect 10796 2446 10824 5034
rect 10888 4049 10916 10764
rect 10980 7993 11008 11290
rect 11072 11121 11100 11290
rect 11058 11112 11114 11121
rect 11058 11047 11114 11056
rect 11072 10674 11100 11047
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 10966 7984 11022 7993
rect 10966 7919 11022 7928
rect 11072 6474 11100 10610
rect 11164 10606 11192 12038
rect 11244 11552 11296 11558
rect 11348 11540 11376 12038
rect 11296 11512 11376 11540
rect 11428 11552 11480 11558
rect 11244 11494 11296 11500
rect 11428 11494 11480 11500
rect 11440 11286 11468 11494
rect 11428 11280 11480 11286
rect 11428 11222 11480 11228
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11348 10742 11376 11154
rect 11428 11008 11480 11014
rect 11428 10950 11480 10956
rect 11440 10742 11468 10950
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 11428 10736 11480 10742
rect 11428 10678 11480 10684
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11348 10470 11376 10678
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11532 9674 11560 12854
rect 11900 12434 11928 14758
rect 12817 14716 13113 14736
rect 12873 14714 12897 14716
rect 12953 14714 12977 14716
rect 13033 14714 13057 14716
rect 12895 14662 12897 14714
rect 12959 14662 12971 14714
rect 13033 14662 13035 14714
rect 12873 14660 12897 14662
rect 12953 14660 12977 14662
rect 13033 14660 13057 14662
rect 12817 14640 13113 14660
rect 13924 14074 13952 16400
rect 14464 14612 14516 14618
rect 14464 14554 14516 14560
rect 13912 14068 13964 14074
rect 13912 14010 13964 14016
rect 12817 13628 13113 13648
rect 12873 13626 12897 13628
rect 12953 13626 12977 13628
rect 13033 13626 13057 13628
rect 12895 13574 12897 13626
rect 12959 13574 12971 13626
rect 13033 13574 13035 13626
rect 12873 13572 12897 13574
rect 12953 13572 12977 13574
rect 13033 13572 13057 13574
rect 12817 13552 13113 13572
rect 14280 13524 14332 13530
rect 14280 13466 14332 13472
rect 12440 12912 12492 12918
rect 12440 12854 12492 12860
rect 12164 12436 12216 12442
rect 11900 12406 12020 12434
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 11808 11082 11836 12242
rect 11900 12209 11928 12242
rect 11886 12200 11942 12209
rect 11886 12135 11942 12144
rect 11992 12102 12020 12406
rect 12164 12378 12216 12384
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 11612 11076 11664 11082
rect 11612 11018 11664 11024
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 11624 10606 11652 11018
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 11716 10674 11744 10950
rect 11992 10810 12020 12038
rect 12072 11824 12124 11830
rect 12072 11766 12124 11772
rect 12084 11558 12112 11766
rect 12176 11626 12204 12378
rect 12256 12368 12308 12374
rect 12308 12328 12388 12356
rect 12256 12310 12308 12316
rect 12164 11620 12216 11626
rect 12164 11562 12216 11568
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11612 10600 11664 10606
rect 11612 10542 11664 10548
rect 11624 10130 11652 10542
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 11624 9722 11652 10066
rect 11440 9646 11560 9674
rect 11612 9716 11664 9722
rect 11612 9658 11664 9664
rect 11150 9480 11206 9489
rect 11150 9415 11206 9424
rect 11164 9382 11192 9415
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 11164 8945 11192 9318
rect 11244 9104 11296 9110
rect 11244 9046 11296 9052
rect 11150 8936 11206 8945
rect 11150 8871 11206 8880
rect 11164 7818 11192 8871
rect 11152 7812 11204 7818
rect 11152 7754 11204 7760
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 10980 6446 11100 6474
rect 10980 6118 11008 6446
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10980 4554 11008 6054
rect 11072 4826 11100 6326
rect 11164 5914 11192 6802
rect 11256 6225 11284 9046
rect 11336 7744 11388 7750
rect 11336 7686 11388 7692
rect 11348 7342 11376 7686
rect 11440 7478 11468 9646
rect 11624 8498 11652 9658
rect 11716 9602 11744 10202
rect 11808 9722 11836 10406
rect 11796 9716 11848 9722
rect 11796 9658 11848 9664
rect 11794 9616 11850 9625
rect 11716 9574 11794 9602
rect 11794 9551 11796 9560
rect 11848 9551 11850 9560
rect 11888 9580 11940 9586
rect 11796 9522 11848 9528
rect 11888 9522 11940 9528
rect 11794 9480 11850 9489
rect 11900 9466 11928 9522
rect 11850 9438 11928 9466
rect 11794 9415 11850 9424
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11716 8498 11744 8910
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11428 7472 11480 7478
rect 11428 7414 11480 7420
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11348 7002 11376 7142
rect 11336 6996 11388 7002
rect 11336 6938 11388 6944
rect 11348 6361 11376 6938
rect 11440 6882 11468 7414
rect 11532 7002 11560 7890
rect 11624 7426 11652 8434
rect 11808 8430 11836 8774
rect 11992 8480 12020 10406
rect 12084 9518 12112 11154
rect 12072 9512 12124 9518
rect 12072 9454 12124 9460
rect 12084 9178 12112 9454
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 12176 9110 12204 11562
rect 12360 11370 12388 12328
rect 12452 11762 12480 12854
rect 12817 12540 13113 12560
rect 12873 12538 12897 12540
rect 12953 12538 12977 12540
rect 13033 12538 13057 12540
rect 12895 12486 12897 12538
rect 12959 12486 12971 12538
rect 13033 12486 13035 12538
rect 12873 12484 12897 12486
rect 12953 12484 12977 12486
rect 13033 12484 13057 12486
rect 12817 12464 13113 12484
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13176 12164 13228 12170
rect 13176 12106 13228 12112
rect 12440 11756 12492 11762
rect 12440 11698 12492 11704
rect 12622 11520 12678 11529
rect 12622 11455 12678 11464
rect 12360 11342 12572 11370
rect 12346 11248 12402 11257
rect 12346 11183 12402 11192
rect 12254 11112 12310 11121
rect 12254 11047 12310 11056
rect 12268 10470 12296 11047
rect 12360 11014 12388 11183
rect 12544 11150 12572 11342
rect 12636 11286 12664 11455
rect 12817 11452 13113 11472
rect 12873 11450 12897 11452
rect 12953 11450 12977 11452
rect 13033 11450 13057 11452
rect 12895 11398 12897 11450
rect 12959 11398 12971 11450
rect 13033 11398 13035 11450
rect 12873 11396 12897 11398
rect 12953 11396 12977 11398
rect 13033 11396 13057 11398
rect 12817 11376 13113 11396
rect 13188 11354 13216 12106
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 13280 11558 13308 12038
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12532 11144 12584 11150
rect 12532 11086 12584 11092
rect 13280 11082 13308 11494
rect 13726 11384 13782 11393
rect 13360 11348 13412 11354
rect 13412 11308 13584 11336
rect 13832 11354 13860 12174
rect 13726 11319 13782 11328
rect 13820 11348 13872 11354
rect 13360 11290 13412 11296
rect 13268 11076 13320 11082
rect 13268 11018 13320 11024
rect 13452 11076 13504 11082
rect 13452 11018 13504 11024
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 13174 10840 13230 10849
rect 13174 10775 13230 10784
rect 13188 10577 13216 10775
rect 13280 10713 13308 11018
rect 13266 10704 13322 10713
rect 13266 10639 13322 10648
rect 13174 10568 13230 10577
rect 12532 10532 12584 10538
rect 13174 10503 13230 10512
rect 12532 10474 12584 10480
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 12544 9926 12572 10474
rect 12817 10364 13113 10384
rect 12873 10362 12897 10364
rect 12953 10362 12977 10364
rect 13033 10362 13057 10364
rect 12895 10310 12897 10362
rect 12959 10310 12971 10362
rect 13033 10310 13035 10362
rect 12873 10308 12897 10310
rect 12953 10308 12977 10310
rect 13033 10308 13057 10310
rect 12817 10288 13113 10308
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 12256 9920 12308 9926
rect 12532 9920 12584 9926
rect 12308 9880 12388 9908
rect 12256 9862 12308 9868
rect 12254 9752 12310 9761
rect 12360 9722 12388 9880
rect 12532 9862 12584 9868
rect 12254 9687 12310 9696
rect 12348 9716 12400 9722
rect 12268 9654 12296 9687
rect 12348 9658 12400 9664
rect 12256 9648 12308 9654
rect 12256 9590 12308 9596
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 12360 9382 12388 9522
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12164 9104 12216 9110
rect 12164 9046 12216 9052
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 12164 8900 12216 8906
rect 12164 8842 12216 8848
rect 12176 8566 12204 8842
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 11992 8452 12112 8480
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11886 8392 11942 8401
rect 11886 8327 11888 8336
rect 11940 8327 11942 8336
rect 11888 8298 11940 8304
rect 12084 7970 12112 8452
rect 12176 8362 12204 8502
rect 12164 8356 12216 8362
rect 12164 8298 12216 8304
rect 12084 7942 12204 7970
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 12072 7880 12124 7886
rect 12072 7822 12124 7828
rect 11808 7528 11836 7822
rect 11888 7540 11940 7546
rect 11808 7500 11888 7528
rect 11888 7482 11940 7488
rect 12084 7426 12112 7822
rect 11624 7410 12112 7426
rect 11612 7404 12112 7410
rect 11664 7398 12112 7404
rect 11612 7346 11664 7352
rect 11888 7268 11940 7274
rect 11808 7228 11888 7256
rect 11520 6996 11572 7002
rect 11520 6938 11572 6944
rect 11808 6934 11836 7228
rect 11888 7210 11940 7216
rect 12176 7154 12204 7942
rect 12268 7206 12296 8978
rect 12360 8430 12388 9114
rect 12544 8566 12572 9862
rect 12636 9586 12664 10066
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12636 9110 12664 9522
rect 13188 9489 13216 10503
rect 13174 9480 13230 9489
rect 13174 9415 13230 9424
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 13176 9376 13228 9382
rect 13176 9318 13228 9324
rect 12624 9104 12676 9110
rect 12624 9046 12676 9052
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12532 8560 12584 8566
rect 12532 8502 12584 8508
rect 12636 8498 12664 8774
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 12728 8430 12756 9318
rect 12817 9276 13113 9296
rect 12873 9274 12897 9276
rect 12953 9274 12977 9276
rect 13033 9274 13057 9276
rect 12895 9222 12897 9274
rect 12959 9222 12971 9274
rect 13033 9222 13035 9274
rect 12873 9220 12897 9222
rect 12953 9220 12977 9222
rect 13033 9220 13057 9222
rect 12817 9200 13113 9220
rect 13188 9178 13216 9318
rect 13280 9217 13308 10639
rect 13360 9648 13412 9654
rect 13464 9625 13492 11018
rect 13556 10266 13584 11308
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13360 9590 13412 9596
rect 13450 9616 13506 9625
rect 13372 9382 13400 9590
rect 13450 9551 13506 9560
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 13266 9208 13322 9217
rect 13176 9172 13228 9178
rect 13266 9143 13322 9152
rect 13176 9114 13228 9120
rect 13358 9072 13414 9081
rect 13358 9007 13360 9016
rect 13412 9007 13414 9016
rect 13360 8978 13412 8984
rect 13176 8968 13228 8974
rect 13176 8910 13228 8916
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13188 8566 13216 8910
rect 13280 8566 13308 8910
rect 13360 8900 13412 8906
rect 13360 8842 13412 8848
rect 13176 8560 13228 8566
rect 13176 8502 13228 8508
rect 13268 8560 13320 8566
rect 13268 8502 13320 8508
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 12716 8424 12768 8430
rect 12716 8366 12768 8372
rect 11900 7126 12204 7154
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 11796 6928 11848 6934
rect 11440 6854 11652 6882
rect 11796 6870 11848 6876
rect 11624 6798 11652 6854
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11428 6724 11480 6730
rect 11428 6666 11480 6672
rect 11334 6352 11390 6361
rect 11334 6287 11390 6296
rect 11242 6216 11298 6225
rect 11242 6151 11298 6160
rect 11348 6118 11376 6287
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 10968 4548 11020 4554
rect 10968 4490 11020 4496
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11072 4282 11100 4422
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 11060 4276 11112 4282
rect 11060 4218 11112 4224
rect 10874 4040 10930 4049
rect 10874 3975 10930 3984
rect 10980 3992 11008 4218
rect 11164 3992 11192 5170
rect 11256 5166 11284 5646
rect 11440 5574 11468 6666
rect 11532 6458 11560 6734
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11520 6180 11572 6186
rect 11520 6122 11572 6128
rect 11336 5568 11388 5574
rect 11336 5510 11388 5516
rect 11428 5568 11480 5574
rect 11428 5510 11480 5516
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 10980 3964 11192 3992
rect 10980 3534 11008 3964
rect 11256 3890 11284 4966
rect 11348 4078 11376 5510
rect 11428 4752 11480 4758
rect 11428 4694 11480 4700
rect 11440 4214 11468 4694
rect 11428 4208 11480 4214
rect 11428 4150 11480 4156
rect 11336 4072 11388 4078
rect 11336 4014 11388 4020
rect 11164 3862 11284 3890
rect 10968 3528 11020 3534
rect 10966 3496 10968 3505
rect 11020 3496 11022 3505
rect 10966 3431 11022 3440
rect 10784 2440 10836 2446
rect 11164 2428 11192 3862
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 11440 2990 11468 3674
rect 11428 2984 11480 2990
rect 11428 2926 11480 2932
rect 11532 2922 11560 6122
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11624 4010 11652 6054
rect 11808 5914 11836 6054
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 11716 5370 11744 5714
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 11716 4690 11744 5306
rect 11808 5234 11836 5510
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11796 5092 11848 5098
rect 11796 5034 11848 5040
rect 11808 4826 11836 5034
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 11704 4684 11756 4690
rect 11704 4626 11756 4632
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 11716 4185 11744 4422
rect 11702 4176 11758 4185
rect 11702 4111 11758 4120
rect 11612 4004 11664 4010
rect 11612 3946 11664 3952
rect 11520 2916 11572 2922
rect 11520 2858 11572 2864
rect 11716 2774 11744 4111
rect 11900 3097 11928 7126
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 11980 6792 12032 6798
rect 12084 6746 12112 6938
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 12032 6740 12112 6746
rect 11980 6734 12112 6740
rect 11992 6718 12112 6734
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11992 5710 12020 6394
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11992 5273 12020 5646
rect 11978 5264 12034 5273
rect 11978 5199 12034 5208
rect 11980 5160 12032 5166
rect 11980 5102 12032 5108
rect 11992 4486 12020 5102
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 11980 3596 12032 3602
rect 11980 3538 12032 3544
rect 11886 3088 11942 3097
rect 11796 3052 11848 3058
rect 11992 3058 12020 3538
rect 11886 3023 11942 3032
rect 11980 3052 12032 3058
rect 11796 2994 11848 3000
rect 11256 2746 11744 2774
rect 11256 2650 11284 2746
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11808 2446 11836 2994
rect 11900 2922 11928 3023
rect 11980 2994 12032 3000
rect 11888 2916 11940 2922
rect 11888 2858 11940 2864
rect 12084 2854 12112 6718
rect 12176 6322 12204 6802
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 12176 5710 12204 6258
rect 12360 5914 12388 8366
rect 12817 8188 13113 8208
rect 12873 8186 12897 8188
rect 12953 8186 12977 8188
rect 13033 8186 13057 8188
rect 12895 8134 12897 8186
rect 12959 8134 12971 8186
rect 13033 8134 13035 8186
rect 12873 8132 12897 8134
rect 12953 8132 12977 8134
rect 13033 8132 13057 8134
rect 12817 8112 13113 8132
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12544 6236 12572 8026
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 12912 7478 12940 7890
rect 12900 7472 12952 7478
rect 12900 7414 12952 7420
rect 13268 7200 13320 7206
rect 13268 7142 13320 7148
rect 12817 7100 13113 7120
rect 12873 7098 12897 7100
rect 12953 7098 12977 7100
rect 13033 7098 13057 7100
rect 12895 7046 12897 7098
rect 12959 7046 12971 7098
rect 13033 7046 13035 7098
rect 12873 7044 12897 7046
rect 12953 7044 12977 7046
rect 13033 7044 13057 7046
rect 12817 7024 13113 7044
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 12728 6390 12756 6802
rect 13084 6792 13136 6798
rect 13136 6752 13216 6780
rect 13084 6734 13136 6740
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12716 6384 12768 6390
rect 12820 6361 12848 6598
rect 12716 6326 12768 6332
rect 12806 6352 12862 6361
rect 12624 6316 12676 6322
rect 12806 6287 12862 6296
rect 12624 6258 12676 6264
rect 12452 6208 12572 6236
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 12452 4690 12480 6208
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12544 4826 12572 6054
rect 12636 5098 12664 6258
rect 12716 6248 12768 6254
rect 12716 6190 12768 6196
rect 12624 5092 12676 5098
rect 12624 5034 12676 5040
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12256 4684 12308 4690
rect 12176 4644 12256 4672
rect 12176 4146 12204 4644
rect 12256 4626 12308 4632
rect 12440 4684 12492 4690
rect 12440 4626 12492 4632
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12256 4480 12308 4486
rect 12544 4457 12572 4558
rect 12256 4422 12308 4428
rect 12530 4448 12586 4457
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 12268 4078 12296 4422
rect 12530 4383 12586 4392
rect 12346 4176 12402 4185
rect 12636 4146 12664 5034
rect 12728 4826 12756 6190
rect 12817 6012 13113 6032
rect 12873 6010 12897 6012
rect 12953 6010 12977 6012
rect 13033 6010 13057 6012
rect 12895 5958 12897 6010
rect 12959 5958 12971 6010
rect 13033 5958 13035 6010
rect 12873 5956 12897 5958
rect 12953 5956 12977 5958
rect 13033 5956 13057 5958
rect 12817 5936 13113 5956
rect 13188 5574 13216 6752
rect 13280 5778 13308 7142
rect 13268 5772 13320 5778
rect 13268 5714 13320 5720
rect 13176 5568 13228 5574
rect 13176 5510 13228 5516
rect 13188 5370 13216 5510
rect 13176 5364 13228 5370
rect 13176 5306 13228 5312
rect 13174 5128 13230 5137
rect 13372 5114 13400 8842
rect 13464 8430 13492 9551
rect 13452 8424 13504 8430
rect 13452 8366 13504 8372
rect 13556 7562 13584 10202
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 13648 9722 13676 9998
rect 13636 9716 13688 9722
rect 13636 9658 13688 9664
rect 13740 9042 13768 11319
rect 13820 11290 13872 11296
rect 13924 11150 13952 12242
rect 14094 11928 14150 11937
rect 14292 11898 14320 13466
rect 14476 12102 14504 14554
rect 16120 14476 16172 14482
rect 16120 14418 16172 14424
rect 15384 14340 15436 14346
rect 15384 14282 15436 14288
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 14556 12708 14608 12714
rect 14556 12650 14608 12656
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14094 11863 14150 11872
rect 14280 11892 14332 11898
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 13464 7534 13584 7562
rect 13464 6458 13492 7534
rect 13544 7472 13596 7478
rect 13544 7414 13596 7420
rect 13556 7002 13584 7414
rect 13544 6996 13596 7002
rect 13544 6938 13596 6944
rect 13542 6760 13598 6769
rect 13542 6695 13598 6704
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13556 6254 13584 6695
rect 13648 6338 13676 8774
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13740 8090 13768 8434
rect 13832 8362 13860 9998
rect 13924 8922 13952 11086
rect 14108 11014 14136 11863
rect 14280 11834 14332 11840
rect 14372 11892 14424 11898
rect 14372 11834 14424 11840
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 14108 9722 14136 10950
rect 14200 9994 14228 11086
rect 14384 10810 14412 11834
rect 14568 11286 14596 12650
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 14844 12306 14872 12582
rect 14832 12300 14884 12306
rect 14832 12242 14884 12248
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14556 11280 14608 11286
rect 14556 11222 14608 11228
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14188 9988 14240 9994
rect 14188 9930 14240 9936
rect 14096 9716 14148 9722
rect 14096 9658 14148 9664
rect 14096 9512 14148 9518
rect 14096 9454 14148 9460
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 14016 9042 14044 9318
rect 14004 9036 14056 9042
rect 14004 8978 14056 8984
rect 13924 8894 14044 8922
rect 13912 8832 13964 8838
rect 13912 8774 13964 8780
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13818 7984 13874 7993
rect 13924 7954 13952 8774
rect 14016 8362 14044 8894
rect 14004 8356 14056 8362
rect 14004 8298 14056 8304
rect 13818 7919 13820 7928
rect 13872 7919 13874 7928
rect 13912 7948 13964 7954
rect 13820 7890 13872 7896
rect 13912 7890 13964 7896
rect 13832 7426 13860 7890
rect 13728 7404 13780 7410
rect 13832 7398 13952 7426
rect 13728 7346 13780 7352
rect 13740 6866 13768 7346
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13728 6724 13780 6730
rect 13728 6666 13780 6672
rect 13740 6458 13768 6666
rect 13832 6474 13860 7142
rect 13924 7002 13952 7398
rect 14108 7342 14136 9454
rect 14200 8974 14228 9930
rect 14280 9648 14332 9654
rect 14280 9590 14332 9596
rect 14292 9518 14320 9590
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14384 9382 14412 10746
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 14648 10124 14700 10130
rect 14648 10066 14700 10072
rect 14464 9920 14516 9926
rect 14464 9862 14516 9868
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 14372 9104 14424 9110
rect 14372 9046 14424 9052
rect 14384 8974 14412 9046
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14280 8356 14332 8362
rect 14280 8298 14332 8304
rect 14292 8265 14320 8298
rect 14278 8256 14334 8265
rect 14278 8191 14334 8200
rect 14384 8090 14412 8910
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14280 7744 14332 7750
rect 14280 7686 14332 7692
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 14016 7041 14044 7142
rect 14002 7032 14058 7041
rect 13912 6996 13964 7002
rect 14002 6967 14058 6976
rect 13912 6938 13964 6944
rect 14016 6633 14044 6967
rect 14002 6624 14058 6633
rect 14002 6559 14058 6568
rect 13728 6452 13780 6458
rect 13832 6446 13952 6474
rect 13728 6394 13780 6400
rect 13648 6310 13860 6338
rect 13544 6248 13596 6254
rect 13636 6248 13688 6254
rect 13544 6190 13596 6196
rect 13634 6216 13636 6225
rect 13688 6216 13690 6225
rect 13452 6112 13504 6118
rect 13450 6080 13452 6089
rect 13504 6080 13506 6089
rect 13450 6015 13506 6024
rect 13230 5086 13400 5114
rect 13174 5063 13230 5072
rect 12817 4924 13113 4944
rect 12873 4922 12897 4924
rect 12953 4922 12977 4924
rect 13033 4922 13057 4924
rect 12895 4870 12897 4922
rect 12959 4870 12971 4922
rect 13033 4870 13035 4922
rect 12873 4868 12897 4870
rect 12953 4868 12977 4870
rect 13033 4868 13057 4870
rect 12817 4848 13113 4868
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 13082 4720 13138 4729
rect 13188 4690 13216 5063
rect 13082 4655 13138 4664
rect 13176 4684 13228 4690
rect 12346 4111 12402 4120
rect 12624 4140 12676 4146
rect 12256 4072 12308 4078
rect 12256 4014 12308 4020
rect 12164 2984 12216 2990
rect 12164 2926 12216 2932
rect 12072 2848 12124 2854
rect 12072 2790 12124 2796
rect 12176 2514 12204 2926
rect 12360 2825 12388 4111
rect 12624 4082 12676 4088
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 12728 3670 12756 4082
rect 13096 4078 13124 4655
rect 13464 4672 13492 6015
rect 13176 4626 13228 4632
rect 13372 4644 13492 4672
rect 13084 4072 13136 4078
rect 13084 4014 13136 4020
rect 13176 3936 13228 3942
rect 13176 3878 13228 3884
rect 12817 3836 13113 3856
rect 12873 3834 12897 3836
rect 12953 3834 12977 3836
rect 13033 3834 13057 3836
rect 12895 3782 12897 3834
rect 12959 3782 12971 3834
rect 13033 3782 13035 3834
rect 12873 3780 12897 3782
rect 12953 3780 12977 3782
rect 13033 3780 13057 3782
rect 12817 3760 13113 3780
rect 12716 3664 12768 3670
rect 12716 3606 12768 3612
rect 12440 3528 12492 3534
rect 12438 3496 12440 3505
rect 12492 3496 12494 3505
rect 12438 3431 12494 3440
rect 13188 3194 13216 3878
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 13372 2990 13400 4644
rect 13556 3942 13584 6190
rect 13634 6151 13690 6160
rect 13728 6180 13780 6186
rect 13728 6122 13780 6128
rect 13634 6080 13690 6089
rect 13634 6015 13690 6024
rect 13648 5846 13676 6015
rect 13636 5840 13688 5846
rect 13636 5782 13688 5788
rect 13648 4826 13676 5782
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13452 3120 13504 3126
rect 13452 3062 13504 3068
rect 13360 2984 13412 2990
rect 13360 2926 13412 2932
rect 12624 2848 12676 2854
rect 12346 2816 12402 2825
rect 12624 2790 12676 2796
rect 12346 2751 12402 2760
rect 12636 2650 12664 2790
rect 12817 2748 13113 2768
rect 12873 2746 12897 2748
rect 12953 2746 12977 2748
rect 13033 2746 13057 2748
rect 12895 2694 12897 2746
rect 12959 2694 12971 2746
rect 13033 2694 13035 2746
rect 12873 2692 12897 2694
rect 12953 2692 12977 2694
rect 13033 2692 13057 2694
rect 12817 2672 13113 2692
rect 12624 2644 12676 2650
rect 12624 2586 12676 2592
rect 13464 2514 13492 3062
rect 13648 2854 13676 4014
rect 13636 2848 13688 2854
rect 13636 2790 13688 2796
rect 13740 2514 13768 6122
rect 13832 6118 13860 6310
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13820 5636 13872 5642
rect 13820 5578 13872 5584
rect 13832 5166 13860 5578
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 13832 4146 13860 4422
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13832 3738 13860 4082
rect 13820 3732 13872 3738
rect 13820 3674 13872 3680
rect 13924 3602 13952 6446
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 14016 6322 14044 6394
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 14016 5710 14044 6258
rect 14108 5914 14136 7278
rect 14188 6792 14240 6798
rect 14188 6734 14240 6740
rect 14200 6322 14228 6734
rect 14188 6316 14240 6322
rect 14188 6258 14240 6264
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 14096 5772 14148 5778
rect 14096 5714 14148 5720
rect 14004 5704 14056 5710
rect 14004 5646 14056 5652
rect 14004 5568 14056 5574
rect 14004 5510 14056 5516
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 13912 3392 13964 3398
rect 13912 3334 13964 3340
rect 13924 3074 13952 3334
rect 13832 3046 13952 3074
rect 12164 2508 12216 2514
rect 12164 2450 12216 2456
rect 13452 2508 13504 2514
rect 13452 2450 13504 2456
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 10784 2382 10836 2388
rect 11072 2400 11192 2428
rect 11796 2440 11848 2446
rect 10600 1896 10652 1902
rect 10600 1838 10652 1844
rect 11072 1834 11100 2400
rect 11796 2382 11848 2388
rect 11244 2372 11296 2378
rect 11244 2314 11296 2320
rect 11152 2304 11204 2310
rect 11152 2246 11204 2252
rect 11164 2106 11192 2246
rect 11152 2100 11204 2106
rect 11152 2042 11204 2048
rect 11060 1828 11112 1834
rect 11060 1770 11112 1776
rect 11256 800 11284 2314
rect 11336 2304 11388 2310
rect 11336 2246 11388 2252
rect 11348 2038 11376 2246
rect 11336 2032 11388 2038
rect 11336 1974 11388 1980
rect 12176 1562 12204 2450
rect 12256 2372 12308 2378
rect 12256 2314 12308 2320
rect 13084 2372 13136 2378
rect 13084 2314 13136 2320
rect 12164 1556 12216 1562
rect 12164 1498 12216 1504
rect 12268 1170 12296 2314
rect 12176 1142 12296 1170
rect 12176 800 12204 1142
rect 13096 800 13124 2314
rect 13832 2310 13860 3046
rect 13912 2848 13964 2854
rect 14016 2825 14044 5510
rect 14108 3398 14136 5714
rect 14200 5574 14228 6054
rect 14188 5568 14240 5574
rect 14188 5510 14240 5516
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 14200 4486 14228 5102
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 14188 3528 14240 3534
rect 14188 3470 14240 3476
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 13912 2790 13964 2796
rect 14002 2816 14058 2825
rect 13924 2650 13952 2790
rect 14002 2751 14058 2760
rect 13912 2644 13964 2650
rect 13912 2586 13964 2592
rect 13912 2372 13964 2378
rect 13912 2314 13964 2320
rect 13820 2304 13872 2310
rect 13820 2246 13872 2252
rect 13924 800 13952 2314
rect 14108 2310 14136 3334
rect 14096 2304 14148 2310
rect 14096 2246 14148 2252
rect 14200 1766 14228 3470
rect 14292 2990 14320 7686
rect 14384 7410 14412 8026
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14384 5846 14412 6734
rect 14372 5840 14424 5846
rect 14372 5782 14424 5788
rect 14370 4584 14426 4593
rect 14370 4519 14372 4528
rect 14424 4519 14426 4528
rect 14372 4490 14424 4496
rect 14370 4176 14426 4185
rect 14370 4111 14426 4120
rect 14384 4078 14412 4111
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 14280 2984 14332 2990
rect 14384 2961 14412 3878
rect 14476 2990 14504 9862
rect 14568 9654 14596 10066
rect 14556 9648 14608 9654
rect 14556 9590 14608 9596
rect 14660 9178 14688 10066
rect 14648 9172 14700 9178
rect 14648 9114 14700 9120
rect 14648 9036 14700 9042
rect 14648 8978 14700 8984
rect 14660 8498 14688 8978
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14554 8392 14610 8401
rect 14752 8378 14780 12038
rect 15028 11898 15056 14010
rect 15292 14000 15344 14006
rect 15292 13942 15344 13948
rect 15304 12986 15332 13942
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15304 12306 15332 12786
rect 15396 12374 15424 14282
rect 15782 14172 16078 14192
rect 15838 14170 15862 14172
rect 15918 14170 15942 14172
rect 15998 14170 16022 14172
rect 15860 14118 15862 14170
rect 15924 14118 15936 14170
rect 15998 14118 16000 14170
rect 15838 14116 15862 14118
rect 15918 14116 15942 14118
rect 15998 14116 16022 14118
rect 15782 14096 16078 14116
rect 16132 13938 16160 14418
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 16224 13870 16252 16487
rect 16486 15736 16542 15745
rect 16486 15671 16542 15680
rect 16500 14482 16528 15671
rect 16946 15464 17002 15473
rect 16946 15399 17002 15408
rect 16960 14482 16988 15399
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 16948 14476 17000 14482
rect 16948 14418 17000 14424
rect 16500 14074 16528 14418
rect 16580 14340 16632 14346
rect 16580 14282 16632 14288
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 16304 13728 16356 13734
rect 16304 13670 16356 13676
rect 15782 13084 16078 13104
rect 15838 13082 15862 13084
rect 15918 13082 15942 13084
rect 15998 13082 16022 13084
rect 15860 13030 15862 13082
rect 15924 13030 15936 13082
rect 15998 13030 16000 13082
rect 15838 13028 15862 13030
rect 15918 13028 15942 13030
rect 15998 13028 16022 13030
rect 15782 13008 16078 13028
rect 16316 12986 16344 13670
rect 16394 13560 16450 13569
rect 16394 13495 16396 13504
rect 16448 13495 16450 13504
rect 16396 13466 16448 13472
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 15568 12980 15620 12986
rect 15568 12922 15620 12928
rect 16304 12980 16356 12986
rect 16304 12922 16356 12928
rect 15384 12368 15436 12374
rect 15384 12310 15436 12316
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15016 11892 15068 11898
rect 15016 11834 15068 11840
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 15028 11694 15056 11834
rect 14924 11688 14976 11694
rect 14924 11630 14976 11636
rect 15016 11688 15068 11694
rect 15016 11630 15068 11636
rect 14936 11354 14964 11630
rect 14924 11348 14976 11354
rect 14924 11290 14976 11296
rect 15016 11076 15068 11082
rect 15016 11018 15068 11024
rect 15028 10606 15056 11018
rect 15120 10849 15148 11834
rect 15304 11626 15332 12242
rect 15292 11620 15344 11626
rect 15292 11562 15344 11568
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15106 10840 15162 10849
rect 15212 10810 15240 11154
rect 15106 10775 15162 10784
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 15016 10600 15068 10606
rect 15016 10542 15068 10548
rect 14924 10532 14976 10538
rect 14924 10474 14976 10480
rect 14936 10062 14964 10474
rect 14924 10056 14976 10062
rect 14924 9998 14976 10004
rect 14924 9648 14976 9654
rect 14924 9590 14976 9596
rect 14832 8560 14884 8566
rect 14832 8502 14884 8508
rect 14554 8327 14610 8336
rect 14660 8350 14780 8378
rect 14568 8294 14596 8327
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14568 7993 14596 8230
rect 14554 7984 14610 7993
rect 14554 7919 14610 7928
rect 14556 7268 14608 7274
rect 14556 7210 14608 7216
rect 14568 6458 14596 7210
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14554 4856 14610 4865
rect 14554 4791 14556 4800
rect 14608 4791 14610 4800
rect 14556 4762 14608 4768
rect 14660 4078 14688 8350
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14752 7342 14780 7686
rect 14740 7336 14792 7342
rect 14740 7278 14792 7284
rect 14738 7168 14794 7177
rect 14738 7103 14794 7112
rect 14752 5914 14780 7103
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 14752 4826 14780 5850
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14740 4276 14792 4282
rect 14740 4218 14792 4224
rect 14648 4072 14700 4078
rect 14554 4040 14610 4049
rect 14648 4014 14700 4020
rect 14554 3975 14610 3984
rect 14568 3602 14596 3975
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14556 3596 14608 3602
rect 14556 3538 14608 3544
rect 14660 3058 14688 3878
rect 14648 3052 14700 3058
rect 14648 2994 14700 3000
rect 14464 2984 14516 2990
rect 14280 2926 14332 2932
rect 14370 2952 14426 2961
rect 14464 2926 14516 2932
rect 14370 2887 14426 2896
rect 14280 2848 14332 2854
rect 14556 2848 14608 2854
rect 14280 2790 14332 2796
rect 14462 2816 14518 2825
rect 14292 2650 14320 2790
rect 14556 2790 14608 2796
rect 14462 2751 14518 2760
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 14188 1760 14240 1766
rect 14188 1702 14240 1708
rect 14292 1630 14320 2246
rect 14476 2106 14504 2751
rect 14568 2582 14596 2790
rect 14556 2576 14608 2582
rect 14556 2518 14608 2524
rect 14752 2514 14780 4218
rect 14844 2990 14872 8502
rect 14936 8362 14964 9590
rect 15028 9110 15056 10542
rect 15212 10062 15240 10746
rect 15304 10266 15332 11562
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 15396 9908 15424 12310
rect 15474 11928 15530 11937
rect 15474 11863 15530 11872
rect 15488 11762 15516 11863
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15476 10532 15528 10538
rect 15476 10474 15528 10480
rect 15120 9880 15424 9908
rect 15120 9518 15148 9880
rect 15488 9761 15516 10474
rect 15474 9752 15530 9761
rect 15292 9716 15344 9722
rect 15474 9687 15530 9696
rect 15292 9658 15344 9664
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 15212 9178 15240 9522
rect 15200 9172 15252 9178
rect 15200 9114 15252 9120
rect 15016 9104 15068 9110
rect 15304 9058 15332 9658
rect 15488 9654 15516 9687
rect 15476 9648 15528 9654
rect 15476 9590 15528 9596
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 15016 9046 15068 9052
rect 15108 9036 15160 9042
rect 15108 8978 15160 8984
rect 15212 9030 15332 9058
rect 15120 8430 15148 8978
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 14924 8356 14976 8362
rect 14924 8298 14976 8304
rect 14924 6860 14976 6866
rect 14924 6802 14976 6808
rect 14936 6390 14964 6802
rect 14924 6384 14976 6390
rect 14924 6326 14976 6332
rect 14922 6216 14978 6225
rect 14922 6151 14978 6160
rect 14936 5778 14964 6151
rect 15108 6112 15160 6118
rect 15108 6054 15160 6060
rect 15120 5914 15148 6054
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 15016 5840 15068 5846
rect 15016 5782 15068 5788
rect 14924 5772 14976 5778
rect 14924 5714 14976 5720
rect 14924 5636 14976 5642
rect 14924 5578 14976 5584
rect 14936 5166 14964 5578
rect 15028 5370 15056 5782
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 15016 5364 15068 5370
rect 15016 5306 15068 5312
rect 15028 5234 15056 5306
rect 15016 5228 15068 5234
rect 15016 5170 15068 5176
rect 14924 5160 14976 5166
rect 14924 5102 14976 5108
rect 15028 4622 15056 5170
rect 15120 4758 15148 5714
rect 15212 5681 15240 9030
rect 15290 8528 15346 8537
rect 15290 8463 15292 8472
rect 15344 8463 15346 8472
rect 15292 8434 15344 8440
rect 15396 7970 15424 9454
rect 15474 9072 15530 9081
rect 15474 9007 15530 9016
rect 15488 7993 15516 9007
rect 15304 7954 15424 7970
rect 15292 7948 15424 7954
rect 15344 7942 15424 7948
rect 15474 7984 15530 7993
rect 15474 7919 15530 7928
rect 15292 7890 15344 7896
rect 15292 7268 15344 7274
rect 15292 7210 15344 7216
rect 15198 5672 15254 5681
rect 15198 5607 15254 5616
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 15212 5166 15240 5510
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15108 4752 15160 4758
rect 15108 4694 15160 4700
rect 15016 4616 15068 4622
rect 15016 4558 15068 4564
rect 15108 4140 15160 4146
rect 15212 4128 15240 4966
rect 15160 4100 15240 4128
rect 15108 4082 15160 4088
rect 14924 3936 14976 3942
rect 14924 3878 14976 3884
rect 14936 3534 14964 3878
rect 14924 3528 14976 3534
rect 14924 3470 14976 3476
rect 14832 2984 14884 2990
rect 14832 2926 14884 2932
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 14936 2582 14964 2790
rect 15120 2650 15148 4082
rect 15304 3754 15332 7210
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 15212 3726 15332 3754
rect 15212 2854 15240 3726
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 15304 3194 15332 3538
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 15396 2990 15424 6054
rect 15488 5166 15516 7919
rect 15580 7274 15608 12922
rect 16408 12434 16436 13262
rect 16488 12640 16540 12646
rect 16488 12582 16540 12588
rect 16316 12406 16436 12434
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15672 10554 15700 12242
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 15782 11996 16078 12016
rect 15838 11994 15862 11996
rect 15918 11994 15942 11996
rect 15998 11994 16022 11996
rect 15860 11942 15862 11994
rect 15924 11942 15936 11994
rect 15998 11942 16000 11994
rect 15838 11940 15862 11942
rect 15918 11940 15942 11942
rect 15998 11940 16022 11942
rect 15782 11920 16078 11940
rect 15782 10908 16078 10928
rect 15838 10906 15862 10908
rect 15918 10906 15942 10908
rect 15998 10906 16022 10908
rect 15860 10854 15862 10906
rect 15924 10854 15936 10906
rect 15998 10854 16000 10906
rect 15838 10852 15862 10854
rect 15918 10852 15942 10854
rect 15998 10852 16022 10854
rect 15782 10832 16078 10852
rect 15672 10526 15792 10554
rect 15660 10464 15712 10470
rect 15660 10406 15712 10412
rect 15672 9466 15700 10406
rect 15764 10033 15792 10526
rect 16132 10130 16160 12038
rect 16212 11688 16264 11694
rect 16212 11630 16264 11636
rect 16120 10124 16172 10130
rect 16120 10066 16172 10072
rect 15750 10024 15806 10033
rect 15750 9959 15806 9968
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 15782 9820 16078 9840
rect 15838 9818 15862 9820
rect 15918 9818 15942 9820
rect 15998 9818 16022 9820
rect 15860 9766 15862 9818
rect 15924 9766 15936 9818
rect 15998 9766 16000 9818
rect 15838 9764 15862 9766
rect 15918 9764 15942 9766
rect 15998 9764 16022 9766
rect 15782 9744 16078 9764
rect 16026 9688 16082 9697
rect 16026 9623 16082 9632
rect 15672 9438 15976 9466
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15764 8945 15792 9318
rect 15948 9110 15976 9438
rect 15844 9104 15896 9110
rect 15844 9046 15896 9052
rect 15936 9104 15988 9110
rect 16040 9081 16068 9623
rect 16132 9586 16160 9862
rect 16120 9580 16172 9586
rect 16120 9522 16172 9528
rect 16224 9518 16252 11630
rect 16212 9512 16264 9518
rect 16212 9454 16264 9460
rect 15936 9046 15988 9052
rect 16026 9072 16082 9081
rect 15856 8974 15884 9046
rect 15844 8968 15896 8974
rect 15750 8936 15806 8945
rect 15844 8910 15896 8916
rect 15750 8871 15806 8880
rect 15660 8832 15712 8838
rect 15948 8820 15976 9046
rect 16026 9007 16082 9016
rect 16212 8832 16264 8838
rect 15948 8792 16160 8820
rect 15660 8774 15712 8780
rect 15672 8362 15700 8774
rect 15782 8732 16078 8752
rect 15838 8730 15862 8732
rect 15918 8730 15942 8732
rect 15998 8730 16022 8732
rect 15860 8678 15862 8730
rect 15924 8678 15936 8730
rect 15998 8678 16000 8730
rect 15838 8676 15862 8678
rect 15918 8676 15942 8678
rect 15998 8676 16022 8678
rect 15782 8656 16078 8676
rect 16132 8616 16160 8792
rect 16212 8774 16264 8780
rect 16040 8588 16160 8616
rect 16040 8498 16068 8588
rect 16028 8492 16080 8498
rect 16028 8434 16080 8440
rect 15936 8424 15988 8430
rect 16224 8378 16252 8774
rect 16316 8650 16344 12406
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16408 11898 16436 12038
rect 16396 11892 16448 11898
rect 16396 11834 16448 11840
rect 16396 11552 16448 11558
rect 16394 11520 16396 11529
rect 16448 11520 16450 11529
rect 16394 11455 16450 11464
rect 16500 11218 16528 12582
rect 16592 12238 16620 14282
rect 16960 14006 16988 14418
rect 16948 14000 17000 14006
rect 16948 13942 17000 13948
rect 17224 14000 17276 14006
rect 17224 13942 17276 13948
rect 17132 13864 17184 13870
rect 17132 13806 17184 13812
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16684 12374 16712 13262
rect 16948 13252 17000 13258
rect 16948 13194 17000 13200
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16764 12640 16816 12646
rect 16764 12582 16816 12588
rect 16672 12368 16724 12374
rect 16672 12310 16724 12316
rect 16580 12232 16632 12238
rect 16580 12174 16632 12180
rect 16578 11928 16634 11937
rect 16578 11863 16634 11872
rect 16592 11762 16620 11863
rect 16684 11830 16712 12310
rect 16672 11824 16724 11830
rect 16672 11766 16724 11772
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16776 11642 16804 12582
rect 16868 11898 16896 12922
rect 16960 12442 16988 13194
rect 17038 12744 17094 12753
rect 17038 12679 17094 12688
rect 17052 12442 17080 12679
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 16960 12170 16988 12378
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16856 11892 16908 11898
rect 16856 11834 16908 11840
rect 16592 11614 16804 11642
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 16592 11098 16620 11614
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16776 11218 16804 11494
rect 16868 11393 16896 11494
rect 16854 11384 16910 11393
rect 16854 11319 16910 11328
rect 16764 11212 16816 11218
rect 16764 11154 16816 11160
rect 16408 11082 16620 11098
rect 16396 11076 16620 11082
rect 16448 11070 16620 11076
rect 16396 11018 16448 11024
rect 16488 11008 16540 11014
rect 16488 10950 16540 10956
rect 16500 10538 16528 10950
rect 16396 10532 16448 10538
rect 16396 10474 16448 10480
rect 16488 10532 16540 10538
rect 16488 10474 16540 10480
rect 16408 9722 16436 10474
rect 16500 9994 16528 10474
rect 16592 10130 16620 11070
rect 16672 11076 16724 11082
rect 16672 11018 16724 11024
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 16488 9988 16540 9994
rect 16488 9930 16540 9936
rect 16580 9920 16632 9926
rect 16486 9888 16542 9897
rect 16580 9862 16632 9868
rect 16486 9823 16542 9832
rect 16396 9716 16448 9722
rect 16396 9658 16448 9664
rect 16500 9217 16528 9823
rect 16592 9518 16620 9862
rect 16580 9512 16632 9518
rect 16580 9454 16632 9460
rect 16684 9450 16712 11018
rect 16672 9444 16724 9450
rect 16672 9386 16724 9392
rect 16486 9208 16542 9217
rect 16486 9143 16542 9152
rect 16500 9024 16528 9143
rect 16500 8996 16620 9024
rect 16316 8622 16436 8650
rect 15988 8372 16252 8378
rect 15936 8366 16252 8372
rect 15660 8356 15712 8362
rect 15948 8350 16252 8366
rect 16302 8392 16358 8401
rect 16302 8327 16358 8336
rect 15660 8298 15712 8304
rect 16118 8256 16174 8265
rect 16118 8191 16174 8200
rect 15782 7644 16078 7664
rect 15838 7642 15862 7644
rect 15918 7642 15942 7644
rect 15998 7642 16022 7644
rect 15860 7590 15862 7642
rect 15924 7590 15936 7642
rect 15998 7590 16000 7642
rect 15838 7588 15862 7590
rect 15918 7588 15942 7590
rect 15998 7588 16022 7590
rect 15782 7568 16078 7588
rect 15660 7336 15712 7342
rect 15660 7278 15712 7284
rect 15568 7268 15620 7274
rect 15568 7210 15620 7216
rect 15672 6934 15700 7278
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 16028 7200 16080 7206
rect 16028 7142 16080 7148
rect 15856 6934 15884 7142
rect 15660 6928 15712 6934
rect 15660 6870 15712 6876
rect 15844 6928 15896 6934
rect 15844 6870 15896 6876
rect 15660 6792 15712 6798
rect 16040 6769 16068 7142
rect 15660 6734 15712 6740
rect 16026 6760 16082 6769
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15580 6322 15608 6598
rect 15568 6316 15620 6322
rect 15568 6258 15620 6264
rect 15672 5846 15700 6734
rect 16026 6695 16082 6704
rect 15782 6556 16078 6576
rect 15838 6554 15862 6556
rect 15918 6554 15942 6556
rect 15998 6554 16022 6556
rect 15860 6502 15862 6554
rect 15924 6502 15936 6554
rect 15998 6502 16000 6554
rect 15838 6500 15862 6502
rect 15918 6500 15942 6502
rect 15998 6500 16022 6502
rect 15782 6480 16078 6500
rect 16132 6338 16160 8191
rect 16212 8084 16264 8090
rect 16212 8026 16264 8032
rect 16224 7993 16252 8026
rect 16210 7984 16266 7993
rect 16316 7954 16344 8327
rect 16210 7919 16266 7928
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16212 7880 16264 7886
rect 16212 7822 16264 7828
rect 16224 7410 16252 7822
rect 16212 7404 16264 7410
rect 16212 7346 16264 7352
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16316 7041 16344 7142
rect 16302 7032 16358 7041
rect 16302 6967 16358 6976
rect 16212 6928 16264 6934
rect 16212 6870 16264 6876
rect 15764 6310 16160 6338
rect 16224 6322 16252 6870
rect 16212 6316 16264 6322
rect 15660 5840 15712 5846
rect 15660 5782 15712 5788
rect 15568 5704 15620 5710
rect 15764 5658 15792 6310
rect 16212 6258 16264 6264
rect 16120 5772 16172 5778
rect 16120 5714 16172 5720
rect 15568 5646 15620 5652
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 15488 3058 15516 4966
rect 15580 3738 15608 5646
rect 15672 5630 15792 5658
rect 15672 5166 15700 5630
rect 15782 5468 16078 5488
rect 15838 5466 15862 5468
rect 15918 5466 15942 5468
rect 15998 5466 16022 5468
rect 15860 5414 15862 5466
rect 15924 5414 15936 5466
rect 15998 5414 16000 5466
rect 15838 5412 15862 5414
rect 15918 5412 15942 5414
rect 15998 5412 16022 5414
rect 15782 5392 16078 5412
rect 15750 5264 15806 5273
rect 15750 5199 15806 5208
rect 15660 5160 15712 5166
rect 15660 5102 15712 5108
rect 15672 4865 15700 5102
rect 15658 4856 15714 4865
rect 15658 4791 15714 4800
rect 15764 4706 15792 5199
rect 15934 5128 15990 5137
rect 15934 5063 15936 5072
rect 15988 5063 15990 5072
rect 15936 5034 15988 5040
rect 15672 4678 15792 4706
rect 15568 3732 15620 3738
rect 15568 3674 15620 3680
rect 15672 3602 15700 4678
rect 15782 4380 16078 4400
rect 15838 4378 15862 4380
rect 15918 4378 15942 4380
rect 15998 4378 16022 4380
rect 15860 4326 15862 4378
rect 15924 4326 15936 4378
rect 15998 4326 16000 4378
rect 15838 4324 15862 4326
rect 15918 4324 15942 4326
rect 15998 4324 16022 4326
rect 15782 4304 16078 4324
rect 16132 3777 16160 5714
rect 16212 5636 16264 5642
rect 16212 5578 16264 5584
rect 16224 5234 16252 5578
rect 16212 5228 16264 5234
rect 16212 5170 16264 5176
rect 16224 4758 16252 5170
rect 16316 5166 16344 6967
rect 16408 5778 16436 8622
rect 16488 8424 16540 8430
rect 16488 8366 16540 8372
rect 16500 8129 16528 8366
rect 16486 8120 16542 8129
rect 16486 8055 16542 8064
rect 16592 7426 16620 8996
rect 16672 8560 16724 8566
rect 16672 8502 16724 8508
rect 16684 8401 16712 8502
rect 16670 8392 16726 8401
rect 16670 8327 16726 8336
rect 16672 7948 16724 7954
rect 16672 7890 16724 7896
rect 16684 7546 16712 7890
rect 16776 7857 16804 11154
rect 16856 11008 16908 11014
rect 16856 10950 16908 10956
rect 16868 9042 16896 10950
rect 16960 10810 16988 12106
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 17052 11694 17080 12038
rect 17144 11937 17172 13806
rect 17236 13530 17264 13942
rect 17328 13802 17356 16895
rect 17866 16400 17922 17200
rect 17774 16144 17830 16153
rect 17774 16079 17830 16088
rect 17682 15056 17738 15065
rect 17682 14991 17738 15000
rect 17500 14816 17552 14822
rect 17500 14758 17552 14764
rect 17512 14550 17540 14758
rect 17696 14550 17724 14991
rect 17500 14544 17552 14550
rect 17500 14486 17552 14492
rect 17684 14544 17736 14550
rect 17684 14486 17736 14492
rect 17500 14340 17552 14346
rect 17500 14282 17552 14288
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17420 13841 17448 14214
rect 17406 13832 17462 13841
rect 17316 13796 17368 13802
rect 17406 13767 17462 13776
rect 17316 13738 17368 13744
rect 17224 13524 17276 13530
rect 17224 13466 17276 13472
rect 17328 13190 17356 13738
rect 17316 13184 17368 13190
rect 17316 13126 17368 13132
rect 17316 12912 17368 12918
rect 17316 12854 17368 12860
rect 17224 12300 17276 12306
rect 17224 12242 17276 12248
rect 17130 11928 17186 11937
rect 17236 11898 17264 12242
rect 17130 11863 17186 11872
rect 17224 11892 17276 11898
rect 17224 11834 17276 11840
rect 17132 11824 17184 11830
rect 17132 11766 17184 11772
rect 17040 11688 17092 11694
rect 17038 11656 17040 11665
rect 17092 11656 17094 11665
rect 17038 11591 17094 11600
rect 17040 11212 17092 11218
rect 17040 11154 17092 11160
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 16960 9518 16988 10542
rect 17052 10470 17080 11154
rect 17040 10464 17092 10470
rect 17040 10406 17092 10412
rect 17052 10266 17080 10406
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 17144 10198 17172 11766
rect 17224 10804 17276 10810
rect 17224 10746 17276 10752
rect 17132 10192 17184 10198
rect 17132 10134 17184 10140
rect 17040 10124 17092 10130
rect 17040 10066 17092 10072
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16960 9178 16988 9454
rect 16948 9172 17000 9178
rect 16948 9114 17000 9120
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 17052 8974 17080 10066
rect 17236 10010 17264 10746
rect 17144 9982 17264 10010
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 17052 8650 17080 8910
rect 16960 8622 17080 8650
rect 16960 8362 16988 8622
rect 17040 8560 17092 8566
rect 17040 8502 17092 8508
rect 16948 8356 17000 8362
rect 16948 8298 17000 8304
rect 16762 7848 16818 7857
rect 16762 7783 16818 7792
rect 16672 7540 16724 7546
rect 16672 7482 16724 7488
rect 16592 7398 16712 7426
rect 16488 6996 16540 7002
rect 16488 6938 16540 6944
rect 16500 5794 16528 6938
rect 16580 6452 16632 6458
rect 16580 6394 16632 6400
rect 16592 6254 16620 6394
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 16396 5772 16448 5778
rect 16500 5766 16620 5794
rect 16396 5714 16448 5720
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16396 5568 16448 5574
rect 16396 5510 16448 5516
rect 16304 5160 16356 5166
rect 16304 5102 16356 5108
rect 16212 4752 16264 4758
rect 16212 4694 16264 4700
rect 16304 4684 16356 4690
rect 16304 4626 16356 4632
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 16224 4078 16252 4422
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16118 3768 16174 3777
rect 16118 3703 16174 3712
rect 16224 3602 16252 4014
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 16212 3596 16264 3602
rect 16212 3538 16264 3544
rect 16316 3466 16344 4626
rect 16408 3754 16436 5510
rect 16500 4146 16528 5646
rect 16592 4690 16620 5766
rect 16684 5234 16712 7398
rect 16776 7002 16804 7783
rect 16856 7744 16908 7750
rect 16856 7686 16908 7692
rect 16948 7744 17000 7750
rect 16948 7686 17000 7692
rect 16764 6996 16816 7002
rect 16764 6938 16816 6944
rect 16868 6322 16896 7686
rect 16960 6322 16988 7686
rect 17052 6390 17080 8502
rect 17144 7206 17172 9982
rect 17224 9444 17276 9450
rect 17224 9386 17276 9392
rect 17236 8838 17264 9386
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 17236 8498 17264 8774
rect 17224 8492 17276 8498
rect 17224 8434 17276 8440
rect 17224 8288 17276 8294
rect 17224 8230 17276 8236
rect 17132 7200 17184 7206
rect 17132 7142 17184 7148
rect 17040 6384 17092 6390
rect 17040 6326 17092 6332
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 17052 6202 17080 6326
rect 16960 6174 17080 6202
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 16672 5228 16724 5234
rect 16672 5170 16724 5176
rect 16672 4752 16724 4758
rect 16672 4694 16724 4700
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 16592 4282 16620 4626
rect 16580 4276 16632 4282
rect 16580 4218 16632 4224
rect 16488 4140 16540 4146
rect 16488 4082 16540 4088
rect 16408 3738 16528 3754
rect 16408 3732 16540 3738
rect 16408 3726 16488 3732
rect 16488 3674 16540 3680
rect 16486 3632 16542 3641
rect 16396 3596 16448 3602
rect 16486 3567 16542 3576
rect 16396 3538 16448 3544
rect 16212 3460 16264 3466
rect 16212 3402 16264 3408
rect 16304 3460 16356 3466
rect 16304 3402 16356 3408
rect 15660 3392 15712 3398
rect 15660 3334 15712 3340
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15476 3052 15528 3058
rect 15476 2994 15528 3000
rect 15384 2984 15436 2990
rect 15384 2926 15436 2932
rect 15476 2916 15528 2922
rect 15476 2858 15528 2864
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 15108 2644 15160 2650
rect 15108 2586 15160 2592
rect 14924 2576 14976 2582
rect 14924 2518 14976 2524
rect 14740 2508 14792 2514
rect 14740 2450 14792 2456
rect 14832 2372 14884 2378
rect 14832 2314 14884 2320
rect 14464 2100 14516 2106
rect 14464 2042 14516 2048
rect 14280 1624 14332 1630
rect 14280 1566 14332 1572
rect 14844 800 14872 2314
rect 3422 776 3478 785
rect 3422 711 3478 720
rect 3974 0 4030 800
rect 4894 0 4950 800
rect 5814 0 5870 800
rect 6734 0 6790 800
rect 7562 0 7618 800
rect 8482 0 8538 800
rect 9402 0 9458 800
rect 10322 0 10378 800
rect 11242 0 11298 800
rect 12162 0 12218 800
rect 13082 0 13138 800
rect 13910 0 13966 800
rect 14830 0 14886 800
rect 15488 241 15516 2858
rect 15580 2854 15608 3130
rect 15672 2990 15700 3334
rect 15782 3292 16078 3312
rect 15838 3290 15862 3292
rect 15918 3290 15942 3292
rect 15998 3290 16022 3292
rect 15860 3238 15862 3290
rect 15924 3238 15936 3290
rect 15998 3238 16000 3290
rect 15838 3236 15862 3238
rect 15918 3236 15942 3238
rect 15998 3236 16022 3238
rect 15782 3216 16078 3236
rect 16224 2990 16252 3402
rect 16408 3058 16436 3538
rect 16500 3058 16528 3567
rect 16684 3534 16712 4694
rect 16960 4690 16988 6174
rect 17040 6112 17092 6118
rect 17040 6054 17092 6060
rect 17052 5914 17080 6054
rect 17040 5908 17092 5914
rect 17040 5850 17092 5856
rect 17040 5772 17092 5778
rect 17040 5714 17092 5720
rect 17052 5370 17080 5714
rect 17040 5364 17092 5370
rect 17040 5306 17092 5312
rect 16948 4684 17000 4690
rect 16948 4626 17000 4632
rect 17144 4622 17172 6190
rect 17236 6118 17264 8230
rect 17224 6112 17276 6118
rect 17224 6054 17276 6060
rect 17328 5114 17356 12854
rect 17512 12782 17540 14282
rect 17696 14090 17724 14486
rect 17604 14062 17724 14090
rect 17604 13530 17632 14062
rect 17788 14006 17816 16079
rect 17880 14618 17908 16400
rect 18142 14648 18198 14657
rect 17868 14612 17920 14618
rect 18142 14583 18198 14592
rect 17868 14554 17920 14560
rect 18156 14482 18184 14583
rect 18144 14476 18196 14482
rect 18144 14418 18196 14424
rect 18420 14476 18472 14482
rect 18420 14418 18472 14424
rect 18156 14074 18184 14418
rect 18328 14272 18380 14278
rect 18432 14249 18460 14418
rect 18512 14340 18564 14346
rect 18512 14282 18564 14288
rect 18328 14214 18380 14220
rect 18418 14240 18474 14249
rect 18144 14068 18196 14074
rect 18144 14010 18196 14016
rect 17776 14000 17828 14006
rect 17776 13942 17828 13948
rect 17684 13932 17736 13938
rect 17684 13874 17736 13880
rect 17592 13524 17644 13530
rect 17592 13466 17644 13472
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17604 12889 17632 13126
rect 17590 12880 17646 12889
rect 17590 12815 17646 12824
rect 17500 12776 17552 12782
rect 17500 12718 17552 12724
rect 17500 12640 17552 12646
rect 17500 12582 17552 12588
rect 17512 12434 17540 12582
rect 17512 12406 17632 12434
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 17420 11218 17448 12038
rect 17512 11937 17540 12174
rect 17498 11928 17554 11937
rect 17498 11863 17554 11872
rect 17512 11694 17540 11863
rect 17500 11688 17552 11694
rect 17500 11630 17552 11636
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17408 11212 17460 11218
rect 17408 11154 17460 11160
rect 17420 10441 17448 11154
rect 17512 10713 17540 11494
rect 17498 10704 17554 10713
rect 17498 10639 17554 10648
rect 17406 10432 17462 10441
rect 17406 10367 17462 10376
rect 17500 10192 17552 10198
rect 17500 10134 17552 10140
rect 17408 9988 17460 9994
rect 17408 9930 17460 9936
rect 17420 8294 17448 9930
rect 17512 8838 17540 10134
rect 17500 8832 17552 8838
rect 17500 8774 17552 8780
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17408 7200 17460 7206
rect 17408 7142 17460 7148
rect 17420 7002 17448 7142
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17408 6792 17460 6798
rect 17408 6734 17460 6740
rect 17420 5302 17448 6734
rect 17408 5296 17460 5302
rect 17408 5238 17460 5244
rect 17236 5086 17356 5114
rect 17132 4616 17184 4622
rect 17132 4558 17184 4564
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 17144 4146 17172 4422
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 16960 3738 16988 3878
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 16764 3460 16816 3466
rect 16764 3402 16816 3408
rect 16672 3392 16724 3398
rect 16672 3334 16724 3340
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 16488 3052 16540 3058
rect 16488 2994 16540 3000
rect 16684 2990 16712 3334
rect 15660 2984 15712 2990
rect 15660 2926 15712 2932
rect 16212 2984 16264 2990
rect 16212 2926 16264 2932
rect 16672 2984 16724 2990
rect 16672 2926 16724 2932
rect 16028 2916 16080 2922
rect 16028 2858 16080 2864
rect 16488 2916 16540 2922
rect 16488 2858 16540 2864
rect 15568 2848 15620 2854
rect 15568 2790 15620 2796
rect 15936 2848 15988 2854
rect 15936 2790 15988 2796
rect 15948 2582 15976 2790
rect 15936 2576 15988 2582
rect 15936 2518 15988 2524
rect 16040 2514 16068 2858
rect 16212 2848 16264 2854
rect 16212 2790 16264 2796
rect 16028 2508 16080 2514
rect 16028 2450 16080 2456
rect 15660 2372 15712 2378
rect 15660 2314 15712 2320
rect 15672 1170 15700 2314
rect 15782 2204 16078 2224
rect 15838 2202 15862 2204
rect 15918 2202 15942 2204
rect 15998 2202 16022 2204
rect 15860 2150 15862 2202
rect 15924 2150 15936 2202
rect 15998 2150 16000 2202
rect 15838 2148 15862 2150
rect 15918 2148 15942 2150
rect 15998 2148 16022 2150
rect 15782 2128 16078 2148
rect 16224 2106 16252 2790
rect 16212 2100 16264 2106
rect 16212 2042 16264 2048
rect 15672 1142 15792 1170
rect 15764 800 15792 1142
rect 15474 232 15530 241
rect 15474 167 15530 176
rect 15750 0 15806 800
rect 16500 513 16528 2858
rect 16580 2848 16632 2854
rect 16580 2790 16632 2796
rect 16592 2446 16620 2790
rect 16580 2440 16632 2446
rect 16580 2382 16632 2388
rect 16776 898 16804 3402
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 16868 2990 16896 3130
rect 16856 2984 16908 2990
rect 16856 2926 16908 2932
rect 17236 2774 17264 5086
rect 17316 5024 17368 5030
rect 17316 4966 17368 4972
rect 17408 5024 17460 5030
rect 17408 4966 17460 4972
rect 17328 4078 17356 4966
rect 17420 4826 17448 4966
rect 17512 4826 17540 8570
rect 17408 4820 17460 4826
rect 17408 4762 17460 4768
rect 17500 4820 17552 4826
rect 17500 4762 17552 4768
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17316 4072 17368 4078
rect 17316 4014 17368 4020
rect 17420 3398 17448 4558
rect 17500 3596 17552 3602
rect 17500 3538 17552 3544
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 16960 2746 17264 2774
rect 16854 2680 16910 2689
rect 16854 2615 16910 2624
rect 16868 2582 16896 2615
rect 16960 2582 16988 2746
rect 16856 2576 16908 2582
rect 16856 2518 16908 2524
rect 16948 2576 17000 2582
rect 16948 2518 17000 2524
rect 17512 2514 17540 3538
rect 17604 2990 17632 12406
rect 17696 11354 17724 13874
rect 17788 13802 17816 13942
rect 17960 13932 18012 13938
rect 17960 13874 18012 13880
rect 17776 13796 17828 13802
rect 17776 13738 17828 13744
rect 17774 13560 17830 13569
rect 17774 13495 17776 13504
rect 17828 13495 17830 13504
rect 17776 13466 17828 13472
rect 17868 12708 17920 12714
rect 17868 12650 17920 12656
rect 17880 12345 17908 12650
rect 17866 12336 17922 12345
rect 17866 12271 17922 12280
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 17684 11348 17736 11354
rect 17684 11290 17736 11296
rect 17776 11280 17828 11286
rect 17776 11222 17828 11228
rect 17684 11076 17736 11082
rect 17684 11018 17736 11024
rect 17696 9110 17724 11018
rect 17788 10130 17816 11222
rect 17880 10554 17908 12038
rect 17972 11257 18000 13874
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 18052 13388 18104 13394
rect 18052 13330 18104 13336
rect 18064 13161 18092 13330
rect 18050 13152 18106 13161
rect 18050 13087 18106 13096
rect 18050 12744 18106 12753
rect 18050 12679 18052 12688
rect 18104 12679 18106 12688
rect 18144 12708 18196 12714
rect 18052 12650 18104 12656
rect 18144 12650 18196 12656
rect 18052 12096 18104 12102
rect 18052 12038 18104 12044
rect 17958 11248 18014 11257
rect 17958 11183 18014 11192
rect 17880 10526 18000 10554
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 17776 9920 17828 9926
rect 17776 9862 17828 9868
rect 17788 9178 17816 9862
rect 17880 9722 17908 10406
rect 17868 9716 17920 9722
rect 17868 9658 17920 9664
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17684 9104 17736 9110
rect 17684 9046 17736 9052
rect 17880 8974 17908 9658
rect 17972 9194 18000 10526
rect 18064 9353 18092 12038
rect 18156 11801 18184 12650
rect 18142 11792 18198 11801
rect 18142 11727 18198 11736
rect 18142 11656 18198 11665
rect 18142 11591 18144 11600
rect 18196 11591 18198 11600
rect 18144 11562 18196 11568
rect 18144 11144 18196 11150
rect 18144 11086 18196 11092
rect 18156 10062 18184 11086
rect 18248 10198 18276 13466
rect 18340 12986 18368 14214
rect 18418 14175 18474 14184
rect 18420 13864 18472 13870
rect 18418 13832 18420 13841
rect 18472 13832 18474 13841
rect 18418 13767 18474 13776
rect 18418 13560 18474 13569
rect 18418 13495 18474 13504
rect 18432 13462 18460 13495
rect 18420 13456 18472 13462
rect 18420 13398 18472 13404
rect 18328 12980 18380 12986
rect 18328 12922 18380 12928
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 18432 12345 18460 12718
rect 18418 12336 18474 12345
rect 18418 12271 18474 12280
rect 18420 12164 18472 12170
rect 18420 12106 18472 12112
rect 18432 11626 18460 12106
rect 18420 11620 18472 11626
rect 18420 11562 18472 11568
rect 18432 10849 18460 11562
rect 18524 11121 18552 14282
rect 18972 11280 19024 11286
rect 18970 11248 18972 11257
rect 19024 11248 19026 11257
rect 18970 11183 19026 11192
rect 18510 11112 18566 11121
rect 18510 11047 18566 11056
rect 18418 10840 18474 10849
rect 18418 10775 18474 10784
rect 18512 10464 18564 10470
rect 18512 10406 18564 10412
rect 18236 10192 18288 10198
rect 18236 10134 18288 10140
rect 18144 10056 18196 10062
rect 18144 9998 18196 10004
rect 18248 9994 18276 10134
rect 18524 10033 18552 10406
rect 18510 10024 18566 10033
rect 18236 9988 18288 9994
rect 18566 9982 18644 10010
rect 18510 9959 18566 9968
rect 18236 9930 18288 9936
rect 18510 9752 18566 9761
rect 18510 9687 18566 9696
rect 18524 9654 18552 9687
rect 18512 9648 18564 9654
rect 18512 9590 18564 9596
rect 18328 9376 18380 9382
rect 18050 9344 18106 9353
rect 18328 9318 18380 9324
rect 18050 9279 18106 9288
rect 17972 9166 18092 9194
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17776 7948 17828 7954
rect 17776 7890 17828 7896
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 17696 7478 17724 7822
rect 17788 7546 17816 7890
rect 17880 7834 17908 8774
rect 17960 8356 18012 8362
rect 17960 8298 18012 8304
rect 17972 8022 18000 8298
rect 17960 8016 18012 8022
rect 17960 7958 18012 7964
rect 17880 7806 18000 7834
rect 17866 7712 17922 7721
rect 17866 7647 17922 7656
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 17684 7472 17736 7478
rect 17684 7414 17736 7420
rect 17880 6866 17908 7647
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 17972 6746 18000 7806
rect 18064 7313 18092 9166
rect 18144 8356 18196 8362
rect 18144 8298 18196 8304
rect 18156 7449 18184 8298
rect 18142 7440 18198 7449
rect 18340 7410 18368 9318
rect 18524 9042 18552 9590
rect 18512 9036 18564 9042
rect 18512 8978 18564 8984
rect 18616 8430 18644 9982
rect 18604 8424 18656 8430
rect 18604 8366 18656 8372
rect 18142 7375 18198 7384
rect 18328 7404 18380 7410
rect 18328 7346 18380 7352
rect 18050 7304 18106 7313
rect 18050 7239 18106 7248
rect 18328 7268 18380 7274
rect 17880 6718 18000 6746
rect 17684 6656 17736 6662
rect 17684 6598 17736 6604
rect 17696 6322 17724 6598
rect 17880 6458 17908 6718
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 17684 6316 17736 6322
rect 17684 6258 17736 6264
rect 17696 5846 17724 6258
rect 17868 6112 17920 6118
rect 17868 6054 17920 6060
rect 17684 5840 17736 5846
rect 17684 5782 17736 5788
rect 17696 5302 17724 5782
rect 17776 5568 17828 5574
rect 17880 5545 17908 6054
rect 17776 5510 17828 5516
rect 17866 5536 17922 5545
rect 17684 5296 17736 5302
rect 17684 5238 17736 5244
rect 17684 5024 17736 5030
rect 17684 4966 17736 4972
rect 17696 3670 17724 4966
rect 17788 4146 17816 5510
rect 17866 5471 17922 5480
rect 17868 5228 17920 5234
rect 17868 5170 17920 5176
rect 17880 4622 17908 5170
rect 18064 5166 18092 7239
rect 18328 7210 18380 7216
rect 18144 7200 18196 7206
rect 18144 7142 18196 7148
rect 18156 5914 18184 7142
rect 18234 7032 18290 7041
rect 18234 6967 18290 6976
rect 18248 6866 18276 6967
rect 18340 6866 18368 7210
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 18328 6860 18380 6866
rect 18328 6802 18380 6808
rect 18512 6724 18564 6730
rect 18512 6666 18564 6672
rect 18524 6633 18552 6666
rect 18510 6624 18566 6633
rect 18510 6559 18566 6568
rect 18510 6216 18566 6225
rect 18510 6151 18512 6160
rect 18564 6151 18566 6160
rect 18512 6122 18564 6128
rect 18510 5944 18566 5953
rect 18144 5908 18196 5914
rect 18510 5879 18566 5888
rect 18144 5850 18196 5856
rect 18524 5846 18552 5879
rect 18512 5840 18564 5846
rect 18512 5782 18564 5788
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 18510 5128 18566 5137
rect 18510 5063 18512 5072
rect 18564 5063 18566 5072
rect 18512 5034 18564 5040
rect 17960 5024 18012 5030
rect 17960 4966 18012 4972
rect 17868 4616 17920 4622
rect 17868 4558 17920 4564
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 17972 3670 18000 4966
rect 18510 4720 18566 4729
rect 18510 4655 18512 4664
rect 18564 4655 18566 4664
rect 18512 4626 18564 4632
rect 18052 4548 18104 4554
rect 18052 4490 18104 4496
rect 18064 4078 18092 4490
rect 18328 4480 18380 4486
rect 18328 4422 18380 4428
rect 18142 4312 18198 4321
rect 18142 4247 18198 4256
rect 18156 4146 18184 4247
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 17684 3664 17736 3670
rect 17684 3606 17736 3612
rect 17960 3664 18012 3670
rect 17960 3606 18012 3612
rect 18142 3632 18198 3641
rect 18142 3567 18144 3576
rect 18196 3567 18198 3576
rect 18144 3538 18196 3544
rect 17960 3392 18012 3398
rect 17960 3334 18012 3340
rect 17684 3120 17736 3126
rect 17684 3062 17736 3068
rect 17592 2984 17644 2990
rect 17592 2926 17644 2932
rect 17696 2514 17724 3062
rect 17972 2990 18000 3334
rect 18340 2990 18368 4422
rect 18510 4040 18566 4049
rect 18510 3975 18512 3984
rect 18564 3975 18566 3984
rect 18512 3946 18564 3952
rect 18512 3460 18564 3466
rect 18512 3402 18564 3408
rect 18524 3233 18552 3402
rect 18510 3224 18566 3233
rect 18510 3159 18566 3168
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 17868 2916 17920 2922
rect 17868 2858 17920 2864
rect 18144 2916 18196 2922
rect 18144 2858 18196 2864
rect 17774 2680 17830 2689
rect 17774 2615 17830 2624
rect 17788 2582 17816 2615
rect 17776 2576 17828 2582
rect 17776 2518 17828 2524
rect 17500 2508 17552 2514
rect 17500 2450 17552 2456
rect 17684 2508 17736 2514
rect 17684 2450 17736 2456
rect 16856 2372 16908 2378
rect 16856 2314 16908 2320
rect 17040 2372 17092 2378
rect 17040 2314 17092 2320
rect 17592 2372 17644 2378
rect 17592 2314 17644 2320
rect 16868 921 16896 2314
rect 17052 1329 17080 2314
rect 17038 1320 17094 1329
rect 17038 1255 17094 1264
rect 16684 870 16804 898
rect 16854 912 16910 921
rect 16684 800 16712 870
rect 16854 847 16910 856
rect 17604 800 17632 2314
rect 17880 1737 17908 2858
rect 18156 2825 18184 2858
rect 18420 2848 18472 2854
rect 18142 2816 18198 2825
rect 18420 2790 18472 2796
rect 18142 2751 18198 2760
rect 18432 2417 18460 2790
rect 19432 2440 19484 2446
rect 18418 2408 18474 2417
rect 19432 2382 19484 2388
rect 18418 2343 18474 2352
rect 18512 2372 18564 2378
rect 18512 2314 18564 2320
rect 18420 2304 18472 2310
rect 18420 2246 18472 2252
rect 17866 1728 17922 1737
rect 17866 1663 17922 1672
rect 18432 1170 18460 2246
rect 18524 2145 18552 2314
rect 18510 2136 18566 2145
rect 18510 2071 18566 2080
rect 18432 1142 18552 1170
rect 18524 800 18552 1142
rect 19444 800 19472 2382
rect 16486 504 16542 513
rect 16486 439 16542 448
rect 16670 0 16726 800
rect 17590 0 17646 800
rect 18510 0 18566 800
rect 19430 0 19486 800
<< via2 >>
rect 3054 16904 3110 16960
rect 1490 15952 1546 16008
rect 1858 15000 1914 15056
rect 2226 14612 2282 14648
rect 2226 14592 2228 14612
rect 2228 14592 2280 14612
rect 2280 14592 2282 14612
rect 1858 14320 1914 14376
rect 2134 13948 2136 13968
rect 2136 13948 2188 13968
rect 2188 13948 2190 13968
rect 2134 13912 2190 13948
rect 2778 13640 2834 13696
rect 3514 16632 3570 16688
rect 17314 16904 17370 16960
rect 16210 16496 16266 16552
rect 3882 16224 3938 16280
rect 4250 15544 4306 15600
rect 4158 15272 4214 15328
rect 3921 14170 3977 14172
rect 4001 14170 4057 14172
rect 4081 14170 4137 14172
rect 4161 14170 4217 14172
rect 3921 14118 3947 14170
rect 3947 14118 3977 14170
rect 4001 14118 4011 14170
rect 4011 14118 4057 14170
rect 4081 14118 4127 14170
rect 4127 14118 4137 14170
rect 4161 14118 4191 14170
rect 4191 14118 4217 14170
rect 3921 14116 3977 14118
rect 4001 14116 4057 14118
rect 4081 14116 4137 14118
rect 4161 14116 4217 14118
rect 1398 13232 1454 13288
rect 2226 12960 2282 13016
rect 1490 12688 1546 12744
rect 6886 14714 6942 14716
rect 6966 14714 7022 14716
rect 7046 14714 7102 14716
rect 7126 14714 7182 14716
rect 6886 14662 6912 14714
rect 6912 14662 6942 14714
rect 6966 14662 6976 14714
rect 6976 14662 7022 14714
rect 7046 14662 7092 14714
rect 7092 14662 7102 14714
rect 7126 14662 7156 14714
rect 7156 14662 7182 14714
rect 6886 14660 6942 14662
rect 6966 14660 7022 14662
rect 7046 14660 7102 14662
rect 7126 14660 7182 14662
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9878 14170
rect 9878 14118 9908 14170
rect 9932 14118 9942 14170
rect 9942 14118 9988 14170
rect 10012 14118 10058 14170
rect 10058 14118 10068 14170
rect 10092 14118 10122 14170
rect 10122 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 6886 13626 6942 13628
rect 6966 13626 7022 13628
rect 7046 13626 7102 13628
rect 7126 13626 7182 13628
rect 6886 13574 6912 13626
rect 6912 13574 6942 13626
rect 6966 13574 6976 13626
rect 6976 13574 7022 13626
rect 7046 13574 7092 13626
rect 7092 13574 7102 13626
rect 7126 13574 7156 13626
rect 7156 13574 7182 13626
rect 6886 13572 6942 13574
rect 6966 13572 7022 13574
rect 7046 13572 7102 13574
rect 7126 13572 7182 13574
rect 3921 13082 3977 13084
rect 4001 13082 4057 13084
rect 4081 13082 4137 13084
rect 4161 13082 4217 13084
rect 3921 13030 3947 13082
rect 3947 13030 3977 13082
rect 4001 13030 4011 13082
rect 4011 13030 4057 13082
rect 4081 13030 4127 13082
rect 4127 13030 4137 13082
rect 4161 13030 4191 13082
rect 4191 13030 4217 13082
rect 3921 13028 3977 13030
rect 4001 13028 4057 13030
rect 4081 13028 4137 13030
rect 4161 13028 4217 13030
rect 1398 12008 1454 12064
rect 1858 12280 1914 12336
rect 1490 11328 1546 11384
rect 1398 10920 1454 10976
rect 1490 9968 1546 10024
rect 1490 8336 1546 8392
rect 1490 8064 1546 8120
rect 1398 7656 1454 7712
rect 1398 7384 1454 7440
rect 1490 6704 1546 6760
rect 1766 11600 1822 11656
rect 1950 11192 2006 11248
rect 1858 10648 1914 10704
rect 1674 10376 1730 10432
rect 1950 9968 2006 10024
rect 1674 7384 1730 7440
rect 1674 5752 1730 5808
rect 1398 4664 1454 4720
rect 1582 4664 1638 4720
rect 1490 4120 1546 4176
rect 1490 3440 1546 3496
rect 2226 10240 2282 10296
rect 3054 9696 3110 9752
rect 3921 11994 3977 11996
rect 4001 11994 4057 11996
rect 4081 11994 4137 11996
rect 4161 11994 4217 11996
rect 3921 11942 3947 11994
rect 3947 11942 3977 11994
rect 4001 11942 4011 11994
rect 4011 11942 4057 11994
rect 4081 11942 4127 11994
rect 4127 11942 4137 11994
rect 4161 11942 4191 11994
rect 4191 11942 4217 11994
rect 3921 11940 3977 11942
rect 4001 11940 4057 11942
rect 4081 11940 4137 11942
rect 4161 11940 4217 11942
rect 3974 11636 3976 11656
rect 3976 11636 4028 11656
rect 4028 11636 4030 11656
rect 3974 11600 4030 11636
rect 2042 5208 2098 5264
rect 3330 8744 3386 8800
rect 3238 8472 3294 8528
rect 2410 6160 2466 6216
rect 2318 5752 2374 5808
rect 2410 5344 2466 5400
rect 1858 3712 1914 3768
rect 2134 4392 2190 4448
rect 2870 6976 2926 7032
rect 2778 6332 2780 6352
rect 2780 6332 2832 6352
rect 2832 6332 2834 6352
rect 2778 6296 2834 6332
rect 2962 5888 3018 5944
rect 2686 5636 2742 5672
rect 2686 5616 2688 5636
rect 2688 5616 2740 5636
rect 2740 5616 2742 5636
rect 3054 5752 3110 5808
rect 2870 5516 2872 5536
rect 2872 5516 2924 5536
rect 2924 5516 2926 5536
rect 2870 5480 2926 5516
rect 2594 4528 2650 4584
rect 2594 3984 2650 4040
rect 3921 10906 3977 10908
rect 4001 10906 4057 10908
rect 4081 10906 4137 10908
rect 4161 10906 4217 10908
rect 3921 10854 3947 10906
rect 3947 10854 3977 10906
rect 4001 10854 4011 10906
rect 4011 10854 4057 10906
rect 4081 10854 4127 10906
rect 4127 10854 4137 10906
rect 4161 10854 4191 10906
rect 4191 10854 4217 10906
rect 3921 10852 3977 10854
rect 4001 10852 4057 10854
rect 4081 10852 4137 10854
rect 4161 10852 4217 10854
rect 3921 9818 3977 9820
rect 4001 9818 4057 9820
rect 4081 9818 4137 9820
rect 4161 9818 4217 9820
rect 3921 9766 3947 9818
rect 3947 9766 3977 9818
rect 4001 9766 4011 9818
rect 4011 9766 4057 9818
rect 4081 9766 4127 9818
rect 4127 9766 4137 9818
rect 4161 9766 4191 9818
rect 4191 9766 4217 9818
rect 3921 9764 3977 9766
rect 4001 9764 4057 9766
rect 4081 9764 4137 9766
rect 4161 9764 4217 9766
rect 4434 9968 4490 10024
rect 3790 9288 3846 9344
rect 4066 9288 4122 9344
rect 3882 9016 3938 9072
rect 4802 12044 4804 12064
rect 4804 12044 4856 12064
rect 4856 12044 4858 12064
rect 4802 12008 4858 12044
rect 5170 11872 5226 11928
rect 4710 10104 4766 10160
rect 4802 9968 4858 10024
rect 4894 9716 4950 9752
rect 4894 9696 4896 9716
rect 4896 9696 4948 9716
rect 4948 9696 4950 9716
rect 4710 9424 4766 9480
rect 4434 9016 4490 9072
rect 4158 8880 4214 8936
rect 3422 7384 3478 7440
rect 3422 5888 3478 5944
rect 3921 8730 3977 8732
rect 4001 8730 4057 8732
rect 4081 8730 4137 8732
rect 4161 8730 4217 8732
rect 3921 8678 3947 8730
rect 3947 8678 3977 8730
rect 4001 8678 4011 8730
rect 4011 8678 4057 8730
rect 4081 8678 4127 8730
rect 4127 8678 4137 8730
rect 4161 8678 4191 8730
rect 4191 8678 4217 8730
rect 3921 8676 3977 8678
rect 4001 8676 4057 8678
rect 4081 8676 4137 8678
rect 4161 8676 4217 8678
rect 3974 8200 4030 8256
rect 3606 6432 3662 6488
rect 3422 5480 3478 5536
rect 3921 7642 3977 7644
rect 4001 7642 4057 7644
rect 4081 7642 4137 7644
rect 4161 7642 4217 7644
rect 3921 7590 3947 7642
rect 3947 7590 3977 7642
rect 4001 7590 4011 7642
rect 4011 7590 4057 7642
rect 4081 7590 4127 7642
rect 4127 7590 4137 7642
rect 4161 7590 4191 7642
rect 4191 7590 4217 7642
rect 3921 7588 3977 7590
rect 4001 7588 4057 7590
rect 4081 7588 4137 7590
rect 4161 7588 4217 7590
rect 4434 8200 4490 8256
rect 3921 6554 3977 6556
rect 4001 6554 4057 6556
rect 4081 6554 4137 6556
rect 4161 6554 4217 6556
rect 3921 6502 3947 6554
rect 3947 6502 3977 6554
rect 4001 6502 4011 6554
rect 4011 6502 4057 6554
rect 4081 6502 4127 6554
rect 4127 6502 4137 6554
rect 4161 6502 4191 6554
rect 4191 6502 4217 6554
rect 3921 6500 3977 6502
rect 4001 6500 4057 6502
rect 4081 6500 4137 6502
rect 4161 6500 4217 6502
rect 4342 6432 4398 6488
rect 3790 6024 3846 6080
rect 4250 5636 4306 5672
rect 4250 5616 4252 5636
rect 4252 5616 4304 5636
rect 4304 5616 4306 5636
rect 3921 5466 3977 5468
rect 4001 5466 4057 5468
rect 4081 5466 4137 5468
rect 4161 5466 4217 5468
rect 3921 5414 3947 5466
rect 3947 5414 3977 5466
rect 4001 5414 4011 5466
rect 4011 5414 4057 5466
rect 4081 5414 4127 5466
rect 4127 5414 4137 5466
rect 4161 5414 4191 5466
rect 4191 5414 4217 5466
rect 3921 5412 3977 5414
rect 4001 5412 4057 5414
rect 4081 5412 4137 5414
rect 4161 5412 4217 5414
rect 3882 5108 3884 5128
rect 3884 5108 3936 5128
rect 3936 5108 3938 5128
rect 3882 5072 3938 5108
rect 3054 4120 3110 4176
rect 2962 3848 3018 3904
rect 2318 2932 2320 2952
rect 2320 2932 2372 2952
rect 2372 2932 2374 2952
rect 2318 2896 2374 2932
rect 2686 2624 2742 2680
rect 3422 3032 3478 3088
rect 2962 1128 3018 1184
rect 3921 4378 3977 4380
rect 4001 4378 4057 4380
rect 4081 4378 4137 4380
rect 4161 4378 4217 4380
rect 3921 4326 3947 4378
rect 3947 4326 3977 4378
rect 4001 4326 4011 4378
rect 4011 4326 4057 4378
rect 4081 4326 4127 4378
rect 4127 4326 4137 4378
rect 4161 4326 4191 4378
rect 4191 4326 4217 4378
rect 3921 4324 3977 4326
rect 4001 4324 4057 4326
rect 4081 4324 4137 4326
rect 4161 4324 4217 4326
rect 4158 3848 4214 3904
rect 3698 3440 3754 3496
rect 3921 3290 3977 3292
rect 4001 3290 4057 3292
rect 4081 3290 4137 3292
rect 4161 3290 4217 3292
rect 3921 3238 3947 3290
rect 3947 3238 3977 3290
rect 4001 3238 4011 3290
rect 4011 3238 4057 3290
rect 4081 3238 4127 3290
rect 4127 3238 4137 3290
rect 4161 3238 4191 3290
rect 4191 3238 4217 3290
rect 3921 3236 3977 3238
rect 4001 3236 4057 3238
rect 4081 3236 4137 3238
rect 4161 3236 4217 3238
rect 3330 2080 3386 2136
rect 3238 1808 3294 1864
rect 3146 1400 3202 1456
rect 2870 448 2926 504
rect 2778 176 2834 232
rect 3790 2760 3846 2816
rect 4894 7928 4950 7984
rect 4894 7384 4950 7440
rect 5078 10260 5134 10296
rect 5078 10240 5080 10260
rect 5080 10240 5132 10260
rect 5132 10240 5134 10260
rect 5078 9288 5134 9344
rect 5354 11872 5410 11928
rect 5354 10104 5410 10160
rect 5170 8200 5226 8256
rect 5722 10512 5778 10568
rect 6886 12538 6942 12540
rect 6966 12538 7022 12540
rect 7046 12538 7102 12540
rect 7126 12538 7182 12540
rect 6886 12486 6912 12538
rect 6912 12486 6942 12538
rect 6966 12486 6976 12538
rect 6976 12486 7022 12538
rect 7046 12486 7092 12538
rect 7092 12486 7102 12538
rect 7126 12486 7156 12538
rect 7156 12486 7182 12538
rect 6886 12484 6942 12486
rect 6966 12484 7022 12486
rect 7046 12484 7102 12486
rect 7126 12484 7182 12486
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9878 13082
rect 9878 13030 9908 13082
rect 9932 13030 9942 13082
rect 9942 13030 9988 13082
rect 10012 13030 10058 13082
rect 10058 13030 10068 13082
rect 10092 13030 10122 13082
rect 10122 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 5906 12280 5962 12336
rect 6182 11736 6238 11792
rect 6090 10920 6146 10976
rect 6274 11056 6330 11112
rect 5906 10648 5962 10704
rect 5538 9696 5594 9752
rect 5630 9580 5686 9616
rect 5630 9560 5632 9580
rect 5632 9560 5684 9580
rect 5684 9560 5686 9580
rect 5538 9016 5594 9072
rect 4618 3984 4674 4040
rect 4618 3884 4620 3904
rect 4620 3884 4672 3904
rect 4672 3884 4674 3904
rect 4618 3848 4674 3884
rect 5262 7928 5318 7984
rect 5354 6160 5410 6216
rect 5814 7928 5870 7984
rect 6090 10140 6092 10160
rect 6092 10140 6144 10160
rect 6144 10140 6146 10160
rect 6090 10104 6146 10140
rect 6182 9696 6238 9752
rect 5722 6432 5778 6488
rect 6550 12144 6606 12200
rect 7838 12180 7840 12200
rect 7840 12180 7892 12200
rect 7892 12180 7894 12200
rect 7838 12144 7894 12180
rect 6642 10240 6698 10296
rect 5354 4664 5410 4720
rect 5262 4392 5318 4448
rect 5170 3440 5226 3496
rect 3698 2352 3754 2408
rect 3921 2202 3977 2204
rect 4001 2202 4057 2204
rect 4081 2202 4137 2204
rect 4161 2202 4217 2204
rect 3921 2150 3947 2202
rect 3947 2150 3977 2202
rect 4001 2150 4011 2202
rect 4011 2150 4057 2202
rect 4081 2150 4127 2202
rect 4127 2150 4137 2202
rect 4161 2150 4191 2202
rect 4191 2150 4217 2202
rect 3921 2148 3977 2150
rect 4001 2148 4057 2150
rect 4081 2148 4137 2150
rect 4161 2148 4217 2150
rect 5998 4528 6054 4584
rect 5814 4392 5870 4448
rect 5630 3032 5686 3088
rect 6458 5108 6460 5128
rect 6460 5108 6512 5128
rect 6512 5108 6514 5128
rect 6458 5072 6514 5108
rect 6366 4528 6422 4584
rect 6886 11450 6942 11452
rect 6966 11450 7022 11452
rect 7046 11450 7102 11452
rect 7126 11450 7182 11452
rect 6886 11398 6912 11450
rect 6912 11398 6942 11450
rect 6966 11398 6976 11450
rect 6976 11398 7022 11450
rect 7046 11398 7092 11450
rect 7092 11398 7102 11450
rect 7126 11398 7156 11450
rect 7156 11398 7182 11450
rect 6886 11396 6942 11398
rect 6966 11396 7022 11398
rect 7046 11396 7102 11398
rect 7126 11396 7182 11398
rect 7378 11328 7434 11384
rect 6886 10362 6942 10364
rect 6966 10362 7022 10364
rect 7046 10362 7102 10364
rect 7126 10362 7182 10364
rect 6886 10310 6912 10362
rect 6912 10310 6942 10362
rect 6966 10310 6976 10362
rect 6976 10310 7022 10362
rect 7046 10310 7092 10362
rect 7092 10310 7102 10362
rect 7126 10310 7156 10362
rect 7156 10310 7182 10362
rect 6886 10308 6942 10310
rect 6966 10308 7022 10310
rect 7046 10308 7102 10310
rect 7126 10308 7182 10310
rect 6826 10104 6882 10160
rect 6918 10004 6920 10024
rect 6920 10004 6972 10024
rect 6972 10004 6974 10024
rect 6918 9968 6974 10004
rect 7286 9968 7342 10024
rect 7470 9580 7526 9616
rect 7470 9560 7472 9580
rect 7472 9560 7524 9580
rect 7524 9560 7526 9580
rect 6886 9274 6942 9276
rect 6966 9274 7022 9276
rect 7046 9274 7102 9276
rect 7126 9274 7182 9276
rect 6886 9222 6912 9274
rect 6912 9222 6942 9274
rect 6966 9222 6976 9274
rect 6976 9222 7022 9274
rect 7046 9222 7092 9274
rect 7092 9222 7102 9274
rect 7126 9222 7156 9274
rect 7156 9222 7182 9274
rect 6886 9220 6942 9222
rect 6966 9220 7022 9222
rect 7046 9220 7102 9222
rect 7126 9220 7182 9222
rect 7286 8472 7342 8528
rect 6886 8186 6942 8188
rect 6966 8186 7022 8188
rect 7046 8186 7102 8188
rect 7126 8186 7182 8188
rect 6886 8134 6912 8186
rect 6912 8134 6942 8186
rect 6966 8134 6976 8186
rect 6976 8134 7022 8186
rect 7046 8134 7092 8186
rect 7092 8134 7102 8186
rect 7126 8134 7156 8186
rect 7156 8134 7182 8186
rect 6886 8132 6942 8134
rect 6966 8132 7022 8134
rect 7046 8132 7102 8134
rect 7126 8132 7182 8134
rect 6886 7098 6942 7100
rect 6966 7098 7022 7100
rect 7046 7098 7102 7100
rect 7126 7098 7182 7100
rect 6886 7046 6912 7098
rect 6912 7046 6942 7098
rect 6966 7046 6976 7098
rect 6976 7046 7022 7098
rect 7046 7046 7092 7098
rect 7092 7046 7102 7098
rect 7126 7046 7156 7098
rect 7156 7046 7182 7098
rect 6886 7044 6942 7046
rect 6966 7044 7022 7046
rect 7046 7044 7102 7046
rect 7126 7044 7182 7046
rect 6886 6010 6942 6012
rect 6966 6010 7022 6012
rect 7046 6010 7102 6012
rect 7126 6010 7182 6012
rect 6886 5958 6912 6010
rect 6912 5958 6942 6010
rect 6966 5958 6976 6010
rect 6976 5958 7022 6010
rect 7046 5958 7092 6010
rect 7092 5958 7102 6010
rect 7126 5958 7156 6010
rect 7156 5958 7182 6010
rect 6886 5956 6942 5958
rect 6966 5956 7022 5958
rect 7046 5956 7102 5958
rect 7126 5956 7182 5958
rect 7102 5208 7158 5264
rect 7562 8880 7618 8936
rect 7470 5616 7526 5672
rect 6734 5072 6790 5128
rect 6274 4392 6330 4448
rect 6090 2896 6146 2952
rect 6550 4428 6552 4448
rect 6552 4428 6604 4448
rect 6604 4428 6606 4448
rect 6550 4392 6606 4428
rect 6886 4922 6942 4924
rect 6966 4922 7022 4924
rect 7046 4922 7102 4924
rect 7126 4922 7182 4924
rect 6886 4870 6912 4922
rect 6912 4870 6942 4922
rect 6966 4870 6976 4922
rect 6976 4870 7022 4922
rect 7046 4870 7092 4922
rect 7092 4870 7102 4922
rect 7126 4870 7156 4922
rect 7156 4870 7182 4922
rect 6886 4868 6942 4870
rect 6966 4868 7022 4870
rect 7046 4868 7102 4870
rect 7126 4868 7182 4870
rect 8114 12144 8170 12200
rect 8022 10104 8078 10160
rect 8206 11464 8262 11520
rect 8206 9968 8262 10024
rect 8758 11464 8814 11520
rect 8758 10412 8760 10432
rect 8760 10412 8812 10432
rect 8812 10412 8814 10432
rect 8758 10376 8814 10412
rect 9218 11872 9274 11928
rect 9126 10920 9182 10976
rect 9034 10104 9090 10160
rect 8482 9968 8538 10024
rect 8206 9560 8262 9616
rect 8574 9832 8630 9888
rect 8206 8880 8262 8936
rect 8482 8880 8538 8936
rect 8298 7928 8354 7984
rect 8850 7964 8852 7984
rect 8852 7964 8904 7984
rect 8904 7964 8906 7984
rect 8850 7928 8906 7964
rect 9126 9968 9182 10024
rect 9494 9968 9550 10024
rect 9034 7248 9090 7304
rect 8666 6296 8722 6352
rect 8022 5208 8078 5264
rect 8022 5108 8024 5128
rect 8024 5108 8076 5128
rect 8076 5108 8078 5128
rect 8022 5072 8078 5108
rect 6734 4156 6736 4176
rect 6736 4156 6788 4176
rect 6788 4156 6790 4176
rect 6734 4120 6790 4156
rect 7654 4120 7710 4176
rect 6458 2624 6514 2680
rect 6886 3834 6942 3836
rect 6966 3834 7022 3836
rect 7046 3834 7102 3836
rect 7126 3834 7182 3836
rect 6886 3782 6912 3834
rect 6912 3782 6942 3834
rect 6966 3782 6976 3834
rect 6976 3782 7022 3834
rect 7046 3782 7092 3834
rect 7092 3782 7102 3834
rect 7126 3782 7156 3834
rect 7156 3782 7182 3834
rect 6886 3780 6942 3782
rect 6966 3780 7022 3782
rect 7046 3780 7102 3782
rect 7126 3780 7182 3782
rect 8114 3576 8170 3632
rect 6734 2932 6736 2952
rect 6736 2932 6788 2952
rect 6788 2932 6790 2952
rect 6734 2896 6790 2932
rect 6886 2746 6942 2748
rect 6966 2746 7022 2748
rect 7046 2746 7102 2748
rect 7126 2746 7182 2748
rect 6886 2694 6912 2746
rect 6912 2694 6942 2746
rect 6966 2694 6976 2746
rect 6976 2694 7022 2746
rect 7046 2694 7092 2746
rect 7092 2694 7102 2746
rect 7126 2694 7156 2746
rect 7156 2694 7182 2746
rect 6886 2692 6942 2694
rect 6966 2692 7022 2694
rect 7046 2692 7102 2694
rect 7126 2692 7182 2694
rect 8298 2508 8354 2544
rect 8298 2488 8300 2508
rect 8300 2488 8352 2508
rect 8352 2488 8354 2508
rect 8574 4684 8630 4720
rect 8574 4664 8576 4684
rect 8576 4664 8628 4684
rect 8628 4664 8630 4684
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9878 11994
rect 9878 11942 9908 11994
rect 9932 11942 9942 11994
rect 9942 11942 9988 11994
rect 10012 11942 10058 11994
rect 10058 11942 10068 11994
rect 10092 11942 10122 11994
rect 10122 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 10598 12280 10654 12336
rect 9954 11464 10010 11520
rect 9862 11192 9918 11248
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9878 10906
rect 9878 10854 9908 10906
rect 9932 10854 9942 10906
rect 9942 10854 9988 10906
rect 10012 10854 10058 10906
rect 10058 10854 10068 10906
rect 10092 10854 10122 10906
rect 10122 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 9862 10532 9918 10568
rect 9862 10512 9864 10532
rect 9864 10512 9916 10532
rect 9916 10512 9918 10532
rect 10046 10240 10102 10296
rect 10506 11736 10562 11792
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9878 9818
rect 9878 9766 9908 9818
rect 9932 9766 9942 9818
rect 9942 9766 9988 9818
rect 10012 9766 10058 9818
rect 10058 9766 10068 9818
rect 10092 9766 10122 9818
rect 10122 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 9218 4428 9220 4448
rect 9220 4428 9272 4448
rect 9272 4428 9274 4448
rect 9218 4392 9274 4428
rect 8850 2796 8852 2816
rect 8852 2796 8904 2816
rect 8904 2796 8906 2816
rect 8850 2760 8906 2796
rect 9218 3596 9274 3632
rect 9218 3576 9220 3596
rect 9220 3576 9272 3596
rect 9272 3576 9274 3596
rect 9402 4684 9458 4720
rect 9402 4664 9404 4684
rect 9404 4664 9456 4684
rect 9456 4664 9458 4684
rect 10414 10512 10470 10568
rect 10506 10240 10562 10296
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9878 8730
rect 9878 8678 9908 8730
rect 9932 8678 9942 8730
rect 9942 8678 9988 8730
rect 10012 8678 10058 8730
rect 10058 8678 10068 8730
rect 10092 8678 10122 8730
rect 10122 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 10506 9016 10562 9072
rect 9862 7828 9864 7848
rect 9864 7828 9916 7848
rect 9916 7828 9918 7848
rect 9862 7792 9918 7828
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9878 7642
rect 9878 7590 9908 7642
rect 9932 7590 9942 7642
rect 9942 7590 9988 7642
rect 10012 7590 10058 7642
rect 10058 7590 10068 7642
rect 10092 7590 10122 7642
rect 10122 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9878 6554
rect 9878 6502 9908 6554
rect 9932 6502 9942 6554
rect 9942 6502 9988 6554
rect 10012 6502 10058 6554
rect 10058 6502 10068 6554
rect 10092 6502 10122 6554
rect 10122 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9878 5466
rect 9878 5414 9908 5466
rect 9932 5414 9942 5466
rect 9942 5414 9988 5466
rect 10012 5414 10058 5466
rect 10058 5414 10068 5466
rect 10092 5414 10122 5466
rect 10122 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 10690 9580 10746 9616
rect 10690 9560 10692 9580
rect 10692 9560 10744 9580
rect 10744 9560 10746 9580
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9878 4378
rect 9878 4326 9908 4378
rect 9932 4326 9942 4378
rect 9942 4326 9988 4378
rect 10012 4326 10058 4378
rect 10058 4326 10068 4378
rect 10092 4326 10122 4378
rect 10122 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 10322 4392 10378 4448
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9878 3290
rect 9878 3238 9908 3290
rect 9932 3238 9942 3290
rect 9942 3238 9988 3290
rect 10012 3238 10058 3290
rect 10058 3238 10068 3290
rect 10092 3238 10122 3290
rect 10122 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 9954 2624 10010 2680
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9878 2202
rect 9878 2150 9908 2202
rect 9932 2150 9942 2202
rect 9942 2150 9988 2202
rect 10012 2150 10058 2202
rect 10058 2150 10068 2202
rect 10092 2150 10122 2202
rect 10122 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 10690 6568 10746 6624
rect 10690 6316 10746 6352
rect 10690 6296 10692 6316
rect 10692 6296 10744 6316
rect 10744 6296 10746 6316
rect 10598 2508 10654 2544
rect 10598 2488 10600 2508
rect 10600 2488 10652 2508
rect 10652 2488 10654 2508
rect 11058 11056 11114 11112
rect 10966 7928 11022 7984
rect 12817 14714 12873 14716
rect 12897 14714 12953 14716
rect 12977 14714 13033 14716
rect 13057 14714 13113 14716
rect 12817 14662 12843 14714
rect 12843 14662 12873 14714
rect 12897 14662 12907 14714
rect 12907 14662 12953 14714
rect 12977 14662 13023 14714
rect 13023 14662 13033 14714
rect 13057 14662 13087 14714
rect 13087 14662 13113 14714
rect 12817 14660 12873 14662
rect 12897 14660 12953 14662
rect 12977 14660 13033 14662
rect 13057 14660 13113 14662
rect 12817 13626 12873 13628
rect 12897 13626 12953 13628
rect 12977 13626 13033 13628
rect 13057 13626 13113 13628
rect 12817 13574 12843 13626
rect 12843 13574 12873 13626
rect 12897 13574 12907 13626
rect 12907 13574 12953 13626
rect 12977 13574 13023 13626
rect 13023 13574 13033 13626
rect 13057 13574 13087 13626
rect 13087 13574 13113 13626
rect 12817 13572 12873 13574
rect 12897 13572 12953 13574
rect 12977 13572 13033 13574
rect 13057 13572 13113 13574
rect 11886 12144 11942 12200
rect 11150 9424 11206 9480
rect 11150 8880 11206 8936
rect 11794 9580 11850 9616
rect 11794 9560 11796 9580
rect 11796 9560 11848 9580
rect 11848 9560 11850 9580
rect 11794 9424 11850 9480
rect 12817 12538 12873 12540
rect 12897 12538 12953 12540
rect 12977 12538 13033 12540
rect 13057 12538 13113 12540
rect 12817 12486 12843 12538
rect 12843 12486 12873 12538
rect 12897 12486 12907 12538
rect 12907 12486 12953 12538
rect 12977 12486 13023 12538
rect 13023 12486 13033 12538
rect 13057 12486 13087 12538
rect 13087 12486 13113 12538
rect 12817 12484 12873 12486
rect 12897 12484 12953 12486
rect 12977 12484 13033 12486
rect 13057 12484 13113 12486
rect 12622 11464 12678 11520
rect 12346 11192 12402 11248
rect 12254 11056 12310 11112
rect 12817 11450 12873 11452
rect 12897 11450 12953 11452
rect 12977 11450 13033 11452
rect 13057 11450 13113 11452
rect 12817 11398 12843 11450
rect 12843 11398 12873 11450
rect 12897 11398 12907 11450
rect 12907 11398 12953 11450
rect 12977 11398 13023 11450
rect 13023 11398 13033 11450
rect 13057 11398 13087 11450
rect 13087 11398 13113 11450
rect 12817 11396 12873 11398
rect 12897 11396 12953 11398
rect 12977 11396 13033 11398
rect 13057 11396 13113 11398
rect 13726 11328 13782 11384
rect 13174 10784 13230 10840
rect 13266 10648 13322 10704
rect 13174 10512 13230 10568
rect 12817 10362 12873 10364
rect 12897 10362 12953 10364
rect 12977 10362 13033 10364
rect 13057 10362 13113 10364
rect 12817 10310 12843 10362
rect 12843 10310 12873 10362
rect 12897 10310 12907 10362
rect 12907 10310 12953 10362
rect 12977 10310 13023 10362
rect 13023 10310 13033 10362
rect 13057 10310 13087 10362
rect 13087 10310 13113 10362
rect 12817 10308 12873 10310
rect 12897 10308 12953 10310
rect 12977 10308 13033 10310
rect 13057 10308 13113 10310
rect 12254 9696 12310 9752
rect 11886 8356 11942 8392
rect 11886 8336 11888 8356
rect 11888 8336 11940 8356
rect 11940 8336 11942 8356
rect 13174 9424 13230 9480
rect 12817 9274 12873 9276
rect 12897 9274 12953 9276
rect 12977 9274 13033 9276
rect 13057 9274 13113 9276
rect 12817 9222 12843 9274
rect 12843 9222 12873 9274
rect 12897 9222 12907 9274
rect 12907 9222 12953 9274
rect 12977 9222 13023 9274
rect 13023 9222 13033 9274
rect 13057 9222 13087 9274
rect 13087 9222 13113 9274
rect 12817 9220 12873 9222
rect 12897 9220 12953 9222
rect 12977 9220 13033 9222
rect 13057 9220 13113 9222
rect 13450 9560 13506 9616
rect 13266 9152 13322 9208
rect 13358 9036 13414 9072
rect 13358 9016 13360 9036
rect 13360 9016 13412 9036
rect 13412 9016 13414 9036
rect 11334 6296 11390 6352
rect 11242 6160 11298 6216
rect 10874 3984 10930 4040
rect 10966 3476 10968 3496
rect 10968 3476 11020 3496
rect 11020 3476 11022 3496
rect 10966 3440 11022 3476
rect 11702 4120 11758 4176
rect 11978 5208 12034 5264
rect 11886 3032 11942 3088
rect 12817 8186 12873 8188
rect 12897 8186 12953 8188
rect 12977 8186 13033 8188
rect 13057 8186 13113 8188
rect 12817 8134 12843 8186
rect 12843 8134 12873 8186
rect 12897 8134 12907 8186
rect 12907 8134 12953 8186
rect 12977 8134 13023 8186
rect 13023 8134 13033 8186
rect 13057 8134 13087 8186
rect 13087 8134 13113 8186
rect 12817 8132 12873 8134
rect 12897 8132 12953 8134
rect 12977 8132 13033 8134
rect 13057 8132 13113 8134
rect 12817 7098 12873 7100
rect 12897 7098 12953 7100
rect 12977 7098 13033 7100
rect 13057 7098 13113 7100
rect 12817 7046 12843 7098
rect 12843 7046 12873 7098
rect 12897 7046 12907 7098
rect 12907 7046 12953 7098
rect 12977 7046 13023 7098
rect 13023 7046 13033 7098
rect 13057 7046 13087 7098
rect 13087 7046 13113 7098
rect 12817 7044 12873 7046
rect 12897 7044 12953 7046
rect 12977 7044 13033 7046
rect 13057 7044 13113 7046
rect 12806 6296 12862 6352
rect 12530 4392 12586 4448
rect 12346 4120 12402 4176
rect 12817 6010 12873 6012
rect 12897 6010 12953 6012
rect 12977 6010 13033 6012
rect 13057 6010 13113 6012
rect 12817 5958 12843 6010
rect 12843 5958 12873 6010
rect 12897 5958 12907 6010
rect 12907 5958 12953 6010
rect 12977 5958 13023 6010
rect 13023 5958 13033 6010
rect 13057 5958 13087 6010
rect 13087 5958 13113 6010
rect 12817 5956 12873 5958
rect 12897 5956 12953 5958
rect 12977 5956 13033 5958
rect 13057 5956 13113 5958
rect 13174 5072 13230 5128
rect 14094 11872 14150 11928
rect 13542 6704 13598 6760
rect 13818 7948 13874 7984
rect 13818 7928 13820 7948
rect 13820 7928 13872 7948
rect 13872 7928 13874 7948
rect 14278 8200 14334 8256
rect 14002 6976 14058 7032
rect 14002 6568 14058 6624
rect 13634 6196 13636 6216
rect 13636 6196 13688 6216
rect 13688 6196 13690 6216
rect 13450 6060 13452 6080
rect 13452 6060 13504 6080
rect 13504 6060 13506 6080
rect 13450 6024 13506 6060
rect 12817 4922 12873 4924
rect 12897 4922 12953 4924
rect 12977 4922 13033 4924
rect 13057 4922 13113 4924
rect 12817 4870 12843 4922
rect 12843 4870 12873 4922
rect 12897 4870 12907 4922
rect 12907 4870 12953 4922
rect 12977 4870 13023 4922
rect 13023 4870 13033 4922
rect 13057 4870 13087 4922
rect 13087 4870 13113 4922
rect 12817 4868 12873 4870
rect 12897 4868 12953 4870
rect 12977 4868 13033 4870
rect 13057 4868 13113 4870
rect 13082 4664 13138 4720
rect 12817 3834 12873 3836
rect 12897 3834 12953 3836
rect 12977 3834 13033 3836
rect 13057 3834 13113 3836
rect 12817 3782 12843 3834
rect 12843 3782 12873 3834
rect 12897 3782 12907 3834
rect 12907 3782 12953 3834
rect 12977 3782 13023 3834
rect 13023 3782 13033 3834
rect 13057 3782 13087 3834
rect 13087 3782 13113 3834
rect 12817 3780 12873 3782
rect 12897 3780 12953 3782
rect 12977 3780 13033 3782
rect 13057 3780 13113 3782
rect 12438 3476 12440 3496
rect 12440 3476 12492 3496
rect 12492 3476 12494 3496
rect 12438 3440 12494 3476
rect 13634 6160 13690 6196
rect 13634 6024 13690 6080
rect 12346 2760 12402 2816
rect 12817 2746 12873 2748
rect 12897 2746 12953 2748
rect 12977 2746 13033 2748
rect 13057 2746 13113 2748
rect 12817 2694 12843 2746
rect 12843 2694 12873 2746
rect 12897 2694 12907 2746
rect 12907 2694 12953 2746
rect 12977 2694 13023 2746
rect 13023 2694 13033 2746
rect 13057 2694 13087 2746
rect 13087 2694 13113 2746
rect 12817 2692 12873 2694
rect 12897 2692 12953 2694
rect 12977 2692 13033 2694
rect 13057 2692 13113 2694
rect 14002 2760 14058 2816
rect 14370 4548 14426 4584
rect 14370 4528 14372 4548
rect 14372 4528 14424 4548
rect 14424 4528 14426 4548
rect 14370 4120 14426 4176
rect 14554 8336 14610 8392
rect 15782 14170 15838 14172
rect 15862 14170 15918 14172
rect 15942 14170 15998 14172
rect 16022 14170 16078 14172
rect 15782 14118 15808 14170
rect 15808 14118 15838 14170
rect 15862 14118 15872 14170
rect 15872 14118 15918 14170
rect 15942 14118 15988 14170
rect 15988 14118 15998 14170
rect 16022 14118 16052 14170
rect 16052 14118 16078 14170
rect 15782 14116 15838 14118
rect 15862 14116 15918 14118
rect 15942 14116 15998 14118
rect 16022 14116 16078 14118
rect 16486 15680 16542 15736
rect 16946 15408 17002 15464
rect 15782 13082 15838 13084
rect 15862 13082 15918 13084
rect 15942 13082 15998 13084
rect 16022 13082 16078 13084
rect 15782 13030 15808 13082
rect 15808 13030 15838 13082
rect 15862 13030 15872 13082
rect 15872 13030 15918 13082
rect 15942 13030 15988 13082
rect 15988 13030 15998 13082
rect 16022 13030 16052 13082
rect 16052 13030 16078 13082
rect 15782 13028 15838 13030
rect 15862 13028 15918 13030
rect 15942 13028 15998 13030
rect 16022 13028 16078 13030
rect 16394 13524 16450 13560
rect 16394 13504 16396 13524
rect 16396 13504 16448 13524
rect 16448 13504 16450 13524
rect 15106 10784 15162 10840
rect 14554 7928 14610 7984
rect 14554 4820 14610 4856
rect 14554 4800 14556 4820
rect 14556 4800 14608 4820
rect 14608 4800 14610 4820
rect 14738 7112 14794 7168
rect 14554 3984 14610 4040
rect 14370 2896 14426 2952
rect 14462 2760 14518 2816
rect 15474 11872 15530 11928
rect 15474 9696 15530 9752
rect 14922 6160 14978 6216
rect 15290 8492 15346 8528
rect 15290 8472 15292 8492
rect 15292 8472 15344 8492
rect 15344 8472 15346 8492
rect 15474 9016 15530 9072
rect 15474 7928 15530 7984
rect 15198 5616 15254 5672
rect 15782 11994 15838 11996
rect 15862 11994 15918 11996
rect 15942 11994 15998 11996
rect 16022 11994 16078 11996
rect 15782 11942 15808 11994
rect 15808 11942 15838 11994
rect 15862 11942 15872 11994
rect 15872 11942 15918 11994
rect 15942 11942 15988 11994
rect 15988 11942 15998 11994
rect 16022 11942 16052 11994
rect 16052 11942 16078 11994
rect 15782 11940 15838 11942
rect 15862 11940 15918 11942
rect 15942 11940 15998 11942
rect 16022 11940 16078 11942
rect 15782 10906 15838 10908
rect 15862 10906 15918 10908
rect 15942 10906 15998 10908
rect 16022 10906 16078 10908
rect 15782 10854 15808 10906
rect 15808 10854 15838 10906
rect 15862 10854 15872 10906
rect 15872 10854 15918 10906
rect 15942 10854 15988 10906
rect 15988 10854 15998 10906
rect 16022 10854 16052 10906
rect 16052 10854 16078 10906
rect 15782 10852 15838 10854
rect 15862 10852 15918 10854
rect 15942 10852 15998 10854
rect 16022 10852 16078 10854
rect 15750 9968 15806 10024
rect 15782 9818 15838 9820
rect 15862 9818 15918 9820
rect 15942 9818 15998 9820
rect 16022 9818 16078 9820
rect 15782 9766 15808 9818
rect 15808 9766 15838 9818
rect 15862 9766 15872 9818
rect 15872 9766 15918 9818
rect 15942 9766 15988 9818
rect 15988 9766 15998 9818
rect 16022 9766 16052 9818
rect 16052 9766 16078 9818
rect 15782 9764 15838 9766
rect 15862 9764 15918 9766
rect 15942 9764 15998 9766
rect 16022 9764 16078 9766
rect 16026 9632 16082 9688
rect 15750 8880 15806 8936
rect 16026 9016 16082 9072
rect 15782 8730 15838 8732
rect 15862 8730 15918 8732
rect 15942 8730 15998 8732
rect 16022 8730 16078 8732
rect 15782 8678 15808 8730
rect 15808 8678 15838 8730
rect 15862 8678 15872 8730
rect 15872 8678 15918 8730
rect 15942 8678 15988 8730
rect 15988 8678 15998 8730
rect 16022 8678 16052 8730
rect 16052 8678 16078 8730
rect 15782 8676 15838 8678
rect 15862 8676 15918 8678
rect 15942 8676 15998 8678
rect 16022 8676 16078 8678
rect 16394 11500 16396 11520
rect 16396 11500 16448 11520
rect 16448 11500 16450 11520
rect 16394 11464 16450 11500
rect 16578 11872 16634 11928
rect 17038 12688 17094 12744
rect 16854 11328 16910 11384
rect 16486 9832 16542 9888
rect 16486 9152 16542 9208
rect 16302 8336 16358 8392
rect 16118 8200 16174 8256
rect 15782 7642 15838 7644
rect 15862 7642 15918 7644
rect 15942 7642 15998 7644
rect 16022 7642 16078 7644
rect 15782 7590 15808 7642
rect 15808 7590 15838 7642
rect 15862 7590 15872 7642
rect 15872 7590 15918 7642
rect 15942 7590 15988 7642
rect 15988 7590 15998 7642
rect 16022 7590 16052 7642
rect 16052 7590 16078 7642
rect 15782 7588 15838 7590
rect 15862 7588 15918 7590
rect 15942 7588 15998 7590
rect 16022 7588 16078 7590
rect 16026 6704 16082 6760
rect 15782 6554 15838 6556
rect 15862 6554 15918 6556
rect 15942 6554 15998 6556
rect 16022 6554 16078 6556
rect 15782 6502 15808 6554
rect 15808 6502 15838 6554
rect 15862 6502 15872 6554
rect 15872 6502 15918 6554
rect 15942 6502 15988 6554
rect 15988 6502 15998 6554
rect 16022 6502 16052 6554
rect 16052 6502 16078 6554
rect 15782 6500 15838 6502
rect 15862 6500 15918 6502
rect 15942 6500 15998 6502
rect 16022 6500 16078 6502
rect 16210 7928 16266 7984
rect 16302 6976 16358 7032
rect 15782 5466 15838 5468
rect 15862 5466 15918 5468
rect 15942 5466 15998 5468
rect 16022 5466 16078 5468
rect 15782 5414 15808 5466
rect 15808 5414 15838 5466
rect 15862 5414 15872 5466
rect 15872 5414 15918 5466
rect 15942 5414 15988 5466
rect 15988 5414 15998 5466
rect 16022 5414 16052 5466
rect 16052 5414 16078 5466
rect 15782 5412 15838 5414
rect 15862 5412 15918 5414
rect 15942 5412 15998 5414
rect 16022 5412 16078 5414
rect 15750 5208 15806 5264
rect 15658 4800 15714 4856
rect 15934 5092 15990 5128
rect 15934 5072 15936 5092
rect 15936 5072 15988 5092
rect 15988 5072 15990 5092
rect 15782 4378 15838 4380
rect 15862 4378 15918 4380
rect 15942 4378 15998 4380
rect 16022 4378 16078 4380
rect 15782 4326 15808 4378
rect 15808 4326 15838 4378
rect 15862 4326 15872 4378
rect 15872 4326 15918 4378
rect 15942 4326 15988 4378
rect 15988 4326 15998 4378
rect 16022 4326 16052 4378
rect 16052 4326 16078 4378
rect 15782 4324 15838 4326
rect 15862 4324 15918 4326
rect 15942 4324 15998 4326
rect 16022 4324 16078 4326
rect 16486 8064 16542 8120
rect 16670 8336 16726 8392
rect 17774 16088 17830 16144
rect 17682 15000 17738 15056
rect 17406 13776 17462 13832
rect 17130 11872 17186 11928
rect 17038 11636 17040 11656
rect 17040 11636 17092 11656
rect 17092 11636 17094 11656
rect 17038 11600 17094 11636
rect 16762 7792 16818 7848
rect 16118 3712 16174 3768
rect 16486 3576 16542 3632
rect 3422 720 3478 776
rect 15782 3290 15838 3292
rect 15862 3290 15918 3292
rect 15942 3290 15998 3292
rect 16022 3290 16078 3292
rect 15782 3238 15808 3290
rect 15808 3238 15838 3290
rect 15862 3238 15872 3290
rect 15872 3238 15918 3290
rect 15942 3238 15988 3290
rect 15988 3238 15998 3290
rect 16022 3238 16052 3290
rect 16052 3238 16078 3290
rect 15782 3236 15838 3238
rect 15862 3236 15918 3238
rect 15942 3236 15998 3238
rect 16022 3236 16078 3238
rect 18142 14592 18198 14648
rect 17590 12824 17646 12880
rect 17498 11872 17554 11928
rect 17498 10648 17554 10704
rect 17406 10376 17462 10432
rect 15782 2202 15838 2204
rect 15862 2202 15918 2204
rect 15942 2202 15998 2204
rect 16022 2202 16078 2204
rect 15782 2150 15808 2202
rect 15808 2150 15838 2202
rect 15862 2150 15872 2202
rect 15872 2150 15918 2202
rect 15942 2150 15988 2202
rect 15988 2150 15998 2202
rect 16022 2150 16052 2202
rect 16052 2150 16078 2202
rect 15782 2148 15838 2150
rect 15862 2148 15918 2150
rect 15942 2148 15998 2150
rect 16022 2148 16078 2150
rect 15474 176 15530 232
rect 16854 2624 16910 2680
rect 17774 13524 17830 13560
rect 17774 13504 17776 13524
rect 17776 13504 17828 13524
rect 17828 13504 17830 13524
rect 17866 12280 17922 12336
rect 18050 13096 18106 13152
rect 18050 12708 18106 12744
rect 18050 12688 18052 12708
rect 18052 12688 18104 12708
rect 18104 12688 18106 12708
rect 17958 11192 18014 11248
rect 18142 11736 18198 11792
rect 18142 11620 18198 11656
rect 18142 11600 18144 11620
rect 18144 11600 18196 11620
rect 18196 11600 18198 11620
rect 18418 14184 18474 14240
rect 18418 13812 18420 13832
rect 18420 13812 18472 13832
rect 18472 13812 18474 13832
rect 18418 13776 18474 13812
rect 18418 13504 18474 13560
rect 18418 12280 18474 12336
rect 18970 11228 18972 11248
rect 18972 11228 19024 11248
rect 19024 11228 19026 11248
rect 18970 11192 19026 11228
rect 18510 11056 18566 11112
rect 18418 10784 18474 10840
rect 18510 9968 18566 10024
rect 18510 9696 18566 9752
rect 18050 9288 18106 9344
rect 17866 7656 17922 7712
rect 18142 7384 18198 7440
rect 18050 7248 18106 7304
rect 17866 5480 17922 5536
rect 18234 6976 18290 7032
rect 18510 6568 18566 6624
rect 18510 6180 18566 6216
rect 18510 6160 18512 6180
rect 18512 6160 18564 6180
rect 18564 6160 18566 6180
rect 18510 5888 18566 5944
rect 18510 5092 18566 5128
rect 18510 5072 18512 5092
rect 18512 5072 18564 5092
rect 18564 5072 18566 5092
rect 18510 4684 18566 4720
rect 18510 4664 18512 4684
rect 18512 4664 18564 4684
rect 18564 4664 18566 4684
rect 18142 4256 18198 4312
rect 18142 3596 18198 3632
rect 18142 3576 18144 3596
rect 18144 3576 18196 3596
rect 18196 3576 18198 3596
rect 18510 4004 18566 4040
rect 18510 3984 18512 4004
rect 18512 3984 18564 4004
rect 18564 3984 18566 4004
rect 18510 3168 18566 3224
rect 17774 2624 17830 2680
rect 17038 1264 17094 1320
rect 16854 856 16910 912
rect 18142 2760 18198 2816
rect 18418 2352 18474 2408
rect 17866 1672 17922 1728
rect 18510 2080 18566 2136
rect 16486 448 16542 504
<< metal3 >>
rect 0 16962 800 16992
rect 3049 16962 3115 16965
rect 0 16960 3115 16962
rect 0 16904 3054 16960
rect 3110 16904 3115 16960
rect 0 16902 3115 16904
rect 0 16872 800 16902
rect 3049 16899 3115 16902
rect 17309 16962 17375 16965
rect 19200 16962 20000 16992
rect 17309 16960 20000 16962
rect 17309 16904 17314 16960
rect 17370 16904 20000 16960
rect 17309 16902 20000 16904
rect 17309 16899 17375 16902
rect 19200 16872 20000 16902
rect 0 16690 800 16720
rect 3509 16690 3575 16693
rect 0 16688 3575 16690
rect 0 16632 3514 16688
rect 3570 16632 3575 16688
rect 0 16630 3575 16632
rect 0 16600 800 16630
rect 3509 16627 3575 16630
rect 16205 16554 16271 16557
rect 19200 16554 20000 16584
rect 16205 16552 20000 16554
rect 16205 16496 16210 16552
rect 16266 16496 20000 16552
rect 16205 16494 20000 16496
rect 16205 16491 16271 16494
rect 19200 16464 20000 16494
rect 0 16282 800 16312
rect 3877 16282 3943 16285
rect 0 16280 3943 16282
rect 0 16224 3882 16280
rect 3938 16224 3943 16280
rect 0 16222 3943 16224
rect 0 16192 800 16222
rect 3877 16219 3943 16222
rect 17769 16146 17835 16149
rect 19200 16146 20000 16176
rect 17769 16144 20000 16146
rect 17769 16088 17774 16144
rect 17830 16088 20000 16144
rect 17769 16086 20000 16088
rect 17769 16083 17835 16086
rect 19200 16056 20000 16086
rect 0 16010 800 16040
rect 1485 16010 1551 16013
rect 0 16008 1551 16010
rect 0 15952 1490 16008
rect 1546 15952 1551 16008
rect 0 15950 1551 15952
rect 0 15920 800 15950
rect 1485 15947 1551 15950
rect 16481 15738 16547 15741
rect 19200 15738 20000 15768
rect 16481 15736 20000 15738
rect 16481 15680 16486 15736
rect 16542 15680 20000 15736
rect 16481 15678 20000 15680
rect 16481 15675 16547 15678
rect 19200 15648 20000 15678
rect 0 15602 800 15632
rect 4245 15602 4311 15605
rect 0 15600 4311 15602
rect 0 15544 4250 15600
rect 4306 15544 4311 15600
rect 0 15542 4311 15544
rect 0 15512 800 15542
rect 4245 15539 4311 15542
rect 16941 15466 17007 15469
rect 19200 15466 20000 15496
rect 16941 15464 20000 15466
rect 16941 15408 16946 15464
rect 17002 15408 20000 15464
rect 16941 15406 20000 15408
rect 16941 15403 17007 15406
rect 19200 15376 20000 15406
rect 0 15330 800 15360
rect 4153 15330 4219 15333
rect 0 15328 4219 15330
rect 0 15272 4158 15328
rect 4214 15272 4219 15328
rect 0 15270 4219 15272
rect 0 15240 800 15270
rect 4153 15267 4219 15270
rect 0 15058 800 15088
rect 1853 15058 1919 15061
rect 0 15056 1919 15058
rect 0 15000 1858 15056
rect 1914 15000 1919 15056
rect 0 14998 1919 15000
rect 0 14968 800 14998
rect 1853 14995 1919 14998
rect 17677 15058 17743 15061
rect 19200 15058 20000 15088
rect 17677 15056 20000 15058
rect 17677 15000 17682 15056
rect 17738 15000 20000 15056
rect 17677 14998 20000 15000
rect 17677 14995 17743 14998
rect 19200 14968 20000 14998
rect 6874 14720 7194 14721
rect 0 14650 800 14680
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7194 14720
rect 6874 14655 7194 14656
rect 12805 14720 13125 14721
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 14655 13125 14656
rect 2221 14650 2287 14653
rect 0 14648 2287 14650
rect 0 14592 2226 14648
rect 2282 14592 2287 14648
rect 0 14590 2287 14592
rect 0 14560 800 14590
rect 2221 14587 2287 14590
rect 18137 14650 18203 14653
rect 19200 14650 20000 14680
rect 18137 14648 20000 14650
rect 18137 14592 18142 14648
rect 18198 14592 20000 14648
rect 18137 14590 20000 14592
rect 18137 14587 18203 14590
rect 19200 14560 20000 14590
rect 0 14378 800 14408
rect 1853 14378 1919 14381
rect 0 14376 1919 14378
rect 0 14320 1858 14376
rect 1914 14320 1919 14376
rect 0 14318 1919 14320
rect 0 14288 800 14318
rect 1853 14315 1919 14318
rect 18413 14242 18479 14245
rect 19200 14242 20000 14272
rect 18413 14240 20000 14242
rect 18413 14184 18418 14240
rect 18474 14184 20000 14240
rect 18413 14182 20000 14184
rect 18413 14179 18479 14182
rect 3909 14176 4229 14177
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 14111 4229 14112
rect 9840 14176 10160 14177
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 14111 10160 14112
rect 15770 14176 16090 14177
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16090 14176
rect 19200 14152 20000 14182
rect 15770 14111 16090 14112
rect 0 13970 800 14000
rect 2129 13970 2195 13973
rect 0 13968 2195 13970
rect 0 13912 2134 13968
rect 2190 13912 2195 13968
rect 0 13910 2195 13912
rect 0 13880 800 13910
rect 2129 13907 2195 13910
rect 17401 13834 17467 13837
rect 17718 13834 17724 13836
rect 17401 13832 17724 13834
rect 17401 13776 17406 13832
rect 17462 13776 17724 13832
rect 17401 13774 17724 13776
rect 17401 13771 17467 13774
rect 17718 13772 17724 13774
rect 17788 13772 17794 13836
rect 18413 13834 18479 13837
rect 19200 13834 20000 13864
rect 18413 13832 20000 13834
rect 18413 13776 18418 13832
rect 18474 13776 20000 13832
rect 18413 13774 20000 13776
rect 18413 13771 18479 13774
rect 19200 13744 20000 13774
rect 0 13698 800 13728
rect 2773 13698 2839 13701
rect 0 13696 2839 13698
rect 0 13640 2778 13696
rect 2834 13640 2839 13696
rect 0 13638 2839 13640
rect 0 13608 800 13638
rect 2773 13635 2839 13638
rect 6874 13632 7194 13633
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7194 13632
rect 6874 13567 7194 13568
rect 12805 13632 13125 13633
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 13567 13125 13568
rect 16389 13562 16455 13565
rect 17769 13562 17835 13565
rect 16389 13560 17835 13562
rect 16389 13504 16394 13560
rect 16450 13504 17774 13560
rect 17830 13504 17835 13560
rect 16389 13502 17835 13504
rect 16389 13499 16455 13502
rect 17769 13499 17835 13502
rect 18413 13562 18479 13565
rect 19200 13562 20000 13592
rect 18413 13560 20000 13562
rect 18413 13504 18418 13560
rect 18474 13504 20000 13560
rect 18413 13502 20000 13504
rect 18413 13499 18479 13502
rect 19200 13472 20000 13502
rect 0 13290 800 13320
rect 1393 13290 1459 13293
rect 0 13288 1459 13290
rect 0 13232 1398 13288
rect 1454 13232 1459 13288
rect 0 13230 1459 13232
rect 0 13200 800 13230
rect 1393 13227 1459 13230
rect 18045 13154 18111 13157
rect 19200 13154 20000 13184
rect 18045 13152 20000 13154
rect 18045 13096 18050 13152
rect 18106 13096 20000 13152
rect 18045 13094 20000 13096
rect 18045 13091 18111 13094
rect 3909 13088 4229 13089
rect 0 13018 800 13048
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 13023 4229 13024
rect 9840 13088 10160 13089
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 13023 10160 13024
rect 15770 13088 16090 13089
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16090 13088
rect 19200 13064 20000 13094
rect 15770 13023 16090 13024
rect 2221 13018 2287 13021
rect 0 13016 2287 13018
rect 0 12960 2226 13016
rect 2282 12960 2287 13016
rect 0 12958 2287 12960
rect 0 12928 800 12958
rect 2221 12955 2287 12958
rect 16982 12820 16988 12884
rect 17052 12882 17058 12884
rect 17585 12882 17651 12885
rect 17052 12880 17651 12882
rect 17052 12824 17590 12880
rect 17646 12824 17651 12880
rect 17052 12822 17651 12824
rect 17052 12820 17058 12822
rect 17585 12819 17651 12822
rect 0 12746 800 12776
rect 1485 12746 1551 12749
rect 0 12744 1551 12746
rect 0 12688 1490 12744
rect 1546 12688 1551 12744
rect 0 12686 1551 12688
rect 0 12656 800 12686
rect 1485 12683 1551 12686
rect 9622 12684 9628 12748
rect 9692 12746 9698 12748
rect 17033 12746 17099 12749
rect 9692 12744 17099 12746
rect 9692 12688 17038 12744
rect 17094 12688 17099 12744
rect 9692 12686 17099 12688
rect 9692 12684 9698 12686
rect 17033 12683 17099 12686
rect 18045 12746 18111 12749
rect 19200 12746 20000 12776
rect 18045 12744 20000 12746
rect 18045 12688 18050 12744
rect 18106 12688 20000 12744
rect 18045 12686 20000 12688
rect 18045 12683 18111 12686
rect 19200 12656 20000 12686
rect 6874 12544 7194 12545
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7194 12544
rect 6874 12479 7194 12480
rect 12805 12544 13125 12545
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 12805 12479 13125 12480
rect 0 12338 800 12368
rect 1853 12338 1919 12341
rect 0 12336 1919 12338
rect 0 12280 1858 12336
rect 1914 12280 1919 12336
rect 0 12278 1919 12280
rect 0 12248 800 12278
rect 1853 12275 1919 12278
rect 5901 12338 5967 12341
rect 10593 12338 10659 12341
rect 17861 12338 17927 12341
rect 5901 12336 17927 12338
rect 5901 12280 5906 12336
rect 5962 12280 10598 12336
rect 10654 12280 17866 12336
rect 17922 12280 17927 12336
rect 5901 12278 17927 12280
rect 5901 12275 5967 12278
rect 10593 12275 10659 12278
rect 17861 12275 17927 12278
rect 18413 12338 18479 12341
rect 19200 12338 20000 12368
rect 18413 12336 20000 12338
rect 18413 12280 18418 12336
rect 18474 12280 20000 12336
rect 18413 12278 20000 12280
rect 18413 12275 18479 12278
rect 19200 12248 20000 12278
rect 6545 12202 6611 12205
rect 7833 12202 7899 12205
rect 6545 12200 7899 12202
rect 6545 12144 6550 12200
rect 6606 12144 7838 12200
rect 7894 12144 7899 12200
rect 6545 12142 7899 12144
rect 6545 12139 6611 12142
rect 7833 12139 7899 12142
rect 8109 12202 8175 12205
rect 11881 12202 11947 12205
rect 8109 12200 11947 12202
rect 8109 12144 8114 12200
rect 8170 12144 11886 12200
rect 11942 12144 11947 12200
rect 8109 12142 11947 12144
rect 8109 12139 8175 12142
rect 11881 12139 11947 12142
rect 0 12066 800 12096
rect 1393 12066 1459 12069
rect 0 12064 1459 12066
rect 0 12008 1398 12064
rect 1454 12008 1459 12064
rect 0 12006 1459 12008
rect 0 11976 800 12006
rect 1393 12003 1459 12006
rect 4797 12066 4863 12069
rect 9622 12066 9628 12068
rect 4797 12064 9628 12066
rect 4797 12008 4802 12064
rect 4858 12008 9628 12064
rect 4797 12006 9628 12008
rect 4797 12003 4863 12006
rect 3909 12000 4229 12001
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 11935 4229 11936
rect 5214 11933 5274 12006
rect 9622 12004 9628 12006
rect 9692 12004 9698 12068
rect 9840 12000 10160 12001
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 11935 10160 11936
rect 15770 12000 16090 12001
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16090 12000
rect 15770 11935 16090 11936
rect 5165 11928 5274 11933
rect 5165 11872 5170 11928
rect 5226 11872 5274 11928
rect 5165 11870 5274 11872
rect 5349 11930 5415 11933
rect 9213 11930 9279 11933
rect 14089 11930 14155 11933
rect 15469 11930 15535 11933
rect 5349 11928 9279 11930
rect 5349 11872 5354 11928
rect 5410 11872 9218 11928
rect 9274 11872 9279 11928
rect 5349 11870 9279 11872
rect 5165 11867 5231 11870
rect 5349 11867 5415 11870
rect 9213 11867 9279 11870
rect 10366 11928 15535 11930
rect 10366 11872 14094 11928
rect 14150 11872 15474 11928
rect 15530 11872 15535 11928
rect 10366 11870 15535 11872
rect 6177 11794 6243 11797
rect 10366 11794 10426 11870
rect 14089 11867 14155 11870
rect 15469 11867 15535 11870
rect 16573 11930 16639 11933
rect 17125 11930 17191 11933
rect 16573 11928 17191 11930
rect 16573 11872 16578 11928
rect 16634 11872 17130 11928
rect 17186 11872 17191 11928
rect 16573 11870 17191 11872
rect 16573 11867 16639 11870
rect 17125 11867 17191 11870
rect 17493 11930 17559 11933
rect 19200 11930 20000 11960
rect 17493 11928 20000 11930
rect 17493 11872 17498 11928
rect 17554 11872 20000 11928
rect 17493 11870 20000 11872
rect 17493 11867 17559 11870
rect 19200 11840 20000 11870
rect 6177 11792 10426 11794
rect 6177 11736 6182 11792
rect 6238 11736 10426 11792
rect 6177 11734 10426 11736
rect 10501 11794 10567 11797
rect 18137 11794 18203 11797
rect 10501 11792 18203 11794
rect 10501 11736 10506 11792
rect 10562 11736 18142 11792
rect 18198 11736 18203 11792
rect 10501 11734 18203 11736
rect 6177 11731 6243 11734
rect 10501 11731 10567 11734
rect 18137 11731 18203 11734
rect 0 11658 800 11688
rect 1761 11658 1827 11661
rect 0 11656 1827 11658
rect 0 11600 1766 11656
rect 1822 11600 1827 11656
rect 0 11598 1827 11600
rect 0 11568 800 11598
rect 1761 11595 1827 11598
rect 3969 11658 4035 11661
rect 16246 11658 16252 11660
rect 3969 11656 16252 11658
rect 3969 11600 3974 11656
rect 4030 11600 16252 11656
rect 3969 11598 16252 11600
rect 3969 11595 4035 11598
rect 16246 11596 16252 11598
rect 16316 11658 16322 11660
rect 17033 11658 17099 11661
rect 16316 11656 17099 11658
rect 16316 11600 17038 11656
rect 17094 11600 17099 11656
rect 16316 11598 17099 11600
rect 16316 11596 16322 11598
rect 17033 11595 17099 11598
rect 18137 11658 18203 11661
rect 19200 11658 20000 11688
rect 18137 11656 20000 11658
rect 18137 11600 18142 11656
rect 18198 11600 20000 11656
rect 18137 11598 20000 11600
rect 18137 11595 18203 11598
rect 19200 11568 20000 11598
rect 8201 11522 8267 11525
rect 8753 11522 8819 11525
rect 8201 11520 8819 11522
rect 8201 11464 8206 11520
rect 8262 11464 8758 11520
rect 8814 11464 8819 11520
rect 8201 11462 8819 11464
rect 8201 11459 8267 11462
rect 8753 11459 8819 11462
rect 9949 11522 10015 11525
rect 12617 11522 12683 11525
rect 9949 11520 12683 11522
rect 9949 11464 9954 11520
rect 10010 11464 12622 11520
rect 12678 11464 12683 11520
rect 9949 11462 12683 11464
rect 9949 11459 10015 11462
rect 12617 11459 12683 11462
rect 16389 11524 16455 11525
rect 16389 11520 16436 11524
rect 16500 11522 16506 11524
rect 16389 11464 16394 11520
rect 16389 11460 16436 11464
rect 16500 11462 16546 11522
rect 16500 11460 16506 11462
rect 16389 11459 16455 11460
rect 6874 11456 7194 11457
rect 0 11386 800 11416
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7194 11456
rect 6874 11391 7194 11392
rect 12805 11456 13125 11457
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 11391 13125 11392
rect 1485 11386 1551 11389
rect 0 11384 1551 11386
rect 0 11328 1490 11384
rect 1546 11328 1551 11384
rect 0 11326 1551 11328
rect 0 11296 800 11326
rect 1485 11323 1551 11326
rect 7373 11386 7439 11389
rect 13721 11386 13787 11389
rect 16849 11386 16915 11389
rect 7373 11384 11346 11386
rect 7373 11328 7378 11384
rect 7434 11328 11346 11384
rect 7373 11326 11346 11328
rect 7373 11323 7439 11326
rect 1945 11250 2011 11253
rect 9857 11250 9923 11253
rect 1945 11248 9923 11250
rect 1945 11192 1950 11248
rect 2006 11192 9862 11248
rect 9918 11192 9923 11248
rect 1945 11190 9923 11192
rect 1945 11187 2011 11190
rect 9857 11187 9923 11190
rect 6269 11114 6335 11117
rect 11053 11114 11119 11117
rect 6269 11112 11119 11114
rect 6269 11056 6274 11112
rect 6330 11056 11058 11112
rect 11114 11056 11119 11112
rect 6269 11054 11119 11056
rect 11286 11114 11346 11326
rect 13721 11384 16915 11386
rect 13721 11328 13726 11384
rect 13782 11328 16854 11384
rect 16910 11328 16915 11384
rect 13721 11326 16915 11328
rect 13721 11323 13787 11326
rect 16849 11323 16915 11326
rect 12341 11250 12407 11253
rect 17953 11250 18019 11253
rect 12341 11248 18019 11250
rect 12341 11192 12346 11248
rect 12402 11192 17958 11248
rect 18014 11192 18019 11248
rect 12341 11190 18019 11192
rect 12341 11187 12407 11190
rect 17953 11187 18019 11190
rect 18965 11250 19031 11253
rect 19200 11250 20000 11280
rect 18965 11248 20000 11250
rect 18965 11192 18970 11248
rect 19026 11192 20000 11248
rect 18965 11190 20000 11192
rect 18965 11187 19031 11190
rect 19200 11160 20000 11190
rect 12249 11114 12315 11117
rect 18505 11114 18571 11117
rect 11286 11112 18571 11114
rect 11286 11056 12254 11112
rect 12310 11056 18510 11112
rect 18566 11056 18571 11112
rect 11286 11054 18571 11056
rect 6269 11051 6335 11054
rect 11053 11051 11119 11054
rect 12249 11051 12315 11054
rect 18505 11051 18571 11054
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 6085 10978 6151 10981
rect 9121 10978 9187 10981
rect 6085 10976 9187 10978
rect 6085 10920 6090 10976
rect 6146 10920 9126 10976
rect 9182 10920 9187 10976
rect 6085 10918 9187 10920
rect 6085 10915 6151 10918
rect 9121 10915 9187 10918
rect 3909 10912 4229 10913
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 10847 4229 10848
rect 9840 10912 10160 10913
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 10847 10160 10848
rect 15770 10912 16090 10913
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16090 10912
rect 15770 10847 16090 10848
rect 13169 10842 13235 10845
rect 15101 10842 15167 10845
rect 13169 10840 15167 10842
rect 13169 10784 13174 10840
rect 13230 10784 15106 10840
rect 15162 10784 15167 10840
rect 13169 10782 15167 10784
rect 13169 10779 13235 10782
rect 15101 10779 15167 10782
rect 18413 10842 18479 10845
rect 19200 10842 20000 10872
rect 18413 10840 20000 10842
rect 18413 10784 18418 10840
rect 18474 10784 20000 10840
rect 18413 10782 20000 10784
rect 18413 10779 18479 10782
rect 19200 10752 20000 10782
rect 0 10706 800 10736
rect 1853 10706 1919 10709
rect 5901 10706 5967 10709
rect 0 10704 1919 10706
rect 0 10648 1858 10704
rect 1914 10648 1919 10704
rect 0 10646 1919 10648
rect 0 10616 800 10646
rect 1853 10643 1919 10646
rect 5766 10704 5967 10706
rect 5766 10648 5906 10704
rect 5962 10648 5967 10704
rect 5766 10646 5967 10648
rect 5766 10573 5826 10646
rect 5901 10643 5967 10646
rect 13261 10706 13327 10709
rect 17493 10706 17559 10709
rect 13261 10704 17559 10706
rect 13261 10648 13266 10704
rect 13322 10648 17498 10704
rect 17554 10648 17559 10704
rect 13261 10646 17559 10648
rect 13261 10643 13327 10646
rect 17493 10643 17559 10646
rect 5717 10568 5826 10573
rect 5717 10512 5722 10568
rect 5778 10512 5826 10568
rect 5717 10510 5826 10512
rect 9857 10570 9923 10573
rect 10409 10570 10475 10573
rect 13169 10570 13235 10573
rect 9857 10568 10475 10570
rect 9857 10512 9862 10568
rect 9918 10512 10414 10568
rect 10470 10512 10475 10568
rect 9857 10510 10475 10512
rect 5717 10507 5783 10510
rect 9857 10507 9923 10510
rect 10409 10507 10475 10510
rect 12574 10568 13235 10570
rect 12574 10512 13174 10568
rect 13230 10512 13235 10568
rect 12574 10510 13235 10512
rect 0 10434 800 10464
rect 1669 10434 1735 10437
rect 0 10432 1735 10434
rect 0 10376 1674 10432
rect 1730 10376 1735 10432
rect 0 10374 1735 10376
rect 0 10344 800 10374
rect 1669 10371 1735 10374
rect 8753 10434 8819 10437
rect 12574 10434 12634 10510
rect 13169 10507 13235 10510
rect 8753 10432 12634 10434
rect 8753 10376 8758 10432
rect 8814 10376 12634 10432
rect 8753 10374 12634 10376
rect 17401 10434 17467 10437
rect 19200 10434 20000 10464
rect 17401 10432 20000 10434
rect 17401 10376 17406 10432
rect 17462 10376 20000 10432
rect 17401 10374 20000 10376
rect 8753 10371 8819 10374
rect 17401 10371 17467 10374
rect 6874 10368 7194 10369
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7194 10368
rect 6874 10303 7194 10304
rect 12805 10368 13125 10369
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 19200 10344 20000 10374
rect 12805 10303 13125 10304
rect 2221 10298 2287 10301
rect 5073 10298 5139 10301
rect 2221 10296 5139 10298
rect 2221 10240 2226 10296
rect 2282 10240 5078 10296
rect 5134 10240 5139 10296
rect 2221 10238 5139 10240
rect 2221 10235 2287 10238
rect 5073 10235 5139 10238
rect 6637 10298 6703 10301
rect 10041 10298 10107 10301
rect 10501 10298 10567 10301
rect 6637 10296 6746 10298
rect 6637 10240 6642 10296
rect 6698 10240 6746 10296
rect 6637 10235 6746 10240
rect 10041 10296 10567 10298
rect 10041 10240 10046 10296
rect 10102 10240 10506 10296
rect 10562 10240 10567 10296
rect 10041 10238 10567 10240
rect 10041 10235 10107 10238
rect 10501 10235 10567 10238
rect 4705 10162 4771 10165
rect 4432 10160 4771 10162
rect 4432 10104 4710 10160
rect 4766 10104 4771 10160
rect 4432 10102 4771 10104
rect 0 10026 800 10056
rect 4432 10029 4492 10102
rect 4705 10099 4771 10102
rect 5349 10162 5415 10165
rect 6085 10162 6151 10165
rect 5349 10160 6151 10162
rect 5349 10104 5354 10160
rect 5410 10104 6090 10160
rect 6146 10104 6151 10160
rect 5349 10102 6151 10104
rect 6686 10162 6746 10235
rect 6821 10162 6887 10165
rect 6686 10160 6887 10162
rect 6686 10104 6826 10160
rect 6882 10104 6887 10160
rect 6686 10102 6887 10104
rect 5349 10099 5415 10102
rect 6085 10099 6151 10102
rect 6821 10099 6887 10102
rect 8017 10162 8083 10165
rect 9029 10162 9095 10165
rect 8017 10160 9095 10162
rect 8017 10104 8022 10160
rect 8078 10104 9034 10160
rect 9090 10104 9095 10160
rect 8017 10102 9095 10104
rect 8017 10099 8083 10102
rect 9029 10099 9095 10102
rect 1485 10026 1551 10029
rect 0 10024 1551 10026
rect 0 9968 1490 10024
rect 1546 9968 1551 10024
rect 0 9966 1551 9968
rect 0 9936 800 9966
rect 1485 9963 1551 9966
rect 1945 10026 2011 10029
rect 1945 10024 4354 10026
rect 1945 9968 1950 10024
rect 2006 9968 4354 10024
rect 1945 9966 4354 9968
rect 1945 9963 2011 9966
rect 4294 9890 4354 9966
rect 4429 10024 4495 10029
rect 4429 9968 4434 10024
rect 4490 9968 4495 10024
rect 4429 9963 4495 9968
rect 4797 10026 4863 10029
rect 6913 10026 6979 10029
rect 7281 10026 7347 10029
rect 8201 10026 8267 10029
rect 4797 10024 8267 10026
rect 4797 9968 4802 10024
rect 4858 9968 6918 10024
rect 6974 9968 7286 10024
rect 7342 9968 8206 10024
rect 8262 9968 8267 10024
rect 4797 9966 8267 9968
rect 4797 9963 4863 9966
rect 6913 9963 6979 9966
rect 7281 9963 7347 9966
rect 8201 9963 8267 9966
rect 8477 10026 8543 10029
rect 9121 10026 9187 10029
rect 9489 10026 9555 10029
rect 8477 10024 9555 10026
rect 8477 9968 8482 10024
rect 8538 9968 9126 10024
rect 9182 9968 9494 10024
rect 9550 9968 9555 10024
rect 8477 9966 9555 9968
rect 8477 9963 8543 9966
rect 9121 9963 9187 9966
rect 9489 9963 9555 9966
rect 15745 10026 15811 10029
rect 18505 10026 18571 10029
rect 19200 10026 20000 10056
rect 15745 10024 16498 10026
rect 15745 9968 15750 10024
rect 15806 9968 16498 10024
rect 15745 9966 16498 9968
rect 15745 9963 15811 9966
rect 16438 9893 16498 9966
rect 18505 10024 20000 10026
rect 18505 9968 18510 10024
rect 18566 9968 20000 10024
rect 18505 9966 20000 9968
rect 18505 9963 18571 9966
rect 19200 9936 20000 9966
rect 8569 9890 8635 9893
rect 4294 9888 8635 9890
rect 4294 9832 8574 9888
rect 8630 9832 8635 9888
rect 4294 9830 8635 9832
rect 16438 9888 16547 9893
rect 16438 9832 16486 9888
rect 16542 9832 16547 9888
rect 16438 9830 16547 9832
rect 8569 9827 8635 9830
rect 16481 9827 16547 9830
rect 3909 9824 4229 9825
rect 0 9754 800 9784
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 9759 4229 9760
rect 9840 9824 10160 9825
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 9759 10160 9760
rect 15770 9824 16090 9825
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16090 9824
rect 15770 9759 16090 9760
rect 3049 9754 3115 9757
rect 0 9752 3115 9754
rect 0 9696 3054 9752
rect 3110 9696 3115 9752
rect 0 9694 3115 9696
rect 0 9664 800 9694
rect 3049 9691 3115 9694
rect 4889 9754 4955 9757
rect 5533 9754 5599 9757
rect 6177 9756 6243 9757
rect 4889 9752 5599 9754
rect 4889 9696 4894 9752
rect 4950 9696 5538 9752
rect 5594 9696 5599 9752
rect 4889 9694 5599 9696
rect 4889 9691 4955 9694
rect 5533 9691 5599 9694
rect 6126 9692 6132 9756
rect 6196 9754 6243 9756
rect 12249 9754 12315 9757
rect 15469 9754 15535 9757
rect 16430 9754 16436 9756
rect 6196 9752 6288 9754
rect 6238 9696 6288 9752
rect 6196 9694 6288 9696
rect 12249 9752 15535 9754
rect 12249 9696 12254 9752
rect 12310 9696 15474 9752
rect 15530 9696 15535 9752
rect 12249 9694 15535 9696
rect 6196 9692 6243 9694
rect 6177 9691 6243 9692
rect 12249 9691 12315 9694
rect 15469 9691 15535 9694
rect 16254 9694 16436 9754
rect 16021 9690 16087 9693
rect 16254 9690 16314 9694
rect 16430 9692 16436 9694
rect 16500 9692 16506 9756
rect 18505 9754 18571 9757
rect 19200 9754 20000 9784
rect 18505 9752 20000 9754
rect 18505 9696 18510 9752
rect 18566 9696 20000 9752
rect 18505 9694 20000 9696
rect 18505 9691 18571 9694
rect 16021 9688 16314 9690
rect 16021 9632 16026 9688
rect 16082 9632 16314 9688
rect 19200 9664 20000 9694
rect 16021 9630 16314 9632
rect 16021 9627 16087 9630
rect 5625 9618 5691 9621
rect 7465 9618 7531 9621
rect 5625 9616 7531 9618
rect 5625 9560 5630 9616
rect 5686 9560 7470 9616
rect 7526 9560 7531 9616
rect 5625 9558 7531 9560
rect 5625 9555 5691 9558
rect 7465 9555 7531 9558
rect 8201 9618 8267 9621
rect 10685 9618 10751 9621
rect 8201 9616 10751 9618
rect 8201 9560 8206 9616
rect 8262 9560 10690 9616
rect 10746 9560 10751 9616
rect 8201 9558 10751 9560
rect 8201 9555 8267 9558
rect 10685 9555 10751 9558
rect 11789 9618 11855 9621
rect 13445 9618 13511 9621
rect 11789 9616 13511 9618
rect 11789 9560 11794 9616
rect 11850 9560 13450 9616
rect 13506 9560 13511 9616
rect 11789 9558 13511 9560
rect 11789 9555 11855 9558
rect 13445 9555 13511 9558
rect 4705 9482 4771 9485
rect 11145 9482 11211 9485
rect 4705 9480 11211 9482
rect 4705 9424 4710 9480
rect 4766 9424 11150 9480
rect 11206 9424 11211 9480
rect 4705 9422 11211 9424
rect 4705 9419 4771 9422
rect 11145 9419 11211 9422
rect 11789 9482 11855 9485
rect 13169 9482 13235 9485
rect 13302 9482 13308 9484
rect 11789 9480 13308 9482
rect 11789 9424 11794 9480
rect 11850 9424 13174 9480
rect 13230 9424 13308 9480
rect 11789 9422 13308 9424
rect 11789 9419 11855 9422
rect 13169 9419 13235 9422
rect 13302 9420 13308 9422
rect 13372 9420 13378 9484
rect 0 9346 800 9376
rect 3785 9346 3851 9349
rect 0 9344 3851 9346
rect 0 9288 3790 9344
rect 3846 9288 3851 9344
rect 0 9286 3851 9288
rect 0 9256 800 9286
rect 3785 9283 3851 9286
rect 4061 9346 4127 9349
rect 5073 9346 5139 9349
rect 4061 9344 5139 9346
rect 4061 9288 4066 9344
rect 4122 9288 5078 9344
rect 5134 9288 5139 9344
rect 4061 9286 5139 9288
rect 4061 9283 4127 9286
rect 5073 9283 5139 9286
rect 18045 9346 18111 9349
rect 19200 9346 20000 9376
rect 18045 9344 20000 9346
rect 18045 9288 18050 9344
rect 18106 9288 20000 9344
rect 18045 9286 20000 9288
rect 18045 9283 18111 9286
rect 6874 9280 7194 9281
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7194 9280
rect 6874 9215 7194 9216
rect 12805 9280 13125 9281
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 19200 9256 20000 9286
rect 12805 9215 13125 9216
rect 13261 9210 13327 9213
rect 13486 9210 13492 9212
rect 13261 9208 13492 9210
rect 13261 9152 13266 9208
rect 13322 9152 13492 9208
rect 13261 9150 13492 9152
rect 13261 9147 13327 9150
rect 13486 9148 13492 9150
rect 13556 9148 13562 9212
rect 16481 9210 16547 9213
rect 13632 9208 16547 9210
rect 13632 9152 16486 9208
rect 16542 9152 16547 9208
rect 13632 9150 16547 9152
rect 0 9074 800 9104
rect 3877 9074 3943 9077
rect 0 9072 3943 9074
rect 0 9016 3882 9072
rect 3938 9016 3943 9072
rect 0 9014 3943 9016
rect 0 8984 800 9014
rect 3877 9011 3943 9014
rect 4429 9076 4495 9077
rect 4429 9072 4476 9076
rect 4540 9074 4546 9076
rect 5533 9074 5599 9077
rect 10501 9074 10567 9077
rect 4429 9016 4434 9072
rect 4429 9012 4476 9016
rect 4540 9014 4586 9074
rect 5533 9072 10567 9074
rect 5533 9016 5538 9072
rect 5594 9016 10506 9072
rect 10562 9016 10567 9072
rect 5533 9014 10567 9016
rect 4540 9012 4546 9014
rect 4429 9011 4495 9012
rect 5533 9011 5599 9014
rect 10501 9011 10567 9014
rect 12566 9012 12572 9076
rect 12636 9074 12642 9076
rect 13353 9074 13419 9077
rect 12636 9072 13419 9074
rect 12636 9016 13358 9072
rect 13414 9016 13419 9072
rect 12636 9014 13419 9016
rect 12636 9012 12642 9014
rect 13353 9011 13419 9014
rect 4153 8938 4219 8941
rect 7557 8938 7623 8941
rect 4153 8936 7623 8938
rect 4153 8880 4158 8936
rect 4214 8880 7562 8936
rect 7618 8880 7623 8936
rect 4153 8878 7623 8880
rect 4153 8875 4219 8878
rect 7557 8875 7623 8878
rect 8201 8938 8267 8941
rect 8477 8938 8543 8941
rect 8201 8936 8543 8938
rect 8201 8880 8206 8936
rect 8262 8880 8482 8936
rect 8538 8880 8543 8936
rect 8201 8878 8543 8880
rect 8201 8875 8267 8878
rect 8477 8875 8543 8878
rect 11145 8938 11211 8941
rect 13632 8938 13692 9150
rect 16481 9147 16547 9150
rect 15469 9074 15535 9077
rect 16021 9074 16087 9077
rect 15469 9072 16087 9074
rect 15469 9016 15474 9072
rect 15530 9016 16026 9072
rect 16082 9016 16087 9072
rect 15469 9014 16087 9016
rect 15469 9011 15535 9014
rect 16021 9011 16087 9014
rect 11145 8936 13692 8938
rect 11145 8880 11150 8936
rect 11206 8880 13692 8936
rect 11145 8878 13692 8880
rect 15745 8938 15811 8941
rect 19200 8938 20000 8968
rect 15745 8936 20000 8938
rect 15745 8880 15750 8936
rect 15806 8880 20000 8936
rect 15745 8878 20000 8880
rect 11145 8875 11211 8878
rect 15745 8875 15811 8878
rect 19200 8848 20000 8878
rect 0 8802 800 8832
rect 3325 8802 3391 8805
rect 0 8800 3391 8802
rect 0 8744 3330 8800
rect 3386 8744 3391 8800
rect 0 8742 3391 8744
rect 0 8712 800 8742
rect 3325 8739 3391 8742
rect 3909 8736 4229 8737
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 8671 4229 8672
rect 9840 8736 10160 8737
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 8671 10160 8672
rect 15770 8736 16090 8737
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16090 8736
rect 15770 8671 16090 8672
rect 3233 8530 3299 8533
rect 7281 8530 7347 8533
rect 3233 8528 7347 8530
rect 3233 8472 3238 8528
rect 3294 8472 7286 8528
rect 7342 8472 7347 8528
rect 3233 8470 7347 8472
rect 3233 8467 3299 8470
rect 7281 8467 7347 8470
rect 15285 8530 15351 8533
rect 19200 8530 20000 8560
rect 15285 8528 20000 8530
rect 15285 8472 15290 8528
rect 15346 8472 20000 8528
rect 15285 8470 20000 8472
rect 15285 8467 15351 8470
rect 19200 8440 20000 8470
rect 0 8394 800 8424
rect 1485 8394 1551 8397
rect 0 8392 1551 8394
rect 0 8336 1490 8392
rect 1546 8336 1551 8392
rect 0 8334 1551 8336
rect 0 8304 800 8334
rect 1485 8331 1551 8334
rect 11881 8394 11947 8397
rect 14549 8394 14615 8397
rect 11881 8392 14615 8394
rect 11881 8336 11886 8392
rect 11942 8336 14554 8392
rect 14610 8336 14615 8392
rect 11881 8334 14615 8336
rect 11881 8331 11947 8334
rect 14549 8331 14615 8334
rect 16297 8394 16363 8397
rect 16665 8394 16731 8397
rect 16297 8392 16731 8394
rect 16297 8336 16302 8392
rect 16358 8336 16670 8392
rect 16726 8336 16731 8392
rect 16297 8334 16731 8336
rect 16297 8331 16363 8334
rect 16665 8331 16731 8334
rect 3969 8258 4035 8261
rect 4429 8258 4495 8261
rect 5165 8258 5231 8261
rect 3969 8256 5231 8258
rect 3969 8200 3974 8256
rect 4030 8200 4434 8256
rect 4490 8200 5170 8256
rect 5226 8200 5231 8256
rect 3969 8198 5231 8200
rect 3969 8195 4035 8198
rect 4429 8195 4495 8198
rect 5165 8195 5231 8198
rect 14038 8196 14044 8260
rect 14108 8258 14114 8260
rect 14273 8258 14339 8261
rect 14108 8256 14339 8258
rect 14108 8200 14278 8256
rect 14334 8200 14339 8256
rect 14108 8198 14339 8200
rect 14108 8196 14114 8198
rect 14273 8195 14339 8198
rect 16113 8258 16179 8261
rect 16246 8258 16252 8260
rect 16113 8256 16252 8258
rect 16113 8200 16118 8256
rect 16174 8200 16252 8256
rect 16113 8198 16252 8200
rect 16113 8195 16179 8198
rect 16246 8196 16252 8198
rect 16316 8196 16322 8260
rect 6874 8192 7194 8193
rect 0 8122 800 8152
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7194 8192
rect 6874 8127 7194 8128
rect 12805 8192 13125 8193
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 12805 8127 13125 8128
rect 1485 8122 1551 8125
rect 0 8120 1551 8122
rect 0 8064 1490 8120
rect 1546 8064 1551 8120
rect 0 8062 1551 8064
rect 0 8032 800 8062
rect 1485 8059 1551 8062
rect 16481 8122 16547 8125
rect 19200 8122 20000 8152
rect 16481 8120 20000 8122
rect 16481 8064 16486 8120
rect 16542 8064 20000 8120
rect 16481 8062 20000 8064
rect 16481 8059 16547 8062
rect 19200 8032 20000 8062
rect 4889 7986 4955 7989
rect 5257 7986 5323 7989
rect 4889 7984 5323 7986
rect 4889 7928 4894 7984
rect 4950 7928 5262 7984
rect 5318 7928 5323 7984
rect 4889 7926 5323 7928
rect 4889 7923 4955 7926
rect 5257 7923 5323 7926
rect 5809 7986 5875 7989
rect 8293 7986 8359 7989
rect 8845 7986 8911 7989
rect 5809 7984 8911 7986
rect 5809 7928 5814 7984
rect 5870 7928 8298 7984
rect 8354 7928 8850 7984
rect 8906 7928 8911 7984
rect 5809 7926 8911 7928
rect 5809 7923 5875 7926
rect 8293 7923 8359 7926
rect 8845 7923 8911 7926
rect 10961 7986 11027 7989
rect 13813 7986 13879 7989
rect 10961 7984 13879 7986
rect 10961 7928 10966 7984
rect 11022 7928 13818 7984
rect 13874 7928 13879 7984
rect 10961 7926 13879 7928
rect 10961 7923 11027 7926
rect 13813 7923 13879 7926
rect 14549 7986 14615 7989
rect 15469 7986 15535 7989
rect 16205 7986 16271 7989
rect 14549 7984 16271 7986
rect 14549 7928 14554 7984
rect 14610 7928 15474 7984
rect 15530 7928 16210 7984
rect 16266 7928 16271 7984
rect 14549 7926 16271 7928
rect 14549 7923 14615 7926
rect 15469 7923 15535 7926
rect 16205 7923 16271 7926
rect 9622 7788 9628 7852
rect 9692 7850 9698 7852
rect 9857 7850 9923 7853
rect 16757 7850 16823 7853
rect 19200 7850 20000 7880
rect 9692 7848 16823 7850
rect 9692 7792 9862 7848
rect 9918 7792 16762 7848
rect 16818 7792 16823 7848
rect 9692 7790 16823 7792
rect 9692 7788 9698 7790
rect 9857 7787 9923 7790
rect 16757 7787 16823 7790
rect 17910 7790 20000 7850
rect 0 7714 800 7744
rect 17910 7717 17970 7790
rect 19200 7760 20000 7790
rect 1393 7714 1459 7717
rect 0 7712 1459 7714
rect 0 7656 1398 7712
rect 1454 7656 1459 7712
rect 0 7654 1459 7656
rect 0 7624 800 7654
rect 1393 7651 1459 7654
rect 17861 7712 17970 7717
rect 17861 7656 17866 7712
rect 17922 7656 17970 7712
rect 17861 7654 17970 7656
rect 17861 7651 17927 7654
rect 3909 7648 4229 7649
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 7583 4229 7584
rect 9840 7648 10160 7649
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 7583 10160 7584
rect 15770 7648 16090 7649
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16090 7648
rect 15770 7583 16090 7584
rect 0 7442 800 7472
rect 1393 7442 1459 7445
rect 0 7440 1459 7442
rect 0 7384 1398 7440
rect 1454 7384 1459 7440
rect 0 7382 1459 7384
rect 0 7352 800 7382
rect 1393 7379 1459 7382
rect 1669 7442 1735 7445
rect 3417 7442 3483 7445
rect 4889 7442 4955 7445
rect 18137 7442 18203 7445
rect 19200 7442 20000 7472
rect 1669 7440 15762 7442
rect 1669 7384 1674 7440
rect 1730 7384 3422 7440
rect 3478 7384 4894 7440
rect 4950 7384 15762 7440
rect 1669 7382 15762 7384
rect 1669 7379 1735 7382
rect 3417 7379 3483 7382
rect 4889 7379 4955 7382
rect 9029 7306 9095 7309
rect 15702 7306 15762 7382
rect 18137 7440 20000 7442
rect 18137 7384 18142 7440
rect 18198 7384 20000 7440
rect 18137 7382 20000 7384
rect 18137 7379 18203 7382
rect 19200 7352 20000 7382
rect 18045 7306 18111 7309
rect 9029 7304 14658 7306
rect 9029 7248 9034 7304
rect 9090 7248 14658 7304
rect 9029 7246 14658 7248
rect 15702 7304 18111 7306
rect 15702 7248 18050 7304
rect 18106 7248 18111 7304
rect 15702 7246 18111 7248
rect 9029 7243 9095 7246
rect 14598 7170 14658 7246
rect 18045 7243 18111 7246
rect 14733 7170 14799 7173
rect 14598 7168 14799 7170
rect 14598 7112 14738 7168
rect 14794 7112 14799 7168
rect 14598 7110 14799 7112
rect 14733 7107 14799 7110
rect 6874 7104 7194 7105
rect 0 7034 800 7064
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7194 7104
rect 6874 7039 7194 7040
rect 12805 7104 13125 7105
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 7039 13125 7040
rect 2865 7034 2931 7037
rect 0 7032 2931 7034
rect 0 6976 2870 7032
rect 2926 6976 2931 7032
rect 0 6974 2931 6976
rect 0 6944 800 6974
rect 2865 6971 2931 6974
rect 13997 7034 14063 7037
rect 16297 7034 16363 7037
rect 13997 7032 16363 7034
rect 13997 6976 14002 7032
rect 14058 6976 16302 7032
rect 16358 6976 16363 7032
rect 13997 6974 16363 6976
rect 13997 6971 14063 6974
rect 16297 6971 16363 6974
rect 18229 7034 18295 7037
rect 19200 7034 20000 7064
rect 18229 7032 20000 7034
rect 18229 6976 18234 7032
rect 18290 6976 20000 7032
rect 18229 6974 20000 6976
rect 18229 6971 18295 6974
rect 19200 6944 20000 6974
rect 0 6762 800 6792
rect 1485 6762 1551 6765
rect 0 6760 1551 6762
rect 0 6704 1490 6760
rect 1546 6704 1551 6760
rect 0 6702 1551 6704
rect 0 6672 800 6702
rect 1485 6699 1551 6702
rect 13302 6700 13308 6764
rect 13372 6762 13378 6764
rect 13537 6762 13603 6765
rect 13372 6760 13603 6762
rect 13372 6704 13542 6760
rect 13598 6704 13603 6760
rect 13372 6702 13603 6704
rect 13372 6700 13378 6702
rect 13537 6699 13603 6702
rect 14038 6700 14044 6764
rect 14108 6762 14114 6764
rect 16021 6762 16087 6765
rect 14108 6760 16087 6762
rect 14108 6704 16026 6760
rect 16082 6704 16087 6760
rect 14108 6702 16087 6704
rect 14108 6700 14114 6702
rect 16021 6699 16087 6702
rect 10685 6626 10751 6629
rect 13997 6626 14063 6629
rect 10685 6624 14063 6626
rect 10685 6568 10690 6624
rect 10746 6568 14002 6624
rect 14058 6568 14063 6624
rect 10685 6566 14063 6568
rect 10685 6563 10751 6566
rect 13997 6563 14063 6566
rect 18505 6626 18571 6629
rect 19200 6626 20000 6656
rect 18505 6624 20000 6626
rect 18505 6568 18510 6624
rect 18566 6568 20000 6624
rect 18505 6566 20000 6568
rect 18505 6563 18571 6566
rect 3909 6560 4229 6561
rect 0 6490 800 6520
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 6495 4229 6496
rect 9840 6560 10160 6561
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 6495 10160 6496
rect 15770 6560 16090 6561
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16090 6560
rect 19200 6536 20000 6566
rect 15770 6495 16090 6496
rect 3601 6490 3667 6493
rect 0 6488 3667 6490
rect 0 6432 3606 6488
rect 3662 6432 3667 6488
rect 0 6430 3667 6432
rect 0 6400 800 6430
rect 3601 6427 3667 6430
rect 4337 6490 4403 6493
rect 5717 6490 5783 6493
rect 4337 6488 5783 6490
rect 4337 6432 4342 6488
rect 4398 6432 5722 6488
rect 5778 6432 5783 6488
rect 4337 6430 5783 6432
rect 4337 6427 4403 6430
rect 5717 6427 5783 6430
rect 2773 6354 2839 6357
rect 8661 6354 8727 6357
rect 2773 6352 8727 6354
rect 2773 6296 2778 6352
rect 2834 6296 8666 6352
rect 8722 6296 8727 6352
rect 2773 6294 8727 6296
rect 2773 6291 2839 6294
rect 8661 6291 8727 6294
rect 10685 6354 10751 6357
rect 10910 6354 10916 6356
rect 10685 6352 10916 6354
rect 10685 6296 10690 6352
rect 10746 6296 10916 6352
rect 10685 6294 10916 6296
rect 10685 6291 10751 6294
rect 10910 6292 10916 6294
rect 10980 6292 10986 6356
rect 11329 6354 11395 6357
rect 12801 6354 12867 6357
rect 11329 6352 13876 6354
rect 11329 6296 11334 6352
rect 11390 6296 12806 6352
rect 12862 6296 13876 6352
rect 11329 6294 13876 6296
rect 11329 6291 11395 6294
rect 12801 6291 12867 6294
rect 2405 6218 2471 6221
rect 5349 6218 5415 6221
rect 2405 6216 5415 6218
rect 2405 6160 2410 6216
rect 2466 6160 5354 6216
rect 5410 6160 5415 6216
rect 2405 6158 5415 6160
rect 2405 6155 2471 6158
rect 5349 6155 5415 6158
rect 10726 6156 10732 6220
rect 10796 6218 10802 6220
rect 11237 6218 11303 6221
rect 13629 6218 13695 6221
rect 10796 6216 13695 6218
rect 10796 6160 11242 6216
rect 11298 6160 13634 6216
rect 13690 6160 13695 6216
rect 10796 6158 13695 6160
rect 13816 6218 13876 6294
rect 14917 6218 14983 6221
rect 13816 6216 14983 6218
rect 13816 6160 14922 6216
rect 14978 6160 14983 6216
rect 13816 6158 14983 6160
rect 10796 6156 10802 6158
rect 11237 6155 11303 6158
rect 13629 6155 13695 6158
rect 14917 6155 14983 6158
rect 18505 6218 18571 6221
rect 19200 6218 20000 6248
rect 18505 6216 20000 6218
rect 18505 6160 18510 6216
rect 18566 6160 20000 6216
rect 18505 6158 20000 6160
rect 18505 6155 18571 6158
rect 19200 6128 20000 6158
rect 0 6082 800 6112
rect 3785 6082 3851 6085
rect 13445 6084 13511 6085
rect 13445 6082 13492 6084
rect 0 6080 3851 6082
rect 0 6024 3790 6080
rect 3846 6024 3851 6080
rect 0 6022 3851 6024
rect 13400 6080 13492 6082
rect 13400 6024 13450 6080
rect 13400 6022 13492 6024
rect 0 5992 800 6022
rect 3785 6019 3851 6022
rect 13445 6020 13492 6022
rect 13556 6020 13562 6084
rect 13629 6082 13695 6085
rect 14038 6082 14044 6084
rect 13629 6080 14044 6082
rect 13629 6024 13634 6080
rect 13690 6024 14044 6080
rect 13629 6022 14044 6024
rect 13445 6019 13511 6020
rect 13629 6019 13695 6022
rect 14038 6020 14044 6022
rect 14108 6020 14114 6084
rect 6874 6016 7194 6017
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7194 6016
rect 6874 5951 7194 5952
rect 12805 6016 13125 6017
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 12805 5951 13125 5952
rect 2957 5946 3023 5949
rect 3417 5946 3483 5949
rect 2957 5944 3483 5946
rect 2957 5888 2962 5944
rect 3018 5888 3422 5944
rect 3478 5888 3483 5944
rect 2957 5886 3483 5888
rect 2957 5883 3023 5886
rect 3417 5883 3483 5886
rect 18505 5946 18571 5949
rect 19200 5946 20000 5976
rect 18505 5944 20000 5946
rect 18505 5888 18510 5944
rect 18566 5888 20000 5944
rect 18505 5886 20000 5888
rect 18505 5883 18571 5886
rect 19200 5856 20000 5886
rect 0 5810 800 5840
rect 1669 5810 1735 5813
rect 0 5808 1735 5810
rect 0 5752 1674 5808
rect 1730 5752 1735 5808
rect 0 5750 1735 5752
rect 0 5720 800 5750
rect 1669 5747 1735 5750
rect 2313 5810 2379 5813
rect 3049 5810 3115 5813
rect 2313 5808 3115 5810
rect 2313 5752 2318 5808
rect 2374 5752 3054 5808
rect 3110 5752 3115 5808
rect 2313 5750 3115 5752
rect 2313 5747 2379 5750
rect 3049 5747 3115 5750
rect 2681 5674 2747 5677
rect 4245 5674 4311 5677
rect 2681 5672 4311 5674
rect 2681 5616 2686 5672
rect 2742 5616 4250 5672
rect 4306 5616 4311 5672
rect 2681 5614 4311 5616
rect 2681 5611 2747 5614
rect 4245 5611 4311 5614
rect 7465 5674 7531 5677
rect 10910 5674 10916 5676
rect 7465 5672 10916 5674
rect 7465 5616 7470 5672
rect 7526 5616 10916 5672
rect 7465 5614 10916 5616
rect 7465 5611 7531 5614
rect 10910 5612 10916 5614
rect 10980 5612 10986 5676
rect 15193 5674 15259 5677
rect 15193 5672 15578 5674
rect 15193 5616 15198 5672
rect 15254 5616 15578 5672
rect 15193 5614 15578 5616
rect 15193 5611 15259 5614
rect 2865 5538 2931 5541
rect 3417 5538 3483 5541
rect 2865 5536 3483 5538
rect 2865 5480 2870 5536
rect 2926 5480 3422 5536
rect 3478 5480 3483 5536
rect 2865 5478 3483 5480
rect 2865 5475 2931 5478
rect 3417 5475 3483 5478
rect 3909 5472 4229 5473
rect 0 5402 800 5432
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 5407 4229 5408
rect 9840 5472 10160 5473
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 5407 10160 5408
rect 2405 5402 2471 5405
rect 0 5400 2471 5402
rect 0 5344 2410 5400
rect 2466 5344 2471 5400
rect 0 5342 2471 5344
rect 0 5312 800 5342
rect 2405 5339 2471 5342
rect 2037 5266 2103 5269
rect 7097 5266 7163 5269
rect 8017 5266 8083 5269
rect 2037 5264 8083 5266
rect 2037 5208 2042 5264
rect 2098 5208 7102 5264
rect 7158 5208 8022 5264
rect 8078 5208 8083 5264
rect 2037 5206 8083 5208
rect 2037 5203 2103 5206
rect 0 5130 800 5160
rect 6732 5133 6792 5206
rect 7097 5203 7163 5206
rect 8017 5203 8083 5206
rect 11973 5266 12039 5269
rect 15518 5266 15578 5614
rect 17861 5538 17927 5541
rect 19200 5538 20000 5568
rect 17861 5536 20000 5538
rect 17861 5480 17866 5536
rect 17922 5480 20000 5536
rect 17861 5478 20000 5480
rect 17861 5475 17927 5478
rect 15770 5472 16090 5473
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16090 5472
rect 19200 5448 20000 5478
rect 15770 5407 16090 5408
rect 15745 5266 15811 5269
rect 11973 5264 13370 5266
rect 11973 5208 11978 5264
rect 12034 5208 13370 5264
rect 11973 5206 13370 5208
rect 15518 5264 15811 5266
rect 15518 5208 15750 5264
rect 15806 5208 15811 5264
rect 15518 5206 15811 5208
rect 11973 5203 12039 5206
rect 3877 5130 3943 5133
rect 6453 5132 6519 5133
rect 6453 5130 6500 5132
rect 0 5128 3943 5130
rect 0 5072 3882 5128
rect 3938 5072 3943 5128
rect 0 5070 3943 5072
rect 6408 5128 6500 5130
rect 6408 5072 6458 5128
rect 6408 5070 6500 5072
rect 0 5040 800 5070
rect 3877 5067 3943 5070
rect 6453 5068 6500 5070
rect 6564 5068 6570 5132
rect 6729 5128 6795 5133
rect 6729 5072 6734 5128
rect 6790 5072 6795 5128
rect 6453 5067 6519 5068
rect 6729 5067 6795 5072
rect 8017 5130 8083 5133
rect 13169 5130 13235 5133
rect 8017 5128 13235 5130
rect 8017 5072 8022 5128
rect 8078 5072 13174 5128
rect 13230 5072 13235 5128
rect 8017 5070 13235 5072
rect 13310 5130 13370 5206
rect 15745 5203 15811 5206
rect 15929 5130 15995 5133
rect 13310 5128 15995 5130
rect 13310 5072 15934 5128
rect 15990 5072 15995 5128
rect 13310 5070 15995 5072
rect 8017 5067 8083 5070
rect 13169 5067 13235 5070
rect 15929 5067 15995 5070
rect 18505 5130 18571 5133
rect 19200 5130 20000 5160
rect 18505 5128 20000 5130
rect 18505 5072 18510 5128
rect 18566 5072 20000 5128
rect 18505 5070 20000 5072
rect 18505 5067 18571 5070
rect 19200 5040 20000 5070
rect 6874 4928 7194 4929
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7194 4928
rect 6874 4863 7194 4864
rect 12805 4928 13125 4929
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12805 4863 13125 4864
rect 14549 4858 14615 4861
rect 15653 4858 15719 4861
rect 14549 4856 15719 4858
rect 14549 4800 14554 4856
rect 14610 4800 15658 4856
rect 15714 4800 15719 4856
rect 14549 4798 15719 4800
rect 14549 4795 14615 4798
rect 15653 4795 15719 4798
rect 0 4722 800 4752
rect 1393 4722 1459 4725
rect 0 4720 1459 4722
rect 0 4664 1398 4720
rect 1454 4664 1459 4720
rect 0 4662 1459 4664
rect 0 4632 800 4662
rect 1393 4659 1459 4662
rect 1577 4722 1643 4725
rect 5349 4722 5415 4725
rect 1577 4720 5415 4722
rect 1577 4664 1582 4720
rect 1638 4664 5354 4720
rect 5410 4664 5415 4720
rect 1577 4662 5415 4664
rect 1577 4659 1643 4662
rect 5349 4659 5415 4662
rect 8569 4722 8635 4725
rect 9397 4722 9463 4725
rect 8569 4720 9463 4722
rect 8569 4664 8574 4720
rect 8630 4664 9402 4720
rect 9458 4664 9463 4720
rect 8569 4662 9463 4664
rect 8569 4659 8635 4662
rect 9397 4659 9463 4662
rect 10910 4660 10916 4724
rect 10980 4722 10986 4724
rect 13077 4722 13143 4725
rect 10980 4720 13143 4722
rect 10980 4664 13082 4720
rect 13138 4664 13143 4720
rect 10980 4662 13143 4664
rect 10980 4660 10986 4662
rect 13077 4659 13143 4662
rect 18505 4722 18571 4725
rect 19200 4722 20000 4752
rect 18505 4720 20000 4722
rect 18505 4664 18510 4720
rect 18566 4664 20000 4720
rect 18505 4662 20000 4664
rect 18505 4659 18571 4662
rect 19200 4632 20000 4662
rect 2589 4586 2655 4589
rect 5993 4586 6059 4589
rect 2589 4584 6059 4586
rect 2589 4528 2594 4584
rect 2650 4528 5998 4584
rect 6054 4528 6059 4584
rect 2589 4526 6059 4528
rect 2589 4523 2655 4526
rect 5993 4523 6059 4526
rect 6361 4586 6427 4589
rect 14365 4586 14431 4589
rect 6361 4584 14431 4586
rect 6361 4528 6366 4584
rect 6422 4528 14370 4584
rect 14426 4528 14431 4584
rect 6361 4526 14431 4528
rect 6361 4523 6427 4526
rect 14365 4523 14431 4526
rect 0 4450 800 4480
rect 2129 4450 2195 4453
rect 0 4448 2195 4450
rect 0 4392 2134 4448
rect 2190 4392 2195 4448
rect 0 4390 2195 4392
rect 0 4360 800 4390
rect 2129 4387 2195 4390
rect 5257 4450 5323 4453
rect 5809 4450 5875 4453
rect 5257 4448 5875 4450
rect 5257 4392 5262 4448
rect 5318 4392 5814 4448
rect 5870 4392 5875 4448
rect 5257 4390 5875 4392
rect 5257 4387 5323 4390
rect 5809 4387 5875 4390
rect 6126 4388 6132 4452
rect 6196 4450 6202 4452
rect 6269 4450 6335 4453
rect 6196 4448 6335 4450
rect 6196 4392 6274 4448
rect 6330 4392 6335 4448
rect 6196 4390 6335 4392
rect 6196 4388 6202 4390
rect 6269 4387 6335 4390
rect 6545 4450 6611 4453
rect 9213 4450 9279 4453
rect 6545 4448 9279 4450
rect 6545 4392 6550 4448
rect 6606 4392 9218 4448
rect 9274 4392 9279 4448
rect 6545 4390 9279 4392
rect 6545 4387 6611 4390
rect 9213 4387 9279 4390
rect 10317 4450 10383 4453
rect 12525 4452 12591 4453
rect 12525 4450 12572 4452
rect 10317 4448 12572 4450
rect 12636 4450 12642 4452
rect 10317 4392 10322 4448
rect 10378 4392 12530 4448
rect 10317 4390 12572 4392
rect 10317 4387 10383 4390
rect 12525 4388 12572 4390
rect 12636 4390 12718 4450
rect 12636 4388 12642 4390
rect 12525 4387 12591 4388
rect 3909 4384 4229 4385
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 4319 4229 4320
rect 9840 4384 10160 4385
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 4319 10160 4320
rect 15770 4384 16090 4385
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16090 4384
rect 15770 4319 16090 4320
rect 18137 4314 18203 4317
rect 19200 4314 20000 4344
rect 18137 4312 20000 4314
rect 18137 4256 18142 4312
rect 18198 4256 20000 4312
rect 18137 4254 20000 4256
rect 18137 4251 18203 4254
rect 19200 4224 20000 4254
rect 0 4178 800 4208
rect 1485 4178 1551 4181
rect 0 4176 1551 4178
rect 0 4120 1490 4176
rect 1546 4120 1551 4176
rect 0 4118 1551 4120
rect 0 4088 800 4118
rect 1485 4115 1551 4118
rect 3049 4178 3115 4181
rect 6729 4178 6795 4181
rect 3049 4176 6795 4178
rect 3049 4120 3054 4176
rect 3110 4120 6734 4176
rect 6790 4120 6795 4176
rect 3049 4118 6795 4120
rect 3049 4115 3115 4118
rect 6729 4115 6795 4118
rect 7649 4178 7715 4181
rect 11697 4178 11763 4181
rect 7649 4176 11763 4178
rect 7649 4120 7654 4176
rect 7710 4120 11702 4176
rect 11758 4120 11763 4176
rect 7649 4118 11763 4120
rect 7649 4115 7715 4118
rect 11697 4115 11763 4118
rect 12341 4178 12407 4181
rect 14365 4178 14431 4181
rect 12341 4176 14431 4178
rect 12341 4120 12346 4176
rect 12402 4120 14370 4176
rect 14426 4120 14431 4176
rect 12341 4118 14431 4120
rect 12341 4115 12407 4118
rect 14365 4115 14431 4118
rect 2589 4042 2655 4045
rect 4613 4042 4679 4045
rect 2589 4040 4679 4042
rect 2589 3984 2594 4040
rect 2650 3984 4618 4040
rect 4674 3984 4679 4040
rect 2589 3982 4679 3984
rect 2589 3979 2655 3982
rect 4613 3979 4679 3982
rect 10869 4042 10935 4045
rect 14549 4042 14615 4045
rect 10869 4040 14615 4042
rect 10869 3984 10874 4040
rect 10930 3984 14554 4040
rect 14610 3984 14615 4040
rect 10869 3982 14615 3984
rect 10869 3979 10935 3982
rect 14549 3979 14615 3982
rect 18505 4042 18571 4045
rect 19200 4042 20000 4072
rect 18505 4040 20000 4042
rect 18505 3984 18510 4040
rect 18566 3984 20000 4040
rect 18505 3982 20000 3984
rect 18505 3979 18571 3982
rect 19200 3952 20000 3982
rect 2957 3906 3023 3909
rect 4153 3906 4219 3909
rect 2957 3904 4219 3906
rect 2957 3848 2962 3904
rect 3018 3848 4158 3904
rect 4214 3848 4219 3904
rect 2957 3846 4219 3848
rect 2957 3843 3023 3846
rect 4153 3843 4219 3846
rect 4470 3844 4476 3908
rect 4540 3906 4546 3908
rect 4613 3906 4679 3909
rect 4540 3904 4679 3906
rect 4540 3848 4618 3904
rect 4674 3848 4679 3904
rect 4540 3846 4679 3848
rect 4540 3844 4546 3846
rect 4613 3843 4679 3846
rect 6874 3840 7194 3841
rect 0 3770 800 3800
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7194 3840
rect 6874 3775 7194 3776
rect 12805 3840 13125 3841
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 3775 13125 3776
rect 1853 3770 1919 3773
rect 0 3768 1919 3770
rect 0 3712 1858 3768
rect 1914 3712 1919 3768
rect 0 3710 1919 3712
rect 0 3680 800 3710
rect 1853 3707 1919 3710
rect 16113 3770 16179 3773
rect 16113 3768 16498 3770
rect 16113 3712 16118 3768
rect 16174 3712 16498 3768
rect 16113 3710 16498 3712
rect 16113 3707 16179 3710
rect 16438 3637 16498 3710
rect 8109 3634 8175 3637
rect 9213 3634 9279 3637
rect 8109 3632 9279 3634
rect 8109 3576 8114 3632
rect 8170 3576 9218 3632
rect 9274 3576 9279 3632
rect 8109 3574 9279 3576
rect 16438 3632 16547 3637
rect 16438 3576 16486 3632
rect 16542 3576 16547 3632
rect 16438 3574 16547 3576
rect 8109 3571 8175 3574
rect 9213 3571 9279 3574
rect 16481 3571 16547 3574
rect 18137 3634 18203 3637
rect 19200 3634 20000 3664
rect 18137 3632 20000 3634
rect 18137 3576 18142 3632
rect 18198 3576 20000 3632
rect 18137 3574 20000 3576
rect 18137 3571 18203 3574
rect 19200 3544 20000 3574
rect 0 3498 800 3528
rect 1485 3498 1551 3501
rect 0 3496 1551 3498
rect 0 3440 1490 3496
rect 1546 3440 1551 3496
rect 0 3438 1551 3440
rect 0 3408 800 3438
rect 1485 3435 1551 3438
rect 3693 3498 3759 3501
rect 5165 3498 5231 3501
rect 3693 3496 5231 3498
rect 3693 3440 3698 3496
rect 3754 3440 5170 3496
rect 5226 3440 5231 3496
rect 3693 3438 5231 3440
rect 3693 3435 3759 3438
rect 5165 3435 5231 3438
rect 10961 3498 11027 3501
rect 12433 3498 12499 3501
rect 10961 3496 12499 3498
rect 10961 3440 10966 3496
rect 11022 3440 12438 3496
rect 12494 3440 12499 3496
rect 10961 3438 12499 3440
rect 10961 3435 11027 3438
rect 12433 3435 12499 3438
rect 3909 3296 4229 3297
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 3231 4229 3232
rect 9840 3296 10160 3297
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 3231 10160 3232
rect 15770 3296 16090 3297
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16090 3296
rect 15770 3231 16090 3232
rect 18505 3226 18571 3229
rect 19200 3226 20000 3256
rect 18505 3224 20000 3226
rect 18505 3168 18510 3224
rect 18566 3168 20000 3224
rect 18505 3166 20000 3168
rect 18505 3163 18571 3166
rect 19200 3136 20000 3166
rect 0 3090 800 3120
rect 3417 3090 3483 3093
rect 0 3088 3483 3090
rect 0 3032 3422 3088
rect 3478 3032 3483 3088
rect 0 3030 3483 3032
rect 0 3000 800 3030
rect 3417 3027 3483 3030
rect 5625 3090 5691 3093
rect 6494 3090 6500 3092
rect 5625 3088 6500 3090
rect 5625 3032 5630 3088
rect 5686 3032 6500 3088
rect 5625 3030 6500 3032
rect 5625 3027 5691 3030
rect 6494 3028 6500 3030
rect 6564 3090 6570 3092
rect 11881 3090 11947 3093
rect 6564 3088 11947 3090
rect 6564 3032 11886 3088
rect 11942 3032 11947 3088
rect 6564 3030 11947 3032
rect 6564 3028 6570 3030
rect 11881 3027 11947 3030
rect 2313 2954 2379 2957
rect 6085 2954 6151 2957
rect 2313 2952 6151 2954
rect 2313 2896 2318 2952
rect 2374 2896 6090 2952
rect 6146 2896 6151 2952
rect 2313 2894 6151 2896
rect 2313 2891 2379 2894
rect 6085 2891 6151 2894
rect 6729 2954 6795 2957
rect 14365 2954 14431 2957
rect 6729 2952 14431 2954
rect 6729 2896 6734 2952
rect 6790 2896 14370 2952
rect 14426 2896 14431 2952
rect 6729 2894 14431 2896
rect 6729 2891 6795 2894
rect 14365 2891 14431 2894
rect 0 2818 800 2848
rect 3785 2818 3851 2821
rect 0 2816 3851 2818
rect 0 2760 3790 2816
rect 3846 2760 3851 2816
rect 0 2758 3851 2760
rect 0 2728 800 2758
rect 3785 2755 3851 2758
rect 8845 2818 8911 2821
rect 12341 2818 12407 2821
rect 8845 2816 12407 2818
rect 8845 2760 8850 2816
rect 8906 2760 12346 2816
rect 12402 2760 12407 2816
rect 8845 2758 12407 2760
rect 8845 2755 8911 2758
rect 12341 2755 12407 2758
rect 13997 2818 14063 2821
rect 14457 2818 14523 2821
rect 13997 2816 14523 2818
rect 13997 2760 14002 2816
rect 14058 2760 14462 2816
rect 14518 2760 14523 2816
rect 13997 2758 14523 2760
rect 13997 2755 14063 2758
rect 14457 2755 14523 2758
rect 18137 2818 18203 2821
rect 19200 2818 20000 2848
rect 18137 2816 20000 2818
rect 18137 2760 18142 2816
rect 18198 2760 20000 2816
rect 18137 2758 20000 2760
rect 18137 2755 18203 2758
rect 6874 2752 7194 2753
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7194 2752
rect 6874 2687 7194 2688
rect 12805 2752 13125 2753
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 19200 2728 20000 2758
rect 12805 2687 13125 2688
rect 2681 2682 2747 2685
rect 6453 2682 6519 2685
rect 2681 2680 6519 2682
rect 2681 2624 2686 2680
rect 2742 2624 6458 2680
rect 6514 2624 6519 2680
rect 2681 2622 6519 2624
rect 2681 2619 2747 2622
rect 6453 2619 6519 2622
rect 9622 2620 9628 2684
rect 9692 2682 9698 2684
rect 9949 2682 10015 2685
rect 9692 2680 10015 2682
rect 9692 2624 9954 2680
rect 10010 2624 10015 2680
rect 9692 2622 10015 2624
rect 9692 2620 9698 2622
rect 9949 2619 10015 2622
rect 16849 2682 16915 2685
rect 17769 2684 17835 2685
rect 16982 2682 16988 2684
rect 16849 2680 16988 2682
rect 16849 2624 16854 2680
rect 16910 2624 16988 2680
rect 16849 2622 16988 2624
rect 16849 2619 16915 2622
rect 16982 2620 16988 2622
rect 17052 2620 17058 2684
rect 17718 2682 17724 2684
rect 17678 2622 17724 2682
rect 17788 2680 17835 2684
rect 17830 2624 17835 2680
rect 17718 2620 17724 2622
rect 17788 2620 17835 2624
rect 17769 2619 17835 2620
rect 4838 2484 4844 2548
rect 4908 2546 4914 2548
rect 8293 2546 8359 2549
rect 4908 2544 8359 2546
rect 4908 2488 8298 2544
rect 8354 2488 8359 2544
rect 4908 2486 8359 2488
rect 4908 2484 4914 2486
rect 8293 2483 8359 2486
rect 10593 2546 10659 2549
rect 10726 2546 10732 2548
rect 10593 2544 10732 2546
rect 10593 2488 10598 2544
rect 10654 2488 10732 2544
rect 10593 2486 10732 2488
rect 10593 2483 10659 2486
rect 10726 2484 10732 2486
rect 10796 2484 10802 2548
rect 0 2410 800 2440
rect 3693 2410 3759 2413
rect 0 2408 3759 2410
rect 0 2352 3698 2408
rect 3754 2352 3759 2408
rect 0 2350 3759 2352
rect 0 2320 800 2350
rect 3693 2347 3759 2350
rect 18413 2410 18479 2413
rect 19200 2410 20000 2440
rect 18413 2408 20000 2410
rect 18413 2352 18418 2408
rect 18474 2352 20000 2408
rect 18413 2350 20000 2352
rect 18413 2347 18479 2350
rect 19200 2320 20000 2350
rect 3909 2208 4229 2209
rect 0 2138 800 2168
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2143 4229 2144
rect 9840 2208 10160 2209
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2143 10160 2144
rect 15770 2208 16090 2209
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16090 2208
rect 15770 2143 16090 2144
rect 3325 2138 3391 2141
rect 0 2136 3391 2138
rect 0 2080 3330 2136
rect 3386 2080 3391 2136
rect 0 2078 3391 2080
rect 0 2048 800 2078
rect 3325 2075 3391 2078
rect 18505 2138 18571 2141
rect 19200 2138 20000 2168
rect 18505 2136 20000 2138
rect 18505 2080 18510 2136
rect 18566 2080 20000 2136
rect 18505 2078 20000 2080
rect 18505 2075 18571 2078
rect 19200 2048 20000 2078
rect 0 1866 800 1896
rect 3233 1866 3299 1869
rect 0 1864 3299 1866
rect 0 1808 3238 1864
rect 3294 1808 3299 1864
rect 0 1806 3299 1808
rect 0 1776 800 1806
rect 3233 1803 3299 1806
rect 17861 1730 17927 1733
rect 19200 1730 20000 1760
rect 17861 1728 20000 1730
rect 17861 1672 17866 1728
rect 17922 1672 20000 1728
rect 17861 1670 20000 1672
rect 17861 1667 17927 1670
rect 19200 1640 20000 1670
rect 0 1458 800 1488
rect 3141 1458 3207 1461
rect 0 1456 3207 1458
rect 0 1400 3146 1456
rect 3202 1400 3207 1456
rect 0 1398 3207 1400
rect 0 1368 800 1398
rect 3141 1395 3207 1398
rect 17033 1322 17099 1325
rect 19200 1322 20000 1352
rect 17033 1320 20000 1322
rect 17033 1264 17038 1320
rect 17094 1264 20000 1320
rect 17033 1262 20000 1264
rect 17033 1259 17099 1262
rect 19200 1232 20000 1262
rect 0 1186 800 1216
rect 2957 1186 3023 1189
rect 0 1184 3023 1186
rect 0 1128 2962 1184
rect 3018 1128 3023 1184
rect 0 1126 3023 1128
rect 0 1096 800 1126
rect 2957 1123 3023 1126
rect 16849 914 16915 917
rect 19200 914 20000 944
rect 16849 912 20000 914
rect 16849 856 16854 912
rect 16910 856 20000 912
rect 16849 854 20000 856
rect 16849 851 16915 854
rect 19200 824 20000 854
rect 0 778 800 808
rect 3417 778 3483 781
rect 0 776 3483 778
rect 0 720 3422 776
rect 3478 720 3483 776
rect 0 718 3483 720
rect 0 688 800 718
rect 3417 715 3483 718
rect 0 506 800 536
rect 2865 506 2931 509
rect 0 504 2931 506
rect 0 448 2870 504
rect 2926 448 2931 504
rect 0 446 2931 448
rect 0 416 800 446
rect 2865 443 2931 446
rect 16481 506 16547 509
rect 19200 506 20000 536
rect 16481 504 20000 506
rect 16481 448 16486 504
rect 16542 448 20000 504
rect 16481 446 20000 448
rect 16481 443 16547 446
rect 19200 416 20000 446
rect 0 234 800 264
rect 2773 234 2839 237
rect 0 232 2839 234
rect 0 176 2778 232
rect 2834 176 2839 232
rect 0 174 2839 176
rect 0 144 800 174
rect 2773 171 2839 174
rect 15469 234 15535 237
rect 19200 234 20000 264
rect 15469 232 20000 234
rect 15469 176 15474 232
rect 15530 176 20000 232
rect 15469 174 20000 176
rect 15469 171 15535 174
rect 19200 144 20000 174
<< via3 >>
rect 6882 14716 6946 14720
rect 6882 14660 6886 14716
rect 6886 14660 6942 14716
rect 6942 14660 6946 14716
rect 6882 14656 6946 14660
rect 6962 14716 7026 14720
rect 6962 14660 6966 14716
rect 6966 14660 7022 14716
rect 7022 14660 7026 14716
rect 6962 14656 7026 14660
rect 7042 14716 7106 14720
rect 7042 14660 7046 14716
rect 7046 14660 7102 14716
rect 7102 14660 7106 14716
rect 7042 14656 7106 14660
rect 7122 14716 7186 14720
rect 7122 14660 7126 14716
rect 7126 14660 7182 14716
rect 7182 14660 7186 14716
rect 7122 14656 7186 14660
rect 12813 14716 12877 14720
rect 12813 14660 12817 14716
rect 12817 14660 12873 14716
rect 12873 14660 12877 14716
rect 12813 14656 12877 14660
rect 12893 14716 12957 14720
rect 12893 14660 12897 14716
rect 12897 14660 12953 14716
rect 12953 14660 12957 14716
rect 12893 14656 12957 14660
rect 12973 14716 13037 14720
rect 12973 14660 12977 14716
rect 12977 14660 13033 14716
rect 13033 14660 13037 14716
rect 12973 14656 13037 14660
rect 13053 14716 13117 14720
rect 13053 14660 13057 14716
rect 13057 14660 13113 14716
rect 13113 14660 13117 14716
rect 13053 14656 13117 14660
rect 3917 14172 3981 14176
rect 3917 14116 3921 14172
rect 3921 14116 3977 14172
rect 3977 14116 3981 14172
rect 3917 14112 3981 14116
rect 3997 14172 4061 14176
rect 3997 14116 4001 14172
rect 4001 14116 4057 14172
rect 4057 14116 4061 14172
rect 3997 14112 4061 14116
rect 4077 14172 4141 14176
rect 4077 14116 4081 14172
rect 4081 14116 4137 14172
rect 4137 14116 4141 14172
rect 4077 14112 4141 14116
rect 4157 14172 4221 14176
rect 4157 14116 4161 14172
rect 4161 14116 4217 14172
rect 4217 14116 4221 14172
rect 4157 14112 4221 14116
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 15778 14172 15842 14176
rect 15778 14116 15782 14172
rect 15782 14116 15838 14172
rect 15838 14116 15842 14172
rect 15778 14112 15842 14116
rect 15858 14172 15922 14176
rect 15858 14116 15862 14172
rect 15862 14116 15918 14172
rect 15918 14116 15922 14172
rect 15858 14112 15922 14116
rect 15938 14172 16002 14176
rect 15938 14116 15942 14172
rect 15942 14116 15998 14172
rect 15998 14116 16002 14172
rect 15938 14112 16002 14116
rect 16018 14172 16082 14176
rect 16018 14116 16022 14172
rect 16022 14116 16078 14172
rect 16078 14116 16082 14172
rect 16018 14112 16082 14116
rect 17724 13772 17788 13836
rect 6882 13628 6946 13632
rect 6882 13572 6886 13628
rect 6886 13572 6942 13628
rect 6942 13572 6946 13628
rect 6882 13568 6946 13572
rect 6962 13628 7026 13632
rect 6962 13572 6966 13628
rect 6966 13572 7022 13628
rect 7022 13572 7026 13628
rect 6962 13568 7026 13572
rect 7042 13628 7106 13632
rect 7042 13572 7046 13628
rect 7046 13572 7102 13628
rect 7102 13572 7106 13628
rect 7042 13568 7106 13572
rect 7122 13628 7186 13632
rect 7122 13572 7126 13628
rect 7126 13572 7182 13628
rect 7182 13572 7186 13628
rect 7122 13568 7186 13572
rect 12813 13628 12877 13632
rect 12813 13572 12817 13628
rect 12817 13572 12873 13628
rect 12873 13572 12877 13628
rect 12813 13568 12877 13572
rect 12893 13628 12957 13632
rect 12893 13572 12897 13628
rect 12897 13572 12953 13628
rect 12953 13572 12957 13628
rect 12893 13568 12957 13572
rect 12973 13628 13037 13632
rect 12973 13572 12977 13628
rect 12977 13572 13033 13628
rect 13033 13572 13037 13628
rect 12973 13568 13037 13572
rect 13053 13628 13117 13632
rect 13053 13572 13057 13628
rect 13057 13572 13113 13628
rect 13113 13572 13117 13628
rect 13053 13568 13117 13572
rect 3917 13084 3981 13088
rect 3917 13028 3921 13084
rect 3921 13028 3977 13084
rect 3977 13028 3981 13084
rect 3917 13024 3981 13028
rect 3997 13084 4061 13088
rect 3997 13028 4001 13084
rect 4001 13028 4057 13084
rect 4057 13028 4061 13084
rect 3997 13024 4061 13028
rect 4077 13084 4141 13088
rect 4077 13028 4081 13084
rect 4081 13028 4137 13084
rect 4137 13028 4141 13084
rect 4077 13024 4141 13028
rect 4157 13084 4221 13088
rect 4157 13028 4161 13084
rect 4161 13028 4217 13084
rect 4217 13028 4221 13084
rect 4157 13024 4221 13028
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 15778 13084 15842 13088
rect 15778 13028 15782 13084
rect 15782 13028 15838 13084
rect 15838 13028 15842 13084
rect 15778 13024 15842 13028
rect 15858 13084 15922 13088
rect 15858 13028 15862 13084
rect 15862 13028 15918 13084
rect 15918 13028 15922 13084
rect 15858 13024 15922 13028
rect 15938 13084 16002 13088
rect 15938 13028 15942 13084
rect 15942 13028 15998 13084
rect 15998 13028 16002 13084
rect 15938 13024 16002 13028
rect 16018 13084 16082 13088
rect 16018 13028 16022 13084
rect 16022 13028 16078 13084
rect 16078 13028 16082 13084
rect 16018 13024 16082 13028
rect 16988 12820 17052 12884
rect 9628 12684 9692 12748
rect 6882 12540 6946 12544
rect 6882 12484 6886 12540
rect 6886 12484 6942 12540
rect 6942 12484 6946 12540
rect 6882 12480 6946 12484
rect 6962 12540 7026 12544
rect 6962 12484 6966 12540
rect 6966 12484 7022 12540
rect 7022 12484 7026 12540
rect 6962 12480 7026 12484
rect 7042 12540 7106 12544
rect 7042 12484 7046 12540
rect 7046 12484 7102 12540
rect 7102 12484 7106 12540
rect 7042 12480 7106 12484
rect 7122 12540 7186 12544
rect 7122 12484 7126 12540
rect 7126 12484 7182 12540
rect 7182 12484 7186 12540
rect 7122 12480 7186 12484
rect 12813 12540 12877 12544
rect 12813 12484 12817 12540
rect 12817 12484 12873 12540
rect 12873 12484 12877 12540
rect 12813 12480 12877 12484
rect 12893 12540 12957 12544
rect 12893 12484 12897 12540
rect 12897 12484 12953 12540
rect 12953 12484 12957 12540
rect 12893 12480 12957 12484
rect 12973 12540 13037 12544
rect 12973 12484 12977 12540
rect 12977 12484 13033 12540
rect 13033 12484 13037 12540
rect 12973 12480 13037 12484
rect 13053 12540 13117 12544
rect 13053 12484 13057 12540
rect 13057 12484 13113 12540
rect 13113 12484 13117 12540
rect 13053 12480 13117 12484
rect 3917 11996 3981 12000
rect 3917 11940 3921 11996
rect 3921 11940 3977 11996
rect 3977 11940 3981 11996
rect 3917 11936 3981 11940
rect 3997 11996 4061 12000
rect 3997 11940 4001 11996
rect 4001 11940 4057 11996
rect 4057 11940 4061 11996
rect 3997 11936 4061 11940
rect 4077 11996 4141 12000
rect 4077 11940 4081 11996
rect 4081 11940 4137 11996
rect 4137 11940 4141 11996
rect 4077 11936 4141 11940
rect 4157 11996 4221 12000
rect 4157 11940 4161 11996
rect 4161 11940 4217 11996
rect 4217 11940 4221 11996
rect 4157 11936 4221 11940
rect 9628 12004 9692 12068
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 15778 11996 15842 12000
rect 15778 11940 15782 11996
rect 15782 11940 15838 11996
rect 15838 11940 15842 11996
rect 15778 11936 15842 11940
rect 15858 11996 15922 12000
rect 15858 11940 15862 11996
rect 15862 11940 15918 11996
rect 15918 11940 15922 11996
rect 15858 11936 15922 11940
rect 15938 11996 16002 12000
rect 15938 11940 15942 11996
rect 15942 11940 15998 11996
rect 15998 11940 16002 11996
rect 15938 11936 16002 11940
rect 16018 11996 16082 12000
rect 16018 11940 16022 11996
rect 16022 11940 16078 11996
rect 16078 11940 16082 11996
rect 16018 11936 16082 11940
rect 16252 11596 16316 11660
rect 16436 11520 16500 11524
rect 16436 11464 16450 11520
rect 16450 11464 16500 11520
rect 16436 11460 16500 11464
rect 6882 11452 6946 11456
rect 6882 11396 6886 11452
rect 6886 11396 6942 11452
rect 6942 11396 6946 11452
rect 6882 11392 6946 11396
rect 6962 11452 7026 11456
rect 6962 11396 6966 11452
rect 6966 11396 7022 11452
rect 7022 11396 7026 11452
rect 6962 11392 7026 11396
rect 7042 11452 7106 11456
rect 7042 11396 7046 11452
rect 7046 11396 7102 11452
rect 7102 11396 7106 11452
rect 7042 11392 7106 11396
rect 7122 11452 7186 11456
rect 7122 11396 7126 11452
rect 7126 11396 7182 11452
rect 7182 11396 7186 11452
rect 7122 11392 7186 11396
rect 12813 11452 12877 11456
rect 12813 11396 12817 11452
rect 12817 11396 12873 11452
rect 12873 11396 12877 11452
rect 12813 11392 12877 11396
rect 12893 11452 12957 11456
rect 12893 11396 12897 11452
rect 12897 11396 12953 11452
rect 12953 11396 12957 11452
rect 12893 11392 12957 11396
rect 12973 11452 13037 11456
rect 12973 11396 12977 11452
rect 12977 11396 13033 11452
rect 13033 11396 13037 11452
rect 12973 11392 13037 11396
rect 13053 11452 13117 11456
rect 13053 11396 13057 11452
rect 13057 11396 13113 11452
rect 13113 11396 13117 11452
rect 13053 11392 13117 11396
rect 3917 10908 3981 10912
rect 3917 10852 3921 10908
rect 3921 10852 3977 10908
rect 3977 10852 3981 10908
rect 3917 10848 3981 10852
rect 3997 10908 4061 10912
rect 3997 10852 4001 10908
rect 4001 10852 4057 10908
rect 4057 10852 4061 10908
rect 3997 10848 4061 10852
rect 4077 10908 4141 10912
rect 4077 10852 4081 10908
rect 4081 10852 4137 10908
rect 4137 10852 4141 10908
rect 4077 10848 4141 10852
rect 4157 10908 4221 10912
rect 4157 10852 4161 10908
rect 4161 10852 4217 10908
rect 4217 10852 4221 10908
rect 4157 10848 4221 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 15778 10908 15842 10912
rect 15778 10852 15782 10908
rect 15782 10852 15838 10908
rect 15838 10852 15842 10908
rect 15778 10848 15842 10852
rect 15858 10908 15922 10912
rect 15858 10852 15862 10908
rect 15862 10852 15918 10908
rect 15918 10852 15922 10908
rect 15858 10848 15922 10852
rect 15938 10908 16002 10912
rect 15938 10852 15942 10908
rect 15942 10852 15998 10908
rect 15998 10852 16002 10908
rect 15938 10848 16002 10852
rect 16018 10908 16082 10912
rect 16018 10852 16022 10908
rect 16022 10852 16078 10908
rect 16078 10852 16082 10908
rect 16018 10848 16082 10852
rect 6882 10364 6946 10368
rect 6882 10308 6886 10364
rect 6886 10308 6942 10364
rect 6942 10308 6946 10364
rect 6882 10304 6946 10308
rect 6962 10364 7026 10368
rect 6962 10308 6966 10364
rect 6966 10308 7022 10364
rect 7022 10308 7026 10364
rect 6962 10304 7026 10308
rect 7042 10364 7106 10368
rect 7042 10308 7046 10364
rect 7046 10308 7102 10364
rect 7102 10308 7106 10364
rect 7042 10304 7106 10308
rect 7122 10364 7186 10368
rect 7122 10308 7126 10364
rect 7126 10308 7182 10364
rect 7182 10308 7186 10364
rect 7122 10304 7186 10308
rect 12813 10364 12877 10368
rect 12813 10308 12817 10364
rect 12817 10308 12873 10364
rect 12873 10308 12877 10364
rect 12813 10304 12877 10308
rect 12893 10364 12957 10368
rect 12893 10308 12897 10364
rect 12897 10308 12953 10364
rect 12953 10308 12957 10364
rect 12893 10304 12957 10308
rect 12973 10364 13037 10368
rect 12973 10308 12977 10364
rect 12977 10308 13033 10364
rect 13033 10308 13037 10364
rect 12973 10304 13037 10308
rect 13053 10364 13117 10368
rect 13053 10308 13057 10364
rect 13057 10308 13113 10364
rect 13113 10308 13117 10364
rect 13053 10304 13117 10308
rect 3917 9820 3981 9824
rect 3917 9764 3921 9820
rect 3921 9764 3977 9820
rect 3977 9764 3981 9820
rect 3917 9760 3981 9764
rect 3997 9820 4061 9824
rect 3997 9764 4001 9820
rect 4001 9764 4057 9820
rect 4057 9764 4061 9820
rect 3997 9760 4061 9764
rect 4077 9820 4141 9824
rect 4077 9764 4081 9820
rect 4081 9764 4137 9820
rect 4137 9764 4141 9820
rect 4077 9760 4141 9764
rect 4157 9820 4221 9824
rect 4157 9764 4161 9820
rect 4161 9764 4217 9820
rect 4217 9764 4221 9820
rect 4157 9760 4221 9764
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 15778 9820 15842 9824
rect 15778 9764 15782 9820
rect 15782 9764 15838 9820
rect 15838 9764 15842 9820
rect 15778 9760 15842 9764
rect 15858 9820 15922 9824
rect 15858 9764 15862 9820
rect 15862 9764 15918 9820
rect 15918 9764 15922 9820
rect 15858 9760 15922 9764
rect 15938 9820 16002 9824
rect 15938 9764 15942 9820
rect 15942 9764 15998 9820
rect 15998 9764 16002 9820
rect 15938 9760 16002 9764
rect 16018 9820 16082 9824
rect 16018 9764 16022 9820
rect 16022 9764 16078 9820
rect 16078 9764 16082 9820
rect 16018 9760 16082 9764
rect 6132 9752 6196 9756
rect 6132 9696 6182 9752
rect 6182 9696 6196 9752
rect 6132 9692 6196 9696
rect 16436 9692 16500 9756
rect 13308 9420 13372 9484
rect 6882 9276 6946 9280
rect 6882 9220 6886 9276
rect 6886 9220 6942 9276
rect 6942 9220 6946 9276
rect 6882 9216 6946 9220
rect 6962 9276 7026 9280
rect 6962 9220 6966 9276
rect 6966 9220 7022 9276
rect 7022 9220 7026 9276
rect 6962 9216 7026 9220
rect 7042 9276 7106 9280
rect 7042 9220 7046 9276
rect 7046 9220 7102 9276
rect 7102 9220 7106 9276
rect 7042 9216 7106 9220
rect 7122 9276 7186 9280
rect 7122 9220 7126 9276
rect 7126 9220 7182 9276
rect 7182 9220 7186 9276
rect 7122 9216 7186 9220
rect 12813 9276 12877 9280
rect 12813 9220 12817 9276
rect 12817 9220 12873 9276
rect 12873 9220 12877 9276
rect 12813 9216 12877 9220
rect 12893 9276 12957 9280
rect 12893 9220 12897 9276
rect 12897 9220 12953 9276
rect 12953 9220 12957 9276
rect 12893 9216 12957 9220
rect 12973 9276 13037 9280
rect 12973 9220 12977 9276
rect 12977 9220 13033 9276
rect 13033 9220 13037 9276
rect 12973 9216 13037 9220
rect 13053 9276 13117 9280
rect 13053 9220 13057 9276
rect 13057 9220 13113 9276
rect 13113 9220 13117 9276
rect 13053 9216 13117 9220
rect 13492 9148 13556 9212
rect 4476 9072 4540 9076
rect 4476 9016 4490 9072
rect 4490 9016 4540 9072
rect 4476 9012 4540 9016
rect 12572 9012 12636 9076
rect 3917 8732 3981 8736
rect 3917 8676 3921 8732
rect 3921 8676 3977 8732
rect 3977 8676 3981 8732
rect 3917 8672 3981 8676
rect 3997 8732 4061 8736
rect 3997 8676 4001 8732
rect 4001 8676 4057 8732
rect 4057 8676 4061 8732
rect 3997 8672 4061 8676
rect 4077 8732 4141 8736
rect 4077 8676 4081 8732
rect 4081 8676 4137 8732
rect 4137 8676 4141 8732
rect 4077 8672 4141 8676
rect 4157 8732 4221 8736
rect 4157 8676 4161 8732
rect 4161 8676 4217 8732
rect 4217 8676 4221 8732
rect 4157 8672 4221 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 15778 8732 15842 8736
rect 15778 8676 15782 8732
rect 15782 8676 15838 8732
rect 15838 8676 15842 8732
rect 15778 8672 15842 8676
rect 15858 8732 15922 8736
rect 15858 8676 15862 8732
rect 15862 8676 15918 8732
rect 15918 8676 15922 8732
rect 15858 8672 15922 8676
rect 15938 8732 16002 8736
rect 15938 8676 15942 8732
rect 15942 8676 15998 8732
rect 15998 8676 16002 8732
rect 15938 8672 16002 8676
rect 16018 8732 16082 8736
rect 16018 8676 16022 8732
rect 16022 8676 16078 8732
rect 16078 8676 16082 8732
rect 16018 8672 16082 8676
rect 14044 8196 14108 8260
rect 16252 8196 16316 8260
rect 6882 8188 6946 8192
rect 6882 8132 6886 8188
rect 6886 8132 6942 8188
rect 6942 8132 6946 8188
rect 6882 8128 6946 8132
rect 6962 8188 7026 8192
rect 6962 8132 6966 8188
rect 6966 8132 7022 8188
rect 7022 8132 7026 8188
rect 6962 8128 7026 8132
rect 7042 8188 7106 8192
rect 7042 8132 7046 8188
rect 7046 8132 7102 8188
rect 7102 8132 7106 8188
rect 7042 8128 7106 8132
rect 7122 8188 7186 8192
rect 7122 8132 7126 8188
rect 7126 8132 7182 8188
rect 7182 8132 7186 8188
rect 7122 8128 7186 8132
rect 12813 8188 12877 8192
rect 12813 8132 12817 8188
rect 12817 8132 12873 8188
rect 12873 8132 12877 8188
rect 12813 8128 12877 8132
rect 12893 8188 12957 8192
rect 12893 8132 12897 8188
rect 12897 8132 12953 8188
rect 12953 8132 12957 8188
rect 12893 8128 12957 8132
rect 12973 8188 13037 8192
rect 12973 8132 12977 8188
rect 12977 8132 13033 8188
rect 13033 8132 13037 8188
rect 12973 8128 13037 8132
rect 13053 8188 13117 8192
rect 13053 8132 13057 8188
rect 13057 8132 13113 8188
rect 13113 8132 13117 8188
rect 13053 8128 13117 8132
rect 9628 7788 9692 7852
rect 3917 7644 3981 7648
rect 3917 7588 3921 7644
rect 3921 7588 3977 7644
rect 3977 7588 3981 7644
rect 3917 7584 3981 7588
rect 3997 7644 4061 7648
rect 3997 7588 4001 7644
rect 4001 7588 4057 7644
rect 4057 7588 4061 7644
rect 3997 7584 4061 7588
rect 4077 7644 4141 7648
rect 4077 7588 4081 7644
rect 4081 7588 4137 7644
rect 4137 7588 4141 7644
rect 4077 7584 4141 7588
rect 4157 7644 4221 7648
rect 4157 7588 4161 7644
rect 4161 7588 4217 7644
rect 4217 7588 4221 7644
rect 4157 7584 4221 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 15778 7644 15842 7648
rect 15778 7588 15782 7644
rect 15782 7588 15838 7644
rect 15838 7588 15842 7644
rect 15778 7584 15842 7588
rect 15858 7644 15922 7648
rect 15858 7588 15862 7644
rect 15862 7588 15918 7644
rect 15918 7588 15922 7644
rect 15858 7584 15922 7588
rect 15938 7644 16002 7648
rect 15938 7588 15942 7644
rect 15942 7588 15998 7644
rect 15998 7588 16002 7644
rect 15938 7584 16002 7588
rect 16018 7644 16082 7648
rect 16018 7588 16022 7644
rect 16022 7588 16078 7644
rect 16078 7588 16082 7644
rect 16018 7584 16082 7588
rect 6882 7100 6946 7104
rect 6882 7044 6886 7100
rect 6886 7044 6942 7100
rect 6942 7044 6946 7100
rect 6882 7040 6946 7044
rect 6962 7100 7026 7104
rect 6962 7044 6966 7100
rect 6966 7044 7022 7100
rect 7022 7044 7026 7100
rect 6962 7040 7026 7044
rect 7042 7100 7106 7104
rect 7042 7044 7046 7100
rect 7046 7044 7102 7100
rect 7102 7044 7106 7100
rect 7042 7040 7106 7044
rect 7122 7100 7186 7104
rect 7122 7044 7126 7100
rect 7126 7044 7182 7100
rect 7182 7044 7186 7100
rect 7122 7040 7186 7044
rect 12813 7100 12877 7104
rect 12813 7044 12817 7100
rect 12817 7044 12873 7100
rect 12873 7044 12877 7100
rect 12813 7040 12877 7044
rect 12893 7100 12957 7104
rect 12893 7044 12897 7100
rect 12897 7044 12953 7100
rect 12953 7044 12957 7100
rect 12893 7040 12957 7044
rect 12973 7100 13037 7104
rect 12973 7044 12977 7100
rect 12977 7044 13033 7100
rect 13033 7044 13037 7100
rect 12973 7040 13037 7044
rect 13053 7100 13117 7104
rect 13053 7044 13057 7100
rect 13057 7044 13113 7100
rect 13113 7044 13117 7100
rect 13053 7040 13117 7044
rect 13308 6700 13372 6764
rect 14044 6700 14108 6764
rect 3917 6556 3981 6560
rect 3917 6500 3921 6556
rect 3921 6500 3977 6556
rect 3977 6500 3981 6556
rect 3917 6496 3981 6500
rect 3997 6556 4061 6560
rect 3997 6500 4001 6556
rect 4001 6500 4057 6556
rect 4057 6500 4061 6556
rect 3997 6496 4061 6500
rect 4077 6556 4141 6560
rect 4077 6500 4081 6556
rect 4081 6500 4137 6556
rect 4137 6500 4141 6556
rect 4077 6496 4141 6500
rect 4157 6556 4221 6560
rect 4157 6500 4161 6556
rect 4161 6500 4217 6556
rect 4217 6500 4221 6556
rect 4157 6496 4221 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 15778 6556 15842 6560
rect 15778 6500 15782 6556
rect 15782 6500 15838 6556
rect 15838 6500 15842 6556
rect 15778 6496 15842 6500
rect 15858 6556 15922 6560
rect 15858 6500 15862 6556
rect 15862 6500 15918 6556
rect 15918 6500 15922 6556
rect 15858 6496 15922 6500
rect 15938 6556 16002 6560
rect 15938 6500 15942 6556
rect 15942 6500 15998 6556
rect 15998 6500 16002 6556
rect 15938 6496 16002 6500
rect 16018 6556 16082 6560
rect 16018 6500 16022 6556
rect 16022 6500 16078 6556
rect 16078 6500 16082 6556
rect 16018 6496 16082 6500
rect 10916 6292 10980 6356
rect 10732 6156 10796 6220
rect 13492 6080 13556 6084
rect 13492 6024 13506 6080
rect 13506 6024 13556 6080
rect 13492 6020 13556 6024
rect 14044 6020 14108 6084
rect 6882 6012 6946 6016
rect 6882 5956 6886 6012
rect 6886 5956 6942 6012
rect 6942 5956 6946 6012
rect 6882 5952 6946 5956
rect 6962 6012 7026 6016
rect 6962 5956 6966 6012
rect 6966 5956 7022 6012
rect 7022 5956 7026 6012
rect 6962 5952 7026 5956
rect 7042 6012 7106 6016
rect 7042 5956 7046 6012
rect 7046 5956 7102 6012
rect 7102 5956 7106 6012
rect 7042 5952 7106 5956
rect 7122 6012 7186 6016
rect 7122 5956 7126 6012
rect 7126 5956 7182 6012
rect 7182 5956 7186 6012
rect 7122 5952 7186 5956
rect 12813 6012 12877 6016
rect 12813 5956 12817 6012
rect 12817 5956 12873 6012
rect 12873 5956 12877 6012
rect 12813 5952 12877 5956
rect 12893 6012 12957 6016
rect 12893 5956 12897 6012
rect 12897 5956 12953 6012
rect 12953 5956 12957 6012
rect 12893 5952 12957 5956
rect 12973 6012 13037 6016
rect 12973 5956 12977 6012
rect 12977 5956 13033 6012
rect 13033 5956 13037 6012
rect 12973 5952 13037 5956
rect 13053 6012 13117 6016
rect 13053 5956 13057 6012
rect 13057 5956 13113 6012
rect 13113 5956 13117 6012
rect 13053 5952 13117 5956
rect 10916 5612 10980 5676
rect 3917 5468 3981 5472
rect 3917 5412 3921 5468
rect 3921 5412 3977 5468
rect 3977 5412 3981 5468
rect 3917 5408 3981 5412
rect 3997 5468 4061 5472
rect 3997 5412 4001 5468
rect 4001 5412 4057 5468
rect 4057 5412 4061 5468
rect 3997 5408 4061 5412
rect 4077 5468 4141 5472
rect 4077 5412 4081 5468
rect 4081 5412 4137 5468
rect 4137 5412 4141 5468
rect 4077 5408 4141 5412
rect 4157 5468 4221 5472
rect 4157 5412 4161 5468
rect 4161 5412 4217 5468
rect 4217 5412 4221 5468
rect 4157 5408 4221 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 15778 5468 15842 5472
rect 15778 5412 15782 5468
rect 15782 5412 15838 5468
rect 15838 5412 15842 5468
rect 15778 5408 15842 5412
rect 15858 5468 15922 5472
rect 15858 5412 15862 5468
rect 15862 5412 15918 5468
rect 15918 5412 15922 5468
rect 15858 5408 15922 5412
rect 15938 5468 16002 5472
rect 15938 5412 15942 5468
rect 15942 5412 15998 5468
rect 15998 5412 16002 5468
rect 15938 5408 16002 5412
rect 16018 5468 16082 5472
rect 16018 5412 16022 5468
rect 16022 5412 16078 5468
rect 16078 5412 16082 5468
rect 16018 5408 16082 5412
rect 6500 5128 6564 5132
rect 6500 5072 6514 5128
rect 6514 5072 6564 5128
rect 6500 5068 6564 5072
rect 6882 4924 6946 4928
rect 6882 4868 6886 4924
rect 6886 4868 6942 4924
rect 6942 4868 6946 4924
rect 6882 4864 6946 4868
rect 6962 4924 7026 4928
rect 6962 4868 6966 4924
rect 6966 4868 7022 4924
rect 7022 4868 7026 4924
rect 6962 4864 7026 4868
rect 7042 4924 7106 4928
rect 7042 4868 7046 4924
rect 7046 4868 7102 4924
rect 7102 4868 7106 4924
rect 7042 4864 7106 4868
rect 7122 4924 7186 4928
rect 7122 4868 7126 4924
rect 7126 4868 7182 4924
rect 7182 4868 7186 4924
rect 7122 4864 7186 4868
rect 12813 4924 12877 4928
rect 12813 4868 12817 4924
rect 12817 4868 12873 4924
rect 12873 4868 12877 4924
rect 12813 4864 12877 4868
rect 12893 4924 12957 4928
rect 12893 4868 12897 4924
rect 12897 4868 12953 4924
rect 12953 4868 12957 4924
rect 12893 4864 12957 4868
rect 12973 4924 13037 4928
rect 12973 4868 12977 4924
rect 12977 4868 13033 4924
rect 13033 4868 13037 4924
rect 12973 4864 13037 4868
rect 13053 4924 13117 4928
rect 13053 4868 13057 4924
rect 13057 4868 13113 4924
rect 13113 4868 13117 4924
rect 13053 4864 13117 4868
rect 10916 4660 10980 4724
rect 6132 4388 6196 4452
rect 12572 4448 12636 4452
rect 12572 4392 12586 4448
rect 12586 4392 12636 4448
rect 12572 4388 12636 4392
rect 3917 4380 3981 4384
rect 3917 4324 3921 4380
rect 3921 4324 3977 4380
rect 3977 4324 3981 4380
rect 3917 4320 3981 4324
rect 3997 4380 4061 4384
rect 3997 4324 4001 4380
rect 4001 4324 4057 4380
rect 4057 4324 4061 4380
rect 3997 4320 4061 4324
rect 4077 4380 4141 4384
rect 4077 4324 4081 4380
rect 4081 4324 4137 4380
rect 4137 4324 4141 4380
rect 4077 4320 4141 4324
rect 4157 4380 4221 4384
rect 4157 4324 4161 4380
rect 4161 4324 4217 4380
rect 4217 4324 4221 4380
rect 4157 4320 4221 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 15778 4380 15842 4384
rect 15778 4324 15782 4380
rect 15782 4324 15838 4380
rect 15838 4324 15842 4380
rect 15778 4320 15842 4324
rect 15858 4380 15922 4384
rect 15858 4324 15862 4380
rect 15862 4324 15918 4380
rect 15918 4324 15922 4380
rect 15858 4320 15922 4324
rect 15938 4380 16002 4384
rect 15938 4324 15942 4380
rect 15942 4324 15998 4380
rect 15998 4324 16002 4380
rect 15938 4320 16002 4324
rect 16018 4380 16082 4384
rect 16018 4324 16022 4380
rect 16022 4324 16078 4380
rect 16078 4324 16082 4380
rect 16018 4320 16082 4324
rect 4476 3844 4540 3908
rect 6882 3836 6946 3840
rect 6882 3780 6886 3836
rect 6886 3780 6942 3836
rect 6942 3780 6946 3836
rect 6882 3776 6946 3780
rect 6962 3836 7026 3840
rect 6962 3780 6966 3836
rect 6966 3780 7022 3836
rect 7022 3780 7026 3836
rect 6962 3776 7026 3780
rect 7042 3836 7106 3840
rect 7042 3780 7046 3836
rect 7046 3780 7102 3836
rect 7102 3780 7106 3836
rect 7042 3776 7106 3780
rect 7122 3836 7186 3840
rect 7122 3780 7126 3836
rect 7126 3780 7182 3836
rect 7182 3780 7186 3836
rect 7122 3776 7186 3780
rect 12813 3836 12877 3840
rect 12813 3780 12817 3836
rect 12817 3780 12873 3836
rect 12873 3780 12877 3836
rect 12813 3776 12877 3780
rect 12893 3836 12957 3840
rect 12893 3780 12897 3836
rect 12897 3780 12953 3836
rect 12953 3780 12957 3836
rect 12893 3776 12957 3780
rect 12973 3836 13037 3840
rect 12973 3780 12977 3836
rect 12977 3780 13033 3836
rect 13033 3780 13037 3836
rect 12973 3776 13037 3780
rect 13053 3836 13117 3840
rect 13053 3780 13057 3836
rect 13057 3780 13113 3836
rect 13113 3780 13117 3836
rect 13053 3776 13117 3780
rect 3917 3292 3981 3296
rect 3917 3236 3921 3292
rect 3921 3236 3977 3292
rect 3977 3236 3981 3292
rect 3917 3232 3981 3236
rect 3997 3292 4061 3296
rect 3997 3236 4001 3292
rect 4001 3236 4057 3292
rect 4057 3236 4061 3292
rect 3997 3232 4061 3236
rect 4077 3292 4141 3296
rect 4077 3236 4081 3292
rect 4081 3236 4137 3292
rect 4137 3236 4141 3292
rect 4077 3232 4141 3236
rect 4157 3292 4221 3296
rect 4157 3236 4161 3292
rect 4161 3236 4217 3292
rect 4217 3236 4221 3292
rect 4157 3232 4221 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 15778 3292 15842 3296
rect 15778 3236 15782 3292
rect 15782 3236 15838 3292
rect 15838 3236 15842 3292
rect 15778 3232 15842 3236
rect 15858 3292 15922 3296
rect 15858 3236 15862 3292
rect 15862 3236 15918 3292
rect 15918 3236 15922 3292
rect 15858 3232 15922 3236
rect 15938 3292 16002 3296
rect 15938 3236 15942 3292
rect 15942 3236 15998 3292
rect 15998 3236 16002 3292
rect 15938 3232 16002 3236
rect 16018 3292 16082 3296
rect 16018 3236 16022 3292
rect 16022 3236 16078 3292
rect 16078 3236 16082 3292
rect 16018 3232 16082 3236
rect 6500 3028 6564 3092
rect 6882 2748 6946 2752
rect 6882 2692 6886 2748
rect 6886 2692 6942 2748
rect 6942 2692 6946 2748
rect 6882 2688 6946 2692
rect 6962 2748 7026 2752
rect 6962 2692 6966 2748
rect 6966 2692 7022 2748
rect 7022 2692 7026 2748
rect 6962 2688 7026 2692
rect 7042 2748 7106 2752
rect 7042 2692 7046 2748
rect 7046 2692 7102 2748
rect 7102 2692 7106 2748
rect 7042 2688 7106 2692
rect 7122 2748 7186 2752
rect 7122 2692 7126 2748
rect 7126 2692 7182 2748
rect 7182 2692 7186 2748
rect 7122 2688 7186 2692
rect 12813 2748 12877 2752
rect 12813 2692 12817 2748
rect 12817 2692 12873 2748
rect 12873 2692 12877 2748
rect 12813 2688 12877 2692
rect 12893 2748 12957 2752
rect 12893 2692 12897 2748
rect 12897 2692 12953 2748
rect 12953 2692 12957 2748
rect 12893 2688 12957 2692
rect 12973 2748 13037 2752
rect 12973 2692 12977 2748
rect 12977 2692 13033 2748
rect 13033 2692 13037 2748
rect 12973 2688 13037 2692
rect 13053 2748 13117 2752
rect 13053 2692 13057 2748
rect 13057 2692 13113 2748
rect 13113 2692 13117 2748
rect 13053 2688 13117 2692
rect 9628 2620 9692 2684
rect 16988 2620 17052 2684
rect 17724 2680 17788 2684
rect 17724 2624 17774 2680
rect 17774 2624 17788 2680
rect 17724 2620 17788 2624
rect 4844 2484 4908 2548
rect 10732 2484 10796 2548
rect 3917 2204 3981 2208
rect 3917 2148 3921 2204
rect 3921 2148 3977 2204
rect 3977 2148 3981 2204
rect 3917 2144 3981 2148
rect 3997 2204 4061 2208
rect 3997 2148 4001 2204
rect 4001 2148 4057 2204
rect 4057 2148 4061 2204
rect 3997 2144 4061 2148
rect 4077 2204 4141 2208
rect 4077 2148 4081 2204
rect 4081 2148 4137 2204
rect 4137 2148 4141 2204
rect 4077 2144 4141 2148
rect 4157 2204 4221 2208
rect 4157 2148 4161 2204
rect 4161 2148 4217 2204
rect 4217 2148 4221 2204
rect 4157 2144 4221 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 15778 2204 15842 2208
rect 15778 2148 15782 2204
rect 15782 2148 15838 2204
rect 15838 2148 15842 2204
rect 15778 2144 15842 2148
rect 15858 2204 15922 2208
rect 15858 2148 15862 2204
rect 15862 2148 15918 2204
rect 15918 2148 15922 2204
rect 15858 2144 15922 2148
rect 15938 2204 16002 2208
rect 15938 2148 15942 2204
rect 15942 2148 15998 2204
rect 15998 2148 16002 2204
rect 15938 2144 16002 2148
rect 16018 2204 16082 2208
rect 16018 2148 16022 2204
rect 16022 2148 16078 2204
rect 16078 2148 16082 2204
rect 16018 2144 16082 2148
<< metal4 >>
rect 3909 14176 4229 14736
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 13088 4229 14112
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 12000 4229 13024
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 10912 4229 11936
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 9824 4229 10848
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 8736 4229 9760
rect 6874 14720 7195 14736
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7195 14720
rect 6874 13632 7195 14656
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7195 13632
rect 6874 12544 7195 13568
rect 9840 14176 10160 14736
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 13088 10160 14112
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9627 12748 9693 12749
rect 9627 12684 9628 12748
rect 9692 12684 9693 12748
rect 9627 12683 9693 12684
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7195 12544
rect 6874 11456 7195 12480
rect 9630 12069 9690 12683
rect 9627 12068 9693 12069
rect 9627 12004 9628 12068
rect 9692 12004 9693 12068
rect 9627 12003 9693 12004
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7195 11456
rect 6874 10368 7195 11392
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7195 10368
rect 6131 9756 6197 9757
rect 6131 9692 6132 9756
rect 6196 9692 6197 9756
rect 6131 9691 6197 9692
rect 4475 9076 4541 9077
rect 4475 9012 4476 9076
rect 4540 9012 4541 9076
rect 4475 9011 4541 9012
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 7648 4229 8672
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 6560 4229 7584
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 5472 4229 6496
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 4384 4229 5408
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 3296 4229 4320
rect 4478 3909 4538 9011
rect 6134 4453 6194 9691
rect 6874 9280 7195 10304
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7195 9280
rect 6874 8192 7195 9216
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7195 8192
rect 6874 7104 7195 8128
rect 9840 12000 10160 13024
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 10912 10160 11936
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 9824 10160 10848
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 8736 10160 9760
rect 12805 14720 13125 14736
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 13632 13125 14656
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 12544 13125 13568
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 12805 11456 13125 12480
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 10368 13125 11392
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 12805 9280 13125 10304
rect 15770 14176 16091 14736
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16091 14176
rect 15770 13088 16091 14112
rect 17723 13836 17789 13837
rect 17723 13772 17724 13836
rect 17788 13772 17789 13836
rect 17723 13771 17789 13772
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16091 13088
rect 15770 12000 16091 13024
rect 16987 12884 17053 12885
rect 16987 12820 16988 12884
rect 17052 12820 17053 12884
rect 16987 12819 17053 12820
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16091 12000
rect 15770 10912 16091 11936
rect 16251 11660 16317 11661
rect 16251 11596 16252 11660
rect 16316 11596 16317 11660
rect 16251 11595 16317 11596
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16091 10912
rect 15770 9824 16091 10848
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16091 9824
rect 13307 9484 13373 9485
rect 13307 9420 13308 9484
rect 13372 9420 13373 9484
rect 13307 9419 13373 9420
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12571 9076 12637 9077
rect 12571 9012 12572 9076
rect 12636 9012 12637 9076
rect 12571 9011 12637 9012
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9627 7852 9693 7853
rect 9627 7788 9628 7852
rect 9692 7788 9693 7852
rect 9627 7787 9693 7788
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7195 7104
rect 6874 6016 7195 7040
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7195 6016
rect 6499 5132 6565 5133
rect 6499 5068 6500 5132
rect 6564 5068 6565 5132
rect 6499 5067 6565 5068
rect 6131 4452 6197 4453
rect 6131 4388 6132 4452
rect 6196 4388 6197 4452
rect 6131 4387 6197 4388
rect 4475 3908 4541 3909
rect 4475 3844 4476 3908
rect 4540 3844 4541 3908
rect 4475 3843 4541 3844
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 2208 4229 3232
rect 4478 2790 4538 3843
rect 6502 3093 6562 5067
rect 6874 4928 7195 5952
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7195 4928
rect 6874 3840 7195 4864
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7195 3840
rect 6499 3092 6565 3093
rect 6499 3028 6500 3092
rect 6564 3028 6565 3092
rect 6499 3027 6565 3028
rect 4478 2730 4906 2790
rect 4846 2549 4906 2730
rect 6874 2752 7195 3776
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7195 2752
rect 4843 2548 4909 2549
rect 4843 2484 4844 2548
rect 4908 2484 4909 2548
rect 4843 2483 4909 2484
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2128 4229 2144
rect 6874 2128 7195 2688
rect 9630 2685 9690 7787
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 6560 10160 7584
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 5472 10160 6496
rect 10915 6356 10981 6357
rect 10915 6292 10916 6356
rect 10980 6292 10981 6356
rect 10915 6291 10981 6292
rect 10731 6220 10797 6221
rect 10731 6156 10732 6220
rect 10796 6156 10797 6220
rect 10731 6155 10797 6156
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 4384 10160 5408
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 3296 10160 4320
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9627 2684 9693 2685
rect 9627 2620 9628 2684
rect 9692 2620 9693 2684
rect 9627 2619 9693 2620
rect 9840 2208 10160 3232
rect 10734 2549 10794 6155
rect 10918 5677 10978 6291
rect 10915 5676 10981 5677
rect 10915 5612 10916 5676
rect 10980 5612 10981 5676
rect 10915 5611 10981 5612
rect 10918 4725 10978 5611
rect 10915 4724 10981 4725
rect 10915 4660 10916 4724
rect 10980 4660 10981 4724
rect 10915 4659 10981 4660
rect 12574 4453 12634 9011
rect 12805 8192 13125 9216
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 12805 7104 13125 8128
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 6016 13125 7040
rect 13310 6765 13370 9419
rect 13491 9212 13557 9213
rect 13491 9148 13492 9212
rect 13556 9148 13557 9212
rect 13491 9147 13557 9148
rect 13307 6764 13373 6765
rect 13307 6700 13308 6764
rect 13372 6700 13373 6764
rect 13307 6699 13373 6700
rect 13494 6085 13554 9147
rect 15770 8736 16091 9760
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16091 8736
rect 14043 8260 14109 8261
rect 14043 8196 14044 8260
rect 14108 8196 14109 8260
rect 14043 8195 14109 8196
rect 14046 6765 14106 8195
rect 15770 7648 16091 8672
rect 16254 8261 16314 11595
rect 16435 11524 16501 11525
rect 16435 11460 16436 11524
rect 16500 11460 16501 11524
rect 16435 11459 16501 11460
rect 16438 9757 16498 11459
rect 16435 9756 16501 9757
rect 16435 9692 16436 9756
rect 16500 9692 16501 9756
rect 16435 9691 16501 9692
rect 16251 8260 16317 8261
rect 16251 8196 16252 8260
rect 16316 8196 16317 8260
rect 16251 8195 16317 8196
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16091 7648
rect 14043 6764 14109 6765
rect 14043 6700 14044 6764
rect 14108 6700 14109 6764
rect 14043 6699 14109 6700
rect 14046 6085 14106 6699
rect 15770 6560 16091 7584
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16091 6560
rect 13491 6084 13557 6085
rect 13491 6020 13492 6084
rect 13556 6020 13557 6084
rect 13491 6019 13557 6020
rect 14043 6084 14109 6085
rect 14043 6020 14044 6084
rect 14108 6020 14109 6084
rect 14043 6019 14109 6020
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 12805 4928 13125 5952
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12571 4452 12637 4453
rect 12571 4388 12572 4452
rect 12636 4388 12637 4452
rect 12571 4387 12637 4388
rect 12805 3840 13125 4864
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 2752 13125 3776
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 10731 2548 10797 2549
rect 10731 2484 10732 2548
rect 10796 2484 10797 2548
rect 10731 2483 10797 2484
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 12805 2128 13125 2688
rect 15770 5472 16091 6496
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16091 5472
rect 15770 4384 16091 5408
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16091 4384
rect 15770 3296 16091 4320
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16091 3296
rect 15770 2208 16091 3232
rect 16990 2685 17050 12819
rect 17726 2685 17786 13771
rect 16987 2684 17053 2685
rect 16987 2620 16988 2684
rect 17052 2620 17053 2684
rect 16987 2619 17053 2620
rect 17723 2684 17789 2685
rect 17723 2620 17724 2684
rect 17788 2620 17789 2684
rect 17723 2619 17789 2620
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16091 2208
rect 15770 2128 16091 2144
use sky130_fd_sc_hd__clkbuf_2  output76 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 1748 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output70
timestamp 1624635492
transform -1 0 1748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1624635492
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output79
timestamp 1624635492
transform -1 0 2116 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output71
timestamp 1624635492
transform -1 0 2116 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output84
timestamp 1624635492
transform -1 0 2484 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output54
timestamp 1624635492
transform -1 0 2484 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 3036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output86
timestamp 1624635492
transform -1 0 3220 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output85
timestamp 1624635492
transform -1 0 2852 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output82
timestamp 1624635492
transform -1 0 2852 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3864 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output88
timestamp 1624635492
transform -1 0 3956 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output87
timestamp 1624635492
transform -1 0 3588 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output83
timestamp 1624635492
transform -1 0 3772 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output61
timestamp 1624635492
transform -1 0 3404 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_31
timestamp 1624635492
transform 1 0 3956 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35
timestamp 1624635492
transform 1 0 4324 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output62
timestamp 1624635492
transform -1 0 4324 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 4416 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1624635492
transform 1 0 4048 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1624635492
transform -1 0 5060 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1624635492
transform -1 0 5796 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output64
timestamp 1624635492
transform -1 0 6164 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output63
timestamp 1624635492
transform -1 0 5612 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1624635492
transform 1 0 5060 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__A0
timestamp 1624635492
transform -1 0 6716 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 6440 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output68
timestamp 1624635492
transform 1 0 6624 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output65
timestamp 1624635492
transform -1 0 7084 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1624635492
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1624635492
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _35_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 6164 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _21_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5888 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1624635492
transform -1 0 9016 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_1_
timestamp 1624635492
transform 1 0 8280 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_0_
timestamp 1624635492
transform 1 0 7452 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l4_in_0_
timestamp 1624635492
transform -1 0 8188 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output66
timestamp 1624635492
transform 1 0 7084 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output67
timestamp 1624635492
transform 1 0 6992 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1624635492
transform 1 0 9844 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1624635492
transform 1 0 10672 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1624635492
transform 1 0 9016 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l1_in_0_
timestamp 1624635492
transform 1 0 10212 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9384 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1624635492
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A0
timestamp 1624635492
transform -1 0 9384 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_2_
timestamp 1624635492
transform -1 0 12696 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_3_
timestamp 1624635492
transform -1 0 12512 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_1_
timestamp 1624635492
transform 1 0 12512 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1624635492
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1624635492
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output55
timestamp 1624635492
transform -1 0 11592 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A0
timestamp 1624635492
transform -1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 11224 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_113
timestamp 1624635492
transform 1 0 11500 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output56
timestamp 1624635492
transform -1 0 13064 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 13340 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output69
timestamp 1624635492
transform -1 0 13800 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output57
timestamp 1624635492
transform -1 0 13432 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_138
timestamp 1624635492
transform 1 0 13800 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output122
timestamp 1624635492
transform 1 0 13524 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output58
timestamp 1624635492
transform -1 0 14260 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 13892 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1624635492
transform -1 0 14444 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 14168 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_145
timestamp 1624635492
transform 1 0 14444 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1624635492
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_153
timestamp 1624635492
transform 1 0 15180 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_149
timestamp 1624635492
transform 1 0 14812 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1624635492
transform -1 0 15364 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output119
timestamp 1624635492
transform 1 0 15364 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output59
timestamp 1624635492
transform -1 0 15180 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_1_
timestamp 1624635492
transform 1 0 15272 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 14904 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 14536 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 14536 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output60
timestamp 1624635492
transform -1 0 16100 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_1_N_FTB01
timestamp 1624635492
transform -1 0 16376 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 16100 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 16376 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output118
timestamp 1624635492
transform 1 0 16376 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output115
timestamp 1624635492
transform 1 0 16744 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1624635492
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_1_S_FTB01
timestamp 1624635492
transform 1 0 16560 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1624635492
transform 1 0 16928 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output120
timestamp 1624635492
transform 1 0 17112 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output112
timestamp 1624635492
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1624635492
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output113
timestamp 1624635492
transform 1 0 17480 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output52
timestamp 1624635492
transform -1 0 17940 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output103
timestamp 1624635492
transform 1 0 17848 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output102
timestamp 1624635492
transform 1 0 18216 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output91
timestamp 1624635492
transform 1 0 18216 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1624635492
transform -1 0 18216 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624635492
transform -1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624635492
transform -1 0 18860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 2852 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1624635492
transform -1 0 3772 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624635492
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_19
timestamp 1624635492
transform 1 0 2852 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 4600 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1624635492
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output89
timestamp 1624635492
transform -1 0 4232 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output90
timestamp 1624635492
transform -1 0 4600 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 6072 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp 1624635492
transform 1 0 7544 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp 1624635492
transform 1 0 7820 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1624635492
transform 1 0 8188 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_76
timestamp 1624635492
transform 1 0 8096 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1624635492
transform -1 0 10948 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 10580 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1624635492
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_103
timestamp 1624635492
transform 1 0 10580 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 10948 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 12420 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 13892 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 14352 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1624635492
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_142
timestamp 1624635492
transform 1 0 14168 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_3_
timestamp 1624635492
transform 1 0 15456 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_0_
timestamp 1624635492
transform 1 0 16284 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l4_in_0_
timestamp 1624635492
transform -1 0 15456 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1624635492
transform -1 0 17848 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1624635492
transform -1 0 17572 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output104
timestamp 1624635492
transform 1 0 18216 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output105
timestamp 1624635492
transform 1 0 17848 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1624635492
transform 1 0 17112 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624635492
transform -1 0 18860 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 2944 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624635492
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output72
timestamp 1624635492
transform -1 0 1748 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output73
timestamp 1624635492
transform -1 0 2116 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output75
timestamp 1624635492
transform -1 0 2484 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output78
timestamp 1624635492
transform -1 0 2852 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_19
timestamp 1624635492
transform 1 0 2852 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1624635492
transform 1 0 4508 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_36
timestamp 1624635492
transform 1 0 4416 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _36_
timestamp 1624635492
transform 1 0 6440 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1624635492
transform 1 0 5336 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1624635492
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 6716 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 6900 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 9844 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _44_
timestamp 1624635492
transform 1 0 9844 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 10120 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1624635492
transform 1 0 10580 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A0
timestamp 1624635492
transform -1 0 10580 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_0_
timestamp 1624635492
transform 1 0 11868 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1624635492
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 11684 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A0
timestamp 1624635492
transform -1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l1_in_0_
timestamp 1624635492
transform -1 0 13524 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_0_
timestamp 1624635492
transform 1 0 13524 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 14352 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 16376 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  prog_clk_3_E_FTB01 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 14904 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1624635492
transform -1 0 16560 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1624635492
transform -1 0 16836 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_0_
timestamp 1624635492
transform 1 0 16928 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1624635492
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output106
timestamp 1624635492
transform 1 0 18216 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output107
timestamp 1624635492
transform 1 0 17848 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_181
timestamp 1624635492
transform 1 0 17756 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624635492
transform -1 0 18860 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1624635492
transform 1 0 2576 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1624635492
transform 1 0 1748 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624635492
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output74
timestamp 1624635492
transform -1 0 1748 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _37_
timestamp 1624635492
transform -1 0 3680 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1624635492
transform 1 0 3864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1624635492
transform 1 0 4140 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1624635492
transform 1 0 4508 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1624635492
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_28
timestamp 1624635492
transform 1 0 3680 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_36
timestamp 1624635492
transform 1 0 4416 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _43_
timestamp 1624635492
transform 1 0 5336 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _45_
timestamp 1624635492
transform 1 0 5612 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _46_
timestamp 1624635492
transform 1 0 5888 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1624635492
transform 1 0 6164 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1624635492
transform -1 0 8188 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1624635492
transform 1 0 6992 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1624635492
transform -1 0 9016 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_73
timestamp 1624635492
transform 1 0 7820 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 9108 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l4_in_0_
timestamp 1624635492
transform -1 0 11224 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1624635492
transform 1 0 9568 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1624635492
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__A0
timestamp 1624635492
transform -1 0 9568 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_2_
timestamp 1624635492
transform -1 0 12880 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_3_
timestamp 1624635492
transform -1 0 12052 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1624635492
transform 1 0 13708 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_1_
timestamp 1624635492
transform 1 0 12880 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1624635492
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1624635492
transform -1 0 14628 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A0
timestamp 1624635492
transform -1 0 14260 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_140
timestamp 1624635492
transform 1 0 13984 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 14996 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1624635492
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1624635492
transform -1 0 18216 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1624635492
transform -1 0 17112 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1624635492
transform -1 0 16836 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_0_
timestamp 1624635492
transform 1 0 17112 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output108
timestamp 1624635492
transform 1 0 18216 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_167
timestamp 1624635492
transform 1 0 16468 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624635492
transform -1 0 18860 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 2392 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1624635492
transform -1 0 2392 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1624635492
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1624635492
transform -1 0 1564 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1624635492
transform 1 0 4232 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 5980 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  output77
timestamp 1624635492
transform -1 0 4232 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _47_
timestamp 1624635492
transform 1 0 6440 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1624635492
transform 1 0 5980 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1624635492
transform 1 0 6716 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1624635492
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_56
timestamp 1624635492
transform 1 0 6256 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1624635492
transform 1 0 7544 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1624635492
transform 1 0 8372 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 11224 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 9200 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 9476 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 13156 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 11224 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1624635492
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_113
timestamp 1624635492
transform 1 0 11500 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 14904 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_top_ipin_0.prog_clk
timestamp 1624635492
transform 1 0 13156 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1624635492
transform -1 0 16560 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1624635492
transform -1 0 15456 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_2_
timestamp 1624635492
transform 1 0 15456 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_top_ipin_0.prog_clk
timestamp 1624635492
transform -1 0 15180 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1624635492
transform 1 0 17940 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1624635492
transform -1 0 16836 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_1_
timestamp 1624635492
transform 1 0 17112 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1624635492
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output109
timestamp 1624635492
transform 1 0 18216 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1624635492
transform -1 0 17112 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1624635492
transform -1 0 18860 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_9
timestamp 1624635492
transform 1 0 1932 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_9
timestamp 1624635492
transform 1 0 1932 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1380 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input5
timestamp 1624635492
transform 1 0 1380 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1624635492
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1624635492
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1624635492
transform -1 0 2852 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1624635492
transform -1 0 2852 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1624635492
transform 1 0 2852 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 4324 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4324 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1624635492
transform 1 0 3864 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1624635492
transform 1 0 4784 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1624635492
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_28
timestamp 1624635492
transform 1 0 3680 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_39
timestamp 1624635492
transform 1 0 4692 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1624635492
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 8004 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1624635492
transform -1 0 6440 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1624635492
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output81
timestamp 1624635492
transform -1 0 6164 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1624635492
transform -1 0 6348 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 6716 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_58
timestamp 1624635492
transform 1 0 6440 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 7820 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1624635492
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1624635492
transform 1 0 6900 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_7_72
timestamp 1624635492
transform 1 0 7728 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1624635492
transform -1 0 9936 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9108 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 9384 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1624635492
transform -1 0 10764 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1624635492
transform -1 0 11408 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1624635492
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_89
timestamp 1624635492
transform 1 0 9292 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1624635492
transform 1 0 11776 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 12236 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_1_
timestamp 1624635492
transform 1 0 12328 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_2_
timestamp 1624635492
transform -1 0 11592 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_3_
timestamp 1624635492
transform 1 0 11408 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 12328 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1624635492
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_115
timestamp 1624635492
transform 1 0 11684 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_0_
timestamp 1624635492
transform -1 0 14812 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_1_
timestamp 1624635492
transform -1 0 15180 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_2_
timestamp 1624635492
transform -1 0 13984 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1624635492
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_top_ipin_0.prog_clk
timestamp 1624635492
transform -1 0 13984 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1624635492
transform 1 0 13984 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_142
timestamp 1624635492
transform 1 0 14168 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1624635492
transform -1 0 15640 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_0_
timestamp 1624635492
transform 1 0 14812 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l4_in_0_
timestamp 1624635492
transform 1 0 15640 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_1_
timestamp 1624635492
transform -1 0 16468 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1624635492
transform 1 0 15180 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_172
timestamp 1624635492
transform 1 0 16928 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1624635492
transform 1 0 16468 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1624635492
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_2_
timestamp 1624635492
transform 1 0 17020 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 1624635492
transform -1 0 16836 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output110
timestamp 1624635492
transform 1 0 17848 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output93
timestamp 1624635492
transform 1 0 18216 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output92
timestamp 1624635492
transform 1 0 18216 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1624635492
transform -1 0 18216 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 16468 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1624635492
transform -1 0 18860 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1624635492
transform -1 0 18860 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 1472 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1624635492
transform 1 0 2944 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1624635492
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1624635492
transform 1 0 1380 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1624635492
transform 1 0 3864 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1624635492
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output80
timestamp 1624635492
transform -1 0 5060 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 6532 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1624635492
transform -1 0 7544 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1624635492
transform -1 0 6716 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1624635492
transform -1 0 8464 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_top_ipin_0.prog_clk
timestamp 1624635492
transform -1 0 8740 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_top_ipin_0.prog_clk
timestamp 1624635492
transform -1 0 9016 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_70
timestamp 1624635492
transform 1 0 7544 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 10580 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1624635492
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 10580 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 13064 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_1_
timestamp 1624635492
transform -1 0 11592 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1624635492
transform -1 0 13432 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 14352 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_1_
timestamp 1624635492
transform 1 0 13432 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1624635492
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_130
timestamp 1624635492
transform 1 0 13064 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 15824 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  output94
timestamp 1624635492
transform 1 0 18216 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output95
timestamp 1624635492
transform 1 0 17848 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output97
timestamp 1624635492
transform 1 0 17480 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A0
timestamp 1624635492
transform -1 0 17480 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1624635492
transform -1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1624635492
transform 1 0 2576 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1624635492
transform -1 0 2576 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1624635492
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1624635492
transform 1 0 4232 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1624635492
transform 1 0 4508 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 6256 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1624635492
transform -1 0 4232 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1624635492
transform 1 0 6440 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1624635492
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_56
timestamp 1624635492
transform 1 0 6256 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _16_
timestamp 1624635492
transform -1 0 7544 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1624635492
transform 1 0 7544 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1624635492
transform -1 0 8648 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1624635492
transform 1 0 8648 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1624635492
transform -1 0 10304 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1624635492
transform -1 0 11132 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 11684 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1624635492
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_top_ipin_0.prog_clk
timestamp 1624635492
transform -1 0 11592 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1624635492
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1624635492
transform -1 0 14444 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 14444 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_0_
timestamp 1624635492
transform 1 0 13156 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_1_
timestamp 1624635492
transform -1 0 16744 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_2_
timestamp 1624635492
transform -1 0 17756 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_3_
timestamp 1624635492
transform 1 0 17756 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1624635492
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_170
timestamp 1624635492
transform 1 0 16744 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1624635492
transform -1 0 18860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1624635492
transform 1 0 1840 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1624635492
transform 1 0 2668 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1624635492
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1624635492
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_7
timestamp 1624635492
transform 1 0 1748 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1624635492
transform -1 0 3772 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1624635492
transform 1 0 3864 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1624635492
transform -1 0 5520 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1624635492
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1624635492
transform -1 0 5796 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1624635492
transform -1 0 6072 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 7544 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1624635492
transform -1 0 8372 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_top_ipin_0.prog_clk
timestamp 1624635492
transform 1 0 8372 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 8648 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1624635492
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_top_ipin_0.prog_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 11500 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 9108 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 9292 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 9476 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 12328 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l4_in_0_
timestamp 1624635492
transform -1 0 12328 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1624635492
transform -1 0 14260 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 15916 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1624635492
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 13800 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_144
timestamp 1624635492
transform 1 0 14352 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_0_
timestamp 1624635492
transform -1 0 16836 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_161
timestamp 1624635492
transform 1 0 15916 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_0_
timestamp 1624635492
transform 1 0 16836 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_1_
timestamp 1624635492
transform 1 0 17664 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1624635492
transform -1 0 18860 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_189
timestamp 1624635492
transform 1 0 18492 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 2944 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 2944 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1624635492
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1624635492
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 4416 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 6440 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1624635492
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_top_ipin_0.prog_clk
timestamp 1624635492
transform 1 0 5888 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1624635492
transform -1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 9476 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_74
timestamp 1624635492
transform 1 0 7912 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 11592 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 9936 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_95
timestamp 1624635492
transform 1 0 9844 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_0_
timestamp 1624635492
transform -1 0 13156 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1624635492
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_115
timestamp 1624635492
transform 1 0 11684 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_0_
timestamp 1624635492
transform 1 0 13156 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_1_
timestamp 1624635492
transform 1 0 13984 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 1624635492
transform -1 0 16468 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l4_in_0_
timestamp 1624635492
transform 1 0 15364 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output99
timestamp 1624635492
transform 1 0 14996 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 14812 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l1_in_0_
timestamp 1624635492
transform 1 0 16928 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1624635492
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input36
timestamp 1624635492
transform -1 0 18584 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output96
timestamp 1624635492
transform 1 0 17848 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output98
timestamp 1624635492
transform 1 0 16468 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_181
timestamp 1624635492
transform 1 0 17756 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1624635492
transform -1 0 18860 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 3220 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1624635492
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1624635492
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1624635492
transform -1 0 4692 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1624635492
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1624635492
transform 1 0 4692 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1624635492
transform 1 0 3220 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1624635492
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4968 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1624635492
transform -1 0 7268 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1624635492
transform 1 0 8188 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1624635492
transform -1 0 8096 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_76
timestamp 1624635492
transform 1 0 8096 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9200 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1624635492
transform 1 0 10672 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1624635492
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_87
timestamp 1624635492
transform 1 0 9108 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_0_
timestamp 1624635492
transform -1 0 12972 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_top_ipin_0.prog_clk
timestamp 1624635492
transform -1 0 12144 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 11684 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 11500 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1624635492
transform -1 0 14260 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 14352 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_2_
timestamp 1624635492
transform 1 0 12972 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1624635492
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1624635492
transform 1 0 13800 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 15824 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_1_
timestamp 1624635492
transform 1 0 17296 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  input25
timestamp 1624635492
transform -1 0 18584 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_185
timestamp 1624635492
transform 1 0 18124 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1624635492
transform -1 0 18860 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1624635492
transform 1 0 1932 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 2852 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1624635492
transform -1 0 3772 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1624635492
transform -1 0 3036 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1624635492
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1624635492
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input18
timestamp 1624635492
transform 1 0 1380 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_19
timestamp 1624635492
transform 1 0 2852 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1624635492
transform 1 0 4324 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1624635492
transform 1 0 4140 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1624635492
transform 1 0 3036 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1624635492
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1624635492
transform 1 0 3864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1624635492
transform 1 0 3864 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_34
timestamp 1624635492
transform 1 0 4232 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 6440 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1624635492
transform 1 0 5152 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1624635492
transform -1 0 5796 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1624635492
transform -1 0 7084 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1624635492
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_top_ipin_0.prog_clk
timestamp 1624635492
transform 1 0 6072 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_top_ipin_0.prog_clk
timestamp 1624635492
transform 1 0 5796 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 5980 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_55
timestamp 1624635492
transform 1 0 6164 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 7912 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1624635492
transform 1 0 7084 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1624635492
transform 1 0 7912 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_top_ipin_0.prog_clk
timestamp 1624635492
transform -1 0 9016 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9384 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 11684 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1624635492
transform -1 0 10212 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1624635492
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 9108 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_89
timestamp 1624635492
transform 1 0 9292 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_113
timestamp 1624635492
transform 1 0 11500 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 10856 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_top_ipin_0.prog_clk
timestamp 1624635492
transform 1 0 11224 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1624635492
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 11684 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 11868 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 12052 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 12236 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_1_
timestamp 1624635492
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 11868 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1624635492
transform -1 0 13708 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_2_
timestamp 1624635492
transform 1 0 13708 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_1_
timestamp 1624635492
transform -1 0 14168 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l4_in_0_
timestamp 1624635492
transform 1 0 14352 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1624635492
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1624635492
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_142
timestamp 1624635492
transform 1 0 14168 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_3_
timestamp 1624635492
transform 1 0 14536 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l1_in_0_
timestamp 1624635492
transform -1 0 16008 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_0_
timestamp 1624635492
transform 1 0 16100 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_0_
timestamp 1624635492
transform 1 0 15916 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output100
timestamp 1624635492
transform 1 0 15548 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A0
timestamp 1624635492
transform -1 0 15548 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_162
timestamp 1624635492
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 16928 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_1_
timestamp 1624635492
transform 1 0 16928 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_2_
timestamp 1624635492
transform 1 0 17756 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1624635492
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_170
timestamp 1624635492
transform 1 0 16744 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1624635492
transform -1 0 18860 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1624635492
transform -1 0 18860 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1624635492
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1624635492
transform 1 0 2300 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1624635492
transform -1 0 2300 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1624635492
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1624635492
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 5520 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1624635492
transform 1 0 3220 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_22
timestamp 1624635492
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 6440 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1624635492
transform -1 0 6348 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1624635492
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1624635492
transform 1 0 7912 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1624635492
transform 1 0 10304 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9476 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 8924 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 12236 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1624635492
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 12052 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 11868 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1624635492
transform 1 0 11500 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 13708 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 16652 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 16928 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1624635492
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1624635492
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1624635492
transform -1 0 18860 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1624635492
transform -1 0 18584 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 3772 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1624635492
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1624635492
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1624635492
transform 1 0 1748 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1624635492
transform -1 0 2300 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1624635492
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1624635492
transform -1 0 4048 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1624635492
transform -1 0 4232 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1624635492
transform -1 0 4416 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1624635492
transform -1 0 4600 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 4784 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 4784 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 6900 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 4968 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_46
timestamp 1624635492
transform 1 0 5336 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1624635492
transform 1 0 7176 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1624635492
transform -1 0 9016 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 8004 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 7084 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_65
timestamp 1624635492
transform 1 0 7084 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 10948 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1624635492
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 9108 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 9292 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1624635492
transform -1 0 11776 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1624635492
transform 1 0 11776 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 12972 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 13156 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 13340 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 13524 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 13708 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 13892 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 14076 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_144
timestamp 1624635492
transform 1 0 14352 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1624635492
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 14444 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 15088 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_top_ipin_0.prog_clk
timestamp 1624635492
transform -1 0 15088 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 14812 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1624635492
transform 1 0 18308 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1624635492
transform 1 0 16836 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp 1624635492
transform 1 0 16560 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_3_
timestamp 1624635492
transform 1 0 17480 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  input37
timestamp 1624635492
transform -1 0 17480 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1624635492
transform -1 0 18860 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1624635492
transform -1 0 2852 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1624635492
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1624635492
transform 1 0 1748 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1624635492
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1624635492
transform 1 0 2852 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1624635492
transform 1 0 3220 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A0
timestamp 1624635492
transform -1 0 3864 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1624635492
transform -1 0 3680 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 3864 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1624635492
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_38
timestamp 1624635492
transform 1 0 4600 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1624635492
transform 1 0 4876 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_43
timestamp 1624635492
transform 1 0 5060 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 5336 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 5152 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 5520 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 5704 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_60
timestamp 1624635492
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_54
timestamp 1624635492
transform 1 0 6072 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1624635492
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1624635492
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1624635492
transform 1 0 6440 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1624635492
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1624635492
transform 1 0 6716 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1624635492
transform 1 0 7636 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 8280 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 7912 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 8096 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_70
timestamp 1624635492
transform 1 0 7544 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1624635492
transform 1 0 9752 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1624635492
transform -1 0 11500 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_103
timestamp 1624635492
transform 1 0 10580 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1624635492
transform 1 0 11684 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1624635492
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 12328 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1624635492
transform 1 0 11500 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_124 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 12512 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 14352 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 13984 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 14168 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_136 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 13616 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 15088 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1624635492
transform 1 0 14904 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1624635492
transform 1 0 16376 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_0__A0
timestamp 1624635492
transform -1 0 16376 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 14536 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 14720 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp 1624635492
transform -1 0 17296 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1624635492
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input38
timestamp 1624635492
transform -1 0 18584 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1624635492
transform -1 0 18032 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1624635492
transform -1 0 17664 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1624635492
transform -1 0 16836 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_168
timestamp 1624635492
transform 1 0 16560 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_172
timestamp 1624635492
transform 1 0 16928 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1624635492
transform -1 0 18860 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1624635492
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1624635492
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1624635492
transform 1 0 1748 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1624635492
transform -1 0 2300 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1624635492
transform -1 0 2484 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1624635492
transform -1 0 2668 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1624635492
transform -1 0 2852 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1624635492
transform -1 0 3036 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1624635492
transform -1 0 3404 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1624635492
transform -1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1624635492
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 3864 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1624635492
transform 1 0 4232 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1624635492
transform 1 0 4416 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_38
timestamp 1624635492
transform 1 0 4600 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 4692 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1624635492
transform -1 0 5060 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1624635492
transform 1 0 5060 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 5428 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 5244 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1624635492
transform 1 0 5612 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_51
timestamp 1624635492
transform 1 0 5796 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A1
timestamp 1624635492
transform -1 0 6072 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1624635492
transform 1 0 6072 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 6440 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1624635492
transform 1 0 6256 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_60
timestamp 1624635492
transform 1 0 6624 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1624635492
transform 1 0 6716 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 7268 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1624635492
transform 1 0 7084 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1624635492
transform 1 0 6900 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_69
timestamp 1624635492
transform 1 0 7452 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1624635492
transform 1 0 8188 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1624635492
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1624635492
transform -1 0 9936 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1624635492
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A0
timestamp 1624635492
transform -1 0 10120 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 10120 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 10304 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1624635492
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1624635492
transform 1 0 8924 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 11224 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_106 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 10856 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_112
timestamp 1624635492
transform 1 0 11408 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_124
timestamp 1624635492
transform 1 0 12512 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1624635492
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_3_E_FTB01_A
timestamp 1624635492
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_136 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 13616 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_142
timestamp 1624635492
transform 1 0 14168 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_144
timestamp 1624635492
transform 1 0 14352 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_147
timestamp 1624635492
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 15180 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 15364 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 15548 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 15732 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_0__A0
timestamp 1624635492
transform -1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_163
timestamp 1624635492
transform 1 0 16100 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1624635492
transform -1 0 16376 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1624635492
transform -1 0 16560 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_168
timestamp 1624635492
transform 1 0 16560 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1624635492
transform -1 0 16836 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1624635492
transform 1 0 16836 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_173
timestamp 1624635492
transform 1 0 17020 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1624635492
transform -1 0 17296 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1624635492
transform -1 0 17480 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1624635492
transform -1 0 17848 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1624635492
transform -1 0 17664 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output101
timestamp 1624635492
transform 1 0 17848 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1624635492
transform -1 0 18584 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1624635492
transform -1 0 18860 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1624635492
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1624635492
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1624635492
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1624635492
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1624635492
transform 1 0 1748 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _32_
timestamp 1624635492
transform 1 0 1748 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1624635492
transform 1 0 2116 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_2_W_FTB01
timestamp 1624635492
transform 1 0 2392 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  prog_clk_2_E_FTB01
timestamp 1624635492
transform 1 0 2024 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1624635492
transform -1 0 3036 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1624635492
transform -1 0 3036 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1624635492
transform -1 0 2852 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1624635492
transform -1 0 2852 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1624635492
transform -1 0 2668 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1624635492
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1624635492
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A0
timestamp 1624635492
transform -1 0 3404 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A0
timestamp 1624635492
transform -1 0 3680 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1624635492
transform -1 0 3864 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_25
timestamp 1624635492
transform 1 0 3404 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_30
timestamp 1624635492
transform 1 0 3864 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3036 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_30
timestamp 1624635492
transform 1 0 3864 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _34_
timestamp 1624635492
transform 1 0 6072 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1624635492
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_42
timestamp 1624635492
transform 1 0 4968 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_54
timestamp 1624635492
transform 1 0 6072 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_58
timestamp 1624635492
transform 1 0 6440 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_42
timestamp 1624635492
transform 1 0 4968 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_57
timestamp 1624635492
transform 1 0 6348 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_70
timestamp 1624635492
transform 1 0 7544 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_82
timestamp 1624635492
transform 1 0 8648 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_69
timestamp 1624635492
transform 1 0 7452 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_81
timestamp 1624635492
transform 1 0 8556 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1624635492
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 9108 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_85
timestamp 1624635492
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_89
timestamp 1624635492
transform 1 0 9292 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_101
timestamp 1624635492
transform 1 0 10396 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 1624635492
transform 1 0 8924 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_87
timestamp 1624635492
transform 1 0 9108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_99
timestamp 1624635492
transform 1 0 10212 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1624635492
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 1624635492
transform 1 0 11500 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_115
timestamp 1624635492
transform 1 0 11684 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_111
timestamp 1624635492
transform 1 0 11316 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_123
timestamp 1624635492
transform 1 0 12420 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1624635492
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_127
timestamp 1624635492
transform 1 0 12788 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_139
timestamp 1624635492
transform 1 0 13892 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_135
timestamp 1624635492
transform 1 0 13524 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_144
timestamp 1624635492
transform 1 0 14352 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_151
timestamp 1624635492
transform 1 0 14996 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_156
timestamp 1624635492
transform 1 0 15456 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_155
timestamp 1624635492
transform 1 0 15364 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_1_S_FTB01_A
timestamp 1624635492
transform 1 0 15456 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_1_N_FTB01_A
timestamp 1624635492
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_162
timestamp 1624635492
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output120_A
timestamp 1624635492
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A1
timestamp 1624635492
transform -1 0 16008 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 16192 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1624635492
transform -1 0 16560 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_168
timestamp 1624635492
transform 1 0 16560 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A0
timestamp 1624635492
transform -1 0 16652 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 16836 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1624635492
transform -1 0 16836 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1624635492
transform -1 0 17020 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1624635492
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1624635492
transform -1 0 17112 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1624635492
transform -1 0 17296 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1624635492
transform -1 0 17204 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1624635492
transform -1 0 17388 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  clk_2_E_FTB01
timestamp 1624635492
transform 1 0 17296 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1624635492
transform -1 0 17572 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  clk_3_E_FTB01
timestamp 1624635492
transform -1 0 17848 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  clk_1_S_FTB01
timestamp 1624635492
transform -1 0 17848 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1624635492
transform -1 0 18216 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1624635492
transform -1 0 18216 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1624635492
transform -1 0 18584 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1624635492
transform -1 0 18584 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1624635492
transform -1 0 18860 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1624635492
transform -1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_2_W_FTB01
timestamp 1624635492
transform 1 0 2484 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_3_W_FTB01
timestamp 1624635492
transform 1 0 2760 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1624635492
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output51
timestamp 1624635492
transform -1 0 1748 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output121
timestamp 1624635492
transform -1 0 2116 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output123
timestamp 1624635492
transform -1 0 2484 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_3_W_FTB01
timestamp 1624635492
transform 1 0 3036 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1624635492
transform -1 0 3496 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1624635492
transform -1 0 3680 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1624635492
transform -1 0 3864 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1624635492
transform -1 0 4048 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_3_W_FTB01_A
timestamp 1624635492
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_34
timestamp 1624635492
transform 1 0 4232 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1624635492
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_46
timestamp 1624635492
transform 1 0 5336 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_54
timestamp 1624635492
transform 1 0 6072 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_58
timestamp 1624635492
transform 1 0 6440 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_70
timestamp 1624635492
transform 1 0 7544 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_82
timestamp 1624635492
transform 1 0 8648 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clk_1_N_FTB01
timestamp 1624635492
transform -1 0 9844 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_90
timestamp 1624635492
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_95
timestamp 1624635492
transform 1 0 9844 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1624635492
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_107
timestamp 1624635492
transform 1 0 10948 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_113
timestamp 1624635492
transform 1 0 11500 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_115
timestamp 1624635492
transform 1 0 11684 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_127
timestamp 1624635492
transform 1 0 12788 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_139
timestamp 1624635492
transform 1 0 13892 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 15548 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1624635492
transform -1 0 16468 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1624635492
transform -1 0 16284 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_W_FTB01_A
timestamp 1624635492
transform 1 0 15364 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_151
timestamp 1624635492
transform 1 0 14996 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1624635492
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1624635492
transform -1 0 18584 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1624635492
transform -1 0 18216 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1624635492
transform -1 0 17848 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1624635492
transform -1 0 17480 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1624635492
transform -1 0 17112 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1624635492
transform -1 0 16836 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1624635492
transform -1 0 16652 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1624635492
transform -1 0 18860 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1624635492
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1624635492
transform 1 0 2484 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1624635492
transform 1 0 2760 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1624635492
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output114
timestamp 1624635492
transform -1 0 2116 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output116
timestamp 1624635492
transform -1 0 2484 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1624635492
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1624635492
transform 1 0 3036 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1624635492
transform -1 0 3588 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1624635492
transform 1 0 3864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1624635492
transform 1 0 4140 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 1624635492
transform -1 0 4692 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1624635492
transform -1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1624635492
transform -1 0 4876 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1624635492
transform -1 0 5060 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1624635492
transform 1 0 6440 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output53
timestamp 1624635492
transform -1 0 6256 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_43
timestamp 1624635492
transform 1 0 5060 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_51
timestamp 1624635492
transform 1 0 5796 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_56
timestamp 1624635492
transform 1 0 6256 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_59
timestamp 1624635492
transform 1 0 6532 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_71
timestamp 1624635492
transform 1 0 7636 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_83
timestamp 1624635492
transform 1 0 8740 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1624635492
transform 1 0 9108 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output111
timestamp 1624635492
transform -1 0 10212 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_88
timestamp 1624635492
transform 1 0 9200 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_94
timestamp 1624635492
transform 1 0 9752 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_99
timestamp 1624635492
transform 1 0 10212 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1624635492
transform 1 0 11776 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_111
timestamp 1624635492
transform 1 0 11316 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_115
timestamp 1624635492
transform 1 0 11684 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_117
timestamp 1624635492
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1624635492
transform 1 0 14444 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_129
timestamp 1624635492
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1624635492
transform 1 0 14076 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1624635492
transform -1 0 16744 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output117
timestamp 1624635492
transform 1 0 16100 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1624635492
transform -1 0 16100 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_146
timestamp 1624635492
transform 1 0 14536 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_158
timestamp 1624635492
transform 1 0 15640 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _33_
timestamp 1624635492
transform 1 0 17204 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1624635492
transform 1 0 17112 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1624635492
transform -1 0 18584 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input29
timestamp 1624635492
transform -1 0 18216 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1624635492
transform -1 0 17848 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1624635492
transform -1 0 17112 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1624635492
transform -1 0 18860 0 -1 14688
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 13608 800 13728 6 REGIN_FEEDTHROUGH
port 0 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 REGOUT_FEEDTHROUGH
port 1 nsew signal tristate
rlabel metal2 s 16670 0 16726 800 6 SC_IN_BOT
port 2 nsew signal input
rlabel metal2 s 1950 16400 2006 17200 6 SC_IN_TOP
port 3 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 SC_OUT_BOT
port 4 nsew signal tristate
rlabel metal2 s 5906 16400 5962 17200 6 SC_OUT_TOP
port 5 nsew signal tristate
rlabel metal2 s 2134 0 2190 800 6 bottom_grid_pin_0_
port 6 nsew signal tristate
rlabel metal2 s 11242 0 11298 800 6 bottom_grid_pin_10_
port 7 nsew signal tristate
rlabel metal2 s 12162 0 12218 800 6 bottom_grid_pin_11_
port 8 nsew signal tristate
rlabel metal2 s 13082 0 13138 800 6 bottom_grid_pin_12_
port 9 nsew signal tristate
rlabel metal2 s 13910 0 13966 800 6 bottom_grid_pin_13_
port 10 nsew signal tristate
rlabel metal2 s 14830 0 14886 800 6 bottom_grid_pin_14_
port 11 nsew signal tristate
rlabel metal2 s 15750 0 15806 800 6 bottom_grid_pin_15_
port 12 nsew signal tristate
rlabel metal2 s 3054 0 3110 800 6 bottom_grid_pin_1_
port 13 nsew signal tristate
rlabel metal2 s 3974 0 4030 800 6 bottom_grid_pin_2_
port 14 nsew signal tristate
rlabel metal2 s 4894 0 4950 800 6 bottom_grid_pin_3_
port 15 nsew signal tristate
rlabel metal2 s 5814 0 5870 800 6 bottom_grid_pin_4_
port 16 nsew signal tristate
rlabel metal2 s 6734 0 6790 800 6 bottom_grid_pin_5_
port 17 nsew signal tristate
rlabel metal2 s 7562 0 7618 800 6 bottom_grid_pin_6_
port 18 nsew signal tristate
rlabel metal2 s 8482 0 8538 800 6 bottom_grid_pin_7_
port 19 nsew signal tristate
rlabel metal2 s 9402 0 9458 800 6 bottom_grid_pin_8_
port 20 nsew signal tristate
rlabel metal2 s 10322 0 10378 800 6 bottom_grid_pin_9_
port 21 nsew signal tristate
rlabel metal2 s 386 0 442 800 6 ccff_head
port 22 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 ccff_tail
port 23 nsew signal tristate
rlabel metal3 s 0 6672 800 6792 6 chanx_left_in[0]
port 24 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 chanx_left_in[10]
port 25 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[11]
port 26 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 chanx_left_in[12]
port 27 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[13]
port 28 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[14]
port 29 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 chanx_left_in[15]
port 30 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 chanx_left_in[16]
port 31 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[17]
port 32 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 chanx_left_in[18]
port 33 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 chanx_left_in[19]
port 34 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 chanx_left_in[1]
port 35 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 chanx_left_in[2]
port 36 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 chanx_left_in[3]
port 37 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[4]
port 38 nsew signal input
rlabel metal3 s 0 8304 800 8424 6 chanx_left_in[5]
port 39 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 chanx_left_in[6]
port 40 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[7]
port 41 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 chanx_left_in[8]
port 42 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 chanx_left_in[9]
port 43 nsew signal input
rlabel metal3 s 0 144 800 264 6 chanx_left_out[0]
port 44 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 chanx_left_out[10]
port 45 nsew signal tristate
rlabel metal3 s 0 3680 800 3800 6 chanx_left_out[11]
port 46 nsew signal tristate
rlabel metal3 s 0 4088 800 4208 6 chanx_left_out[12]
port 47 nsew signal tristate
rlabel metal3 s 0 4360 800 4480 6 chanx_left_out[13]
port 48 nsew signal tristate
rlabel metal3 s 0 4632 800 4752 6 chanx_left_out[14]
port 49 nsew signal tristate
rlabel metal3 s 0 5040 800 5160 6 chanx_left_out[15]
port 50 nsew signal tristate
rlabel metal3 s 0 5312 800 5432 6 chanx_left_out[16]
port 51 nsew signal tristate
rlabel metal3 s 0 5720 800 5840 6 chanx_left_out[17]
port 52 nsew signal tristate
rlabel metal3 s 0 5992 800 6112 6 chanx_left_out[18]
port 53 nsew signal tristate
rlabel metal3 s 0 6400 800 6520 6 chanx_left_out[19]
port 54 nsew signal tristate
rlabel metal3 s 0 416 800 536 6 chanx_left_out[1]
port 55 nsew signal tristate
rlabel metal3 s 0 688 800 808 6 chanx_left_out[2]
port 56 nsew signal tristate
rlabel metal3 s 0 1096 800 1216 6 chanx_left_out[3]
port 57 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 chanx_left_out[4]
port 58 nsew signal tristate
rlabel metal3 s 0 1776 800 1896 6 chanx_left_out[5]
port 59 nsew signal tristate
rlabel metal3 s 0 2048 800 2168 6 chanx_left_out[6]
port 60 nsew signal tristate
rlabel metal3 s 0 2320 800 2440 6 chanx_left_out[7]
port 61 nsew signal tristate
rlabel metal3 s 0 2728 800 2848 6 chanx_left_out[8]
port 62 nsew signal tristate
rlabel metal3 s 0 3000 800 3120 6 chanx_left_out[9]
port 63 nsew signal tristate
rlabel metal3 s 19200 9664 20000 9784 6 chanx_right_in[0]
port 64 nsew signal input
rlabel metal3 s 19200 13472 20000 13592 6 chanx_right_in[10]
port 65 nsew signal input
rlabel metal3 s 19200 13744 20000 13864 6 chanx_right_in[11]
port 66 nsew signal input
rlabel metal3 s 19200 14152 20000 14272 6 chanx_right_in[12]
port 67 nsew signal input
rlabel metal3 s 19200 14560 20000 14680 6 chanx_right_in[13]
port 68 nsew signal input
rlabel metal3 s 19200 14968 20000 15088 6 chanx_right_in[14]
port 69 nsew signal input
rlabel metal3 s 19200 15376 20000 15496 6 chanx_right_in[15]
port 70 nsew signal input
rlabel metal3 s 19200 15648 20000 15768 6 chanx_right_in[16]
port 71 nsew signal input
rlabel metal3 s 19200 16056 20000 16176 6 chanx_right_in[17]
port 72 nsew signal input
rlabel metal3 s 19200 16464 20000 16584 6 chanx_right_in[18]
port 73 nsew signal input
rlabel metal3 s 19200 16872 20000 16992 6 chanx_right_in[19]
port 74 nsew signal input
rlabel metal3 s 19200 9936 20000 10056 6 chanx_right_in[1]
port 75 nsew signal input
rlabel metal3 s 19200 10344 20000 10464 6 chanx_right_in[2]
port 76 nsew signal input
rlabel metal3 s 19200 10752 20000 10872 6 chanx_right_in[3]
port 77 nsew signal input
rlabel metal3 s 19200 11160 20000 11280 6 chanx_right_in[4]
port 78 nsew signal input
rlabel metal3 s 19200 11568 20000 11688 6 chanx_right_in[5]
port 79 nsew signal input
rlabel metal3 s 19200 11840 20000 11960 6 chanx_right_in[6]
port 80 nsew signal input
rlabel metal3 s 19200 12248 20000 12368 6 chanx_right_in[7]
port 81 nsew signal input
rlabel metal3 s 19200 12656 20000 12776 6 chanx_right_in[8]
port 82 nsew signal input
rlabel metal3 s 19200 13064 20000 13184 6 chanx_right_in[9]
port 83 nsew signal input
rlabel metal3 s 19200 2048 20000 2168 6 chanx_right_out[0]
port 84 nsew signal tristate
rlabel metal3 s 19200 5856 20000 5976 6 chanx_right_out[10]
port 85 nsew signal tristate
rlabel metal3 s 19200 6128 20000 6248 6 chanx_right_out[11]
port 86 nsew signal tristate
rlabel metal3 s 19200 6536 20000 6656 6 chanx_right_out[12]
port 87 nsew signal tristate
rlabel metal3 s 19200 6944 20000 7064 6 chanx_right_out[13]
port 88 nsew signal tristate
rlabel metal3 s 19200 7352 20000 7472 6 chanx_right_out[14]
port 89 nsew signal tristate
rlabel metal3 s 19200 7760 20000 7880 6 chanx_right_out[15]
port 90 nsew signal tristate
rlabel metal3 s 19200 8032 20000 8152 6 chanx_right_out[16]
port 91 nsew signal tristate
rlabel metal3 s 19200 8440 20000 8560 6 chanx_right_out[17]
port 92 nsew signal tristate
rlabel metal3 s 19200 8848 20000 8968 6 chanx_right_out[18]
port 93 nsew signal tristate
rlabel metal3 s 19200 9256 20000 9376 6 chanx_right_out[19]
port 94 nsew signal tristate
rlabel metal3 s 19200 2320 20000 2440 6 chanx_right_out[1]
port 95 nsew signal tristate
rlabel metal3 s 19200 2728 20000 2848 6 chanx_right_out[2]
port 96 nsew signal tristate
rlabel metal3 s 19200 3136 20000 3256 6 chanx_right_out[3]
port 97 nsew signal tristate
rlabel metal3 s 19200 3544 20000 3664 6 chanx_right_out[4]
port 98 nsew signal tristate
rlabel metal3 s 19200 3952 20000 4072 6 chanx_right_out[5]
port 99 nsew signal tristate
rlabel metal3 s 19200 4224 20000 4344 6 chanx_right_out[6]
port 100 nsew signal tristate
rlabel metal3 s 19200 4632 20000 4752 6 chanx_right_out[7]
port 101 nsew signal tristate
rlabel metal3 s 19200 5040 20000 5160 6 chanx_right_out[8]
port 102 nsew signal tristate
rlabel metal3 s 19200 5448 20000 5568 6 chanx_right_out[9]
port 103 nsew signal tristate
rlabel metal2 s 9862 16400 9918 17200 6 clk_1_N_out
port 104 nsew signal tristate
rlabel metal2 s 18510 0 18566 800 6 clk_1_S_out
port 105 nsew signal tristate
rlabel metal3 s 0 16872 800 16992 6 clk_1_W_in
port 106 nsew signal input
rlabel metal3 s 19200 1640 20000 1760 6 clk_2_E_out
port 107 nsew signal tristate
rlabel metal3 s 0 16600 800 16720 6 clk_2_W_in
port 108 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 clk_2_W_out
port 109 nsew signal tristate
rlabel metal3 s 19200 1232 20000 1352 6 clk_3_E_out
port 110 nsew signal tristate
rlabel metal3 s 0 16192 800 16312 6 clk_3_W_in
port 111 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 clk_3_W_out
port 112 nsew signal tristate
rlabel metal2 s 13910 16400 13966 17200 6 prog_clk_0_N_in
port 113 nsew signal input
rlabel metal2 s 17866 16400 17922 17200 6 prog_clk_0_W_out
port 114 nsew signal tristate
rlabel metal3 s 19200 824 20000 944 6 prog_clk_1_N_out
port 115 nsew signal tristate
rlabel metal2 s 19430 0 19486 800 6 prog_clk_1_S_out
port 116 nsew signal tristate
rlabel metal3 s 0 15920 800 16040 6 prog_clk_1_W_in
port 117 nsew signal input
rlabel metal3 s 19200 416 20000 536 6 prog_clk_2_E_out
port 118 nsew signal tristate
rlabel metal3 s 0 15512 800 15632 6 prog_clk_2_W_in
port 119 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 prog_clk_2_W_out
port 120 nsew signal tristate
rlabel metal3 s 19200 144 20000 264 6 prog_clk_3_E_out
port 121 nsew signal tristate
rlabel metal3 s 0 15240 800 15360 6 prog_clk_3_W_in
port 122 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 prog_clk_3_W_out
port 123 nsew signal tristate
rlabel metal4 s 15771 2128 16091 14736 6 VPWR
port 124 nsew power bidirectional
rlabel metal4 s 9840 2128 10160 14736 6 VPWR
port 125 nsew power bidirectional
rlabel metal4 s 3909 2128 4229 14736 6 VPWR
port 126 nsew power bidirectional
rlabel metal4 s 12805 2128 13125 14736 6 VGND
port 127 nsew ground bidirectional
rlabel metal4 s 6875 2128 7195 14736 6 VGND
port 128 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 17200
<< end >>
