* NGSPICE file created from left_tile.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

.subckt left_tile VGND VPWR ccff_head ccff_head_0 ccff_tail ccff_tail_0 chanx_right_in[0]
+ chanx_right_in[10] chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14]
+ chanx_right_in[15] chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19]
+ chanx_right_in[1] chanx_right_in[20] chanx_right_in[21] chanx_right_in[22] chanx_right_in[23]
+ chanx_right_in[24] chanx_right_in[25] chanx_right_in[26] chanx_right_in[27] chanx_right_in[28]
+ chanx_right_in[29] chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5]
+ chanx_right_in[6] chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0]
+ chanx_right_out[10] chanx_right_out[11] chanx_right_out[12] chanx_right_out[13]
+ chanx_right_out[14] chanx_right_out[15] chanx_right_out[16] chanx_right_out[17]
+ chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[20] chanx_right_out[21]
+ chanx_right_out[22] chanx_right_out[23] chanx_right_out[24] chanx_right_out[25]
+ chanx_right_out[26] chanx_right_out[27] chanx_right_out[28] chanx_right_out[29]
+ chanx_right_out[2] chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6]
+ chanx_right_out[7] chanx_right_out[8] chanx_right_out[9] chany_bottom_in[0] chany_bottom_in[10]
+ chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14]
+ chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18]
+ chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[20] chany_bottom_in[21] chany_bottom_in[22]
+ chany_bottom_in[23] chany_bottom_in[24] chany_bottom_in[25] chany_bottom_in[26]
+ chany_bottom_in[27] chany_bottom_in[28] chany_bottom_in[29] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[20] chany_bottom_out[21] chany_bottom_out[22]
+ chany_bottom_out[23] chany_bottom_out[24] chany_bottom_out[25] chany_bottom_out[26]
+ chany_bottom_out[27] chany_bottom_out[28] chany_bottom_out[29] chany_bottom_out[2]
+ chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6]
+ chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9] chany_top_in_0[0] chany_top_in_0[10]
+ chany_top_in_0[11] chany_top_in_0[12] chany_top_in_0[13] chany_top_in_0[14] chany_top_in_0[15]
+ chany_top_in_0[16] chany_top_in_0[17] chany_top_in_0[18] chany_top_in_0[19] chany_top_in_0[1]
+ chany_top_in_0[20] chany_top_in_0[21] chany_top_in_0[22] chany_top_in_0[23] chany_top_in_0[24]
+ chany_top_in_0[25] chany_top_in_0[26] chany_top_in_0[27] chany_top_in_0[28] chany_top_in_0[29]
+ chany_top_in_0[2] chany_top_in_0[3] chany_top_in_0[4] chany_top_in_0[5] chany_top_in_0[6]
+ chany_top_in_0[7] chany_top_in_0[8] chany_top_in_0[9] chany_top_out_0[0] chany_top_out_0[10]
+ chany_top_out_0[11] chany_top_out_0[12] chany_top_out_0[13] chany_top_out_0[14]
+ chany_top_out_0[15] chany_top_out_0[16] chany_top_out_0[17] chany_top_out_0[18]
+ chany_top_out_0[19] chany_top_out_0[1] chany_top_out_0[20] chany_top_out_0[21] chany_top_out_0[22]
+ chany_top_out_0[23] chany_top_out_0[24] chany_top_out_0[25] chany_top_out_0[26]
+ chany_top_out_0[27] chany_top_out_0[28] chany_top_out_0[29] chany_top_out_0[2] chany_top_out_0[3]
+ chany_top_out_0[4] chany_top_out_0[5] chany_top_out_0[6] chany_top_out_0[7] chany_top_out_0[8]
+ chany_top_out_0[9] gfpga_pad_io_soc_dir[0] gfpga_pad_io_soc_dir[1] gfpga_pad_io_soc_dir[2]
+ gfpga_pad_io_soc_dir[3] gfpga_pad_io_soc_in[0] gfpga_pad_io_soc_in[1] gfpga_pad_io_soc_in[2]
+ gfpga_pad_io_soc_in[3] gfpga_pad_io_soc_out[0] gfpga_pad_io_soc_out[1] gfpga_pad_io_soc_out[2]
+ gfpga_pad_io_soc_out[3] isol_n prog_clk prog_reset_bottom_in prog_reset_bottom_out
+ prog_reset_left_in prog_reset_right_out prog_reset_top_in prog_reset_top_out reset_bottom_in
+ reset_bottom_out reset_right_in reset_top_in reset_top_out right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_ right_width_0_height_0_subtile_0__pin_inpad_0_
+ right_width_0_height_0_subtile_1__pin_inpad_0_ right_width_0_height_0_subtile_2__pin_inpad_0_
+ right_width_0_height_0_subtile_3__pin_inpad_0_ test_enable_bottom_in test_enable_bottom_out
+ test_enable_right_in test_enable_top_in test_enable_top_out top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
+ top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_ top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
+ top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4_ net65 net34 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l4_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X cby_0__1_.cby_0__1_.mem_right_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xcby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_74_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_9_0_prog_clk sb_0__1_.mem_right_track_22.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_22.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_14.out sky130_fd_sc_hd__clkbuf_1
XFILLER_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput220 net220 VGND VGND VPWR VPWR prog_reset_top_out sky130_fd_sc_hd__buf_12
XFILLER_59_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk sb_0__1_.mem_right_track_54.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_54.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_90_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__272 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__272/HI
+ net272 sky130_fd_sc_hd__conb_1
X_200_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_131_ sb_0__1_.mux_right_track_12.out VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_8.mux_l1_in_0_ net73 net80 sb_0__1_.mem_right_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_2_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l3_in_1_ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_11.mux_l1_in_0_ net88 net73 sb_0__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_37_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_114_ sb_0__1_.mux_right_track_46.out VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_right_track_14.mux_l3_in_0_ sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_right_track_14.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_56.mux_l1_in_0_ net54 net110 sb_0__1_.mem_right_track_56.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_57_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2_ net57 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_45.mux_l2_in_1__227 VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_45.mux_l2_in_1__227/HI
+ net227 sky130_fd_sc_hd__conb_1
XANTENNA_5 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_45.out sky130_fd_sc_hd__clkbuf_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_5_0_prog_clk sb_0__1_.mem_top_track_10.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_95_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_14.mux_l2_in_1_ net234 net39 sb_0__1_.mem_right_track_14.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3_ net71 net40 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_24.mux_l1_in_1__240 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_24.mux_l1_in_1__240/HI
+ net240 sky130_fd_sc_hd__conb_1
XFILLER_77_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_6.mux_l2_in_1__257 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_6.mux_l2_in_1__257/HI
+ net257 sky130_fd_sc_hd__conb_1
XFILLER_67_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_1_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_1.ccff_tail net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_55_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk sb_0__1_.mem_right_track_22.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_22.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_6_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_6_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_12.mux_l3_in_0_ sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_top_track_12.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_20_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput210 net210 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[0] sky130_fd_sc_hd__buf_12
Xoutput221 net221 VGND VGND VPWR VPWR reset_bottom_out sky130_fd_sc_hd__buf_12
XFILLER_58_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk sb_0__1_.mem_right_track_52.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_54.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_130_ sb_0__1_.mux_right_track_14.out VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_top_track_6.mux_l1_in_3_ net269 net59 sb_0__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_7_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_36.out sky130_fd_sc_hd__clkbuf_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l3_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_93_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_36.mux_l2_in_1__265 VGND VGND VPWR VPWR sb_0__1_.mux_top_track_36.mux_l2_in_1__265/HI
+ net265 sky130_fd_sc_hd__conb_1
XFILLER_85_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_113_ sb_0__1_.mux_right_track_48.out VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_12.mux_l2_in_1_ net261 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_top_track_12.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_66_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_1_ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_6 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_6.mux_l3_in_0_ sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X
+ sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X sb_0__1_.mem_top_track_10.ccff_head
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_89_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_12.mux_l1_in_2_ net56 net42 sb_0__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_0__1_.mem_top_track_10.ccff_head
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xinput110 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_ VGND VGND VPWR
+ VPWR net110 sky130_fd_sc_hd__buf_2
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_14.mux_l2_in_0_ net105 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_14.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_3.out sky130_fd_sc_hd__clkbuf_1
XFILLER_79_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2_ net78 net47 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_top_track_6.mux_l2_in_1_ sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_95_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk sb_0__1_.mem_right_track_20.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_22.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput200 net200 VGND VGND VPWR VPWR chany_top_out_0[28] sky130_fd_sc_hd__buf_12
Xoutput222 net222 VGND VGND VPWR VPWR reset_top_out sky130_fd_sc_hd__buf_12
Xoutput211 net211 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[1] sky130_fd_sc_hd__buf_12
XFILLER_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_6.mux_l1_in_2_ net46 net26 sb_0__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_189_ net47 VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_2
XFILLER_89_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_112_ sb_0__1_.mux_right_track_50.out VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk sb_0__1_.mem_right_track_28.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_78_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_top_track_12.mux_l2_in_0_ sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_93_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_7 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_12.mux_l1_in_1_ net14 net6 sb_0__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput100 prog_reset_top_in VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
XFILLER_95_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput111 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_ VGND VGND VPWR
+ VPWR net111 sky130_fd_sc_hd__buf_2
XFILLER_76_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_9_0_prog_clk sb_0__1_.mem_bottom_track_11.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_ net81 net50 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_top_track_6.mux_l2_in_0_ sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_10_0_prog_clk sb_0__1_.mem_bottom_track_5.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_58_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_14.mux_l1_in_0_ net69 net70 sb_0__1_.mem_right_track_14.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xleft_tile_270 VGND VGND VPWR VPWR left_tile_270/HI chanx_right_out[0] sky130_fd_sc_hd__conb_1
XFILLER_46_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_26.mux_l2_in_0_ sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_26.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_76_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput201 net201 VGND VGND VPWR VPWR chany_top_out_0[29] sky130_fd_sc_hd__buf_12
Xoutput223 net223 VGND VGND VPWR VPWR test_enable_bottom_out sky130_fd_sc_hd__buf_12
Xoutput212 net212 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[2] sky130_fd_sc_hd__buf_12
XFILLER_74_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_top_track_6.mux_l1_in_1_ net8 net20 sb_0__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_11_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_188_ net46 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_2
XFILLER_89_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_3.mux_l3_in_0_ sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_bottom_track_3.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_83_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_111_ sb_0__1_.mux_right_track_52.out VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_26.mux_l1_in_1_ net241 net60 sb_0__1_.mem_right_track_26.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_50_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_6_0_prog_clk sb_0__1_.mem_right_track_26.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_3_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_8 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_bottom_track_3.mux_l2_in_1_ net225 right_width_0_height_0_subtile_1__pin_inpad_0_
+ sb_0__1_.mem_bottom_track_3.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk sb_0__1_.mem_right_track_40.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_40.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_21_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_top_track_12.mux_l1_in_0_ net18 net115 sb_0__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_5_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput101 reset_bottom_in VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__buf_2
Xinput112 test_enable_bottom_in VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__buf_2
XFILLER_48_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk sb_0__1_.mem_bottom_track_11.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_ sb_0__1_.mux_bottom_track_3.out
+ net53 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_36.mux_l3_in_0_ sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_top_track_36.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_89_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net94 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR right_width_0_height_0_subtile_2__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_10_0_prog_clk sb_0__1_.mem_bottom_track_5.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_top_track_36.mux_l2_in_1_ net265 net38 sb_0__1_.mem_top_track_36.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_32_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput224 net224 VGND VGND VPWR VPWR test_enable_top_out sky130_fd_sc_hd__buf_12
Xoutput202 net202 VGND VGND VPWR VPWR chany_top_out_0[2] sky130_fd_sc_hd__buf_12
Xoutput213 net213 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[3] sky130_fd_sc_hd__buf_12
XFILLER_87_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_6.mux_l1_in_0_ net117 net115 sb_0__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_11_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ net119 net97 VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
XFILLER_80_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_187_ sb_0__1_.mux_top_track_20.out VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_4.mux_l3_in_0_ sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_right_track_4.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_5_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_5_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_51_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_110_ sb_0__1_.mux_right_track_54.out VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_2
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_26.mux_l1_in_0_ net111 net90 sb_0__1_.mem_right_track_26.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_38.mux_l2_in_0_ net247 sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_38.ccff_tail VGND VGND VPWR VPWR sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_40.mux_l2_in_0_ net249 sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_40.ccff_tail VGND VGND VPWR VPWR sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_9 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_4.mux_l2_in_1_ net248 net47 sb_0__1_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_62_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
Xsb_0__1_.mux_bottom_track_3.mux_l2_in_0_ sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk sb_0__1_.mem_right_track_38.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_40.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput102 reset_right_in VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_1
Xinput113 test_enable_right_in VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk sb_0__1_.mem_bottom_track_11.ccff_head
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_right_track_36.mux_l2_in_1__246 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_36.mux_l2_in_1__246/HI
+ net246 sky130_fd_sc_hd__conb_1
XFILLER_50_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_13_0_prog_clk sb_0__1_.mem_right_track_14.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_14.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_49_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_3.mux_l1_in_1_ net4 net16 sb_0__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_32_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_20.out sky130_fd_sc_hd__clkbuf_1
XFILLER_94_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_3_0_prog_clk sb_0__1_.mem_bottom_track_3.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk sb_0__1_.mem_right_track_46.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_46.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_78_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_36.mux_l2_in_0_ net32 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_top_track_36.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput203 net203 VGND VGND VPWR VPWR chany_top_out_0[3] sky130_fd_sc_hd__buf_12
Xoutput214 net214 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[0] sky130_fd_sc_hd__buf_12
XFILLER_87_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_186_ net43 VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_2
XFILLER_37_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_169_ net55 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_2
XFILLER_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail net97 VGND
+ VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_11_0_prog_clk sb_0__1_.mem_right_track_0.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_15_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_4.mux_l2_in_0_ sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput114 test_enable_top_in VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_1
Xinput103 reset_top_in VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_38.mux_l1_in_0_ net57 net109 sb_0__1_.mem_right_track_38.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_44_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_40.mux_l1_in_0_ net61 net110 sb_0__1_.mem_right_track_40.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_52.mux_l2_in_0_ net254 sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_52.ccff_tail VGND VGND VPWR VPWR sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_4.mux_l1_in_1_ net109 net106 sb_0__1_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_67_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_14.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_14.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_29_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_3.mux_l1_in_0_ net92 net78 sb_0__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_17_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk sb_0__1_.mem_right_track_44.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_46.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_68_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_4_0_prog_clk cby_0__1_.cby_0__1_.ccff_tail net98 VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput204 net204 VGND VGND VPWR VPWR chany_top_out_0[4] sky130_fd_sc_hd__buf_12
Xoutput215 net215 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[1] sky130_fd_sc_hd__buf_12
XFILLER_87_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_13.out sky130_fd_sc_hd__clkbuf_2
XFILLER_95_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_185_ net42 VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_36.mux_l1_in_0_ net15 net118 sb_0__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_56.mux_l2_in_0__256 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_56.mux_l2_in_0__256/HI
+ net256 sky130_fd_sc_hd__conb_1
XFILLER_59_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_168_ net44 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_12_0_prog_clk sb_0__1_.mem_top_track_52.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_0.ccff_head sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_36.out sky130_fd_sc_hd__clkbuf_1
XFILLER_69_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_10.out sky130_fd_sc_hd__clkbuf_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_11_0_prog_clk sb_0__1_.mem_right_track_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_20.mux_l2_in_1__263 VGND VGND VPWR VPWR sb_0__1_.mux_top_track_20.mux_l2_in_1__263/HI
+ net263 sky130_fd_sc_hd__conb_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput104 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ VGND VGND VPWR
+ VPWR net104 sky130_fd_sc_hd__buf_2
Xinput115 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND VPWR
+ VPWR net115 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3_ net273 sb_0__1_.mux_bottom_track_53.out
+ cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_12.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_14.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_right_track_4.mux_l1_in_0_ net77 net83 sb_0__1_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_67_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_12_0_prog_clk sb_0__1_.mem_top_track_4.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_91_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_6.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_6.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_bottom_track_29.mux_l3_in_0_ sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_bottom_track_29.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4_ net64 net62 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput205 net205 VGND VGND VPWR VPWR chany_top_out_0[5] sky130_fd_sc_hd__buf_12
Xoutput216 net216 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[2] sky130_fd_sc_hd__buf_12
Xsb_0__1_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_8.out sky130_fd_sc_hd__clkbuf_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_52.mux_l1_in_0_ net52 net108 sb_0__1_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_10.mux_l3_in_0_ sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_right_track_10.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_63_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_184_ net41 VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_2
XFILLER_89_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l4_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cby_0__1_.cby_0__1_.mem_right_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_5_0_prog_clk sb_0__1_.mem_top_track_20.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_20.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_92_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_29.mux_l2_in_1_ net279 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_bottom_track_29.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_18.mux_l2_in_1__236 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_18.mux_l2_in_1__236/HI
+ net236 sky130_fd_sc_hd__conb_1
XFILLER_87_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_167_ sb_0__1_.mux_bottom_track_1.out VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_10.mux_l2_in_1_ net232 net42 sb_0__1_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk sb_0__1_.mem_top_track_52.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_52.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_69_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l3_in_1_ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_29.mux_l1_in_2_ right_width_0_height_0_subtile_2__pin_inpad_0_
+ net28 sb_0__1_.mem_bottom_track_29.mem_out\[0\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_0.ccff_head
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_4_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_4_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_29.out sky130_fd_sc_hd__clkbuf_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput105 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_ VGND VGND VPWR
+ VPWR net105 sky130_fd_sc_hd__buf_2
Xinput116 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_ VGND VGND VPWR
+ VPWR net116 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_32.out sky130_fd_sc_hd__clkbuf_1
XFILLER_44_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2_ net56 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk sb_0__1_.mem_top_track_4.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_91_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_4.mux_l2_in_1__266 VGND VGND VPWR VPWR sb_0__1_.mux_top_track_4.mux_l2_in_1__266/HI
+ net266 sky130_fd_sc_hd__conb_1
XFILLER_23_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_26.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_26.out sky130_fd_sc_hd__clkbuf_1
XFILLER_31_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_6.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3_ sb_0__1_.mux_bottom_track_29.out
+ net39 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xoutput206 net206 VGND VGND VPWR VPWR chany_top_out_0[6] sky130_fd_sc_hd__buf_12
Xoutput217 net217 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[3] sky130_fd_sc_hd__buf_12
XFILLER_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_183_ sb_0__1_.mux_top_track_28.out VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_7_0_prog_clk sb_0__1_.mem_top_track_20.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_20.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_77_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_29.mux_l2_in_0_ sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_92_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_top_track_2.mux_l3_in_0_ sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_top_track_2.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_87_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_166_ sb_0__1_.mux_bottom_track_3.out VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_10.mux_l2_in_0_ sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_13_0_prog_clk sb_0__1_.mem_top_track_44.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_52.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_22.mux_l3_in_0_ sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_right_track_22.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_16_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l3_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_29.mux_l1_in_1_ net10 net22 sb_0__1_.mem_bottom_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_7_0_prog_clk sb_0__1_.mem_right_track_32.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_32.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_2.mux_l2_in_1_ net262 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_top_track_2.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_218_ net112 VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_2
X_149_ sb_0__1_.mux_bottom_track_37.out VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput117 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_ VGND VGND VPWR
+ VPWR net117 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput106 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_ VGND VGND VPWR
+ VPWR net106 sky130_fd_sc_hd__buf_2
XFILLER_88_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_10.mux_l1_in_1_ net109 net106 sb_0__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_22.mux_l2_in_1_ net239 net34 sb_0__1_.mem_right_track_22.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_30_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1_ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_2.mux_l1_in_2_ net62 net48 sb_0__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_1_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk sb_0__1_.mem_top_track_2.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_76_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_54.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_54.out sky130_fd_sc_hd__clkbuf_1
XFILLER_12_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_4.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_22.mux_l2_in_1__239 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_22.mux_l2_in_1__239/HI
+ net239 sky130_fd_sc_hd__conb_1
XFILLER_1_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2_ net77 net46 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput207 net207 VGND VGND VPWR VPWR chany_top_out_0[7] sky130_fd_sc_hd__buf_12
Xoutput218 net218 VGND VGND VPWR VPWR prog_reset_bottom_out sky130_fd_sc_hd__buf_12
XFILLER_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_20.mux_l3_in_0_ sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_top_track_20.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_48.out sky130_fd_sc_hd__clkbuf_1
XFILLER_48_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_182_ net39 VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_2
XFILLER_89_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_9_0_prog_clk sb_0__1_.mem_top_track_12.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_20.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_92_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_165_ sb_0__1_.mux_bottom_track_5.out VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_20.mux_l2_in_1_ net263 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_top_track_20.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_29.mux_l1_in_0_ net74 net69 sb_0__1_.mem_bottom_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_6_0_prog_clk sb_0__1_.mem_right_track_30.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_32.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_2.mux_l2_in_0_ sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_74_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_217_ net112 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_1
X_148_ net65 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_2
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput118 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_ VGND VGND VPWR
+ VPWR net118 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput107 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_ VGND VGND VPWR
+ VPWR net107 sky130_fd_sc_hd__buf_2
XFILLER_56_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_10.mux_l1_in_0_ net72 net79 sb_0__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_top_track_20.mux_l1_in_2_ net55 net41 sb_0__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_4_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_1_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[2\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_22.mux_l2_in_0_ net109 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_22.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_top_track_52.mux_l2_in_1__268 VGND VGND VPWR VPWR sb_0__1_.mux_top_track_52.mux_l2_in_1__268/HI
+ net268 sky130_fd_sc_hd__conb_1
XFILLER_85_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_2.mux_l1_in_1_ net28 net10 sb_0__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_88_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_38.mux_l2_in_0__247 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_38.mux_l2_in_0__247/HI
+ net247 sky130_fd_sc_hd__conb_1
XFILLER_17_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_4.mux_l2_in_1__248 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_4.mux_l2_in_1__248/HI
+ net248 sky130_fd_sc_hd__conb_1
XFILLER_12_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk sb_0__1_.mem_right_track_38.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_38.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_75_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_ sb_0__1_.mux_bottom_track_11.out
+ net49 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput208 net208 VGND VGND VPWR VPWR chany_top_out_0[8] sky130_fd_sc_hd__buf_12
Xoutput219 net219 VGND VGND VPWR VPWR prog_reset_right_out sky130_fd_sc_hd__buf_12
XFILLER_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_181_ net38 VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_10_0_prog_clk sb_0__1_.mem_bottom_track_21.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_21.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_164_ sb_0__1_.mux_bottom_track_7.out VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_20.mux_l2_in_0_ sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_4.out sky130_fd_sc_hd__clkbuf_1
XFILLER_45_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk sb_0__1_.mem_bottom_track_53.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dfrtp_4
XFILLER_56_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_216_ net112 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_1
X_147_ net64 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_2
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput108 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ VGND VGND VPWR
+ VPWR net108 sky130_fd_sc_hd__buf_2
XFILLER_84_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_20.mux_l1_in_1_ net3 net5 sb_0__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_1_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput90 chany_top_in_0[7] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_top_track_2.mux_l1_in_0_ net22 net116 sb_0__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_3_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_3_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_72_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_0_0_prog_clk sb_0__1_.mem_right_track_36.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_38.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_57_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_494 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_top_track_2.mux_l2_in_1__262 VGND VGND VPWR VPWR sb_0__1_.mux_top_track_2.mux_l2_in_1__262/HI
+ net262 sky130_fd_sc_hd__conb_1
XFILLER_7_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_0.mux_l3_in_0_ sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_right_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_54_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_22.mux_l1_in_0_ net63 net64 sb_0__1_.mem_right_track_22.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_ sb_0__1_.mux_bottom_track_5.out
+ net52 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput209 net209 VGND VGND VPWR VPWR chany_top_out_0[9] sky130_fd_sc_hd__buf_12
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_34.mux_l2_in_0_ sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_34.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_67_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_180_ net37 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_10_0_prog_clk sb_0__1_.mem_right_track_50.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_50.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_1_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_0.mux_l2_in_1_ net231 net51 sb_0__1_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_11_0_prog_clk sb_0__1_.mem_bottom_track_21.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_21.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_48_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_163_ net81 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_34.mux_l1_in_1_ net245 net55 sb_0__1_.mem_right_track_34.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_49_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk sb_0__1_.mem_bottom_track_45.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_53.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_56_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_215_ net112 VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_2
X_146_ net92 VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_2
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput109 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_ VGND VGND VPWR
+ VPWR net109 sky130_fd_sc_hd__clkbuf_4
XFILLER_29_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_20.mux_l1_in_0_ net17 net116 sb_0__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.out sky130_fd_sc_hd__clkbuf_1
XFILLER_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_129_ sb_0__1_.mux_right_track_16.out VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_2
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput80 chany_top_in_0[25] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_1
Xinput91 chany_top_in_0[8] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_5_0_prog_clk sb_0__1_.mem_top_track_12.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_86_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk sb_0__1_.mem_right_track_48.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_50.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_89_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_0.mux_l2_in_0_ sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_5_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk sb_0__1_.mem_bottom_track_13.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_21.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_83_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk sb_0__1_.mem_top_track_44.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_bottom_track_13.mux_l3_in_0_ sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_bottom_track_13.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_54.mux_l2_in_0__255 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_54.mux_l2_in_0__255/HI
+ net255 sky130_fd_sc_hd__conb_1
XFILLER_39_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_10.mux_l1_in_3__260 VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.mux_l1_in_3__260/HI
+ net260 sky130_fd_sc_hd__conb_1
XFILLER_10_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_162_ sb_0__1_.mux_bottom_track_11.out VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_34.mux_l1_in_0_ net107 net85 sb_0__1_.mem_right_track_34.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_40_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_46.mux_l2_in_0_ net251 sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_46.ccff_tail VGND VGND VPWR VPWR sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_0.mux_l1_in_3__259 VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.mux_l1_in_3__259/HI
+ net259 sky130_fd_sc_hd__conb_1
Xinput1 ccff_head VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_68_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_prog_clk prog_clk VGND VGND VPWR VPWR clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_0.mux_l1_in_1_ net110 net107 sb_0__1_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_214_ net101 VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_2
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_145_ sb_0__1_.mux_bottom_track_45.out VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_2
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_13.mux_l2_in_1_ net277 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_bottom_track_13.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk sb_0__1_.mem_right_track_56.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_1.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_38_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_29_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_4_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_0.ccff_tail net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_79_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput190 net190 VGND VGND VPWR VPWR chany_top_out_0[19] sky130_fd_sc_hd__buf_12
XFILLER_87_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_128_ sb_0__1_.mux_right_track_18.out VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_2
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput81 chany_top_in_0[26] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_4
Xinput70 chany_top_in_0[16] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_1
Xinput92 chany_top_in_0[9] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_2
XFILLER_69_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_0_0_prog_clk cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
+ net98 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dfrtp_4
XFILLER_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_13.mux_l1_in_2_ right_width_0_height_0_subtile_0__pin_inpad_0_
+ net26 sb_0__1_.mem_bottom_track_13.mem_out\[0\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_44.mux_l2_in_0_ sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_44.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_23_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_5_0_prog_clk sb_0__1_.mem_top_track_12.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_16.mux_l2_in_1__235 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_16.mux_l2_in_1__235/HI
+ net235 sky130_fd_sc_hd__conb_1
XFILLER_79_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_13_0_prog_clk sb_0__1_.mem_top_track_36.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_86_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_161_ sb_0__1_.mux_bottom_track_13.out VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_44.mux_l1_in_1_ net267 net37 sb_0__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_7_0_prog_clk sb_0__1_.mem_right_track_24.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_24.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput2 ccff_head_0 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_0.mux_l1_in_0_ net104 net81 sb_0__1_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_213_ net101 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_1
X_144_ net90 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_2
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_13.mux_l2_in_0_ sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_4.out sky130_fd_sc_hd__clkbuf_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk sb_0__1_.mem_right_track_54.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_56.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_40 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput191 net191 VGND VGND VPWR VPWR chany_top_out_0[1] sky130_fd_sc_hd__buf_12
Xoutput180 net180 VGND VGND VPWR VPWR chany_top_out_0[0] sky130_fd_sc_hd__buf_12
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_46.mux_l1_in_0_ net45 net105 sb_0__1_.mem_right_track_46.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_46_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_127_ sb_0__1_.mux_right_track_20.out VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_2
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput82 chany_top_in_0[27] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_1
Xinput71 chany_top_in_0[17] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_2
Xinput60 chany_bottom_in[7] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_4
Xinput93 gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_bottom_track_13.mux_l1_in_1_ net8 net20 sb_0__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_40_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_3_0_prog_clk sb_0__1_.mem_bottom_track_1.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3_ net274 net86 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_0__1_.mem_top_track_10.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_83_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_2_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_2_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_11_0_prog_clk sb_0__1_.mem_bottom_track_45.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_45.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_86_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_160_ net78 VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_44.mux_l1_in_0_ net31 net13 sb_0__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4_ net92 net61 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_9_0_prog_clk sb_0__1_.mem_right_track_22.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_24.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_73_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_22.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_22.out sky130_fd_sc_hd__clkbuf_1
XFILLER_5_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput3 chanx_right_in[0] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l4_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X cby_0__1_.cby_0__1_.ccff_tail
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_212_ net101 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_143_ net89 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_41 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_30 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput170 net170 VGND VGND VPWR VPWR chany_bottom_out[28] sky130_fd_sc_hd__buf_12
XFILLER_79_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput181 net181 VGND VGND VPWR VPWR chany_top_out_0[10] sky130_fd_sc_hd__buf_12
Xoutput192 net192 VGND VGND VPWR VPWR chany_top_out_0[20] sky130_fd_sc_hd__buf_12
Xsb_0__1_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_16.out sky130_fd_sc_hd__clkbuf_1
XFILLER_87_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_15_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_15_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_75_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_126_ sb_0__1_.mux_right_track_22.out VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_2
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_37.mux_l2_in_1__226 VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_37.mux_l2_in_1__226/HI
+ net226 sky130_fd_sc_hd__conb_1
XFILLER_34_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput72 chany_top_in_0[18] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_2
Xinput50 chany_bottom_in[25] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput61 chany_bottom_in[8] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_2
Xinput83 chany_top_in_0[28] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_1
Xinput94 gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l3_in_1_ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_bottom_track_13.mux_l1_in_0_ net86 net72 sb_0__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_40_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_109_ sb_0__1_.mux_right_track_56.out VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_37.mux_l3_in_0_ sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_bottom_track_37.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_right_track_20.mux_l2_in_1__238 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_20.mux_l2_in_1__238/HI
+ net238 sky130_fd_sc_hd__conb_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_53.out sky130_fd_sc_hd__clkbuf_2
XFILLER_69_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk sb_0__1_.mem_bottom_track_1.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_16.mux_l3_in_0_ sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_right_track_16.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_4_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2_ net55 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_8_0_prog_clk sb_0__1_.mem_bottom_track_13.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_22_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_bottom_track_37.mux_l2_in_1_ net226 right_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_0__1_.mem_bottom_track_37.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_11_0_prog_clk sb_0__1_.mem_bottom_track_45.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_45.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_16.mux_l2_in_1_ net235 net38 sb_0__1_.mem_right_track_16.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_50.out sky130_fd_sc_hd__clkbuf_1
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3_ net69 net38 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_10_0_prog_clk sb_0__1_.mem_bottom_track_7.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput4 chanx_right_in[10] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_28.mux_l2_in_1__264 VGND VGND VPWR VPWR sb_0__1_.mux_top_track_28.mux_l2_in_1__264/HI
+ net264 sky130_fd_sc_hd__conb_1
XFILLER_70_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_211_ net101 VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_142_ net88 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_2
XFILLER_51_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__273 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__273/HI
+ net273 sky130_fd_sc_hd__conb_1
Xsb_0__1_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_44.out sky130_fd_sc_hd__clkbuf_1
XFILLER_37_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_20 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_31 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput160 net160 VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_12
Xoutput193 net193 VGND VGND VPWR VPWR chany_top_out_0[21] sky130_fd_sc_hd__buf_12
Xoutput182 net182 VGND VGND VPWR VPWR chany_top_out_0[11] sky130_fd_sc_hd__buf_12
Xoutput171 net171 VGND VGND VPWR VPWR chany_bottom_out[29] sky130_fd_sc_hd__buf_12
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_125_ sb_0__1_.mux_right_track_24.out VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_2
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput40 chany_bottom_in[16] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_2
Xinput73 chany_top_in_0[19] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_2
Xinput51 chany_bottom_in[26] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_4
Xinput62 chany_bottom_in[9] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_4
Xinput84 chany_top_in_0[29] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_1
Xinput95 gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l3_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_38.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_38.out sky130_fd_sc_hd__clkbuf_1
XFILLER_16_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_10.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_73_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk sb_0__1_.mem_bottom_track_1.ccff_head
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1_ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk sb_0__1_.mem_bottom_track_13.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_13.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_22_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_5_0_prog_clk sb_0__1_.mem_top_track_36.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_36.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_89_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net95 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR right_width_0_height_0_subtile_1__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_37.mux_l2_in_0_ sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_37.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk sb_0__1_.mem_bottom_track_37.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_45.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_67_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_16.mux_l2_in_0_ net106 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_16.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2_ net76 net45 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk sb_0__1_.mem_bottom_track_7.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_68_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_5.out sky130_fd_sc_hd__clkbuf_1
XFILLER_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput5 chanx_right_in[11] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_210_ net98 VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__clkbuf_1
XFILLER_23_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_141_ sb_0__1_.mux_bottom_track_53.out VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_37.mux_l1_in_1_ net29 net11 sb_0__1_.mem_bottom_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_2_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_10 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput150 net150 VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_12
Xoutput161 net161 VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_12
Xoutput194 net194 VGND VGND VPWR VPWR chany_top_out_0[22] sky130_fd_sc_hd__buf_12
Xoutput183 net183 VGND VGND VPWR VPWR chany_top_out_0[12] sky130_fd_sc_hd__buf_12
Xoutput172 net172 VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_12
XFILLER_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_124_ sb_0__1_.mux_right_track_26.out VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_2
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput30 chanx_right_in[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
Xinput63 chany_top_in_0[0] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_1
Xinput52 chany_bottom_in[27] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput41 chany_bottom_in[17] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_4
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
Xinput85 chany_top_in_0[2] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_2
Xinput74 chany_top_in_0[1] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_2
Xinput96 gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_2.mux_l2_in_1__237 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_2.mux_l2_in_1__237/HI
+ net237 sky130_fd_sc_hd__conb_1
XFILLER_87_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.out sky130_fd_sc_hd__clkbuf_1
XFILLER_16_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_10.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk sb_0__1_.mem_bottom_track_11.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_54_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk sb_0__1_.mem_top_track_36.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_36.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_13_0_prog_clk sb_0__1_.mem_right_track_16.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_16.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_ sb_0__1_.mux_bottom_track_7.out
+ net51 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_1_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_1_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_73_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk sb_0__1_.mem_bottom_track_5.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_49_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput6 chanx_right_in[12] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_10_0_prog_clk sb_0__1_.mem_right_track_48.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_48.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_140_ net86 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_37.mux_l1_in_0_ net23 net68 sb_0__1_.mem_bottom_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_2_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_48.mux_l2_in_0__252 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_48.mux_l2_in_0__252/HI
+ net252 sky130_fd_sc_hd__conb_1
XFILLER_33_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_41_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_40.mux_l2_in_0__249 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_40.mux_l2_in_0__249/HI
+ net249 sky130_fd_sc_hd__conb_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_16.mux_l1_in_0_ net66 net68 sb_0__1_.mem_right_track_16.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_69_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_11 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_33 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput151 net151 VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_12
Xoutput140 net140 VGND VGND VPWR VPWR chanx_right_out[28] sky130_fd_sc_hd__buf_12
Xoutput195 net195 VGND VGND VPWR VPWR chany_top_out_0[23] sky130_fd_sc_hd__buf_12
Xoutput184 net184 VGND VGND VPWR VPWR chany_top_out_0[13] sky130_fd_sc_hd__buf_12
Xoutput173 net173 VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_12
Xoutput162 net162 VGND VGND VPWR VPWR chany_bottom_out[20] sky130_fd_sc_hd__buf_12
Xsb_0__1_.mux_right_track_28.mux_l2_in_0_ sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_28.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_123_ sb_0__1_.mux_right_track_28.out VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_30.mux_l2_in_0_ sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_30.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_61_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput31 chanx_right_in[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput20 chanx_right_in[25] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput64 chany_top_in_0[10] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_2
Xinput53 chany_bottom_in[28] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput42 chany_bottom_in[18] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_2
Xinput86 chany_top_in_0[3] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_2
Xinput75 chany_top_in_0[20] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_1
Xinput97 isol_n VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_2
XFILLER_29_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_0.mux_l2_in_1__231 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_0.mux_l2_in_1__231/HI
+ net231 sky130_fd_sc_hd__conb_1
XFILLER_0_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_10.ccff_head
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_31_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_13_0_prog_clk sb_0__1_.mem_top_track_0.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_bottom_track_5.mux_l3_in_0_ sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_bottom_track_5.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_14_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_14_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_30_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_28.mux_l1_in_1_ net242 net59 sb_0__1_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_89_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_2.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_84_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_30.mux_l1_in_1_ net243 net58 sb_0__1_.mem_right_track_30.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_48_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_0__1_.mem_top_track_28.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_36.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_bottom_track_5.mux_l2_in_1_ net228 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_bottom_track_5.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_16.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_16.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_86_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_52.mux_l2_in_0__254 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_52.mux_l2_in_0__254/HI
+ net254 sky130_fd_sc_hd__conb_1
XFILLER_6_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_ sb_0__1_.mux_bottom_track_1.out
+ net54 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput7 chanx_right_in[13] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk sb_0__1_.mem_right_track_46.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_48.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_5.mux_l1_in_2_ right_width_0_height_0_subtile_2__pin_inpad_0_
+ net3 sb_0__1_.mem_bottom_track_5.mem_out\[0\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_199_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_12 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput152 net152 VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_12
Xoutput130 net130 VGND VGND VPWR VPWR chanx_right_out[19] sky130_fd_sc_hd__buf_12
Xoutput141 net141 VGND VGND VPWR VPWR chanx_right_out[29] sky130_fd_sc_hd__buf_12
Xoutput185 net185 VGND VGND VPWR VPWR chany_top_out_0[14] sky130_fd_sc_hd__buf_12
Xoutput174 net174 VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_12
Xoutput163 net163 VGND VGND VPWR VPWR chany_bottom_out[21] sky130_fd_sc_hd__buf_12
Xoutput196 net196 VGND VGND VPWR VPWR chany_top_out_0[24] sky130_fd_sc_hd__buf_12
XFILLER_28_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_122_ sb_0__1_.mux_right_track_30.out VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
XFILLER_3_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput10 chanx_right_in[16] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
Xinput21 chanx_right_in[26] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput43 chany_bottom_in[19] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_2
Xinput54 chany_bottom_in[29] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput32 chanx_right_in[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput76 chany_top_in_0[21] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_2
Xinput65 chany_top_in_0[11] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_2
Xinput87 chany_top_in_0[4] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_1
Xinput98 prog_reset_bottom_in VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_16
XFILLER_57_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk sb_0__1_.mem_top_track_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_6.mux_l3_in_0_ sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_right_track_6.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_28.mux_l1_in_0_ net104 net89 sb_0__1_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_2.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_30.mux_l1_in_0_ net105 net88 sb_0__1_.mem_right_track_30.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_bottom_track_21.mux_l2_in_1__278 VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_21.mux_l2_in_1__278/HI
+ net278 sky130_fd_sc_hd__conb_1
XFILLER_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_6.mux_l2_in_1_ net257 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_right_track_6.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_9_0_prog_clk sb_0__1_.mem_bottom_track_37.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_37.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_bottom_track_5.mux_l2_in_0_ sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_14.mux_l2_in_1__234 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_14.mux_l2_in_1__234/HI
+ net234 sky130_fd_sc_hd__conb_1
XFILLER_63_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_14.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_16.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_12_0_prog_clk sb_0__1_.mem_top_track_6.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_8.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 chanx_right_in[14] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_6.mux_l1_in_2_ net46 net110 sb_0__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_34.mux_l1_in_1__245 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_34.mux_l1_in_1__245/HI
+ net245 sky130_fd_sc_hd__conb_1
XFILLER_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_5.mux_l1_in_1_ net5 net17 sb_0__1_.mem_bottom_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_67_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_198_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_13 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_24 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_35 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput120 net120 VGND VGND VPWR VPWR ccff_tail_0 sky130_fd_sc_hd__buf_12
Xoutput142 net142 VGND VGND VPWR VPWR chanx_right_out[2] sky130_fd_sc_hd__buf_12
Xoutput131 net131 VGND VGND VPWR VPWR chanx_right_out[1] sky130_fd_sc_hd__buf_12
Xoutput186 net186 VGND VGND VPWR VPWR chany_top_out_0[15] sky130_fd_sc_hd__buf_12
Xoutput175 net175 VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_12
Xoutput153 net153 VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_12
Xoutput164 net164 VGND VGND VPWR VPWR chany_bottom_out[22] sky130_fd_sc_hd__buf_12
Xoutput197 net197 VGND VGND VPWR VPWR chany_top_out_0[25] sky130_fd_sc_hd__buf_12
XFILLER_28_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_121_ sb_0__1_.mux_right_track_32.out VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput11 chanx_right_in[17] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput22 chanx_right_in[27] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput33 chany_bottom_in[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
Xinput44 chany_bottom_in[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_2
Xinput55 chany_bottom_in[2] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_4
Xinput77 chany_top_in_0[22] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_2
Xinput88 chany_top_in_0[5] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_2
Xinput66 chany_top_in_0[12] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_1
Xinput99 prog_reset_left_in VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_12.mux_l2_in_1__261 VGND VGND VPWR VPWR sb_0__1_.mux_top_track_12.mux_l2_in_1__261/HI
+ net261 sky130_fd_sc_hd__conb_1
XFILLER_37_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_52.mux_l3_in_0_ sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_right_track_0.ccff_head
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_57_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk net1 net98
+ VGND VGND VPWR VPWR sb_0__1_.mem_top_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk sb_0__1_.mem_right_track_0.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_27_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_0.out sky130_fd_sc_hd__clkbuf_1
XFILLER_75_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_top_track_52.mux_l2_in_1_ net268 net35 sb_0__1_.mem_top_track_52.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_6.mux_l2_in_0_ sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_13_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk sb_0__1_.mem_bottom_track_37.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_37.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_21_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk sb_0__1_.mem_top_track_6.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_79_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_21.mux_l3_in_0_ sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_bottom_track_21.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_50_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_8.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_8.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput9 chanx_right_in[15] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_54.mux_l2_in_0_ net255 sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_54.ccff_tail VGND VGND VPWR VPWR sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_6.mux_l1_in_1_ net107 net104 sb_0__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_87_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_5.mux_l1_in_0_ net90 net77 sb_0__1_.mem_bottom_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_82_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_21.out sky130_fd_sc_hd__clkbuf_1
XFILLER_73_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_197_ sb_0__1_.mux_top_track_0.out VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mux_bottom_track_21.mux_l2_in_1_ net278 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_bottom_track_21.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__271 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__271/HI
+ net271 sky130_fd_sc_hd__conb_1
XFILLER_2_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_14 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_25 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_36 sb_0__1_.mem_bottom_track_53.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_0_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_0_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xoutput121 net121 VGND VGND VPWR VPWR chanx_right_out[10] sky130_fd_sc_hd__buf_12
Xoutput143 net143 VGND VGND VPWR VPWR chanx_right_out[3] sky130_fd_sc_hd__buf_12
Xoutput132 net132 VGND VGND VPWR VPWR chanx_right_out[20] sky130_fd_sc_hd__buf_12
Xoutput176 net176 VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_12
Xoutput154 net154 VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_12
Xoutput165 net165 VGND VGND VPWR VPWR chany_bottom_out[23] sky130_fd_sc_hd__buf_12
Xoutput198 net198 VGND VGND VPWR VPWR chany_top_out_0[26] sky130_fd_sc_hd__buf_12
Xoutput187 net187 VGND VGND VPWR VPWR chany_top_out_0[16] sky130_fd_sc_hd__buf_12
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_120_ sb_0__1_.mux_right_track_34.out VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput12 chanx_right_in[18] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
Xinput45 chany_bottom_in[20] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_2
Xinput34 chany_bottom_in[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_4
Xinput23 chanx_right_in[28] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput78 chany_top_in_0[23] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__buf_2
Xinput67 chany_top_in_0[13] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_2
Xinput89 chany_top_in_0[6] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_2
Xinput56 chany_bottom_in[3] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_4
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_44.out sky130_fd_sc_hd__clkbuf_1
XFILLER_57_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_bottom_track_21.mux_l1_in_2_ right_width_0_height_0_subtile_1__pin_inpad_0_
+ net27 sb_0__1_.mem_bottom_track_21.mem_out\[0\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_4_0_prog_clk sb_0__1_.mem_right_track_34.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_34.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_5_0_prog_clk sb_0__1_.mem_top_track_28.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_75_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_top_track_52.mux_l2_in_0_ net30 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_top_track_52.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_12.out sky130_fd_sc_hd__clkbuf_1
XFILLER_54_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk sb_0__1_.mem_bottom_track_29.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_37.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_21_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_13_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_13_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk sb_0__1_.mem_top_track_4.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_39_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_6.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_8.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_81_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_4_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[2\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_6.mux_l1_in_0_ net76 net82 sb_0__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_87_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_196_ sb_0__1_.mux_top_track_2.out VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_21.mux_l2_in_0_ sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_15 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_37 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput122 net122 VGND VGND VPWR VPWR chanx_right_out[11] sky130_fd_sc_hd__buf_12
Xoutput133 net133 VGND VGND VPWR VPWR chanx_right_out[21] sky130_fd_sc_hd__buf_12
Xoutput144 net144 VGND VGND VPWR VPWR chanx_right_out[4] sky130_fd_sc_hd__buf_12
Xoutput177 net177 VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_12
Xoutput155 net155 VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_12
Xoutput166 net166 VGND VGND VPWR VPWR chany_bottom_out[24] sky130_fd_sc_hd__buf_12
Xoutput199 net199 VGND VGND VPWR VPWR chany_top_out_0[27] sky130_fd_sc_hd__buf_12
Xoutput188 net188 VGND VGND VPWR VPWR chany_top_out_0[17] sky130_fd_sc_hd__buf_12
XFILLER_28_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_12.mux_l3_in_0_ sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_right_track_12.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_54.mux_l1_in_0_ net53 net109 sb_0__1_.mem_right_track_54.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput13 chanx_right_in[19] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
Xinput46 chany_bottom_in[21] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_4
Xinput35 chany_bottom_in[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_4
Xinput24 chanx_right_in[29] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
Xinput79 chany_top_in_0[24] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_1
Xinput68 chany_top_in_0[14] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_2
X_179_ sb_0__1_.mux_top_track_36.out VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_2
Xinput57 chany_bottom_in[4] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_21.mux_l1_in_1_ net9 net21 sb_0__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_7_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk sb_0__1_.mem_right_track_32.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_34.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_10.mux_l1_in_3_ net260 net58 sb_0__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_right_track_50.mux_l1_in_1__253 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_50.mux_l1_in_1__253/HI
+ net253 sky130_fd_sc_hd__conb_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_12.mux_l2_in_1_ net233 net41 sb_0__1_.mem_right_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_37.out sky130_fd_sc_hd__clkbuf_1
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_5_0_prog_clk sb_0__1_.mem_top_track_28.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_28.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_75_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_right_track_40.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_40.out sky130_fd_sc_hd__clkbuf_1
XFILLER_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_4_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[2\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_34.out sky130_fd_sc_hd__clkbuf_1
XFILLER_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_10.mux_l3_in_0_ sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X
+ sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X sb_0__1_.mem_top_track_10.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_top_track_52.mux_l1_in_0_ net12 net24 sb_0__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_4_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_1_0_prog_clk cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
+ net98 VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_195_ sb_0__1_.mux_top_track_4.out VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_16 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_27 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput123 net123 VGND VGND VPWR VPWR chanx_right_out[12] sky130_fd_sc_hd__buf_12
Xoutput134 net134 VGND VGND VPWR VPWR chanx_right_out[22] sky130_fd_sc_hd__buf_12
Xoutput145 net145 VGND VGND VPWR VPWR chanx_right_out[5] sky130_fd_sc_hd__buf_12
Xoutput167 net167 VGND VGND VPWR VPWR chany_bottom_out[25] sky130_fd_sc_hd__buf_12
Xoutput156 net156 VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_12
Xsb_0__1_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_28.out sky130_fd_sc_hd__clkbuf_1
Xoutput189 net189 VGND VGND VPWR VPWR chany_top_out_0[18] sky130_fd_sc_hd__buf_12
Xoutput178 net178 VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_12
XFILLER_87_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_top_track_10.mux_l2_in_1_ sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput36 chany_bottom_in[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
Xinput14 chanx_right_in[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput25 chanx_right_in[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput69 chany_top_in_0[15] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_2
Xinput47 chany_bottom_in[22] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_4
Xinput58 chany_bottom_in[5] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_4
X_178_ net35 VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail net97 VGND
+ VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XFILLER_33_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_bottom_track_21.mux_l1_in_0_ net85 net71 sb_0__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_top_track_4.mux_l3_in_0_ sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_top_track_4.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_1.out sky130_fd_sc_hd__clkbuf_2
XFILLER_62_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_10.mux_l1_in_2_ net43 net25 sb_0__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_45.mux_l3_in_0_ sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_bottom_track_45.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_12.mux_l2_in_0_ net104 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_12.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_4_0_prog_clk sb_0__1_.mem_top_track_20.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_83_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_4_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_top_track_4.mux_l2_in_1_ net266 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_top_track_4.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_bottom_track_45.mux_l2_in_1_ net227 net30 sb_0__1_.mem_bottom_track_45.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_35_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_55_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_4.mux_l1_in_2_ net60 net47 sb_0__1_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_12_0_prog_clk sb_0__1_.mem_right_track_20.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_20.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_67_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_194_ sb_0__1_.mux_top_track_6.out VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_right_track_46.mux_l2_in_0__251 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_46.mux_l2_in_0__251/HI
+ net251 sky130_fd_sc_hd__conb_1
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_56.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_56.out sky130_fd_sc_hd__clkbuf_1
XFILLER_49_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_10_0_prog_clk sb_0__1_.mem_right_track_52.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_52.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_28 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_17 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput124 net124 VGND VGND VPWR VPWR chanx_right_out[13] sky130_fd_sc_hd__buf_12
Xoutput146 net146 VGND VGND VPWR VPWR chanx_right_out[6] sky130_fd_sc_hd__buf_12
Xoutput168 net168 VGND VGND VPWR VPWR chany_bottom_out[26] sky130_fd_sc_hd__buf_12
Xoutput157 net157 VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_12
Xoutput135 net135 VGND VGND VPWR VPWR chanx_right_out[23] sky130_fd_sc_hd__buf_12
XFILLER_87_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput179 net179 VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_12
XFILLER_87_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_top_track_10.mux_l2_in_0_ sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_55_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput37 chany_bottom_in[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_2
Xinput26 chanx_right_in[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput15 chanx_right_in[20] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput48 chany_bottom_in[23] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_4
Xinput59 chany_bottom_in[6] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_4
X_177_ net34 VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_top_track_10.mux_l1_in_1_ net7 net19 sb_0__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail net97 VGND
+ VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_9_0_prog_clk sb_0__1_.mem_bottom_track_29.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_29.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_88_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_top_track_4.mux_l2_in_0_ sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_45.mux_l2_in_0_ net12 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_bottom_track_45.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_12.mux_l1_in_0_ net71 net75 sb_0__1_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_47_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_24.mux_l2_in_0_ sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_24.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_81_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_0_0_prog_clk
+ net2 net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xsb_0__1_.mux_right_track_36.mux_l3_in_0_ sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_right_track_36.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_top_track_4.mux_l1_in_1_ net27 net9 sb_0__1_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk sb_0__1_.mem_right_track_20.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_20.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_63_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_12_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_12_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_50_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_193_ net51 VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_2
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_1.mux_l3_in_0_ sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_bottom_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk sb_0__1_.mem_right_track_50.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_52.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_18 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_29 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput125 net125 VGND VGND VPWR VPWR chanx_right_out[14] sky130_fd_sc_hd__buf_12
Xoutput147 net147 VGND VGND VPWR VPWR chanx_right_out[7] sky130_fd_sc_hd__buf_12
Xoutput158 net158 VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_12
Xoutput136 net136 VGND VGND VPWR VPWR chanx_right_out[24] sky130_fd_sc_hd__buf_12
Xsb_0__1_.mux_right_track_24.mux_l1_in_1_ net240 net62 sb_0__1_.mem_right_track_24.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_87_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput169 net169 VGND VGND VPWR VPWR chany_bottom_out[27] sky130_fd_sc_hd__buf_12
XFILLER_55_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_36.mux_l2_in_1_ net246 net33 sb_0__1_.mem_right_track_36.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_28.mux_l1_in_1__242 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_28.mux_l1_in_1__242/HI
+ net242 sky130_fd_sc_hd__conb_1
XFILLER_19_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput27 chanx_right_in[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
Xinput16 chanx_right_in[21] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput49 chany_bottom_in[24] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput38 chany_bottom_in[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_4
X_176_ net62 VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_bottom_track_1.mux_l2_in_1_ net275 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_bottom_track_1.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_159_ net77 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_top_track_10.mux_l1_in_0_ net118 net116 sb_0__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_11_0_prog_clk sb_0__1_.mem_bottom_track_29.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_29.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_94_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_0_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_2.ccff_tail net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.out sky130_fd_sc_hd__clkbuf_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_1.mux_l1_in_2_ right_width_0_height_0_subtile_3__pin_inpad_0_
+ right_width_0_height_0_subtile_0__pin_inpad_0_ sb_0__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_12.mux_l2_in_1__233 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_12.mux_l2_in_1__233/HI
+ net233 sky130_fd_sc_hd__conb_1
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_top_track_4.mux_l1_in_0_ net21 net117 sb_0__1_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_13_0_prog_clk sb_0__1_.mem_right_track_18.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_20.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_32.mux_l1_in_1__244 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_32.mux_l1_in_1__244/HI
+ net244 sky130_fd_sc_hd__conb_1
XFILLER_63_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_192_ sb_0__1_.mux_top_track_10.out VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_bottom_track_45.mux_l1_in_0_ net24 net67 sb_0__1_.mem_bottom_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_2.mux_l3_in_0_ sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_right_track_2.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_77_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_19 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput148 net148 VGND VGND VPWR VPWR chanx_right_out[8] sky130_fd_sc_hd__buf_12
Xoutput159 net159 VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_12
Xoutput126 net126 VGND VGND VPWR VPWR chanx_right_out[15] sky130_fd_sc_hd__buf_12
Xoutput137 net137 VGND VGND VPWR VPWR chanx_right_out[25] sky130_fd_sc_hd__buf_12
Xsb_0__1_.mux_right_track_24.mux_l1_in_0_ net110 net92 sb_0__1_.mem_right_track_24.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_36.mux_l2_in_0_ net44 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_36.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput28 chanx_right_in[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
Xinput17 chanx_right_in[22] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dlymetal6s2s_1
X_175_ sb_0__1_.mux_top_track_44.out VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput39 chany_bottom_in[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_4
XFILLER_6_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_11.mux_l1_in_3__276 VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.mux_l1_in_3__276/HI
+ net276 sky130_fd_sc_hd__conb_1
Xsb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk sb_0__1_.mem_right_track_26.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_26.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_56_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_2.mux_l2_in_1_ net237 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_right_track_2.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_bottom_track_1.mux_l2_in_0_ sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_86_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_158_ net76 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk sb_0__1_.mem_bottom_track_21.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_29.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_94_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_right_track_2.mux_l1_in_2_ net48 net111 sb_0__1_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_1.mux_l1_in_1_ net32 net15 sb_0__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_79_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_12.out sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mux_top_track_6.mux_l1_in_3__269 VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.mux_l1_in_3__269/HI
+ net269 sky130_fd_sc_hd__conb_1
XFILLER_91_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_3_0_prog_clk sb_0__1_.mem_bottom_track_3.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_90_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_191_ sb_0__1_.mux_top_track_12.out VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_2
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_89_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput149 net149 VGND VGND VPWR VPWR chanx_right_out[9] sky130_fd_sc_hd__buf_12
Xoutput127 net127 VGND VGND VPWR VPWR chanx_right_out[16] sky130_fd_sc_hd__buf_12
Xoutput138 net138 VGND VGND VPWR VPWR chanx_right_out[26] sky130_fd_sc_hd__buf_12
XFILLER_95_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput18 chanx_right_in[23] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput29 chanx_right_in[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlymetal6s2s_1
X_174_ net60 VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk sb_0__1_.mem_right_track_24.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_26.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_2.mux_l2_in_0_ sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_3_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_157_ sb_0__1_.mux_bottom_track_21.out VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_36.mux_l1_in_0_ net108 net74 sb_0__1_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_48.mux_l2_in_0_ net252 sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_48.ccff_tail VGND VGND VPWR VPWR sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_209_ net98 VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_50.mux_l2_in_0_ sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_50.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_right_track_2.mux_l1_in_1_ net108 net105 sb_0__1_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_93_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_9_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_9_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_bottom_track_1.mux_l1_in_0_ net64 net81 sb_0__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_80_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.out sky130_fd_sc_hd__clkbuf_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net93 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR right_width_0_height_0_subtile_3__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_50.mux_l1_in_1_ net253 net50 sb_0__1_.mem_right_track_50.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_72_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk sb_0__1_.mem_bottom_track_3.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_90_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_190_ net48 VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_5.mux_l2_in_1__228 VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_5.mux_l2_in_1__228/HI
+ net228 sky130_fd_sc_hd__conb_1
XFILLER_20_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput128 net128 VGND VGND VPWR VPWR chanx_right_out[17] sky130_fd_sc_hd__buf_12
Xoutput139 net139 VGND VGND VPWR VPWR chanx_right_out[27] sky130_fd_sc_hd__buf_12
XFILLER_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_173_ net59 VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_2
Xinput19 chanx_right_in[24] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_11_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_11_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_28.out sky130_fd_sc_hd__clkbuf_1
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_156_ net73 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_29.mux_l2_in_1__279 VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_29.mux_l2_in_1__279/HI
+ net279 sky130_fd_sc_hd__conb_1
XFILLER_56_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3_ net271 net89 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_208_ net98 VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_139_ net85 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_2
XFILLER_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_right_track_2.mux_l1_in_0_ net78 net84 sb_0__1_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_93_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_6.out sky130_fd_sc_hd__clkbuf_1
XFILLER_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_48.mux_l1_in_0_ net49 net106 sb_0__1_.mem_right_track_48.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_12.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4_ sb_0__1_.mux_bottom_track_37.out
+ net35 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_50.mux_l1_in_0_ net111 net107 sb_0__1_.mem_right_track_50.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_71_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_6_0_prog_clk sb_0__1_.mem_bottom_track_1.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_75_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk sb_0__1_.mem_right_track_44.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l4_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cby_0__1_.cby_0__1_.mem_right_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput129 net129 VGND VGND VPWR VPWR chanx_right_out[18] sky130_fd_sc_hd__buf_12
XFILLER_68_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net96 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_23_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_172_ net58 VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l3_in_1_ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_30.out sky130_fd_sc_hd__clkbuf_1
XFILLER_3_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_155_ net72 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2_ net58 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_207_ net98 VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_1
X_138_ net74 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_top_track_0.mux_l1_in_3_ net259 net34 sb_0__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_24.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_24.out sky130_fd_sc_hd__clkbuf_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_12.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_93_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3_ net72 net41 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_18.out sky130_fd_sc_hd__clkbuf_1
XFILLER_40_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk sb_0__1_.mem_right_track_40.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_0.mux_l3_in_0_ sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
+ sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X sb_0__1_.mem_top_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_49_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_44.mux_l2_in_0__250 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_44.mux_l2_in_0__250/HI
+ net250 sky130_fd_sc_hd__conb_1
XFILLER_77_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput119 net119 VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_12
XFILLER_95_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_right_track_18.mux_l3_in_0_ sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_right_track_18.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_171_ sb_0__1_.mux_top_track_52.out VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_13_0_prog_clk sb_0__1_.mem_right_track_18.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_18.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_10_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_20.mux_l3_in_0_ sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_right_track_20.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l3_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_top_track_0.mux_l2_in_1_ sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_154_ net71 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_18.mux_l2_in_1_ net236 net37 sb_0__1_.mem_right_track_18.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_20.mux_l2_in_1_ net238 net35 sb_0__1_.mem_right_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_3_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_52.out sky130_fd_sc_hd__clkbuf_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_1_ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_206_ net98 VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__clkbuf_1
X_137_ sb_0__1_.mux_right_track_0.out VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_top_track_0.mux_l1_in_2_ net51 net29 sb_0__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_10.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_93_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_13_0_prog_clk sb_0__1_.mem_top_track_2.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_46.out sky130_fd_sc_hd__clkbuf_1
XFILLER_30_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2_ sb_0__1_.mux_bottom_track_13.out
+ net48 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_8_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_8_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_4_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_4.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_67_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_26.mux_l1_in_1__241 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_26.mux_l1_in_1__241/HI
+ net241 sky130_fd_sc_hd__conb_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_170_ net56 VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk sb_0__1_.mem_right_track_18.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_18.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_10_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_8.mux_l2_in_1__258 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_8.mux_l2_in_1__258/HI
+ net258 sky130_fd_sc_hd__conb_1
XFILLER_5_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_0.mux_l2_in_0_ sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_51_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_153_ sb_0__1_.mux_bottom_track_29.out VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_18.mux_l2_in_0_ net107 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_18.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_10_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_10_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_0__1_.mux_right_track_20.mux_l2_in_0_ net108 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_20.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__274 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__274/HI
+ net274 sky130_fd_sc_hd__conb_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_205_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__clkbuf_1
X_136_ sb_0__1_.mux_right_track_2.out VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_2
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_top_track_0.mux_l1_in_1_ net11 net23 sb_0__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_38_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.out sky130_fd_sc_hd__clkbuf_2
XFILLER_69_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_10.mux_l2_in_1__232 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_10.mux_l2_in_1__232/HI
+ net232 sky130_fd_sc_hd__conb_1
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_119_ sb_0__1_.mux_right_track_36.out VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_2
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk sb_0__1_.mem_top_track_2.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_22_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_ sb_0__1_.mux_bottom_track_7.out
+ net51 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_4.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_4_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_30.mux_l1_in_1__243 VGND VGND VPWR VPWR sb_0__1_.mux_right_track_30.mux_l1_in_1__243/HI
+ net243 sky130_fd_sc_hd__conb_1
XFILLER_77_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_3.mux_l2_in_1__225 VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_3.mux_l2_in_1__225/HI
+ net225 sky130_fd_sc_hd__conb_1
XFILLER_31_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_2.out sky130_fd_sc_hd__clkbuf_1
XFILLER_95_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_28.mux_l3_in_0_ sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_top_track_28.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_59_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_16.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_18.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_152_ net69 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_top_track_28.mux_l2_in_1_ net264 net44 sb_0__1_.mem_top_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_bottom_track_53.mux_l1_in_1__229 VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_53.mux_l1_in_1__229/HI
+ net229 sky130_fd_sc_hd__conb_1
XFILLER_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk sb_0__1_.mem_right_track_30.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_30.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_68_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_204_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_1
XFILLER_23_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_135_ sb_0__1_.mux_right_track_4.out VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_1
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_top_track_0.mux_l1_in_0_ net118 net115 sb_0__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_bottom_track_7.mux_l1_in_3_ net230 right_width_0_height_0_subtile_2__pin_inpad_0_
+ sb_0__1_.mem_bottom_track_7.mem_out\[0\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_18.mux_l1_in_0_ net91 net67 sb_0__1_.mem_right_track_18.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_79_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_4_0_prog_clk cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail
+ net98 VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_118_ sb_0__1_.mux_right_track_38.out VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_2
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_bottom_track_53.mux_l2_in_0_ sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X net120 VGND VGND VPWR VPWR
+ sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_20.mux_l1_in_0_ net87 net65 sb_0__1_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_13_0_prog_clk sb_0__1_.mem_top_track_0.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_ sb_0__1_.mux_bottom_track_1.out
+ net54 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_32.mux_l2_in_0_ sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_32.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_55_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_0_0_prog_clk sb_0__1_.mem_right_track_36.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_36.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_40_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_2.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1 chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_7.mux_l3_in_0_ sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X
+ sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X sb_0__1_.mem_bottom_track_11.ccff_head
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_1_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_53.mux_l1_in_1_ net229 net31 sb_0__1_.mem_bottom_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_5_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_32.mux_l1_in_1_ net244 net56 sb_0__1_.mem_right_track_32.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_59_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_44.mux_l1_in_1__267 VGND VGND VPWR VPWR sb_0__1_.mux_top_track_44.mux_l1_in_1__267/HI
+ net267 sky130_fd_sc_hd__conb_1
XFILLER_93_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_7.mux_l2_in_1_ sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_151_ net68 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_2
XFILLER_50_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_28.mux_l2_in_0_ sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_6_0_prog_clk sb_0__1_.mem_right_track_28.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_30.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_203_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_2
X_134_ sb_0__1_.mux_right_track_6.out VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_2
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_7.mux_l1_in_2_ right_width_0_height_0_subtile_0__pin_inpad_0_
+ net14 sb_0__1_.mem_bottom_track_7.mem_out\[0\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_bottom_track_11.mux_l1_in_3_ net276 right_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_0__1_.mem_bottom_track_11.mem_out\[0\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_28.mux_l1_in_1_ net39 net4 sb_0__1_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_13.mux_l2_in_1__277 VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_13.mux_l2_in_1__277/HI
+ net277 sky130_fd_sc_hd__conb_1
XFILLER_34_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_117_ sb_0__1_.mux_right_track_40.out VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk sb_0__1_.mem_right_track_36.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_36.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_71_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_2 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_8.mux_l3_in_0_ sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_right_track_10.ccff_head
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_11.mux_l3_in_0_ sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X
+ sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X sb_0__1_.mem_bottom_track_11.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_40_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_53.mux_l1_in_0_ net13 net65 sb_0__1_.mem_bottom_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_bottom_track_1.mux_l2_in_1__275 VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_1.mux_l2_in_1__275/HI
+ net275 sky130_fd_sc_hd__conb_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_32.mux_l1_in_0_ net106 net86 sb_0__1_.mem_right_track_32.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_7_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_7_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_44.mux_l2_in_0_ net250 sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_44.ccff_tail VGND VGND VPWR VPWR sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_8.mux_l2_in_1_ net258 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_right_track_8.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_bottom_track_7.mux_l2_in_0_ sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_0_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[2\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_bottom_track_11.mux_l2_in_1_ sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_150_ net67 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_2
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_202_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_2
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_133_ sb_0__1_.mux_right_track_8.out VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_right_track_8.mux_l1_in_2_ net43 net111 sb_0__1_.mem_right_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_7.mux_l1_in_1_ net6 net18 sb_0__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_7.mux_l1_in_3__230 VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.mux_l1_in_3__230/HI
+ net230 sky130_fd_sc_hd__conb_1
XFILLER_65_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_bottom_track_11.mux_l1_in_2_ right_width_0_height_0_subtile_1__pin_inpad_0_
+ net25 sb_0__1_.mem_bottom_track_11.mem_out\[0\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_28.mux_l1_in_0_ net16 net117 sb_0__1_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_69_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_116_ net36 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_2
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk sb_0__1_.mem_right_track_34.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_36.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_3 chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_2.out sky130_fd_sc_hd__clkbuf_1
XFILLER_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_8.mux_l2_in_0_ sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_8.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_64_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_11.mux_l2_in_0_ sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xcby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_0_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_77_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_44.mux_l1_in_0_ net40 net104 sb_0__1_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_32_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_56.mux_l2_in_0_ net256 sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_bottom_track_1.ccff_head VGND VGND VPWR VPWR sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
X_201_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_2
X_132_ sb_0__1_.mux_right_track_10.out VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_8.mux_l1_in_1_ net108 net105 sb_0__1_.mem_right_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_2_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_7.mux_l1_in_0_ net89 net76 sb_0__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_78_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_bottom_track_11.mux_l1_in_1_ net7 net19 sb_0__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_29_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_115_ sb_0__1_.mux_right_track_44.out VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_2
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_52.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_52.out sky130_fd_sc_hd__clkbuf_1
XFILLER_78_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3_ net272 net88 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_4 right_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_5_0_prog_clk sb_0__1_.mem_top_track_10.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_95_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_20.out sky130_fd_sc_hd__clkbuf_1
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
.ends

