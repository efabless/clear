magic
tech sky130A
magscale 1 2
timestamp 1625784757
<< locali >>
rect 20913 19159 20947 19261
rect 19717 18615 19751 18785
rect 14749 17527 14783 17629
rect 17233 17595 17267 17833
rect 14289 17119 14323 17289
rect 6653 16643 6687 16745
rect 22017 15215 22051 15929
rect 19717 14263 19751 14433
rect 8309 12699 8343 12801
rect 22017 12495 22051 13345
rect 3249 12087 3283 12325
rect 17969 12155 18003 12393
rect 19257 11611 19291 11849
rect 6469 10999 6503 11305
rect 22017 11067 22051 12257
rect 13461 9367 13495 9605
rect 14197 9027 14231 9129
rect 14105 8823 14139 8925
rect 12633 7735 12667 7905
rect 9965 7191 9999 7429
rect 10333 7259 10367 7361
rect 14197 7327 14231 7497
rect 16313 7191 16347 7361
rect 22017 6919 22051 7905
rect 4721 6103 4755 6205
rect 11529 6171 11563 6409
rect 7481 5015 7515 5321
rect 16681 5151 16715 5253
rect 10517 5015 10551 5117
rect 5733 3927 5767 4029
rect 4445 3383 4479 3553
rect 10977 3519 11011 3689
rect 12541 3383 12575 3621
rect 9597 2839 9631 3009
rect 12173 2975 12207 3145
rect 5641 2431 5675 2601
<< viali >>
rect 2237 20553 2271 20587
rect 2697 20485 2731 20519
rect 3249 20485 3283 20519
rect 4077 20485 4111 20519
rect 17417 20485 17451 20519
rect 18429 20485 18463 20519
rect 18981 20485 19015 20519
rect 19533 20485 19567 20519
rect 1593 20349 1627 20383
rect 1777 20349 1811 20383
rect 4813 20349 4847 20383
rect 5089 20349 5123 20383
rect 5733 20349 5767 20383
rect 6561 20349 6595 20383
rect 18245 20349 18279 20383
rect 20269 20349 20303 20383
rect 2329 20281 2363 20315
rect 2881 20281 2915 20315
rect 3433 20281 3467 20315
rect 4261 20281 4295 20315
rect 17601 20281 17635 20315
rect 18797 20281 18831 20315
rect 19349 20281 19383 20315
rect 20637 20281 20671 20315
rect 20821 20281 20855 20315
rect 21189 20281 21223 20315
rect 21373 20281 21407 20315
rect 4629 20213 4663 20247
rect 5917 20213 5951 20247
rect 8125 20213 8159 20247
rect 20085 20213 20119 20247
rect 2329 20009 2363 20043
rect 2973 20009 3007 20043
rect 3433 20009 3467 20043
rect 8125 20009 8159 20043
rect 20085 20009 20119 20043
rect 20729 20009 20763 20043
rect 10578 19941 10612 19975
rect 19809 19941 19843 19975
rect 1777 19873 1811 19907
rect 2513 19873 2547 19907
rect 2789 19873 2823 19907
rect 3249 19873 3283 19907
rect 4077 19873 4111 19907
rect 4344 19873 4378 19907
rect 19257 19873 19291 19907
rect 20269 19873 20303 19907
rect 20637 19873 20671 19907
rect 21189 19873 21223 19907
rect 8217 19805 8251 19839
rect 8309 19805 8343 19839
rect 10333 19805 10367 19839
rect 1593 19737 1627 19771
rect 5733 19737 5767 19771
rect 21373 19737 21407 19771
rect 5457 19669 5491 19703
rect 7757 19669 7791 19703
rect 11713 19669 11747 19703
rect 2145 19465 2179 19499
rect 2605 19465 2639 19499
rect 9689 19465 9723 19499
rect 20177 19465 20211 19499
rect 20637 19465 20671 19499
rect 19441 19397 19475 19431
rect 7941 19329 7975 19363
rect 1593 19261 1627 19295
rect 2329 19261 2363 19295
rect 2789 19261 2823 19295
rect 4445 19261 4479 19295
rect 5089 19261 5123 19295
rect 7665 19261 7699 19295
rect 8309 19261 8343 19295
rect 13277 19261 13311 19295
rect 19257 19261 19291 19295
rect 19901 19261 19935 19295
rect 20361 19261 20395 19295
rect 20821 19261 20855 19295
rect 20913 19261 20947 19295
rect 1777 19193 1811 19227
rect 4200 19193 4234 19227
rect 4721 19193 4755 19227
rect 8554 19193 8588 19227
rect 13522 19193 13556 19227
rect 18613 19193 18647 19227
rect 21189 19193 21223 19227
rect 21373 19193 21407 19227
rect 3065 19125 3099 19159
rect 7297 19125 7331 19159
rect 7757 19125 7791 19159
rect 14657 19125 14691 19159
rect 18153 19125 18187 19159
rect 18981 19125 19015 19159
rect 19717 19125 19751 19159
rect 20913 19125 20947 19159
rect 2145 18921 2179 18955
rect 2605 18921 2639 18955
rect 3065 18921 3099 18955
rect 4721 18921 4755 18955
rect 19257 18921 19291 18955
rect 20361 18921 20395 18955
rect 20821 18921 20855 18955
rect 12234 18853 12268 18887
rect 1593 18785 1627 18819
rect 1777 18785 1811 18819
rect 2329 18785 2363 18819
rect 2789 18785 2823 18819
rect 3249 18785 3283 18819
rect 4353 18785 4387 18819
rect 5264 18785 5298 18819
rect 7564 18785 7598 18819
rect 11989 18785 12023 18819
rect 14913 18785 14947 18819
rect 19073 18785 19107 18819
rect 19717 18785 19751 18819
rect 20177 18785 20211 18819
rect 20637 18785 20671 18819
rect 21189 18785 21223 18819
rect 4997 18717 5031 18751
rect 7297 18717 7331 18751
rect 14657 18717 14691 18751
rect 21373 18649 21407 18683
rect 3985 18581 4019 18615
rect 6377 18581 6411 18615
rect 8677 18581 8711 18615
rect 13369 18581 13403 18615
rect 16037 18581 16071 18615
rect 18705 18581 18739 18615
rect 19717 18581 19751 18615
rect 19809 18581 19843 18615
rect 2237 18377 2271 18411
rect 7481 18377 7515 18411
rect 17141 18377 17175 18411
rect 20361 18377 20395 18411
rect 20821 18377 20855 18411
rect 2697 18309 2731 18343
rect 12633 18309 12667 18343
rect 3341 18241 3375 18275
rect 4813 18241 4847 18275
rect 8125 18241 8159 18275
rect 9045 18241 9079 18275
rect 12081 18241 12115 18275
rect 14565 18241 14599 18275
rect 17693 18241 17727 18275
rect 19349 18241 19383 18275
rect 2881 18173 2915 18207
rect 19717 18173 19751 18207
rect 20177 18173 20211 18207
rect 20637 18173 20671 18207
rect 1777 18105 1811 18139
rect 2329 18105 2363 18139
rect 3433 18105 3467 18139
rect 4537 18105 4571 18139
rect 7849 18105 7883 18139
rect 12265 18105 12299 18139
rect 17509 18105 17543 18139
rect 18153 18105 18187 18139
rect 21189 18105 21223 18139
rect 21373 18105 21407 18139
rect 1685 18037 1719 18071
rect 3525 18037 3559 18071
rect 3893 18037 3927 18071
rect 4169 18037 4203 18071
rect 4629 18037 4663 18071
rect 5181 18037 5215 18071
rect 7941 18037 7975 18071
rect 8493 18037 8527 18071
rect 8861 18037 8895 18071
rect 8953 18037 8987 18071
rect 9505 18037 9539 18071
rect 12173 18037 12207 18071
rect 14657 18037 14691 18071
rect 14749 18037 14783 18071
rect 15117 18037 15151 18071
rect 15393 18037 15427 18071
rect 17601 18037 17635 18071
rect 18981 18037 19015 18071
rect 19901 18037 19935 18071
rect 2145 17833 2179 17867
rect 3525 17833 3559 17867
rect 4353 17833 4387 17867
rect 7849 17833 7883 17867
rect 12909 17833 12943 17867
rect 13553 17833 13587 17867
rect 14841 17833 14875 17867
rect 15209 17833 15243 17867
rect 16589 17833 16623 17867
rect 17233 17833 17267 17867
rect 17417 17833 17451 17867
rect 19257 17833 19291 17867
rect 20269 17833 20303 17867
rect 3065 17765 3099 17799
rect 5908 17765 5942 17799
rect 1777 17697 1811 17731
rect 2329 17697 2363 17731
rect 3157 17697 3191 17731
rect 4721 17697 4755 17731
rect 8033 17697 8067 17731
rect 9577 17697 9611 17731
rect 11244 17697 11278 17731
rect 16221 17697 16255 17731
rect 2973 17629 3007 17663
rect 4813 17629 4847 17663
rect 4905 17629 4939 17663
rect 5641 17629 5675 17663
rect 9321 17629 9355 17663
rect 10977 17629 11011 17663
rect 13369 17629 13403 17663
rect 13461 17629 13495 17663
rect 14749 17629 14783 17663
rect 15301 17629 15335 17663
rect 15485 17629 15519 17663
rect 15945 17629 15979 17663
rect 16129 17629 16163 17663
rect 18530 17697 18564 17731
rect 19073 17697 19107 17731
rect 20085 17697 20119 17731
rect 20637 17697 20671 17731
rect 21189 17697 21223 17731
rect 18797 17629 18831 17663
rect 17233 17561 17267 17595
rect 20821 17561 20855 17595
rect 21373 17561 21407 17595
rect 1685 17493 1719 17527
rect 3985 17493 4019 17527
rect 7021 17493 7055 17527
rect 8401 17493 8435 17527
rect 10701 17493 10735 17527
rect 12357 17493 12391 17527
rect 13921 17493 13955 17527
rect 14473 17493 14507 17527
rect 14749 17493 14783 17527
rect 19717 17493 19751 17527
rect 2605 17289 2639 17323
rect 3801 17289 3835 17323
rect 4997 17289 5031 17323
rect 6929 17289 6963 17323
rect 9137 17289 9171 17323
rect 11345 17289 11379 17323
rect 13461 17289 13495 17323
rect 14289 17289 14323 17323
rect 14933 17289 14967 17323
rect 17877 17289 17911 17323
rect 18153 17289 18187 17323
rect 20361 17289 20395 17323
rect 20821 17289 20855 17323
rect 12633 17221 12667 17255
rect 3249 17153 3283 17187
rect 4077 17153 4111 17187
rect 5641 17153 5675 17187
rect 7481 17153 7515 17187
rect 9689 17153 9723 17187
rect 10701 17153 10735 17187
rect 10885 17153 10919 17187
rect 12081 17153 12115 17187
rect 12173 17153 12207 17187
rect 14105 17153 14139 17187
rect 15945 17153 15979 17187
rect 17325 17153 17359 17187
rect 1593 17085 1627 17119
rect 2329 17085 2363 17119
rect 2789 17085 2823 17119
rect 3341 17085 3375 17119
rect 13921 17085 13955 17119
rect 14289 17085 14323 17119
rect 19533 17085 19567 17119
rect 20177 17085 20211 17119
rect 20637 17085 20671 17119
rect 1777 17017 1811 17051
rect 3433 17017 3467 17051
rect 5365 17017 5399 17051
rect 7297 17017 7331 17051
rect 9505 17017 9539 17051
rect 12265 17017 12299 17051
rect 12909 17017 12943 17051
rect 13829 17017 13863 17051
rect 14473 17017 14507 17051
rect 15761 17017 15795 17051
rect 17509 17017 17543 17051
rect 19266 17017 19300 17051
rect 21189 17017 21223 17051
rect 2145 16949 2179 16983
rect 4537 16949 4571 16983
rect 5457 16949 5491 16983
rect 7389 16949 7423 16983
rect 9597 16949 9631 16983
rect 10241 16949 10275 16983
rect 10977 16949 11011 16983
rect 15393 16949 15427 16983
rect 15853 16949 15887 16983
rect 16589 16949 16623 16983
rect 17417 16949 17451 16983
rect 19809 16949 19843 16983
rect 21281 16949 21315 16983
rect 2145 16745 2179 16779
rect 3065 16745 3099 16779
rect 5457 16745 5491 16779
rect 5825 16745 5859 16779
rect 6561 16745 6595 16779
rect 6653 16745 6687 16779
rect 6929 16745 6963 16779
rect 8585 16745 8619 16779
rect 11989 16745 12023 16779
rect 14013 16745 14047 16779
rect 14841 16745 14875 16779
rect 16221 16745 16255 16779
rect 16589 16745 16623 16779
rect 17233 16745 17267 16779
rect 19257 16745 19291 16779
rect 20361 16745 20395 16779
rect 20821 16745 20855 16779
rect 1777 16677 1811 16711
rect 4721 16677 4755 16711
rect 8125 16677 8159 16711
rect 11253 16677 11287 16711
rect 11345 16677 11379 16711
rect 12357 16677 12391 16711
rect 14933 16677 14967 16711
rect 1593 16609 1627 16643
rect 2329 16609 2363 16643
rect 2789 16609 2823 16643
rect 3249 16609 3283 16643
rect 4353 16609 4387 16643
rect 6653 16609 6687 16643
rect 8217 16609 8251 16643
rect 10701 16609 10735 16643
rect 13553 16609 13587 16643
rect 13645 16609 13679 16643
rect 16681 16609 16715 16643
rect 17601 16609 17635 16643
rect 19073 16609 19107 16643
rect 20177 16609 20211 16643
rect 20637 16609 20671 16643
rect 21189 16609 21223 16643
rect 21373 16609 21407 16643
rect 5917 16541 5951 16575
rect 6009 16541 6043 16575
rect 8033 16541 8067 16575
rect 11161 16541 11195 16575
rect 12449 16541 12483 16575
rect 12541 16541 12575 16575
rect 13369 16541 13403 16575
rect 14657 16541 14691 16575
rect 16773 16541 16807 16575
rect 17693 16541 17727 16575
rect 17785 16541 17819 16575
rect 2605 16473 2639 16507
rect 11713 16473 11747 16507
rect 15301 16473 15335 16507
rect 3893 16405 3927 16439
rect 19809 16405 19843 16439
rect 3065 16201 3099 16235
rect 3525 16201 3559 16235
rect 5733 16201 5767 16235
rect 7941 16201 7975 16235
rect 8585 16201 8619 16235
rect 19901 16201 19935 16235
rect 3985 16133 4019 16167
rect 19441 16133 19475 16167
rect 1593 16065 1627 16099
rect 7389 16065 7423 16099
rect 2329 15997 2363 16031
rect 2789 15997 2823 16031
rect 3249 15997 3283 16031
rect 3709 15997 3743 16031
rect 4353 15997 4387 16031
rect 6837 15997 6871 16031
rect 7481 15997 7515 16031
rect 9965 15997 9999 16031
rect 19257 15997 19291 16031
rect 19717 15997 19751 16031
rect 20177 15997 20211 16031
rect 20637 15997 20671 16031
rect 1777 15929 1811 15963
rect 4598 15929 4632 15963
rect 6561 15929 6595 15963
rect 7573 15929 7607 15963
rect 9720 15929 9754 15963
rect 21189 15929 21223 15963
rect 21373 15929 21407 15963
rect 22017 15929 22051 15963
rect 2145 15861 2179 15895
rect 2605 15861 2639 15895
rect 11713 15861 11747 15895
rect 13093 15861 13127 15895
rect 17049 15861 17083 15895
rect 17417 15861 17451 15895
rect 18613 15861 18647 15895
rect 18889 15861 18923 15895
rect 20361 15861 20395 15895
rect 20821 15861 20855 15895
rect 4077 15657 4111 15691
rect 15301 15657 15335 15691
rect 20269 15657 20303 15691
rect 1777 15589 1811 15623
rect 2145 15589 2179 15623
rect 2329 15589 2363 15623
rect 12366 15589 12400 15623
rect 15844 15589 15878 15623
rect 20637 15589 20671 15623
rect 21189 15589 21223 15623
rect 3065 15521 3099 15555
rect 5190 15521 5224 15555
rect 7674 15521 7708 15555
rect 9321 15521 9355 15555
rect 12633 15521 12667 15555
rect 14933 15521 14967 15555
rect 17960 15521 17994 15555
rect 20085 15521 20119 15555
rect 20821 15521 20855 15555
rect 2881 15453 2915 15487
rect 2973 15453 3007 15487
rect 5457 15453 5491 15487
rect 7941 15453 7975 15487
rect 14657 15453 14691 15487
rect 14841 15453 14875 15487
rect 15577 15453 15611 15487
rect 17693 15453 17727 15487
rect 1685 15317 1719 15351
rect 3433 15317 3467 15351
rect 6561 15317 6595 15351
rect 9505 15317 9539 15351
rect 11253 15317 11287 15351
rect 16957 15317 16991 15351
rect 19073 15317 19107 15351
rect 19625 15317 19659 15351
rect 21281 15317 21315 15351
rect 22017 15181 22051 15215
rect 4169 15113 4203 15147
rect 9965 15113 9999 15147
rect 14749 15113 14783 15147
rect 9689 15045 9723 15079
rect 18521 15045 18555 15079
rect 3801 14977 3835 15011
rect 13093 14977 13127 15011
rect 15301 14977 15335 15011
rect 17969 14977 18003 15011
rect 19349 14977 19383 15011
rect 20361 14977 20395 15011
rect 8033 14909 8067 14943
rect 8309 14909 8343 14943
rect 11345 14909 11379 14943
rect 13360 14909 13394 14943
rect 20177 14909 20211 14943
rect 1777 14841 1811 14875
rect 3556 14841 3590 14875
rect 7766 14841 7800 14875
rect 8554 14841 8588 14875
rect 11078 14841 11112 14875
rect 15117 14841 15151 14875
rect 18153 14841 18187 14875
rect 21189 14841 21223 14875
rect 21373 14841 21407 14875
rect 1685 14773 1719 14807
rect 2421 14773 2455 14807
rect 6653 14773 6687 14807
rect 14473 14773 14507 14807
rect 15209 14773 15243 14807
rect 15761 14773 15795 14807
rect 18061 14773 18095 14807
rect 18797 14773 18831 14807
rect 19165 14773 19199 14807
rect 19257 14773 19291 14807
rect 19809 14773 19843 14807
rect 20269 14773 20303 14807
rect 3157 14569 3191 14603
rect 3525 14569 3559 14603
rect 4077 14569 4111 14603
rect 5733 14569 5767 14603
rect 6193 14569 6227 14603
rect 6745 14569 6779 14603
rect 7757 14569 7791 14603
rect 8309 14569 8343 14603
rect 10701 14569 10735 14603
rect 13185 14569 13219 14603
rect 13645 14569 13679 14603
rect 15301 14569 15335 14603
rect 18613 14569 18647 14603
rect 19257 14569 19291 14603
rect 19809 14569 19843 14603
rect 14933 14501 14967 14535
rect 15844 14501 15878 14535
rect 1777 14433 1811 14467
rect 2789 14433 2823 14467
rect 4445 14433 4479 14467
rect 6101 14433 6135 14467
rect 7113 14433 7147 14467
rect 7941 14433 7975 14467
rect 9588 14433 9622 14467
rect 11805 14433 11839 14467
rect 12061 14433 12095 14467
rect 13829 14433 13863 14467
rect 14841 14433 14875 14467
rect 17489 14433 17523 14467
rect 19717 14433 19751 14467
rect 20177 14433 20211 14467
rect 21189 14433 21223 14467
rect 2513 14365 2547 14399
rect 2697 14365 2731 14399
rect 4537 14365 4571 14399
rect 4629 14365 4663 14399
rect 6377 14365 6411 14399
rect 7205 14365 7239 14399
rect 7297 14365 7331 14399
rect 9321 14365 9355 14399
rect 14657 14365 14691 14399
rect 15577 14365 15611 14399
rect 17233 14365 17267 14399
rect 20269 14365 20303 14399
rect 20361 14365 20395 14399
rect 21373 14297 21407 14331
rect 1685 14229 1719 14263
rect 16957 14229 16991 14263
rect 19717 14229 19751 14263
rect 2973 14025 3007 14059
rect 4169 14025 4203 14059
rect 7113 14025 7147 14059
rect 8309 14025 8343 14059
rect 10701 14025 10735 14059
rect 14381 14025 14415 14059
rect 18613 14025 18647 14059
rect 20361 14025 20395 14059
rect 20821 14025 20855 14059
rect 3709 13957 3743 13991
rect 9321 13957 9355 13991
rect 12633 13957 12667 13991
rect 18889 13957 18923 13991
rect 2421 13889 2455 13923
rect 4721 13889 4755 13923
rect 5733 13889 5767 13923
rect 7665 13889 7699 13923
rect 8769 13889 8803 13923
rect 8953 13889 8987 13923
rect 9873 13889 9907 13923
rect 11989 13889 12023 13923
rect 13737 13889 13771 13923
rect 14749 13889 14783 13923
rect 17969 13889 18003 13923
rect 18153 13889 18187 13923
rect 19441 13889 19475 13923
rect 1593 13821 1627 13855
rect 3893 13821 3927 13855
rect 5641 13821 5675 13855
rect 11345 13821 11379 13855
rect 12265 13821 12299 13855
rect 16221 13821 16255 13855
rect 17509 13821 17543 13855
rect 20177 13821 20211 13855
rect 20637 13821 20671 13855
rect 21189 13821 21223 13855
rect 21373 13821 21407 13855
rect 1777 13753 1811 13787
rect 4537 13753 4571 13787
rect 7573 13753 7607 13787
rect 14013 13753 14047 13787
rect 19257 13753 19291 13787
rect 2513 13685 2547 13719
rect 2605 13685 2639 13719
rect 3249 13685 3283 13719
rect 4629 13685 4663 13719
rect 5181 13685 5215 13719
rect 5549 13685 5583 13719
rect 7481 13685 7515 13719
rect 8677 13685 8711 13719
rect 9689 13685 9723 13719
rect 9781 13685 9815 13719
rect 12173 13685 12207 13719
rect 13921 13685 13955 13719
rect 16405 13685 16439 13719
rect 18245 13685 18279 13719
rect 19349 13685 19383 13719
rect 2421 13481 2455 13515
rect 2881 13481 2915 13515
rect 4077 13481 4111 13515
rect 4813 13481 4847 13515
rect 5273 13481 5307 13515
rect 5825 13481 5859 13515
rect 6193 13481 6227 13515
rect 6837 13481 6871 13515
rect 7941 13481 7975 13515
rect 8769 13481 8803 13515
rect 9689 13481 9723 13515
rect 11713 13481 11747 13515
rect 14841 13481 14875 13515
rect 16589 13481 16623 13515
rect 19257 13481 19291 13515
rect 19809 13481 19843 13515
rect 20269 13481 20303 13515
rect 2789 13413 2823 13447
rect 5181 13413 5215 13447
rect 11253 13413 11287 13447
rect 1777 13345 1811 13379
rect 4261 13345 4295 13379
rect 6285 13345 6319 13379
rect 7205 13345 7239 13379
rect 8585 13345 8619 13379
rect 10057 13345 10091 13379
rect 10149 13345 10183 13379
rect 11345 13345 11379 13379
rect 12449 13345 12483 13379
rect 15209 13345 15243 13379
rect 16221 13345 16255 13379
rect 17509 13345 17543 13379
rect 18613 13345 18647 13379
rect 19073 13345 19107 13379
rect 20177 13345 20211 13379
rect 21281 13345 21315 13379
rect 22017 13345 22051 13379
rect 3065 13277 3099 13311
rect 5365 13277 5399 13311
rect 6469 13277 6503 13311
rect 7297 13277 7331 13311
rect 7481 13277 7515 13311
rect 10333 13277 10367 13311
rect 11161 13277 11195 13311
rect 12265 13277 12299 13311
rect 12357 13277 12391 13311
rect 15301 13277 15335 13311
rect 15393 13277 15427 13311
rect 16037 13277 16071 13311
rect 16129 13277 16163 13311
rect 17233 13277 17267 13311
rect 20453 13277 20487 13311
rect 1593 13209 1627 13243
rect 17969 13209 18003 13243
rect 18797 13209 18831 13243
rect 21097 13209 21131 13243
rect 3433 13141 3467 13175
rect 12817 13141 12851 13175
rect 18337 13141 18371 13175
rect 2145 12937 2179 12971
rect 2605 12937 2639 12971
rect 4353 12937 4387 12971
rect 6009 12937 6043 12971
rect 7389 12937 7423 12971
rect 9045 12937 9079 12971
rect 10609 12937 10643 12971
rect 14749 12937 14783 12971
rect 15393 12937 15427 12971
rect 16405 12937 16439 12971
rect 18337 12937 18371 12971
rect 1593 12869 1627 12903
rect 18061 12869 18095 12903
rect 21097 12869 21131 12903
rect 3709 12801 3743 12835
rect 5181 12801 5215 12835
rect 7941 12801 7975 12835
rect 8309 12801 8343 12835
rect 8493 12801 8527 12835
rect 9689 12801 9723 12835
rect 15853 12801 15887 12835
rect 17601 12801 17635 12835
rect 18889 12801 18923 12835
rect 19901 12801 19935 12835
rect 1409 12733 1443 12767
rect 2329 12733 2363 12767
rect 2789 12733 2823 12767
rect 5641 12733 5675 12767
rect 7849 12733 7883 12767
rect 12817 12733 12851 12767
rect 14565 12733 14599 12767
rect 17233 12733 17267 12767
rect 17877 12733 17911 12767
rect 20637 12733 20671 12767
rect 3893 12665 3927 12699
rect 5089 12665 5123 12699
rect 7757 12665 7791 12699
rect 8309 12665 8343 12699
rect 13062 12665 13096 12699
rect 16037 12665 16071 12699
rect 18705 12665 18739 12699
rect 19809 12665 19843 12699
rect 21281 12665 21315 12699
rect 3065 12597 3099 12631
rect 3985 12597 4019 12631
rect 4629 12597 4663 12631
rect 4997 12597 5031 12631
rect 9413 12597 9447 12631
rect 9505 12597 9539 12631
rect 14197 12597 14231 12631
rect 15945 12597 15979 12631
rect 18797 12597 18831 12631
rect 19349 12597 19383 12631
rect 19717 12597 19751 12631
rect 20729 12597 20763 12631
rect 22017 12461 22051 12495
rect 2697 12393 2731 12427
rect 2789 12393 2823 12427
rect 5733 12393 5767 12427
rect 7205 12393 7239 12427
rect 9413 12393 9447 12427
rect 9873 12393 9907 12427
rect 12449 12393 12483 12427
rect 15945 12393 15979 12427
rect 17969 12393 18003 12427
rect 18429 12393 18463 12427
rect 19809 12393 19843 12427
rect 20177 12393 20211 12427
rect 1685 12325 1719 12359
rect 3249 12325 3283 12359
rect 14810 12325 14844 12359
rect 17610 12325 17644 12359
rect 2605 12189 2639 12223
rect 3157 12121 3191 12155
rect 4353 12257 4387 12291
rect 5089 12257 5123 12291
rect 5181 12257 5215 12291
rect 7573 12257 7607 12291
rect 7665 12257 7699 12291
rect 9781 12257 9815 12291
rect 11069 12257 11103 12291
rect 11336 12257 11370 12291
rect 13553 12257 13587 12291
rect 5273 12189 5307 12223
rect 7757 12189 7791 12223
rect 9965 12189 9999 12223
rect 12909 12189 12943 12223
rect 13277 12189 13311 12223
rect 13461 12189 13495 12223
rect 14565 12189 14599 12223
rect 17877 12189 17911 12223
rect 19257 12325 19291 12359
rect 18521 12257 18555 12291
rect 20269 12257 20303 12291
rect 21281 12257 21315 12291
rect 22017 12257 22051 12291
rect 18245 12189 18279 12223
rect 20361 12189 20395 12223
rect 4721 12121 4755 12155
rect 17969 12121 18003 12155
rect 1777 12053 1811 12087
rect 3249 12053 3283 12087
rect 3433 12053 3467 12087
rect 3985 12053 4019 12087
rect 13921 12053 13955 12087
rect 16497 12053 16531 12087
rect 18889 12053 18923 12087
rect 21189 12053 21223 12087
rect 3709 11849 3743 11883
rect 3985 11849 4019 11883
rect 9229 11849 9263 11883
rect 9505 11849 9539 11883
rect 11253 11849 11287 11883
rect 12633 11849 12667 11883
rect 12909 11849 12943 11883
rect 16129 11849 16163 11883
rect 18429 11849 18463 11883
rect 19257 11849 19291 11883
rect 19441 11849 19475 11883
rect 1869 11781 1903 11815
rect 7757 11781 7791 11815
rect 14657 11781 14691 11815
rect 15853 11781 15887 11815
rect 4537 11713 4571 11747
rect 5089 11713 5123 11747
rect 8677 11713 8711 11747
rect 10057 11713 10091 11747
rect 10701 11713 10735 11747
rect 11989 11713 12023 11747
rect 13553 11713 13587 11747
rect 14013 11713 14047 11747
rect 14197 11713 14231 11747
rect 15301 11713 15335 11747
rect 17049 11713 17083 11747
rect 17601 11713 17635 11747
rect 18981 11713 19015 11747
rect 1685 11645 1719 11679
rect 2329 11645 2363 11679
rect 8769 11645 8803 11679
rect 10885 11645 10919 11679
rect 13277 11645 13311 11679
rect 14289 11645 14323 11679
rect 17785 11645 17819 11679
rect 20085 11713 20119 11747
rect 21005 11713 21039 11747
rect 21097 11713 21131 11747
rect 19901 11645 19935 11679
rect 20913 11645 20947 11679
rect 2596 11577 2630 11611
rect 18797 11577 18831 11611
rect 19257 11577 19291 11611
rect 4353 11509 4387 11543
rect 4445 11509 4479 11543
rect 5457 11509 5491 11543
rect 7297 11509 7331 11543
rect 8861 11509 8895 11543
rect 9873 11509 9907 11543
rect 9965 11509 9999 11543
rect 10793 11509 10827 11543
rect 12173 11509 12207 11543
rect 12265 11509 12299 11543
rect 13369 11509 13403 11543
rect 15393 11509 15427 11543
rect 15485 11509 15519 11543
rect 16589 11509 16623 11543
rect 17693 11509 17727 11543
rect 18153 11509 18187 11543
rect 18889 11509 18923 11543
rect 19809 11509 19843 11543
rect 20545 11509 20579 11543
rect 3157 11305 3191 11339
rect 4445 11305 4479 11339
rect 6285 11305 6319 11339
rect 6469 11305 6503 11339
rect 9413 11305 9447 11339
rect 13921 11305 13955 11339
rect 16957 11305 16991 11339
rect 1685 11237 1719 11271
rect 3433 11237 3467 11271
rect 2789 11169 2823 11203
rect 5569 11169 5603 11203
rect 5825 11169 5859 11203
rect 2605 11101 2639 11135
rect 2697 11101 2731 11135
rect 1869 11033 1903 11067
rect 7021 11237 7055 11271
rect 8033 11237 8067 11271
rect 20260 11237 20294 11271
rect 6929 11169 6963 11203
rect 8125 11169 8159 11203
rect 10057 11169 10091 11203
rect 11713 11169 11747 11203
rect 13461 11169 13495 11203
rect 13737 11169 13771 11203
rect 17969 11169 18003 11203
rect 18797 11169 18831 11203
rect 19073 11169 19107 11203
rect 19993 11169 20027 11203
rect 6837 11101 6871 11135
rect 8217 11101 8251 11135
rect 11345 11101 11379 11135
rect 16497 11101 16531 11135
rect 18061 11101 18095 11135
rect 18245 11101 18279 11135
rect 9873 11033 9907 11067
rect 14933 11033 14967 11067
rect 15669 11033 15703 11067
rect 17601 11033 17635 11067
rect 19257 11033 19291 11067
rect 19717 11033 19751 11067
rect 22017 11033 22051 11067
rect 3893 10965 3927 10999
rect 6469 10965 6503 10999
rect 7389 10965 7423 10999
rect 7665 10965 7699 10999
rect 16037 10965 16071 10999
rect 17233 10965 17267 10999
rect 21373 10965 21407 10999
rect 2145 10761 2179 10795
rect 3065 10761 3099 10795
rect 5273 10761 5307 10795
rect 6561 10761 6595 10795
rect 16497 10761 16531 10795
rect 18153 10761 18187 10795
rect 20637 10761 20671 10795
rect 1869 10693 1903 10727
rect 3525 10625 3559 10659
rect 5641 10625 5675 10659
rect 9689 10625 9723 10659
rect 11069 10625 11103 10659
rect 12817 10625 12851 10659
rect 14473 10625 14507 10659
rect 17601 10625 17635 10659
rect 2329 10557 2363 10591
rect 2789 10557 2823 10591
rect 3249 10557 3283 10591
rect 3893 10557 3927 10591
rect 8401 10557 8435 10591
rect 14729 10557 14763 10591
rect 17693 10557 17727 10591
rect 19257 10557 19291 10591
rect 21097 10557 21131 10591
rect 1685 10489 1719 10523
rect 4160 10489 4194 10523
rect 8134 10489 8168 10523
rect 9873 10489 9907 10523
rect 10517 10489 10551 10523
rect 17785 10489 17819 10523
rect 19502 10489 19536 10523
rect 21281 10489 21315 10523
rect 2605 10421 2639 10455
rect 6009 10421 6043 10455
rect 7021 10421 7055 10455
rect 8677 10421 8711 10455
rect 9045 10421 9079 10455
rect 9781 10421 9815 10455
rect 10241 10421 10275 10455
rect 13645 10421 13679 10455
rect 15853 10421 15887 10455
rect 17049 10421 17083 10455
rect 18429 10421 18463 10455
rect 18889 10421 18923 10455
rect 3065 10217 3099 10251
rect 4905 10217 4939 10251
rect 5365 10217 5399 10251
rect 5917 10217 5951 10251
rect 6929 10217 6963 10251
rect 8125 10217 8159 10251
rect 9137 10217 9171 10251
rect 11345 10217 11379 10251
rect 11805 10217 11839 10251
rect 14565 10217 14599 10251
rect 15301 10217 15335 10251
rect 17049 10217 17083 10251
rect 17141 10217 17175 10251
rect 19165 10217 19199 10251
rect 20637 10217 20671 10251
rect 3893 10149 3927 10183
rect 5273 10149 5307 10183
rect 7389 10149 7423 10183
rect 9934 10149 9968 10183
rect 14013 10149 14047 10183
rect 1685 10081 1719 10115
rect 2697 10081 2731 10115
rect 3341 10081 3375 10115
rect 4261 10081 4295 10115
rect 6285 10081 6319 10115
rect 7297 10081 7331 10115
rect 8585 10081 8619 10115
rect 12265 10081 12299 10115
rect 12532 10081 12566 10115
rect 15209 10081 15243 10115
rect 15853 10081 15887 10115
rect 18052 10081 18086 10115
rect 20545 10081 20579 10115
rect 21189 10081 21223 10115
rect 2421 10013 2455 10047
rect 2605 10013 2639 10047
rect 5457 10013 5491 10047
rect 6377 10013 6411 10047
rect 6561 10013 6595 10047
rect 7481 10013 7515 10047
rect 9689 10013 9723 10047
rect 15393 10013 15427 10047
rect 16957 10013 16991 10047
rect 17785 10013 17819 10047
rect 20821 10013 20855 10047
rect 3525 9945 3559 9979
rect 11069 9945 11103 9979
rect 16497 9945 16531 9979
rect 1777 9877 1811 9911
rect 8401 9877 8435 9911
rect 13645 9877 13679 9911
rect 14841 9877 14875 9911
rect 16037 9877 16071 9911
rect 17509 9877 17543 9911
rect 19625 9877 19659 9911
rect 20177 9877 20211 9911
rect 18521 9673 18555 9707
rect 3433 9605 3467 9639
rect 7757 9605 7791 9639
rect 9137 9605 9171 9639
rect 13461 9605 13495 9639
rect 19349 9605 19383 9639
rect 21097 9605 21131 9639
rect 7205 9537 7239 9571
rect 7389 9537 7423 9571
rect 8309 9537 8343 9571
rect 10149 9537 10183 9571
rect 1593 9469 1627 9503
rect 2053 9469 2087 9503
rect 3709 9469 3743 9503
rect 4445 9469 4479 9503
rect 6101 9469 6135 9503
rect 10333 9469 10367 9503
rect 11897 9469 11931 9503
rect 2298 9401 2332 9435
rect 4813 9401 4847 9435
rect 7113 9401 7147 9435
rect 8217 9401 8251 9435
rect 12142 9401 12176 9435
rect 15209 9537 15243 9571
rect 16221 9537 16255 9571
rect 16313 9537 16347 9571
rect 17141 9537 17175 9571
rect 20269 9537 20303 9571
rect 20453 9537 20487 9571
rect 13553 9469 13587 9503
rect 19533 9469 19567 9503
rect 20177 9469 20211 9503
rect 13798 9401 13832 9435
rect 17408 9401 17442 9435
rect 19073 9401 19107 9435
rect 21281 9401 21315 9435
rect 1685 9333 1719 9367
rect 4077 9333 4111 9367
rect 5181 9333 5215 9367
rect 5549 9333 5583 9367
rect 5917 9333 5951 9367
rect 6745 9333 6779 9367
rect 8125 9333 8159 9367
rect 8769 9333 8803 9367
rect 9689 9333 9723 9367
rect 10241 9333 10275 9367
rect 10701 9333 10735 9367
rect 11069 9333 11103 9367
rect 13277 9333 13311 9367
rect 13461 9333 13495 9367
rect 14933 9333 14967 9367
rect 15761 9333 15795 9367
rect 16129 9333 16163 9367
rect 19809 9333 19843 9367
rect 2513 9129 2547 9163
rect 2789 9129 2823 9163
rect 5457 9129 5491 9163
rect 7113 9129 7147 9163
rect 7757 9129 7791 9163
rect 10333 9129 10367 9163
rect 11621 9129 11655 9163
rect 12081 9129 12115 9163
rect 13553 9129 13587 9163
rect 13645 9129 13679 9163
rect 14013 9129 14047 9163
rect 14197 9129 14231 9163
rect 14841 9129 14875 9163
rect 15301 9129 15335 9163
rect 15853 9129 15887 9163
rect 16313 9129 16347 9163
rect 18981 9129 19015 9163
rect 4322 9061 4356 9095
rect 14933 9061 14967 9095
rect 18889 9061 18923 9095
rect 20922 9061 20956 9095
rect 2145 8993 2179 9027
rect 3157 8993 3191 9027
rect 5733 8993 5767 9027
rect 6000 8993 6034 9027
rect 9689 8993 9723 9027
rect 10701 8993 10735 9027
rect 11713 8993 11747 9027
rect 12449 8993 12483 9027
rect 14197 8993 14231 9027
rect 15945 8993 15979 9027
rect 16589 8993 16623 9027
rect 1869 8925 1903 8959
rect 2053 8925 2087 8959
rect 3249 8925 3283 8959
rect 3341 8925 3375 8959
rect 4077 8925 4111 8959
rect 7849 8925 7883 8959
rect 7941 8925 7975 8959
rect 9413 8925 9447 8959
rect 9597 8925 9631 8959
rect 10793 8925 10827 8959
rect 10885 8925 10919 8959
rect 11437 8925 11471 8959
rect 13461 8925 13495 8959
rect 14105 8925 14139 8959
rect 14657 8925 14691 8959
rect 15669 8925 15703 8959
rect 17509 8925 17543 8959
rect 19165 8925 19199 8959
rect 21189 8925 21223 8959
rect 8677 8857 8711 8891
rect 10057 8857 10091 8891
rect 17141 8857 17175 8891
rect 19809 8857 19843 8891
rect 1409 8789 1443 8823
rect 7389 8789 7423 8823
rect 12817 8789 12851 8823
rect 14105 8789 14139 8823
rect 16773 8789 16807 8823
rect 17877 8789 17911 8823
rect 18153 8789 18187 8823
rect 18521 8789 18555 8823
rect 3893 8585 3927 8619
rect 6653 8585 6687 8619
rect 12449 8585 12483 8619
rect 21189 8585 21223 8619
rect 1869 8517 1903 8551
rect 5365 8517 5399 8551
rect 8493 8517 8527 8551
rect 10149 8517 10183 8551
rect 12725 8517 12759 8551
rect 14565 8517 14599 8551
rect 16589 8517 16623 8551
rect 18337 8517 18371 8551
rect 4537 8449 4571 8483
rect 7113 8449 7147 8483
rect 7297 8449 7331 8483
rect 7941 8449 7975 8483
rect 8033 8449 8067 8483
rect 10793 8449 10827 8483
rect 17693 8449 17727 8483
rect 18797 8449 18831 8483
rect 3249 8381 3283 8415
rect 3617 8381 3651 8415
rect 4353 8381 4387 8415
rect 5089 8381 5123 8415
rect 5733 8381 5767 8415
rect 7021 8381 7055 8415
rect 8125 8381 8159 8415
rect 8769 8381 8803 8415
rect 9036 8381 9070 8415
rect 13838 8381 13872 8415
rect 14105 8381 14139 8415
rect 15209 8381 15243 8415
rect 17601 8381 17635 8415
rect 18521 8381 18555 8415
rect 19064 8381 19098 8415
rect 20545 8381 20579 8415
rect 21281 8381 21315 8415
rect 3004 8313 3038 8347
rect 10885 8313 10919 8347
rect 10977 8313 11011 8347
rect 11897 8313 11931 8347
rect 14841 8313 14875 8347
rect 15476 8313 15510 8347
rect 20729 8313 20763 8347
rect 1593 8245 1627 8279
rect 4261 8245 4295 8279
rect 4905 8245 4939 8279
rect 11345 8245 11379 8279
rect 17141 8245 17175 8279
rect 17509 8245 17543 8279
rect 20177 8245 20211 8279
rect 2421 8041 2455 8075
rect 2789 8041 2823 8075
rect 4261 8041 4295 8075
rect 10333 8041 10367 8075
rect 16589 8041 16623 8075
rect 16957 8041 16991 8075
rect 17325 8041 17359 8075
rect 17785 8041 17819 8075
rect 1685 7973 1719 8007
rect 3433 7973 3467 8007
rect 4169 7973 4203 8007
rect 6469 7973 6503 8007
rect 9137 7973 9171 8007
rect 11814 7973 11848 8007
rect 13277 7973 13311 8007
rect 14832 7973 14866 8007
rect 16497 7973 16531 8007
rect 20729 7973 20763 8007
rect 2881 7905 2915 7939
rect 5457 7905 5491 7939
rect 7941 7905 7975 7939
rect 8493 7905 8527 7939
rect 12541 7905 12575 7939
rect 12633 7905 12667 7939
rect 13185 7905 13219 7939
rect 14013 7905 14047 7939
rect 17693 7905 17727 7939
rect 18337 7905 18371 7939
rect 19073 7905 19107 7939
rect 19809 7905 19843 7939
rect 20085 7905 20119 7939
rect 21281 7905 21315 7939
rect 22017 7905 22051 7939
rect 3065 7837 3099 7871
rect 4629 7837 4663 7871
rect 5181 7837 5215 7871
rect 5365 7837 5399 7871
rect 7573 7837 7607 7871
rect 9505 7837 9539 7871
rect 12081 7837 12115 7871
rect 1869 7769 1903 7803
rect 5825 7769 5859 7803
rect 9965 7769 9999 7803
rect 13369 7837 13403 7871
rect 14565 7837 14599 7871
rect 16405 7837 16439 7871
rect 17877 7837 17911 7871
rect 20545 7837 20579 7871
rect 21097 7769 21131 7803
rect 6101 7701 6135 7735
rect 6929 7701 6963 7735
rect 7205 7701 7239 7735
rect 8677 7701 8711 7735
rect 10701 7701 10735 7735
rect 12633 7701 12667 7735
rect 12817 7701 12851 7735
rect 13829 7701 13863 7735
rect 15945 7701 15979 7735
rect 19257 7701 19291 7735
rect 20269 7701 20303 7735
rect 2329 7497 2363 7531
rect 3525 7497 3559 7531
rect 5273 7497 5307 7531
rect 9137 7497 9171 7531
rect 10885 7497 10919 7531
rect 14013 7497 14047 7531
rect 14197 7497 14231 7531
rect 14381 7497 14415 7531
rect 16221 7497 16255 7531
rect 18521 7497 18555 7531
rect 20821 7497 20855 7531
rect 1869 7429 1903 7463
rect 9505 7429 9539 7463
rect 9965 7429 9999 7463
rect 13645 7429 13679 7463
rect 2789 7361 2823 7395
rect 2973 7361 3007 7395
rect 4445 7361 4479 7395
rect 4537 7361 4571 7395
rect 5825 7361 5859 7395
rect 2697 7293 2731 7327
rect 4629 7293 4663 7327
rect 5733 7293 5767 7327
rect 7757 7293 7791 7327
rect 1685 7225 1719 7259
rect 3433 7225 3467 7259
rect 6837 7225 6871 7259
rect 8002 7225 8036 7259
rect 10333 7361 10367 7395
rect 12817 7361 12851 7395
rect 12909 7361 12943 7395
rect 21097 7429 21131 7463
rect 15117 7361 15151 7395
rect 16313 7361 16347 7395
rect 16589 7361 16623 7395
rect 20269 7361 20303 7395
rect 11253 7293 11287 7327
rect 14197 7293 14231 7327
rect 15485 7293 15519 7327
rect 10149 7225 10183 7259
rect 10333 7225 10367 7259
rect 17141 7293 17175 7327
rect 19073 7293 19107 7327
rect 21281 7293 21315 7327
rect 17386 7225 17420 7259
rect 20177 7225 20211 7259
rect 3893 7157 3927 7191
rect 4997 7157 5031 7191
rect 5641 7157 5675 7191
rect 6469 7157 6503 7191
rect 7297 7157 7331 7191
rect 9781 7157 9815 7191
rect 9965 7157 9999 7191
rect 10609 7157 10643 7191
rect 11713 7157 11747 7191
rect 12357 7157 12391 7191
rect 12725 7157 12759 7191
rect 14657 7157 14691 7191
rect 15853 7157 15887 7191
rect 16313 7157 16347 7191
rect 18889 7157 18923 7191
rect 19349 7157 19383 7191
rect 19717 7157 19751 7191
rect 20085 7157 20119 7191
rect 2789 6953 2823 6987
rect 5825 6953 5859 6987
rect 7757 6953 7791 6987
rect 8401 6953 8435 6987
rect 12357 6953 12391 6987
rect 16681 6953 16715 6987
rect 17601 6953 17635 6987
rect 19257 6953 19291 6987
rect 1961 6885 1995 6919
rect 4690 6885 4724 6919
rect 20076 6885 20110 6919
rect 22017 6885 22051 6919
rect 2697 6817 2731 6851
rect 3349 6817 3383 6851
rect 6377 6817 6411 6851
rect 6644 6817 6678 6851
rect 9505 6817 9539 6851
rect 10241 6817 10275 6851
rect 10508 6817 10542 6851
rect 12265 6817 12299 6851
rect 14657 6817 14691 6851
rect 15568 6817 15602 6851
rect 17785 6817 17819 6851
rect 18061 6817 18095 6851
rect 18889 6817 18923 6851
rect 19809 6817 19843 6851
rect 2053 6749 2087 6783
rect 2237 6749 2271 6783
rect 4445 6749 4479 6783
rect 8125 6749 8159 6783
rect 8309 6749 8343 6783
rect 9873 6749 9907 6783
rect 12449 6749 12483 6783
rect 15301 6749 15335 6783
rect 17233 6749 17267 6783
rect 18705 6749 18739 6783
rect 18797 6749 18831 6783
rect 3157 6681 3191 6715
rect 8769 6681 8803 6715
rect 1593 6613 1627 6647
rect 3893 6613 3927 6647
rect 9137 6613 9171 6647
rect 11621 6613 11655 6647
rect 11897 6613 11931 6647
rect 13185 6613 13219 6647
rect 13645 6613 13679 6647
rect 15025 6613 15059 6647
rect 18245 6613 18279 6647
rect 21189 6613 21223 6647
rect 3985 6409 4019 6443
rect 4905 6409 4939 6443
rect 6101 6409 6135 6443
rect 11529 6409 11563 6443
rect 19993 6409 20027 6443
rect 4445 6341 4479 6375
rect 1685 6273 1719 6307
rect 3065 6273 3099 6307
rect 3525 6273 3559 6307
rect 5549 6273 5583 6307
rect 7297 6273 7331 6307
rect 1869 6205 1903 6239
rect 2881 6205 2915 6239
rect 4169 6205 4203 6239
rect 4629 6205 4663 6239
rect 4721 6205 4755 6239
rect 5089 6205 5123 6239
rect 7021 6205 7055 6239
rect 7113 6205 7147 6239
rect 9689 6205 9723 6239
rect 1777 6137 1811 6171
rect 18337 6341 18371 6375
rect 13369 6273 13403 6307
rect 14749 6273 14783 6307
rect 16037 6273 16071 6307
rect 17601 6273 17635 6307
rect 17693 6273 17727 6307
rect 19533 6273 19567 6307
rect 13461 6205 13495 6239
rect 14657 6205 14691 6239
rect 17509 6205 17543 6239
rect 18153 6205 18187 6239
rect 18797 6205 18831 6239
rect 19257 6205 19291 6239
rect 21106 6205 21140 6239
rect 21373 6205 21407 6239
rect 5641 6137 5675 6171
rect 9422 6137 9456 6171
rect 11529 6137 11563 6171
rect 13553 6137 13587 6171
rect 16221 6137 16255 6171
rect 2237 6069 2271 6103
rect 2513 6069 2547 6103
rect 2973 6069 3007 6103
rect 4721 6069 4755 6103
rect 5733 6069 5767 6103
rect 6653 6069 6687 6103
rect 7665 6069 7699 6103
rect 8309 6069 8343 6103
rect 9965 6069 9999 6103
rect 10333 6069 10367 6103
rect 10793 6069 10827 6103
rect 11253 6069 11287 6103
rect 11805 6069 11839 6103
rect 12265 6069 12299 6103
rect 12725 6069 12759 6103
rect 13921 6069 13955 6103
rect 14197 6069 14231 6103
rect 14565 6069 14599 6103
rect 15577 6069 15611 6103
rect 16129 6069 16163 6103
rect 16589 6069 16623 6103
rect 17141 6069 17175 6103
rect 18613 6069 18647 6103
rect 19073 6069 19107 6103
rect 3525 5865 3559 5899
rect 5457 5865 5491 5899
rect 6101 5865 6135 5899
rect 6561 5865 6595 5899
rect 7389 5865 7423 5899
rect 8769 5865 8803 5899
rect 9689 5865 9723 5899
rect 14565 5865 14599 5899
rect 15485 5865 15519 5899
rect 16497 5865 16531 5899
rect 21189 5865 21223 5899
rect 1685 5797 1719 5831
rect 4322 5797 4356 5831
rect 11560 5797 11594 5831
rect 16037 5797 16071 5831
rect 18153 5797 18187 5831
rect 18245 5797 18279 5831
rect 20269 5797 20303 5831
rect 2145 5729 2179 5763
rect 2412 5729 2446 5763
rect 4077 5729 4111 5763
rect 6469 5729 6503 5763
rect 7573 5729 7607 5763
rect 8401 5729 8435 5763
rect 9781 5729 9815 5763
rect 12900 5729 12934 5763
rect 15301 5729 15335 5763
rect 16129 5729 16163 5763
rect 16773 5729 16807 5763
rect 17233 5729 17267 5763
rect 19073 5729 19107 5763
rect 20177 5729 20211 5763
rect 21281 5729 21315 5763
rect 6653 5661 6687 5695
rect 8217 5661 8251 5695
rect 8309 5661 8343 5695
rect 9873 5661 9907 5695
rect 11805 5661 11839 5695
rect 12081 5661 12115 5695
rect 12633 5661 12667 5695
rect 15853 5661 15887 5695
rect 17969 5661 18003 5695
rect 20361 5661 20395 5695
rect 9321 5593 9355 5627
rect 16957 5593 16991 5627
rect 1777 5525 1811 5559
rect 5825 5525 5859 5559
rect 10425 5525 10459 5559
rect 14013 5525 14047 5559
rect 17417 5525 17451 5559
rect 18613 5525 18647 5559
rect 19257 5525 19291 5559
rect 19809 5525 19843 5559
rect 7481 5321 7515 5355
rect 7757 5321 7791 5355
rect 9137 5321 9171 5355
rect 13277 5321 13311 5355
rect 16129 5321 16163 5355
rect 4445 5253 4479 5287
rect 5733 5253 5767 5287
rect 7297 5253 7331 5287
rect 2881 5185 2915 5219
rect 3065 5185 3099 5219
rect 3985 5185 4019 5219
rect 1409 5117 1443 5151
rect 1869 5117 1903 5151
rect 4629 5117 4663 5151
rect 5089 5117 5123 5151
rect 5549 5117 5583 5151
rect 7113 5117 7147 5151
rect 2789 5049 2823 5083
rect 3893 5049 3927 5083
rect 6009 5049 6043 5083
rect 10333 5253 10367 5287
rect 16681 5253 16715 5287
rect 8585 5185 8619 5219
rect 8769 5185 8803 5219
rect 9781 5185 9815 5219
rect 11253 5185 11287 5219
rect 11897 5185 11931 5219
rect 14013 5185 14047 5219
rect 14105 5185 14139 5219
rect 14841 5185 14875 5219
rect 19165 5185 19199 5219
rect 20821 5185 20855 5219
rect 7573 5117 7607 5151
rect 9321 5117 9355 5151
rect 10517 5117 10551 5151
rect 11069 5117 11103 5151
rect 12153 5117 12187 5151
rect 14933 5117 14967 5151
rect 15945 5117 15979 5151
rect 16405 5117 16439 5151
rect 16681 5117 16715 5151
rect 17509 5117 17543 5151
rect 17765 5117 17799 5151
rect 19432 5117 19466 5151
rect 9873 5049 9907 5083
rect 13921 5049 13955 5083
rect 1593 4981 1627 5015
rect 2053 4981 2087 5015
rect 2421 4981 2455 5015
rect 3433 4981 3467 5015
rect 3801 4981 3835 5015
rect 5273 4981 5307 5015
rect 6837 4981 6871 5015
rect 7481 4981 7515 5015
rect 8125 4981 8159 5015
rect 8493 4981 8527 5015
rect 9965 4981 9999 5015
rect 10517 4981 10551 5015
rect 10609 4981 10643 5015
rect 10977 4981 11011 5015
rect 13553 4981 13587 5015
rect 15025 4981 15059 5015
rect 15393 4981 15427 5015
rect 16589 4981 16623 5015
rect 17049 4981 17083 5015
rect 18889 4981 18923 5015
rect 20545 4981 20579 5015
rect 21373 4981 21407 5015
rect 2513 4777 2547 4811
rect 2973 4777 3007 4811
rect 3433 4777 3467 4811
rect 5181 4777 5215 4811
rect 6285 4777 6319 4811
rect 8217 4777 8251 4811
rect 9781 4777 9815 4811
rect 10977 4777 11011 4811
rect 11345 4777 11379 4811
rect 13553 4777 13587 4811
rect 15117 4777 15151 4811
rect 18245 4777 18279 4811
rect 20177 4777 20211 4811
rect 1685 4709 1719 4743
rect 6193 4709 6227 4743
rect 7205 4709 7239 4743
rect 8309 4709 8343 4743
rect 11989 4709 12023 4743
rect 18337 4709 18371 4743
rect 21281 4709 21315 4743
rect 2605 4641 2639 4675
rect 3249 4641 3283 4675
rect 4077 4641 4111 4675
rect 9965 4641 9999 4675
rect 12909 4641 12943 4675
rect 13369 4641 13403 4675
rect 13829 4641 13863 4675
rect 14657 4641 14691 4675
rect 14933 4641 14967 4675
rect 15393 4641 15427 4675
rect 15853 4641 15887 4675
rect 16120 4641 16154 4675
rect 17693 4641 17727 4675
rect 19073 4641 19107 4675
rect 2329 4573 2363 4607
rect 4997 4573 5031 4607
rect 5089 4573 5123 4607
rect 6377 4573 6411 4607
rect 7297 4573 7331 4607
rect 7389 4573 7423 4607
rect 8125 4573 8159 4607
rect 9321 4573 9355 4607
rect 10241 4573 10275 4607
rect 11437 4573 11471 4607
rect 11621 4573 11655 4607
rect 18153 4573 18187 4607
rect 20269 4573 20303 4607
rect 20453 4573 20487 4607
rect 12357 4505 12391 4539
rect 13093 4505 13127 4539
rect 14013 4505 14047 4539
rect 17233 4505 17267 4539
rect 18705 4505 18739 4539
rect 21097 4505 21131 4539
rect 1777 4437 1811 4471
rect 4261 4437 4295 4471
rect 5549 4437 5583 4471
rect 5825 4437 5859 4471
rect 6837 4437 6871 4471
rect 8677 4437 8711 4471
rect 10609 4437 10643 4471
rect 15577 4437 15611 4471
rect 17509 4437 17543 4471
rect 19257 4437 19291 4471
rect 19809 4437 19843 4471
rect 1501 4233 1535 4267
rect 3157 4233 3191 4267
rect 10057 4233 10091 4267
rect 12081 4233 12115 4267
rect 12357 4233 12391 4267
rect 4353 4165 4387 4199
rect 18153 4165 18187 4199
rect 3709 4097 3743 4131
rect 5457 4097 5491 4131
rect 7389 4097 7423 4131
rect 15301 4097 15335 4131
rect 15393 4097 15427 4131
rect 21097 4097 21131 4131
rect 2881 4029 2915 4063
rect 4169 4029 4203 4063
rect 5365 4029 5399 4063
rect 5733 4029 5767 4063
rect 6101 4029 6135 4063
rect 6653 4029 6687 4063
rect 8309 4029 8343 4063
rect 10241 4029 10275 4063
rect 10701 4029 10735 4063
rect 11161 4029 11195 4063
rect 11897 4029 11931 4063
rect 12541 4029 12575 4063
rect 12817 4029 12851 4063
rect 13461 4029 13495 4063
rect 13728 4029 13762 4063
rect 17877 4029 17911 4063
rect 18337 4029 18371 4063
rect 18889 4029 18923 4063
rect 19349 4029 19383 4063
rect 20830 4029 20864 4063
rect 2614 3961 2648 3995
rect 5273 3961 5307 3995
rect 7573 3961 7607 3995
rect 7665 3961 7699 3995
rect 8576 3961 8610 3995
rect 15485 3961 15519 3995
rect 17141 3961 17175 3995
rect 17325 3961 17359 3995
rect 3525 3893 3559 3927
rect 3617 3893 3651 3927
rect 4905 3893 4939 3927
rect 5733 3893 5767 3927
rect 5917 3893 5951 3927
rect 6837 3893 6871 3927
rect 8033 3893 8067 3927
rect 9689 3893 9723 3927
rect 10517 3893 10551 3927
rect 10977 3893 11011 3927
rect 13001 3893 13035 3927
rect 14841 3893 14875 3927
rect 15853 3893 15887 3927
rect 16405 3893 16439 3927
rect 17693 3893 17727 3927
rect 18705 3893 18739 3927
rect 19165 3893 19199 3927
rect 19717 3893 19751 3927
rect 1685 3689 1719 3723
rect 4261 3689 4295 3723
rect 5733 3689 5767 3723
rect 6377 3689 6411 3723
rect 8401 3689 8435 3723
rect 10977 3689 11011 3723
rect 11345 3689 11379 3723
rect 16221 3689 16255 3723
rect 16865 3689 16899 3723
rect 18061 3689 18095 3723
rect 19717 3689 19751 3723
rect 8309 3621 8343 3655
rect 10517 3621 10551 3655
rect 2798 3553 2832 3587
rect 3341 3553 3375 3587
rect 4077 3553 4111 3587
rect 4445 3553 4479 3587
rect 4537 3553 4571 3587
rect 5641 3553 5675 3587
rect 7501 3553 7535 3587
rect 9781 3553 9815 3587
rect 10609 3553 10643 3587
rect 3065 3485 3099 3519
rect 3525 3417 3559 3451
rect 12541 3621 12575 3655
rect 17693 3621 17727 3655
rect 20177 3621 20211 3655
rect 11161 3553 11195 3587
rect 11621 3553 11655 3587
rect 12173 3553 12207 3587
rect 5825 3485 5859 3519
rect 7757 3485 7791 3519
rect 8217 3485 8251 3519
rect 10793 3485 10827 3519
rect 10977 3485 11011 3519
rect 9137 3417 9171 3451
rect 9597 3417 9631 3451
rect 11805 3417 11839 3451
rect 12633 3553 12667 3587
rect 13369 3553 13403 3587
rect 13645 3553 13679 3587
rect 14841 3553 14875 3587
rect 15108 3553 15142 3587
rect 18245 3553 18279 3587
rect 18705 3553 18739 3587
rect 19165 3553 19199 3587
rect 20821 3553 20855 3587
rect 16957 3485 16991 3519
rect 17049 3485 17083 3519
rect 20545 3485 20579 3519
rect 14381 3417 14415 3451
rect 17509 3417 17543 3451
rect 19993 3417 20027 3451
rect 4445 3349 4479 3383
rect 4721 3349 4755 3383
rect 5273 3349 5307 3383
rect 8769 3349 8803 3383
rect 10149 3349 10183 3383
rect 12357 3349 12391 3383
rect 12541 3349 12575 3383
rect 12817 3349 12851 3383
rect 13185 3349 13219 3383
rect 13829 3349 13863 3383
rect 16497 3349 16531 3383
rect 18521 3349 18555 3383
rect 18981 3349 19015 3383
rect 1777 3145 1811 3179
rect 6653 3145 6687 3179
rect 8033 3145 8067 3179
rect 12173 3145 12207 3179
rect 15393 3145 15427 3179
rect 17785 3145 17819 3179
rect 7665 3077 7699 3111
rect 7205 3009 7239 3043
rect 9597 3009 9631 3043
rect 10609 3009 10643 3043
rect 10793 3009 10827 3043
rect 2237 2941 2271 2975
rect 4169 2941 4203 2975
rect 5825 2941 5859 2975
rect 7021 2941 7055 2975
rect 9157 2941 9191 2975
rect 9413 2941 9447 2975
rect 1685 2873 1719 2907
rect 2421 2873 2455 2907
rect 3924 2873 3958 2907
rect 5580 2873 5614 2907
rect 12541 3077 12575 3111
rect 13093 3077 13127 3111
rect 16589 3077 16623 3111
rect 15853 3009 15887 3043
rect 16037 3009 16071 3043
rect 9689 2941 9723 2975
rect 11161 2941 11195 2975
rect 11897 2941 11931 2975
rect 12173 2941 12207 2975
rect 12357 2941 12391 2975
rect 12909 2941 12943 2975
rect 13553 2941 13587 2975
rect 13829 2941 13863 2975
rect 15761 2941 15795 2975
rect 16405 2941 16439 2975
rect 17877 2941 17911 2975
rect 18613 2941 18647 2975
rect 19274 2941 19308 2975
rect 19809 2941 19843 2975
rect 21097 2941 21131 2975
rect 10517 2873 10551 2907
rect 14565 2873 14599 2907
rect 14749 2873 14783 2907
rect 17325 2873 17359 2907
rect 19073 2873 19107 2907
rect 19625 2873 19659 2907
rect 20453 2873 20487 2907
rect 2789 2805 2823 2839
rect 4445 2805 4479 2839
rect 7113 2805 7147 2839
rect 9597 2805 9631 2839
rect 9873 2805 9907 2839
rect 10149 2805 10183 2839
rect 11345 2805 11379 2839
rect 12081 2805 12115 2839
rect 13369 2805 13403 2839
rect 14013 2805 14047 2839
rect 17233 2805 17267 2839
rect 18705 2805 18739 2839
rect 2881 2601 2915 2635
rect 3341 2601 3375 2635
rect 5457 2601 5491 2635
rect 5641 2601 5675 2635
rect 5917 2601 5951 2635
rect 7389 2601 7423 2635
rect 8493 2601 8527 2635
rect 8861 2601 8895 2635
rect 10057 2601 10091 2635
rect 10609 2601 10643 2635
rect 20085 2601 20119 2635
rect 1685 2533 1719 2567
rect 1869 2533 1903 2567
rect 2421 2533 2455 2567
rect 4169 2533 4203 2567
rect 5089 2533 5123 2567
rect 2237 2465 2271 2499
rect 2697 2465 2731 2499
rect 3157 2465 3191 2499
rect 4353 2465 4387 2499
rect 9965 2533 9999 2567
rect 12357 2533 12391 2567
rect 13001 2533 13035 2567
rect 14105 2533 14139 2567
rect 16129 2533 16163 2567
rect 17601 2533 17635 2567
rect 18153 2533 18187 2567
rect 18797 2533 18831 2567
rect 19441 2533 19475 2567
rect 5733 2465 5767 2499
rect 6745 2465 6779 2499
rect 7205 2465 7239 2499
rect 7849 2465 7883 2499
rect 10793 2465 10827 2499
rect 11345 2465 11379 2499
rect 13553 2465 13587 2499
rect 15025 2465 15059 2499
rect 15577 2465 15611 2499
rect 16681 2465 16715 2499
rect 19257 2465 19291 2499
rect 20269 2465 20303 2499
rect 20821 2465 20855 2499
rect 4813 2397 4847 2431
rect 4997 2397 5031 2431
rect 5641 2397 5675 2431
rect 8217 2397 8251 2431
rect 8401 2397 8435 2431
rect 10149 2397 10183 2431
rect 11897 2397 11931 2431
rect 15761 2397 15795 2431
rect 20545 2397 20579 2431
rect 7665 2329 7699 2363
rect 9597 2329 9631 2363
rect 11529 2329 11563 2363
rect 12817 2329 12851 2363
rect 13369 2329 13403 2363
rect 13921 2329 13955 2363
rect 15209 2329 15243 2363
rect 16313 2329 16347 2363
rect 17417 2329 17451 2363
rect 17969 2329 18003 2363
rect 18981 2329 19015 2363
rect 6929 2261 6963 2295
rect 9229 2261 9263 2295
rect 12449 2261 12483 2295
rect 14565 2261 14599 2295
rect 16773 2261 16807 2295
<< metal1 >>
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 2222 20584 2228 20596
rect 2183 20556 2228 20584
rect 2222 20544 2228 20556
rect 2280 20544 2286 20596
rect 2685 20519 2743 20525
rect 2685 20485 2697 20519
rect 2731 20516 2743 20519
rect 2774 20516 2780 20528
rect 2731 20488 2780 20516
rect 2731 20485 2743 20488
rect 2685 20479 2743 20485
rect 2774 20476 2780 20488
rect 2832 20476 2838 20528
rect 3234 20516 3240 20528
rect 3195 20488 3240 20516
rect 3234 20476 3240 20488
rect 3292 20476 3298 20528
rect 4062 20516 4068 20528
rect 4023 20488 4068 20516
rect 4062 20476 4068 20488
rect 4120 20476 4126 20528
rect 17218 20476 17224 20528
rect 17276 20516 17282 20528
rect 17405 20519 17463 20525
rect 17405 20516 17417 20519
rect 17276 20488 17417 20516
rect 17276 20476 17282 20488
rect 17405 20485 17417 20488
rect 17451 20485 17463 20519
rect 17405 20479 17463 20485
rect 18417 20519 18475 20525
rect 18417 20485 18429 20519
rect 18463 20516 18475 20519
rect 18598 20516 18604 20528
rect 18463 20488 18604 20516
rect 18463 20485 18475 20488
rect 18417 20479 18475 20485
rect 18598 20476 18604 20488
rect 18656 20476 18662 20528
rect 18966 20516 18972 20528
rect 18927 20488 18972 20516
rect 18966 20476 18972 20488
rect 19024 20476 19030 20528
rect 19518 20516 19524 20528
rect 19479 20488 19524 20516
rect 19518 20476 19524 20488
rect 19576 20476 19582 20528
rect 1578 20380 1584 20392
rect 1539 20352 1584 20380
rect 1578 20340 1584 20352
rect 1636 20340 1642 20392
rect 1765 20383 1823 20389
rect 1765 20349 1777 20383
rect 1811 20380 1823 20383
rect 2590 20380 2596 20392
rect 1811 20352 2596 20380
rect 1811 20349 1823 20352
rect 1765 20343 1823 20349
rect 2590 20340 2596 20352
rect 2648 20340 2654 20392
rect 4154 20340 4160 20392
rect 4212 20380 4218 20392
rect 4801 20383 4859 20389
rect 4801 20380 4813 20383
rect 4212 20352 4813 20380
rect 4212 20340 4218 20352
rect 4801 20349 4813 20352
rect 4847 20380 4859 20383
rect 5077 20383 5135 20389
rect 5077 20380 5089 20383
rect 4847 20352 5089 20380
rect 4847 20349 4859 20352
rect 4801 20343 4859 20349
rect 5077 20349 5089 20352
rect 5123 20349 5135 20383
rect 5718 20380 5724 20392
rect 5679 20352 5724 20380
rect 5077 20343 5135 20349
rect 5718 20340 5724 20352
rect 5776 20380 5782 20392
rect 6549 20383 6607 20389
rect 6549 20380 6561 20383
rect 5776 20352 6561 20380
rect 5776 20340 5782 20352
rect 6549 20349 6561 20352
rect 6595 20349 6607 20383
rect 6549 20343 6607 20349
rect 18233 20383 18291 20389
rect 18233 20349 18245 20383
rect 18279 20380 18291 20383
rect 19702 20380 19708 20392
rect 18279 20352 19708 20380
rect 18279 20349 18291 20352
rect 18233 20343 18291 20349
rect 19702 20340 19708 20352
rect 19760 20340 19766 20392
rect 20254 20380 20260 20392
rect 20215 20352 20260 20380
rect 20254 20340 20260 20352
rect 20312 20340 20318 20392
rect 2314 20312 2320 20324
rect 2275 20284 2320 20312
rect 2314 20272 2320 20284
rect 2372 20272 2378 20324
rect 2866 20312 2872 20324
rect 2827 20284 2872 20312
rect 2866 20272 2872 20284
rect 2924 20272 2930 20324
rect 2958 20272 2964 20324
rect 3016 20312 3022 20324
rect 3421 20315 3479 20321
rect 3421 20312 3433 20315
rect 3016 20284 3433 20312
rect 3016 20272 3022 20284
rect 3421 20281 3433 20284
rect 3467 20281 3479 20315
rect 4246 20312 4252 20324
rect 4207 20284 4252 20312
rect 3421 20275 3479 20281
rect 4246 20272 4252 20284
rect 4304 20272 4310 20324
rect 9674 20272 9680 20324
rect 9732 20312 9738 20324
rect 17589 20315 17647 20321
rect 17589 20312 17601 20315
rect 9732 20284 17601 20312
rect 9732 20272 9738 20284
rect 17589 20281 17601 20284
rect 17635 20281 17647 20315
rect 18782 20312 18788 20324
rect 18743 20284 18788 20312
rect 17589 20275 17647 20281
rect 18782 20272 18788 20284
rect 18840 20272 18846 20324
rect 19334 20312 19340 20324
rect 19295 20284 19340 20312
rect 19334 20272 19340 20284
rect 19392 20272 19398 20324
rect 20622 20312 20628 20324
rect 20583 20284 20628 20312
rect 20622 20272 20628 20284
rect 20680 20272 20686 20324
rect 20806 20312 20812 20324
rect 20767 20284 20812 20312
rect 20806 20272 20812 20284
rect 20864 20272 20870 20324
rect 21177 20315 21235 20321
rect 21177 20281 21189 20315
rect 21223 20281 21235 20315
rect 21177 20275 21235 20281
rect 21361 20315 21419 20321
rect 21361 20281 21373 20315
rect 21407 20312 21419 20315
rect 21450 20312 21456 20324
rect 21407 20284 21456 20312
rect 21407 20281 21419 20284
rect 21361 20275 21419 20281
rect 4617 20247 4675 20253
rect 4617 20213 4629 20247
rect 4663 20244 4675 20247
rect 4982 20244 4988 20256
rect 4663 20216 4988 20244
rect 4663 20213 4675 20216
rect 4617 20207 4675 20213
rect 4982 20204 4988 20216
rect 5040 20204 5046 20256
rect 5902 20244 5908 20256
rect 5863 20216 5908 20244
rect 5902 20204 5908 20216
rect 5960 20204 5966 20256
rect 8113 20247 8171 20253
rect 8113 20213 8125 20247
rect 8159 20244 8171 20247
rect 8202 20244 8208 20256
rect 8159 20216 8208 20244
rect 8159 20213 8171 20216
rect 8113 20207 8171 20213
rect 8202 20204 8208 20216
rect 8260 20204 8266 20256
rect 19518 20204 19524 20256
rect 19576 20244 19582 20256
rect 20073 20247 20131 20253
rect 20073 20244 20085 20247
rect 19576 20216 20085 20244
rect 19576 20204 19582 20216
rect 20073 20213 20085 20216
rect 20119 20213 20131 20247
rect 20073 20207 20131 20213
rect 20254 20204 20260 20256
rect 20312 20244 20318 20256
rect 21192 20244 21220 20275
rect 21450 20272 21456 20284
rect 21508 20272 21514 20324
rect 20312 20216 21220 20244
rect 20312 20204 20318 20216
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 2314 20040 2320 20052
rect 2275 20012 2320 20040
rect 2314 20000 2320 20012
rect 2372 20000 2378 20052
rect 2958 20040 2964 20052
rect 2919 20012 2964 20040
rect 2958 20000 2964 20012
rect 3016 20000 3022 20052
rect 3421 20043 3479 20049
rect 3421 20009 3433 20043
rect 3467 20040 3479 20043
rect 4246 20040 4252 20052
rect 3467 20012 4252 20040
rect 3467 20009 3479 20012
rect 3421 20003 3479 20009
rect 4246 20000 4252 20012
rect 4304 20000 4310 20052
rect 8113 20043 8171 20049
rect 8113 20009 8125 20043
rect 8159 20040 8171 20043
rect 8202 20040 8208 20052
rect 8159 20012 8208 20040
rect 8159 20009 8171 20012
rect 8113 20003 8171 20009
rect 8202 20000 8208 20012
rect 8260 20000 8266 20052
rect 18782 20000 18788 20052
rect 18840 20040 18846 20052
rect 20073 20043 20131 20049
rect 20073 20040 20085 20043
rect 18840 20012 20085 20040
rect 18840 20000 18846 20012
rect 20073 20009 20085 20012
rect 20119 20009 20131 20043
rect 20073 20003 20131 20009
rect 20530 20000 20536 20052
rect 20588 20040 20594 20052
rect 20717 20043 20775 20049
rect 20717 20040 20729 20043
rect 20588 20012 20729 20040
rect 20588 20000 20594 20012
rect 20717 20009 20729 20012
rect 20763 20009 20775 20043
rect 20717 20003 20775 20009
rect 5074 19972 5080 19984
rect 3252 19944 5080 19972
rect 1762 19904 1768 19916
rect 1723 19876 1768 19904
rect 1762 19864 1768 19876
rect 1820 19864 1826 19916
rect 3252 19913 3280 19944
rect 5074 19932 5080 19944
rect 5132 19932 5138 19984
rect 5902 19932 5908 19984
rect 5960 19972 5966 19984
rect 10566 19975 10624 19981
rect 10566 19972 10578 19975
rect 5960 19944 10578 19972
rect 5960 19932 5966 19944
rect 10566 19941 10578 19944
rect 10612 19941 10624 19975
rect 10566 19935 10624 19941
rect 19797 19975 19855 19981
rect 19797 19941 19809 19975
rect 19843 19972 19855 19975
rect 20162 19972 20168 19984
rect 19843 19944 20168 19972
rect 19843 19941 19855 19944
rect 19797 19935 19855 19941
rect 20162 19932 20168 19944
rect 20220 19932 20226 19984
rect 2501 19907 2559 19913
rect 2501 19873 2513 19907
rect 2547 19873 2559 19907
rect 2501 19867 2559 19873
rect 2777 19907 2835 19913
rect 2777 19873 2789 19907
rect 2823 19904 2835 19907
rect 3237 19907 3295 19913
rect 2823 19876 3188 19904
rect 2823 19873 2835 19876
rect 2777 19867 2835 19873
rect 2516 19836 2544 19867
rect 3050 19836 3056 19848
rect 2516 19808 3056 19836
rect 3050 19796 3056 19808
rect 3108 19796 3114 19848
rect 1578 19768 1584 19780
rect 1539 19740 1584 19768
rect 1578 19728 1584 19740
rect 1636 19728 1642 19780
rect 3160 19700 3188 19876
rect 3237 19873 3249 19907
rect 3283 19873 3295 19907
rect 3237 19867 3295 19873
rect 4065 19907 4123 19913
rect 4065 19873 4077 19907
rect 4111 19904 4123 19907
rect 4154 19904 4160 19916
rect 4111 19876 4160 19904
rect 4111 19873 4123 19876
rect 4065 19867 4123 19873
rect 4154 19864 4160 19876
rect 4212 19864 4218 19916
rect 4338 19913 4344 19916
rect 4332 19904 4344 19913
rect 4299 19876 4344 19904
rect 4332 19867 4344 19876
rect 4338 19864 4344 19867
rect 4396 19864 4402 19916
rect 17954 19864 17960 19916
rect 18012 19904 18018 19916
rect 19245 19907 19303 19913
rect 19245 19904 19257 19907
rect 18012 19876 19257 19904
rect 18012 19864 18018 19876
rect 19245 19873 19257 19876
rect 19291 19904 19303 19907
rect 20257 19907 20315 19913
rect 20257 19904 20269 19907
rect 19291 19876 20269 19904
rect 19291 19873 19303 19876
rect 19245 19867 19303 19873
rect 20257 19873 20269 19876
rect 20303 19873 20315 19907
rect 20257 19867 20315 19873
rect 20346 19864 20352 19916
rect 20404 19904 20410 19916
rect 20625 19907 20683 19913
rect 20625 19904 20637 19907
rect 20404 19876 20637 19904
rect 20404 19864 20410 19876
rect 20625 19873 20637 19876
rect 20671 19873 20683 19907
rect 21174 19904 21180 19916
rect 21135 19876 21180 19904
rect 20625 19867 20683 19873
rect 21174 19864 21180 19876
rect 21232 19864 21238 19916
rect 7650 19796 7656 19848
rect 7708 19836 7714 19848
rect 8205 19839 8263 19845
rect 8205 19836 8217 19839
rect 7708 19808 8217 19836
rect 7708 19796 7714 19808
rect 8205 19805 8217 19808
rect 8251 19805 8263 19839
rect 8205 19799 8263 19805
rect 8297 19839 8355 19845
rect 8297 19805 8309 19839
rect 8343 19805 8355 19839
rect 10318 19836 10324 19848
rect 10279 19808 10324 19836
rect 8297 19799 8355 19805
rect 5721 19771 5779 19777
rect 5721 19768 5733 19771
rect 5184 19740 5733 19768
rect 5184 19700 5212 19740
rect 5721 19737 5733 19740
rect 5767 19768 5779 19771
rect 7834 19768 7840 19780
rect 5767 19740 7840 19768
rect 5767 19737 5779 19740
rect 5721 19731 5779 19737
rect 7834 19728 7840 19740
rect 7892 19728 7898 19780
rect 8312 19768 8340 19799
rect 10318 19796 10324 19808
rect 10376 19796 10382 19848
rect 21358 19768 21364 19780
rect 8220 19740 8340 19768
rect 21319 19740 21364 19768
rect 8220 19712 8248 19740
rect 21358 19728 21364 19740
rect 21416 19728 21422 19780
rect 3160 19672 5212 19700
rect 5258 19660 5264 19712
rect 5316 19700 5322 19712
rect 5445 19703 5503 19709
rect 5445 19700 5457 19703
rect 5316 19672 5457 19700
rect 5316 19660 5322 19672
rect 5445 19669 5457 19672
rect 5491 19669 5503 19703
rect 7742 19700 7748 19712
rect 7703 19672 7748 19700
rect 5445 19663 5503 19669
rect 7742 19660 7748 19672
rect 7800 19660 7806 19712
rect 8202 19660 8208 19712
rect 8260 19660 8266 19712
rect 11698 19700 11704 19712
rect 11659 19672 11704 19700
rect 11698 19660 11704 19672
rect 11756 19660 11762 19712
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 1762 19456 1768 19508
rect 1820 19496 1826 19508
rect 2133 19499 2191 19505
rect 2133 19496 2145 19499
rect 1820 19468 2145 19496
rect 1820 19456 1826 19468
rect 2133 19465 2145 19468
rect 2179 19465 2191 19499
rect 2590 19496 2596 19508
rect 2551 19468 2596 19496
rect 2133 19459 2191 19465
rect 2590 19456 2596 19468
rect 2648 19456 2654 19508
rect 4154 19456 4160 19508
rect 4212 19496 4218 19508
rect 9674 19496 9680 19508
rect 4212 19468 4476 19496
rect 4212 19456 4218 19468
rect 1578 19292 1584 19304
rect 1539 19264 1584 19292
rect 1578 19252 1584 19264
rect 1636 19252 1642 19304
rect 2317 19295 2375 19301
rect 2317 19261 2329 19295
rect 2363 19261 2375 19295
rect 2317 19255 2375 19261
rect 2777 19295 2835 19301
rect 2777 19261 2789 19295
rect 2823 19292 2835 19295
rect 3878 19292 3884 19304
rect 2823 19264 3884 19292
rect 2823 19261 2835 19264
rect 2777 19255 2835 19261
rect 1762 19224 1768 19236
rect 1723 19196 1768 19224
rect 1762 19184 1768 19196
rect 1820 19184 1826 19236
rect 2332 19224 2360 19255
rect 3878 19252 3884 19264
rect 3936 19252 3942 19304
rect 4448 19301 4476 19468
rect 7944 19468 9680 19496
rect 7944 19369 7972 19468
rect 9674 19456 9680 19468
rect 9732 19456 9738 19508
rect 19334 19456 19340 19508
rect 19392 19496 19398 19508
rect 20165 19499 20223 19505
rect 20165 19496 20177 19499
rect 19392 19468 20177 19496
rect 19392 19456 19398 19468
rect 20165 19465 20177 19468
rect 20211 19465 20223 19499
rect 20622 19496 20628 19508
rect 20583 19468 20628 19496
rect 20165 19459 20223 19465
rect 20622 19456 20628 19468
rect 20680 19456 20686 19508
rect 19429 19431 19487 19437
rect 19429 19397 19441 19431
rect 19475 19428 19487 19431
rect 20346 19428 20352 19440
rect 19475 19400 20352 19428
rect 19475 19397 19487 19400
rect 19429 19391 19487 19397
rect 20346 19388 20352 19400
rect 20404 19388 20410 19440
rect 7929 19363 7987 19369
rect 7929 19329 7941 19363
rect 7975 19329 7987 19363
rect 7929 19323 7987 19329
rect 4433 19295 4491 19301
rect 4080 19264 4384 19292
rect 4080 19224 4108 19264
rect 4246 19233 4252 19236
rect 2332 19196 4108 19224
rect 4188 19227 4252 19233
rect 4188 19193 4200 19227
rect 4234 19193 4252 19227
rect 4188 19187 4252 19193
rect 4246 19184 4252 19187
rect 4304 19184 4310 19236
rect 4356 19224 4384 19264
rect 4433 19261 4445 19295
rect 4479 19292 4491 19295
rect 4522 19292 4528 19304
rect 4479 19264 4528 19292
rect 4479 19261 4491 19264
rect 4433 19255 4491 19261
rect 4522 19252 4528 19264
rect 4580 19252 4586 19304
rect 5074 19292 5080 19304
rect 5035 19264 5080 19292
rect 5074 19252 5080 19264
rect 5132 19252 5138 19304
rect 7653 19295 7711 19301
rect 7653 19261 7665 19295
rect 7699 19292 7711 19295
rect 7742 19292 7748 19304
rect 7699 19264 7748 19292
rect 7699 19261 7711 19264
rect 7653 19255 7711 19261
rect 7742 19252 7748 19264
rect 7800 19252 7806 19304
rect 8297 19295 8355 19301
rect 8297 19261 8309 19295
rect 8343 19292 8355 19295
rect 9490 19292 9496 19304
rect 8343 19264 9496 19292
rect 8343 19261 8355 19264
rect 8297 19255 8355 19261
rect 9490 19252 9496 19264
rect 9548 19292 9554 19304
rect 10318 19292 10324 19304
rect 9548 19264 10324 19292
rect 9548 19252 9554 19264
rect 10318 19252 10324 19264
rect 10376 19252 10382 19304
rect 13265 19295 13323 19301
rect 13265 19261 13277 19295
rect 13311 19292 13323 19295
rect 13354 19292 13360 19304
rect 13311 19264 13360 19292
rect 13311 19261 13323 19264
rect 13265 19255 13323 19261
rect 13354 19252 13360 19264
rect 13412 19252 13418 19304
rect 19245 19295 19303 19301
rect 19245 19292 19257 19295
rect 18156 19264 19257 19292
rect 4709 19227 4767 19233
rect 4709 19224 4721 19227
rect 4356 19196 4721 19224
rect 4709 19193 4721 19196
rect 4755 19193 4767 19227
rect 5092 19224 5120 19252
rect 5092 19196 8156 19224
rect 4709 19187 4767 19193
rect 3053 19159 3111 19165
rect 3053 19125 3065 19159
rect 3099 19156 3111 19159
rect 4338 19156 4344 19168
rect 3099 19128 4344 19156
rect 3099 19125 3111 19128
rect 3053 19119 3111 19125
rect 4338 19116 4344 19128
rect 4396 19116 4402 19168
rect 4724 19156 4752 19187
rect 5810 19156 5816 19168
rect 4724 19128 5816 19156
rect 5810 19116 5816 19128
rect 5868 19116 5874 19168
rect 7282 19156 7288 19168
rect 7243 19128 7288 19156
rect 7282 19116 7288 19128
rect 7340 19116 7346 19168
rect 7466 19116 7472 19168
rect 7524 19156 7530 19168
rect 7745 19159 7803 19165
rect 7745 19156 7757 19159
rect 7524 19128 7757 19156
rect 7524 19116 7530 19128
rect 7745 19125 7757 19128
rect 7791 19125 7803 19159
rect 8128 19156 8156 19196
rect 8202 19184 8208 19236
rect 8260 19224 8266 19236
rect 8542 19227 8600 19233
rect 8542 19224 8554 19227
rect 8260 19196 8554 19224
rect 8260 19184 8266 19196
rect 8542 19193 8554 19196
rect 8588 19193 8600 19227
rect 8542 19187 8600 19193
rect 13446 19184 13452 19236
rect 13504 19233 13510 19236
rect 13504 19227 13568 19233
rect 13504 19193 13522 19227
rect 13556 19193 13568 19227
rect 13504 19187 13568 19193
rect 13504 19184 13510 19187
rect 10134 19156 10140 19168
rect 8128 19128 10140 19156
rect 7745 19119 7803 19125
rect 10134 19116 10140 19128
rect 10192 19116 10198 19168
rect 14550 19116 14556 19168
rect 14608 19156 14614 19168
rect 14645 19159 14703 19165
rect 14645 19156 14657 19159
rect 14608 19128 14657 19156
rect 14608 19116 14614 19128
rect 14645 19125 14657 19128
rect 14691 19125 14703 19159
rect 14645 19119 14703 19125
rect 18046 19116 18052 19168
rect 18104 19156 18110 19168
rect 18156 19165 18184 19264
rect 19245 19261 19257 19264
rect 19291 19261 19303 19295
rect 19889 19295 19947 19301
rect 19889 19292 19901 19295
rect 19245 19255 19303 19261
rect 19352 19264 19901 19292
rect 18598 19224 18604 19236
rect 18511 19196 18604 19224
rect 18598 19184 18604 19196
rect 18656 19224 18662 19236
rect 19352 19224 19380 19264
rect 19889 19261 19901 19264
rect 19935 19261 19947 19295
rect 19889 19255 19947 19261
rect 19978 19252 19984 19304
rect 20036 19292 20042 19304
rect 20349 19295 20407 19301
rect 20349 19292 20361 19295
rect 20036 19264 20361 19292
rect 20036 19252 20042 19264
rect 20349 19261 20361 19264
rect 20395 19261 20407 19295
rect 20349 19255 20407 19261
rect 20809 19295 20867 19301
rect 20809 19261 20821 19295
rect 20855 19292 20867 19295
rect 20901 19295 20959 19301
rect 20901 19292 20913 19295
rect 20855 19264 20913 19292
rect 20855 19261 20867 19264
rect 20809 19255 20867 19261
rect 20901 19261 20913 19264
rect 20947 19261 20959 19295
rect 20901 19255 20959 19261
rect 18656 19196 19380 19224
rect 19536 19196 20392 19224
rect 18656 19184 18662 19196
rect 18141 19159 18199 19165
rect 18141 19156 18153 19159
rect 18104 19128 18153 19156
rect 18104 19116 18110 19128
rect 18141 19125 18153 19128
rect 18187 19125 18199 19159
rect 18141 19119 18199 19125
rect 18969 19159 19027 19165
rect 18969 19125 18981 19159
rect 19015 19156 19027 19159
rect 19334 19156 19340 19168
rect 19015 19128 19340 19156
rect 19015 19125 19027 19128
rect 18969 19119 19027 19125
rect 19334 19116 19340 19128
rect 19392 19156 19398 19168
rect 19536 19156 19564 19196
rect 19702 19156 19708 19168
rect 19392 19128 19564 19156
rect 19663 19128 19708 19156
rect 19392 19116 19398 19128
rect 19702 19116 19708 19128
rect 19760 19116 19766 19168
rect 20364 19156 20392 19196
rect 20438 19184 20444 19236
rect 20496 19224 20502 19236
rect 21177 19227 21235 19233
rect 21177 19224 21189 19227
rect 20496 19196 21189 19224
rect 20496 19184 20502 19196
rect 21177 19193 21189 19196
rect 21223 19193 21235 19227
rect 21358 19224 21364 19236
rect 21319 19196 21364 19224
rect 21177 19187 21235 19193
rect 21358 19184 21364 19196
rect 21416 19184 21422 19236
rect 20901 19159 20959 19165
rect 20901 19156 20913 19159
rect 20364 19128 20913 19156
rect 20901 19125 20913 19128
rect 20947 19125 20959 19159
rect 20901 19119 20959 19125
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 1762 18912 1768 18964
rect 1820 18952 1826 18964
rect 2133 18955 2191 18961
rect 2133 18952 2145 18955
rect 1820 18924 2145 18952
rect 1820 18912 1826 18924
rect 2133 18921 2145 18924
rect 2179 18921 2191 18955
rect 2133 18915 2191 18921
rect 2593 18955 2651 18961
rect 2593 18921 2605 18955
rect 2639 18952 2651 18955
rect 2866 18952 2872 18964
rect 2639 18924 2872 18952
rect 2639 18921 2651 18924
rect 2593 18915 2651 18921
rect 2866 18912 2872 18924
rect 2924 18912 2930 18964
rect 3050 18952 3056 18964
rect 3011 18924 3056 18952
rect 3050 18912 3056 18924
rect 3108 18912 3114 18964
rect 4709 18955 4767 18961
rect 4709 18952 4721 18955
rect 3160 18924 4721 18952
rect 1578 18816 1584 18828
rect 1539 18788 1584 18816
rect 1578 18776 1584 18788
rect 1636 18776 1642 18828
rect 1762 18816 1768 18828
rect 1723 18788 1768 18816
rect 1762 18776 1768 18788
rect 1820 18776 1826 18828
rect 2317 18819 2375 18825
rect 2317 18785 2329 18819
rect 2363 18785 2375 18819
rect 2317 18779 2375 18785
rect 2777 18819 2835 18825
rect 2777 18785 2789 18819
rect 2823 18816 2835 18819
rect 3160 18816 3188 18924
rect 4709 18921 4721 18924
rect 4755 18952 4767 18955
rect 6546 18952 6552 18964
rect 4755 18924 6552 18952
rect 4755 18921 4767 18924
rect 4709 18915 4767 18921
rect 6546 18912 6552 18924
rect 6604 18912 6610 18964
rect 19245 18955 19303 18961
rect 19245 18921 19257 18955
rect 19291 18952 19303 18955
rect 19978 18952 19984 18964
rect 19291 18924 19984 18952
rect 19291 18921 19303 18924
rect 19245 18915 19303 18921
rect 19978 18912 19984 18924
rect 20036 18912 20042 18964
rect 20254 18912 20260 18964
rect 20312 18952 20318 18964
rect 20349 18955 20407 18961
rect 20349 18952 20361 18955
rect 20312 18924 20361 18952
rect 20312 18912 20318 18924
rect 20349 18921 20361 18924
rect 20395 18921 20407 18955
rect 20349 18915 20407 18921
rect 20809 18955 20867 18961
rect 20809 18921 20821 18955
rect 20855 18952 20867 18955
rect 21174 18952 21180 18964
rect 20855 18924 21180 18952
rect 20855 18921 20867 18924
rect 20809 18915 20867 18921
rect 21174 18912 21180 18924
rect 21232 18912 21238 18964
rect 7282 18884 7288 18896
rect 3252 18856 7288 18884
rect 3252 18825 3280 18856
rect 7282 18844 7288 18856
rect 7340 18844 7346 18896
rect 11698 18844 11704 18896
rect 11756 18884 11762 18896
rect 12222 18887 12280 18893
rect 12222 18884 12234 18887
rect 11756 18856 12234 18884
rect 11756 18844 11762 18856
rect 12222 18853 12234 18856
rect 12268 18884 12280 18887
rect 13998 18884 14004 18896
rect 12268 18856 14004 18884
rect 12268 18853 12280 18856
rect 12222 18847 12280 18853
rect 13998 18844 14004 18856
rect 14056 18844 14062 18896
rect 2823 18788 3188 18816
rect 3237 18819 3295 18825
rect 2823 18785 2835 18788
rect 2777 18779 2835 18785
rect 3237 18785 3249 18819
rect 3283 18785 3295 18819
rect 3237 18779 3295 18785
rect 2332 18748 2360 18779
rect 4154 18776 4160 18828
rect 4212 18816 4218 18828
rect 4341 18819 4399 18825
rect 4341 18816 4353 18819
rect 4212 18788 4353 18816
rect 4212 18776 4218 18788
rect 4341 18785 4353 18788
rect 4387 18816 4399 18819
rect 5074 18816 5080 18828
rect 4387 18788 5080 18816
rect 4387 18785 4399 18788
rect 4341 18779 4399 18785
rect 5074 18776 5080 18788
rect 5132 18776 5138 18828
rect 5258 18825 5264 18828
rect 5252 18816 5264 18825
rect 5219 18788 5264 18816
rect 5252 18779 5264 18788
rect 5258 18776 5264 18779
rect 5316 18776 5322 18828
rect 7552 18819 7610 18825
rect 7552 18785 7564 18819
rect 7598 18816 7610 18819
rect 9030 18816 9036 18828
rect 7598 18788 9036 18816
rect 7598 18785 7610 18788
rect 7552 18779 7610 18785
rect 9030 18776 9036 18788
rect 9088 18776 9094 18828
rect 11977 18819 12035 18825
rect 11977 18785 11989 18819
rect 12023 18816 12035 18819
rect 12618 18816 12624 18828
rect 12023 18788 12624 18816
rect 12023 18785 12035 18788
rect 11977 18779 12035 18785
rect 12618 18776 12624 18788
rect 12676 18816 12682 18828
rect 12676 18788 13400 18816
rect 12676 18776 12682 18788
rect 13372 18760 13400 18788
rect 14550 18776 14556 18828
rect 14608 18816 14614 18828
rect 14901 18819 14959 18825
rect 14901 18816 14913 18819
rect 14608 18788 14913 18816
rect 14608 18776 14614 18788
rect 14901 18785 14913 18788
rect 14947 18785 14959 18819
rect 14901 18779 14959 18785
rect 19061 18819 19119 18825
rect 19061 18785 19073 18819
rect 19107 18785 19119 18819
rect 19061 18779 19119 18785
rect 19705 18819 19763 18825
rect 19705 18785 19717 18819
rect 19751 18816 19763 18819
rect 20165 18819 20223 18825
rect 20165 18816 20177 18819
rect 19751 18788 20177 18816
rect 19751 18785 19763 18788
rect 19705 18779 19763 18785
rect 20165 18785 20177 18788
rect 20211 18785 20223 18819
rect 20165 18779 20223 18785
rect 20625 18819 20683 18825
rect 20625 18785 20637 18819
rect 20671 18785 20683 18819
rect 21174 18816 21180 18828
rect 21135 18788 21180 18816
rect 20625 18779 20683 18785
rect 2332 18720 2774 18748
rect 2746 18612 2774 18720
rect 4522 18708 4528 18760
rect 4580 18748 4586 18760
rect 4985 18751 5043 18757
rect 4985 18748 4997 18751
rect 4580 18720 4997 18748
rect 4580 18708 4586 18720
rect 4985 18717 4997 18720
rect 5031 18717 5043 18751
rect 7285 18751 7343 18757
rect 7285 18748 7297 18751
rect 4985 18711 5043 18717
rect 6012 18720 7297 18748
rect 3970 18612 3976 18624
rect 2746 18584 3976 18612
rect 3970 18572 3976 18584
rect 4028 18572 4034 18624
rect 5000 18612 5028 18711
rect 5350 18612 5356 18624
rect 5000 18584 5356 18612
rect 5350 18572 5356 18584
rect 5408 18612 5414 18624
rect 6012 18612 6040 18720
rect 7285 18717 7297 18720
rect 7331 18717 7343 18751
rect 7285 18711 7343 18717
rect 13354 18708 13360 18760
rect 13412 18748 13418 18760
rect 14645 18751 14703 18757
rect 14645 18748 14657 18751
rect 13412 18720 14657 18748
rect 13412 18708 13418 18720
rect 14645 18717 14657 18720
rect 14691 18717 14703 18751
rect 19076 18748 19104 18779
rect 20530 18748 20536 18760
rect 19076 18720 20536 18748
rect 14645 18711 14703 18717
rect 20530 18708 20536 18720
rect 20588 18708 20594 18760
rect 20640 18680 20668 18779
rect 21174 18776 21180 18788
rect 21232 18776 21238 18828
rect 21358 18680 21364 18692
rect 19812 18652 20668 18680
rect 21319 18652 21364 18680
rect 19812 18624 19840 18652
rect 21358 18640 21364 18652
rect 21416 18640 21422 18692
rect 5408 18584 6040 18612
rect 6365 18615 6423 18621
rect 5408 18572 5414 18584
rect 6365 18581 6377 18615
rect 6411 18612 6423 18615
rect 7558 18612 7564 18624
rect 6411 18584 7564 18612
rect 6411 18581 6423 18584
rect 6365 18575 6423 18581
rect 7558 18572 7564 18584
rect 7616 18572 7622 18624
rect 8202 18572 8208 18624
rect 8260 18612 8266 18624
rect 8665 18615 8723 18621
rect 8665 18612 8677 18615
rect 8260 18584 8677 18612
rect 8260 18572 8266 18584
rect 8665 18581 8677 18584
rect 8711 18581 8723 18615
rect 13354 18612 13360 18624
rect 13315 18584 13360 18612
rect 8665 18575 8723 18581
rect 13354 18572 13360 18584
rect 13412 18572 13418 18624
rect 15930 18572 15936 18624
rect 15988 18612 15994 18624
rect 16025 18615 16083 18621
rect 16025 18612 16037 18615
rect 15988 18584 16037 18612
rect 15988 18572 15994 18584
rect 16025 18581 16037 18584
rect 16071 18581 16083 18615
rect 18690 18612 18696 18624
rect 18651 18584 18696 18612
rect 16025 18575 16083 18581
rect 18690 18572 18696 18584
rect 18748 18612 18754 18624
rect 19705 18615 19763 18621
rect 19705 18612 19717 18615
rect 18748 18584 19717 18612
rect 18748 18572 18754 18584
rect 19705 18581 19717 18584
rect 19751 18581 19763 18615
rect 19705 18575 19763 18581
rect 19794 18572 19800 18624
rect 19852 18612 19858 18624
rect 19852 18584 19897 18612
rect 19852 18572 19858 18584
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 2222 18408 2228 18420
rect 2183 18380 2228 18408
rect 2222 18368 2228 18380
rect 2280 18368 2286 18420
rect 3970 18368 3976 18420
rect 4028 18408 4034 18420
rect 7466 18408 7472 18420
rect 4028 18380 5028 18408
rect 7427 18380 7472 18408
rect 4028 18368 4034 18380
rect 1762 18300 1768 18352
rect 1820 18340 1826 18352
rect 2685 18343 2743 18349
rect 2685 18340 2697 18343
rect 1820 18312 2697 18340
rect 1820 18300 1826 18312
rect 2685 18309 2697 18312
rect 2731 18309 2743 18343
rect 4338 18340 4344 18352
rect 2685 18303 2743 18309
rect 3344 18312 4344 18340
rect 3344 18281 3372 18312
rect 4338 18300 4344 18312
rect 4396 18340 4402 18352
rect 4890 18340 4896 18352
rect 4396 18312 4896 18340
rect 4396 18300 4402 18312
rect 4890 18300 4896 18312
rect 4948 18300 4954 18352
rect 5000 18340 5028 18380
rect 7466 18368 7472 18380
rect 7524 18368 7530 18420
rect 10870 18368 10876 18420
rect 10928 18408 10934 18420
rect 17129 18411 17187 18417
rect 17129 18408 17141 18411
rect 10928 18380 17141 18408
rect 10928 18368 10934 18380
rect 17129 18377 17141 18380
rect 17175 18377 17187 18411
rect 17129 18371 17187 18377
rect 20349 18411 20407 18417
rect 20349 18377 20361 18411
rect 20395 18408 20407 18411
rect 20438 18408 20444 18420
rect 20395 18380 20444 18408
rect 20395 18377 20407 18380
rect 20349 18371 20407 18377
rect 20438 18368 20444 18380
rect 20496 18368 20502 18420
rect 20809 18411 20867 18417
rect 20809 18377 20821 18411
rect 20855 18408 20867 18411
rect 21174 18408 21180 18420
rect 20855 18380 21180 18408
rect 20855 18377 20867 18380
rect 20809 18371 20867 18377
rect 21174 18368 21180 18380
rect 21232 18368 21238 18420
rect 10686 18340 10692 18352
rect 5000 18312 10692 18340
rect 10686 18300 10692 18312
rect 10744 18300 10750 18352
rect 12621 18343 12679 18349
rect 12621 18309 12633 18343
rect 12667 18340 12679 18343
rect 18874 18340 18880 18352
rect 12667 18312 18880 18340
rect 12667 18309 12679 18312
rect 12621 18303 12679 18309
rect 18874 18300 18880 18312
rect 18932 18300 18938 18352
rect 3329 18275 3387 18281
rect 3329 18241 3341 18275
rect 3375 18241 3387 18275
rect 3329 18235 3387 18241
rect 4801 18275 4859 18281
rect 4801 18241 4813 18275
rect 4847 18272 4859 18275
rect 5258 18272 5264 18284
rect 4847 18244 5264 18272
rect 4847 18241 4859 18244
rect 4801 18235 4859 18241
rect 5258 18232 5264 18244
rect 5316 18232 5322 18284
rect 8113 18275 8171 18281
rect 8113 18241 8125 18275
rect 8159 18272 8171 18275
rect 8202 18272 8208 18284
rect 8159 18244 8208 18272
rect 8159 18241 8171 18244
rect 8113 18235 8171 18241
rect 8202 18232 8208 18244
rect 8260 18232 8266 18284
rect 9030 18272 9036 18284
rect 8991 18244 9036 18272
rect 9030 18232 9036 18244
rect 9088 18272 9094 18284
rect 9582 18272 9588 18284
rect 9088 18244 9588 18272
rect 9088 18232 9094 18244
rect 9582 18232 9588 18244
rect 9640 18232 9646 18284
rect 12069 18275 12127 18281
rect 12069 18241 12081 18275
rect 12115 18272 12127 18275
rect 12342 18272 12348 18284
rect 12115 18244 12348 18272
rect 12115 18241 12127 18244
rect 12069 18235 12127 18241
rect 12342 18232 12348 18244
rect 12400 18232 12406 18284
rect 14550 18272 14556 18284
rect 14511 18244 14556 18272
rect 14550 18232 14556 18244
rect 14608 18232 14614 18284
rect 17678 18272 17684 18284
rect 17639 18244 17684 18272
rect 17678 18232 17684 18244
rect 17736 18232 17742 18284
rect 19337 18275 19395 18281
rect 19337 18241 19349 18275
rect 19383 18272 19395 18275
rect 19383 18244 20484 18272
rect 19383 18241 19395 18244
rect 19337 18235 19395 18241
rect 20456 18216 20484 18244
rect 2869 18207 2927 18213
rect 2869 18173 2881 18207
rect 2915 18204 2927 18207
rect 6822 18204 6828 18216
rect 2915 18176 6828 18204
rect 2915 18173 2927 18176
rect 2869 18167 2927 18173
rect 6822 18164 6828 18176
rect 6880 18164 6886 18216
rect 19426 18164 19432 18216
rect 19484 18204 19490 18216
rect 19705 18207 19763 18213
rect 19705 18204 19717 18207
rect 19484 18176 19717 18204
rect 19484 18164 19490 18176
rect 19705 18173 19717 18176
rect 19751 18173 19763 18207
rect 20165 18207 20223 18213
rect 20165 18204 20177 18207
rect 19705 18167 19763 18173
rect 19904 18176 20177 18204
rect 1762 18136 1768 18148
rect 1723 18108 1768 18136
rect 1762 18096 1768 18108
rect 1820 18096 1826 18148
rect 2314 18136 2320 18148
rect 2275 18108 2320 18136
rect 2314 18096 2320 18108
rect 2372 18096 2378 18148
rect 3418 18136 3424 18148
rect 3379 18108 3424 18136
rect 3418 18096 3424 18108
rect 3476 18096 3482 18148
rect 4525 18139 4583 18145
rect 4525 18136 4537 18139
rect 3896 18108 4537 18136
rect 1670 18068 1676 18080
rect 1631 18040 1676 18068
rect 1670 18028 1676 18040
rect 1728 18028 1734 18080
rect 3510 18068 3516 18080
rect 3471 18040 3516 18068
rect 3510 18028 3516 18040
rect 3568 18028 3574 18080
rect 3896 18077 3924 18108
rect 4525 18105 4537 18108
rect 4571 18105 4583 18139
rect 4525 18099 4583 18105
rect 7837 18139 7895 18145
rect 7837 18105 7849 18139
rect 7883 18136 7895 18139
rect 9122 18136 9128 18148
rect 7883 18108 9128 18136
rect 7883 18105 7895 18108
rect 7837 18099 7895 18105
rect 9122 18096 9128 18108
rect 9180 18096 9186 18148
rect 11974 18096 11980 18148
rect 12032 18136 12038 18148
rect 12253 18139 12311 18145
rect 12253 18136 12265 18139
rect 12032 18108 12265 18136
rect 12032 18096 12038 18108
rect 12253 18105 12265 18108
rect 12299 18105 12311 18139
rect 17494 18136 17500 18148
rect 17407 18108 17500 18136
rect 12253 18099 12311 18105
rect 17494 18096 17500 18108
rect 17552 18136 17558 18148
rect 18141 18139 18199 18145
rect 18141 18136 18153 18139
rect 17552 18108 18153 18136
rect 17552 18096 17558 18108
rect 18141 18105 18153 18108
rect 18187 18105 18199 18139
rect 18141 18099 18199 18105
rect 3881 18071 3939 18077
rect 3881 18037 3893 18071
rect 3927 18037 3939 18071
rect 4154 18068 4160 18080
rect 4115 18040 4160 18068
rect 3881 18031 3939 18037
rect 4154 18028 4160 18040
rect 4212 18028 4218 18080
rect 4614 18068 4620 18080
rect 4575 18040 4620 18068
rect 4614 18028 4620 18040
rect 4672 18028 4678 18080
rect 5166 18068 5172 18080
rect 5127 18040 5172 18068
rect 5166 18028 5172 18040
rect 5224 18028 5230 18080
rect 7929 18071 7987 18077
rect 7929 18037 7941 18071
rect 7975 18068 7987 18071
rect 8481 18071 8539 18077
rect 8481 18068 8493 18071
rect 7975 18040 8493 18068
rect 7975 18037 7987 18040
rect 7929 18031 7987 18037
rect 8481 18037 8493 18040
rect 8527 18037 8539 18071
rect 8846 18068 8852 18080
rect 8807 18040 8852 18068
rect 8481 18031 8539 18037
rect 8846 18028 8852 18040
rect 8904 18028 8910 18080
rect 8938 18028 8944 18080
rect 8996 18068 9002 18080
rect 9398 18068 9404 18080
rect 8996 18040 9404 18068
rect 8996 18028 9002 18040
rect 9398 18028 9404 18040
rect 9456 18068 9462 18080
rect 9493 18071 9551 18077
rect 9493 18068 9505 18071
rect 9456 18040 9505 18068
rect 9456 18028 9462 18040
rect 9493 18037 9505 18040
rect 9539 18037 9551 18071
rect 9493 18031 9551 18037
rect 11698 18028 11704 18080
rect 11756 18068 11762 18080
rect 12161 18071 12219 18077
rect 12161 18068 12173 18071
rect 11756 18040 12173 18068
rect 11756 18028 11762 18040
rect 12161 18037 12173 18040
rect 12207 18037 12219 18071
rect 14642 18068 14648 18080
rect 14603 18040 14648 18068
rect 12161 18031 12219 18037
rect 14642 18028 14648 18040
rect 14700 18028 14706 18080
rect 14734 18028 14740 18080
rect 14792 18068 14798 18080
rect 15105 18071 15163 18077
rect 14792 18040 14837 18068
rect 14792 18028 14798 18040
rect 15105 18037 15117 18071
rect 15151 18068 15163 18071
rect 15194 18068 15200 18080
rect 15151 18040 15200 18068
rect 15151 18037 15163 18040
rect 15105 18031 15163 18037
rect 15194 18028 15200 18040
rect 15252 18028 15258 18080
rect 15378 18068 15384 18080
rect 15339 18040 15384 18068
rect 15378 18028 15384 18040
rect 15436 18028 15442 18080
rect 17586 18028 17592 18080
rect 17644 18068 17650 18080
rect 18966 18068 18972 18080
rect 17644 18040 17689 18068
rect 18927 18040 18972 18068
rect 17644 18028 17650 18040
rect 18966 18028 18972 18040
rect 19024 18028 19030 18080
rect 19904 18077 19932 18176
rect 20165 18173 20177 18176
rect 20211 18173 20223 18207
rect 20165 18167 20223 18173
rect 20438 18164 20444 18216
rect 20496 18204 20502 18216
rect 20625 18207 20683 18213
rect 20625 18204 20637 18207
rect 20496 18176 20637 18204
rect 20496 18164 20502 18176
rect 20625 18173 20637 18176
rect 20671 18173 20683 18207
rect 20625 18167 20683 18173
rect 20254 18096 20260 18148
rect 20312 18136 20318 18148
rect 21177 18139 21235 18145
rect 21177 18136 21189 18139
rect 20312 18108 21189 18136
rect 20312 18096 20318 18108
rect 21177 18105 21189 18108
rect 21223 18105 21235 18139
rect 21358 18136 21364 18148
rect 21319 18108 21364 18136
rect 21177 18099 21235 18105
rect 21358 18096 21364 18108
rect 21416 18096 21422 18148
rect 19889 18071 19947 18077
rect 19889 18037 19901 18071
rect 19935 18037 19947 18071
rect 19889 18031 19947 18037
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 2133 17867 2191 17873
rect 2133 17833 2145 17867
rect 2179 17864 2191 17867
rect 2314 17864 2320 17876
rect 2179 17836 2320 17864
rect 2179 17833 2191 17836
rect 2133 17827 2191 17833
rect 2314 17824 2320 17836
rect 2372 17824 2378 17876
rect 3510 17864 3516 17876
rect 3471 17836 3516 17864
rect 3510 17824 3516 17836
rect 3568 17824 3574 17876
rect 4341 17867 4399 17873
rect 4341 17833 4353 17867
rect 4387 17864 4399 17867
rect 4614 17864 4620 17876
rect 4387 17836 4620 17864
rect 4387 17833 4399 17836
rect 4341 17827 4399 17833
rect 4614 17824 4620 17836
rect 4672 17824 4678 17876
rect 6822 17824 6828 17876
rect 6880 17864 6886 17876
rect 7837 17867 7895 17873
rect 7837 17864 7849 17867
rect 6880 17836 7849 17864
rect 6880 17824 6886 17836
rect 7837 17833 7849 17836
rect 7883 17833 7895 17867
rect 7837 17827 7895 17833
rect 9398 17824 9404 17876
rect 9456 17864 9462 17876
rect 10318 17864 10324 17876
rect 9456 17836 10324 17864
rect 9456 17824 9462 17836
rect 10318 17824 10324 17836
rect 10376 17824 10382 17876
rect 10594 17824 10600 17876
rect 10652 17864 10658 17876
rect 12897 17867 12955 17873
rect 12897 17864 12909 17867
rect 10652 17836 12909 17864
rect 10652 17824 10658 17836
rect 12897 17833 12909 17836
rect 12943 17864 12955 17867
rect 13541 17867 13599 17873
rect 13541 17864 13553 17867
rect 12943 17836 13553 17864
rect 12943 17833 12955 17836
rect 12897 17827 12955 17833
rect 13541 17833 13553 17836
rect 13587 17833 13599 17867
rect 13541 17827 13599 17833
rect 14734 17824 14740 17876
rect 14792 17864 14798 17876
rect 14829 17867 14887 17873
rect 14829 17864 14841 17867
rect 14792 17836 14841 17864
rect 14792 17824 14798 17836
rect 14829 17833 14841 17836
rect 14875 17833 14887 17867
rect 14829 17827 14887 17833
rect 15197 17867 15255 17873
rect 15197 17833 15209 17867
rect 15243 17864 15255 17867
rect 15378 17864 15384 17876
rect 15243 17836 15384 17864
rect 15243 17833 15255 17836
rect 15197 17827 15255 17833
rect 15378 17824 15384 17836
rect 15436 17824 15442 17876
rect 16577 17867 16635 17873
rect 16577 17833 16589 17867
rect 16623 17833 16635 17867
rect 16577 17827 16635 17833
rect 17221 17867 17279 17873
rect 17221 17833 17233 17867
rect 17267 17864 17279 17867
rect 17405 17867 17463 17873
rect 17405 17864 17417 17867
rect 17267 17836 17417 17864
rect 17267 17833 17279 17836
rect 17221 17827 17279 17833
rect 17405 17833 17417 17836
rect 17451 17864 17463 17867
rect 17678 17864 17684 17876
rect 17451 17836 17684 17864
rect 17451 17833 17463 17836
rect 17405 17827 17463 17833
rect 3053 17799 3111 17805
rect 3053 17765 3065 17799
rect 3099 17796 3111 17799
rect 5166 17796 5172 17808
rect 3099 17768 5172 17796
rect 3099 17765 3111 17768
rect 3053 17759 3111 17765
rect 4356 17740 4384 17768
rect 5166 17756 5172 17768
rect 5224 17756 5230 17808
rect 5896 17799 5954 17805
rect 5896 17765 5908 17799
rect 5942 17796 5954 17799
rect 5994 17796 6000 17808
rect 5942 17768 6000 17796
rect 5942 17765 5954 17768
rect 5896 17759 5954 17765
rect 5994 17756 6000 17768
rect 6052 17756 6058 17808
rect 6546 17756 6552 17808
rect 6604 17796 6610 17808
rect 11054 17796 11060 17808
rect 6604 17768 11060 17796
rect 6604 17756 6610 17768
rect 11054 17756 11060 17768
rect 11112 17756 11118 17808
rect 15470 17796 15476 17808
rect 13372 17768 15476 17796
rect 1765 17731 1823 17737
rect 1765 17697 1777 17731
rect 1811 17697 1823 17731
rect 1765 17691 1823 17697
rect 2317 17731 2375 17737
rect 2317 17697 2329 17731
rect 2363 17728 2375 17731
rect 3145 17731 3203 17737
rect 2363 17700 2774 17728
rect 2363 17697 2375 17700
rect 2317 17691 2375 17697
rect 1780 17660 1808 17691
rect 2590 17660 2596 17672
rect 1780 17632 2596 17660
rect 2590 17620 2596 17632
rect 2648 17620 2654 17672
rect 1670 17524 1676 17536
rect 1631 17496 1676 17524
rect 1670 17484 1676 17496
rect 1728 17484 1734 17536
rect 2746 17524 2774 17700
rect 3145 17697 3157 17731
rect 3191 17728 3203 17731
rect 4062 17728 4068 17740
rect 3191 17700 4068 17728
rect 3191 17697 3203 17700
rect 3145 17691 3203 17697
rect 4062 17688 4068 17700
rect 4120 17688 4126 17740
rect 4338 17688 4344 17740
rect 4396 17688 4402 17740
rect 4709 17731 4767 17737
rect 4709 17697 4721 17731
rect 4755 17728 4767 17731
rect 6914 17728 6920 17740
rect 4755 17700 6920 17728
rect 4755 17697 4767 17700
rect 4709 17691 4767 17697
rect 6914 17688 6920 17700
rect 6972 17688 6978 17740
rect 8021 17731 8079 17737
rect 8021 17697 8033 17731
rect 8067 17728 8079 17731
rect 8294 17728 8300 17740
rect 8067 17700 8300 17728
rect 8067 17697 8079 17700
rect 8021 17691 8079 17697
rect 8294 17688 8300 17700
rect 8352 17688 8358 17740
rect 9398 17688 9404 17740
rect 9456 17728 9462 17740
rect 11238 17737 11244 17740
rect 9565 17731 9623 17737
rect 9565 17728 9577 17731
rect 9456 17700 9577 17728
rect 9456 17688 9462 17700
rect 9565 17697 9577 17700
rect 9611 17697 9623 17731
rect 11232 17728 11244 17737
rect 11199 17700 11244 17728
rect 9565 17691 9623 17697
rect 11232 17691 11244 17700
rect 11238 17688 11244 17691
rect 11296 17688 11302 17740
rect 13372 17672 13400 17768
rect 15470 17756 15476 17768
rect 15528 17756 15534 17808
rect 15562 17756 15568 17808
rect 15620 17796 15626 17808
rect 16592 17796 16620 17827
rect 17678 17824 17684 17836
rect 17736 17824 17742 17876
rect 19245 17867 19303 17873
rect 19245 17833 19257 17867
rect 19291 17864 19303 17867
rect 19978 17864 19984 17876
rect 19291 17836 19984 17864
rect 19291 17833 19303 17836
rect 19245 17827 19303 17833
rect 19978 17824 19984 17836
rect 20036 17824 20042 17876
rect 20254 17864 20260 17876
rect 20215 17836 20260 17864
rect 20254 17824 20260 17836
rect 20312 17824 20318 17876
rect 15620 17768 16344 17796
rect 16592 17768 19104 17796
rect 15620 17756 15626 17768
rect 13722 17688 13728 17740
rect 13780 17728 13786 17740
rect 15102 17728 15108 17740
rect 13780 17700 15108 17728
rect 13780 17688 13786 17700
rect 15102 17688 15108 17700
rect 15160 17688 15166 17740
rect 15194 17688 15200 17740
rect 15252 17728 15258 17740
rect 16209 17731 16267 17737
rect 16209 17728 16221 17731
rect 15252 17700 16221 17728
rect 15252 17688 15258 17700
rect 16209 17697 16221 17700
rect 16255 17697 16267 17731
rect 16316 17728 16344 17768
rect 16482 17728 16488 17740
rect 16316 17700 16488 17728
rect 16209 17691 16267 17697
rect 16482 17688 16488 17700
rect 16540 17728 16546 17740
rect 17954 17728 17960 17740
rect 16540 17700 17960 17728
rect 16540 17688 16546 17700
rect 17954 17688 17960 17700
rect 18012 17688 18018 17740
rect 18138 17688 18144 17740
rect 18196 17728 18202 17740
rect 19076 17737 19104 17768
rect 18518 17731 18576 17737
rect 18518 17728 18530 17731
rect 18196 17700 18530 17728
rect 18196 17688 18202 17700
rect 18518 17697 18530 17700
rect 18564 17697 18576 17731
rect 18518 17691 18576 17697
rect 19061 17731 19119 17737
rect 19061 17697 19073 17731
rect 19107 17697 19119 17731
rect 19061 17691 19119 17697
rect 20073 17731 20131 17737
rect 20073 17697 20085 17731
rect 20119 17697 20131 17731
rect 20073 17691 20131 17697
rect 2958 17660 2964 17672
rect 2919 17632 2964 17660
rect 2958 17620 2964 17632
rect 3016 17620 3022 17672
rect 4798 17660 4804 17672
rect 4759 17632 4804 17660
rect 4798 17620 4804 17632
rect 4856 17620 4862 17672
rect 4890 17620 4896 17672
rect 4948 17660 4954 17672
rect 4948 17632 4993 17660
rect 4948 17620 4954 17632
rect 5350 17620 5356 17672
rect 5408 17660 5414 17672
rect 5629 17663 5687 17669
rect 5629 17660 5641 17663
rect 5408 17632 5641 17660
rect 5408 17620 5414 17632
rect 5629 17629 5641 17632
rect 5675 17629 5687 17663
rect 5629 17623 5687 17629
rect 9309 17663 9367 17669
rect 9309 17629 9321 17663
rect 9355 17629 9367 17663
rect 9309 17623 9367 17629
rect 10965 17663 11023 17669
rect 10965 17629 10977 17663
rect 11011 17629 11023 17663
rect 10965 17623 11023 17629
rect 8938 17592 8944 17604
rect 6886 17564 8944 17592
rect 3973 17527 4031 17533
rect 3973 17524 3985 17527
rect 2746 17496 3985 17524
rect 3973 17493 3985 17496
rect 4019 17524 4031 17527
rect 6886 17524 6914 17564
rect 8938 17552 8944 17564
rect 8996 17552 9002 17604
rect 7006 17524 7012 17536
rect 4019 17496 6914 17524
rect 6967 17496 7012 17524
rect 4019 17493 4031 17496
rect 3973 17487 4031 17493
rect 7006 17484 7012 17496
rect 7064 17484 7070 17536
rect 8389 17527 8447 17533
rect 8389 17493 8401 17527
rect 8435 17524 8447 17527
rect 8846 17524 8852 17536
rect 8435 17496 8852 17524
rect 8435 17493 8447 17496
rect 8389 17487 8447 17493
rect 8846 17484 8852 17496
rect 8904 17484 8910 17536
rect 9324 17524 9352 17623
rect 10980 17592 11008 17623
rect 12066 17620 12072 17672
rect 12124 17660 12130 17672
rect 13354 17660 13360 17672
rect 12124 17632 13216 17660
rect 13267 17632 13360 17660
rect 12124 17620 12130 17632
rect 10336 17564 11008 17592
rect 13188 17592 13216 17632
rect 13354 17620 13360 17632
rect 13412 17620 13418 17672
rect 13449 17663 13507 17669
rect 13449 17629 13461 17663
rect 13495 17660 13507 17663
rect 13538 17660 13544 17672
rect 13495 17632 13544 17660
rect 13495 17629 13507 17632
rect 13449 17623 13507 17629
rect 13538 17620 13544 17632
rect 13596 17620 13602 17672
rect 14737 17663 14795 17669
rect 14737 17629 14749 17663
rect 14783 17660 14795 17663
rect 15289 17663 15347 17669
rect 15289 17660 15301 17663
rect 14783 17632 15301 17660
rect 14783 17629 14795 17632
rect 14737 17623 14795 17629
rect 15289 17629 15301 17632
rect 15335 17629 15347 17663
rect 15470 17660 15476 17672
rect 15431 17632 15476 17660
rect 15289 17623 15347 17629
rect 15470 17620 15476 17632
rect 15528 17620 15534 17672
rect 15930 17660 15936 17672
rect 15891 17632 15936 17660
rect 15930 17620 15936 17632
rect 15988 17620 15994 17672
rect 16114 17660 16120 17672
rect 16075 17632 16120 17660
rect 16114 17620 16120 17632
rect 16172 17620 16178 17672
rect 18782 17660 18788 17672
rect 18743 17632 18788 17660
rect 18782 17620 18788 17632
rect 18840 17620 18846 17672
rect 18966 17620 18972 17672
rect 19024 17660 19030 17672
rect 20088 17660 20116 17691
rect 20346 17688 20352 17740
rect 20404 17728 20410 17740
rect 20625 17731 20683 17737
rect 20625 17728 20637 17731
rect 20404 17700 20637 17728
rect 20404 17688 20410 17700
rect 20625 17697 20637 17700
rect 20671 17697 20683 17731
rect 21174 17728 21180 17740
rect 21135 17700 21180 17728
rect 20625 17691 20683 17697
rect 21174 17688 21180 17700
rect 21232 17688 21238 17740
rect 19024 17632 20116 17660
rect 19024 17620 19030 17632
rect 17221 17595 17279 17601
rect 17221 17592 17233 17595
rect 13188 17564 17233 17592
rect 9490 17524 9496 17536
rect 9324 17496 9496 17524
rect 9490 17484 9496 17496
rect 9548 17524 9554 17536
rect 10336 17524 10364 17564
rect 17221 17561 17233 17564
rect 17267 17561 17279 17595
rect 19794 17592 19800 17604
rect 17221 17555 17279 17561
rect 19168 17564 19800 17592
rect 9548 17496 10364 17524
rect 9548 17484 9554 17496
rect 10502 17484 10508 17536
rect 10560 17524 10566 17536
rect 10689 17527 10747 17533
rect 10689 17524 10701 17527
rect 10560 17496 10701 17524
rect 10560 17484 10566 17496
rect 10689 17493 10701 17496
rect 10735 17524 10747 17527
rect 11238 17524 11244 17536
rect 10735 17496 11244 17524
rect 10735 17493 10747 17496
rect 10689 17487 10747 17493
rect 11238 17484 11244 17496
rect 11296 17524 11302 17536
rect 12158 17524 12164 17536
rect 11296 17496 12164 17524
rect 11296 17484 11302 17496
rect 12158 17484 12164 17496
rect 12216 17484 12222 17536
rect 12342 17524 12348 17536
rect 12303 17496 12348 17524
rect 12342 17484 12348 17496
rect 12400 17484 12406 17536
rect 13906 17524 13912 17536
rect 13867 17496 13912 17524
rect 13906 17484 13912 17496
rect 13964 17484 13970 17536
rect 14090 17484 14096 17536
rect 14148 17524 14154 17536
rect 14461 17527 14519 17533
rect 14461 17524 14473 17527
rect 14148 17496 14473 17524
rect 14148 17484 14154 17496
rect 14461 17493 14473 17496
rect 14507 17524 14519 17527
rect 14737 17527 14795 17533
rect 14737 17524 14749 17527
rect 14507 17496 14749 17524
rect 14507 17493 14519 17496
rect 14461 17487 14519 17493
rect 14737 17493 14749 17496
rect 14783 17524 14795 17527
rect 19168 17524 19196 17564
rect 19794 17552 19800 17564
rect 19852 17552 19858 17604
rect 20806 17592 20812 17604
rect 20767 17564 20812 17592
rect 20806 17552 20812 17564
rect 20864 17552 20870 17604
rect 21358 17592 21364 17604
rect 21319 17564 21364 17592
rect 21358 17552 21364 17564
rect 21416 17552 21422 17604
rect 19702 17524 19708 17536
rect 14783 17496 19196 17524
rect 19663 17496 19708 17524
rect 14783 17493 14795 17496
rect 14737 17487 14795 17493
rect 19702 17484 19708 17496
rect 19760 17484 19766 17536
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 1762 17280 1768 17332
rect 1820 17320 1826 17332
rect 2593 17323 2651 17329
rect 2593 17320 2605 17323
rect 1820 17292 2605 17320
rect 1820 17280 1826 17292
rect 2593 17289 2605 17292
rect 2639 17289 2651 17323
rect 2593 17283 2651 17289
rect 3418 17280 3424 17332
rect 3476 17320 3482 17332
rect 3789 17323 3847 17329
rect 3789 17320 3801 17323
rect 3476 17292 3801 17320
rect 3476 17280 3482 17292
rect 3789 17289 3801 17292
rect 3835 17289 3847 17323
rect 3789 17283 3847 17289
rect 4798 17280 4804 17332
rect 4856 17320 4862 17332
rect 4985 17323 5043 17329
rect 4985 17320 4997 17323
rect 4856 17292 4997 17320
rect 4856 17280 4862 17292
rect 4985 17289 4997 17292
rect 5031 17289 5043 17323
rect 6914 17320 6920 17332
rect 6875 17292 6920 17320
rect 4985 17283 5043 17289
rect 6914 17280 6920 17292
rect 6972 17280 6978 17332
rect 9122 17320 9128 17332
rect 9083 17292 9128 17320
rect 9122 17280 9128 17292
rect 9180 17280 9186 17332
rect 11238 17320 11244 17332
rect 9416 17292 11244 17320
rect 2958 17212 2964 17264
rect 3016 17252 3022 17264
rect 4246 17252 4252 17264
rect 3016 17224 4252 17252
rect 3016 17212 3022 17224
rect 3252 17193 3280 17224
rect 4246 17212 4252 17224
rect 4304 17252 4310 17264
rect 4304 17224 5672 17252
rect 4304 17212 4310 17224
rect 3237 17187 3295 17193
rect 3237 17153 3249 17187
rect 3283 17153 3295 17187
rect 4062 17184 4068 17196
rect 4023 17156 4068 17184
rect 3237 17147 3295 17153
rect 4062 17144 4068 17156
rect 4120 17144 4126 17196
rect 5644 17193 5672 17224
rect 8846 17212 8852 17264
rect 8904 17252 8910 17264
rect 9416 17252 9444 17292
rect 11238 17280 11244 17292
rect 11296 17280 11302 17332
rect 11333 17323 11391 17329
rect 11333 17289 11345 17323
rect 11379 17320 11391 17323
rect 11698 17320 11704 17332
rect 11379 17292 11704 17320
rect 11379 17289 11391 17292
rect 11333 17283 11391 17289
rect 11698 17280 11704 17292
rect 11756 17280 11762 17332
rect 13449 17323 13507 17329
rect 13449 17289 13461 17323
rect 13495 17320 13507 17323
rect 13538 17320 13544 17332
rect 13495 17292 13544 17320
rect 13495 17289 13507 17292
rect 13449 17283 13507 17289
rect 13538 17280 13544 17292
rect 13596 17280 13602 17332
rect 14277 17323 14335 17329
rect 14277 17289 14289 17323
rect 14323 17320 14335 17323
rect 14921 17323 14979 17329
rect 14921 17320 14933 17323
rect 14323 17292 14933 17320
rect 14323 17289 14335 17292
rect 14277 17283 14335 17289
rect 14921 17289 14933 17292
rect 14967 17320 14979 17323
rect 15654 17320 15660 17332
rect 14967 17292 15660 17320
rect 14967 17289 14979 17292
rect 14921 17283 14979 17289
rect 15654 17280 15660 17292
rect 15712 17320 15718 17332
rect 17494 17320 17500 17332
rect 15712 17292 17500 17320
rect 15712 17280 15718 17292
rect 17494 17280 17500 17292
rect 17552 17280 17558 17332
rect 17586 17280 17592 17332
rect 17644 17320 17650 17332
rect 17865 17323 17923 17329
rect 17865 17320 17877 17323
rect 17644 17292 17877 17320
rect 17644 17280 17650 17292
rect 17865 17289 17877 17292
rect 17911 17289 17923 17323
rect 18138 17320 18144 17332
rect 18099 17292 18144 17320
rect 17865 17283 17923 17289
rect 18138 17280 18144 17292
rect 18196 17280 18202 17332
rect 20346 17320 20352 17332
rect 20307 17292 20352 17320
rect 20346 17280 20352 17292
rect 20404 17280 20410 17332
rect 20809 17323 20867 17329
rect 20809 17289 20821 17323
rect 20855 17320 20867 17323
rect 21174 17320 21180 17332
rect 20855 17292 21180 17320
rect 20855 17289 20867 17292
rect 20809 17283 20867 17289
rect 21174 17280 21180 17292
rect 21232 17280 21238 17332
rect 8904 17224 9444 17252
rect 8904 17212 8910 17224
rect 10502 17212 10508 17264
rect 10560 17252 10566 17264
rect 12621 17255 12679 17261
rect 10560 17224 10640 17252
rect 10560 17212 10566 17224
rect 5629 17187 5687 17193
rect 5629 17153 5641 17187
rect 5675 17184 5687 17187
rect 7006 17184 7012 17196
rect 5675 17156 7012 17184
rect 5675 17153 5687 17156
rect 5629 17147 5687 17153
rect 7006 17144 7012 17156
rect 7064 17184 7070 17196
rect 7469 17187 7527 17193
rect 7469 17184 7481 17187
rect 7064 17156 7481 17184
rect 7064 17144 7070 17156
rect 7469 17153 7481 17156
rect 7515 17153 7527 17187
rect 7469 17147 7527 17153
rect 9582 17144 9588 17196
rect 9640 17184 9646 17196
rect 9677 17187 9735 17193
rect 9677 17184 9689 17187
rect 9640 17156 9689 17184
rect 9640 17144 9646 17156
rect 9677 17153 9689 17156
rect 9723 17153 9735 17187
rect 10612 17184 10640 17224
rect 12621 17221 12633 17255
rect 12667 17252 12679 17255
rect 12710 17252 12716 17264
rect 12667 17224 12716 17252
rect 12667 17221 12679 17224
rect 12621 17215 12679 17221
rect 12710 17212 12716 17224
rect 12768 17212 12774 17264
rect 13998 17212 14004 17264
rect 14056 17252 14062 17264
rect 14056 17224 14136 17252
rect 14056 17212 14062 17224
rect 10689 17187 10747 17193
rect 10689 17184 10701 17187
rect 10612 17156 10701 17184
rect 9677 17147 9735 17153
rect 10689 17153 10701 17156
rect 10735 17153 10747 17187
rect 10870 17184 10876 17196
rect 10831 17156 10876 17184
rect 10689 17147 10747 17153
rect 10870 17144 10876 17156
rect 10928 17144 10934 17196
rect 11422 17144 11428 17196
rect 11480 17184 11486 17196
rect 12066 17184 12072 17196
rect 11480 17156 12072 17184
rect 11480 17144 11486 17156
rect 12066 17144 12072 17156
rect 12124 17144 12130 17196
rect 12161 17187 12219 17193
rect 12161 17153 12173 17187
rect 12207 17184 12219 17187
rect 12250 17184 12256 17196
rect 12207 17156 12256 17184
rect 12207 17153 12219 17156
rect 12161 17147 12219 17153
rect 12250 17144 12256 17156
rect 12308 17184 12314 17196
rect 13722 17184 13728 17196
rect 12308 17156 13728 17184
rect 12308 17144 12314 17156
rect 13722 17144 13728 17156
rect 13780 17144 13786 17196
rect 14108 17193 14136 17224
rect 14093 17187 14151 17193
rect 14093 17153 14105 17187
rect 14139 17153 14151 17187
rect 14093 17147 14151 17153
rect 15470 17144 15476 17196
rect 15528 17184 15534 17196
rect 15933 17187 15991 17193
rect 15933 17184 15945 17187
rect 15528 17156 15945 17184
rect 15528 17144 15534 17156
rect 15933 17153 15945 17156
rect 15979 17153 15991 17187
rect 15933 17147 15991 17153
rect 17313 17187 17371 17193
rect 17313 17153 17325 17187
rect 17359 17184 17371 17187
rect 18156 17184 18184 17280
rect 17359 17156 18184 17184
rect 17359 17153 17371 17156
rect 17313 17147 17371 17153
rect 1578 17116 1584 17128
rect 1539 17088 1584 17116
rect 1578 17076 1584 17088
rect 1636 17076 1642 17128
rect 2314 17116 2320 17128
rect 2275 17088 2320 17116
rect 2314 17076 2320 17088
rect 2372 17076 2378 17128
rect 2777 17119 2835 17125
rect 2777 17085 2789 17119
rect 2823 17085 2835 17119
rect 2777 17079 2835 17085
rect 3329 17119 3387 17125
rect 3329 17085 3341 17119
rect 3375 17116 3387 17119
rect 4982 17116 4988 17128
rect 3375 17088 4988 17116
rect 3375 17085 3387 17088
rect 3329 17079 3387 17085
rect 1765 17051 1823 17057
rect 1765 17017 1777 17051
rect 1811 17048 1823 17051
rect 2038 17048 2044 17060
rect 1811 17020 2044 17048
rect 1811 17017 1823 17020
rect 1765 17011 1823 17017
rect 2038 17008 2044 17020
rect 2096 17008 2102 17060
rect 1854 16940 1860 16992
rect 1912 16980 1918 16992
rect 2133 16983 2191 16989
rect 2133 16980 2145 16983
rect 1912 16952 2145 16980
rect 1912 16940 1918 16952
rect 2133 16949 2145 16952
rect 2179 16949 2191 16983
rect 2792 16980 2820 17079
rect 4982 17076 4988 17088
rect 5040 17076 5046 17128
rect 10502 17116 10508 17128
rect 5276 17088 10508 17116
rect 2866 17008 2872 17060
rect 2924 17048 2930 17060
rect 3421 17051 3479 17057
rect 3421 17048 3433 17051
rect 2924 17020 3433 17048
rect 2924 17008 2930 17020
rect 3421 17017 3433 17020
rect 3467 17017 3479 17051
rect 3421 17011 3479 17017
rect 4525 16983 4583 16989
rect 4525 16980 4537 16983
rect 2792 16952 4537 16980
rect 2133 16943 2191 16949
rect 4525 16949 4537 16952
rect 4571 16980 4583 16983
rect 5276 16980 5304 17088
rect 10502 17076 10508 17088
rect 10560 17076 10566 17128
rect 12986 17116 12992 17128
rect 11164 17088 12992 17116
rect 5353 17051 5411 17057
rect 5353 17017 5365 17051
rect 5399 17048 5411 17051
rect 5902 17048 5908 17060
rect 5399 17020 5908 17048
rect 5399 17017 5411 17020
rect 5353 17011 5411 17017
rect 5902 17008 5908 17020
rect 5960 17008 5966 17060
rect 7285 17051 7343 17057
rect 7285 17017 7297 17051
rect 7331 17048 7343 17051
rect 9214 17048 9220 17060
rect 7331 17020 9220 17048
rect 7331 17017 7343 17020
rect 7285 17011 7343 17017
rect 9214 17008 9220 17020
rect 9272 17008 9278 17060
rect 9493 17051 9551 17057
rect 9493 17017 9505 17051
rect 9539 17048 9551 17051
rect 11164 17048 11192 17088
rect 12986 17076 12992 17088
rect 13044 17076 13050 17128
rect 13909 17119 13967 17125
rect 13909 17085 13921 17119
rect 13955 17116 13967 17119
rect 14277 17119 14335 17125
rect 14277 17116 14289 17119
rect 13955 17088 14289 17116
rect 13955 17085 13967 17088
rect 13909 17079 13967 17085
rect 14277 17085 14289 17088
rect 14323 17085 14335 17119
rect 14277 17079 14335 17085
rect 18782 17076 18788 17128
rect 18840 17116 18846 17128
rect 19521 17119 19579 17125
rect 19521 17116 19533 17119
rect 18840 17088 19533 17116
rect 18840 17076 18846 17088
rect 19521 17085 19533 17088
rect 19567 17116 19579 17119
rect 20070 17116 20076 17128
rect 19567 17088 20076 17116
rect 19567 17085 19579 17088
rect 19521 17079 19579 17085
rect 20070 17076 20076 17088
rect 20128 17076 20134 17128
rect 20165 17119 20223 17125
rect 20165 17085 20177 17119
rect 20211 17085 20223 17119
rect 20622 17116 20628 17128
rect 20583 17088 20628 17116
rect 20165 17079 20223 17085
rect 9539 17020 11192 17048
rect 9539 17017 9551 17020
rect 9493 17011 9551 17017
rect 11238 17008 11244 17060
rect 11296 17048 11302 17060
rect 12253 17051 12311 17057
rect 11296 17020 12204 17048
rect 11296 17008 11302 17020
rect 4571 16952 5304 16980
rect 4571 16949 4583 16952
rect 4525 16943 4583 16949
rect 5442 16940 5448 16992
rect 5500 16980 5506 16992
rect 5500 16952 5545 16980
rect 5500 16940 5506 16952
rect 5626 16940 5632 16992
rect 5684 16980 5690 16992
rect 7098 16980 7104 16992
rect 5684 16952 7104 16980
rect 5684 16940 5690 16952
rect 7098 16940 7104 16952
rect 7156 16940 7162 16992
rect 7377 16983 7435 16989
rect 7377 16949 7389 16983
rect 7423 16980 7435 16983
rect 8386 16980 8392 16992
rect 7423 16952 8392 16980
rect 7423 16949 7435 16952
rect 7377 16943 7435 16949
rect 8386 16940 8392 16952
rect 8444 16940 8450 16992
rect 9585 16983 9643 16989
rect 9585 16949 9597 16983
rect 9631 16980 9643 16983
rect 10229 16983 10287 16989
rect 10229 16980 10241 16983
rect 9631 16952 10241 16980
rect 9631 16949 9643 16952
rect 9585 16943 9643 16949
rect 10229 16949 10241 16952
rect 10275 16980 10287 16983
rect 10594 16980 10600 16992
rect 10275 16952 10600 16980
rect 10275 16949 10287 16952
rect 10229 16943 10287 16949
rect 10594 16940 10600 16952
rect 10652 16940 10658 16992
rect 10962 16980 10968 16992
rect 10923 16952 10968 16980
rect 10962 16940 10968 16952
rect 11020 16940 11026 16992
rect 12176 16980 12204 17020
rect 12253 17017 12265 17051
rect 12299 17048 12311 17051
rect 12897 17051 12955 17057
rect 12897 17048 12909 17051
rect 12299 17020 12909 17048
rect 12299 17017 12311 17020
rect 12253 17011 12311 17017
rect 12897 17017 12909 17020
rect 12943 17017 12955 17051
rect 13817 17051 13875 17057
rect 13817 17048 13829 17051
rect 12897 17011 12955 17017
rect 13004 17020 13829 17048
rect 13004 16980 13032 17020
rect 13817 17017 13829 17020
rect 13863 17048 13875 17051
rect 14461 17051 14519 17057
rect 14461 17048 14473 17051
rect 13863 17020 14473 17048
rect 13863 17017 13875 17020
rect 13817 17011 13875 17017
rect 14461 17017 14473 17020
rect 14507 17017 14519 17051
rect 14461 17011 14519 17017
rect 15749 17051 15807 17057
rect 15749 17017 15761 17051
rect 15795 17048 15807 17051
rect 17218 17048 17224 17060
rect 15795 17020 17224 17048
rect 15795 17017 15807 17020
rect 15749 17011 15807 17017
rect 17218 17008 17224 17020
rect 17276 17008 17282 17060
rect 17310 17008 17316 17060
rect 17368 17048 17374 17060
rect 17497 17051 17555 17057
rect 17497 17048 17509 17051
rect 17368 17020 17509 17048
rect 17368 17008 17374 17020
rect 17497 17017 17509 17020
rect 17543 17017 17555 17051
rect 17497 17011 17555 17017
rect 19058 17008 19064 17060
rect 19116 17048 19122 17060
rect 19254 17051 19312 17057
rect 19254 17048 19266 17051
rect 19116 17020 19266 17048
rect 19116 17008 19122 17020
rect 19254 17017 19266 17020
rect 19300 17017 19312 17051
rect 19254 17011 19312 17017
rect 19702 17008 19708 17060
rect 19760 17048 19766 17060
rect 20180 17048 20208 17079
rect 20622 17076 20628 17088
rect 20680 17076 20686 17128
rect 19760 17020 20208 17048
rect 19760 17008 19766 17020
rect 20346 17008 20352 17060
rect 20404 17048 20410 17060
rect 21177 17051 21235 17057
rect 21177 17048 21189 17051
rect 20404 17020 21189 17048
rect 20404 17008 20410 17020
rect 21177 17017 21189 17020
rect 21223 17017 21235 17051
rect 21177 17011 21235 17017
rect 15378 16980 15384 16992
rect 12176 16952 13032 16980
rect 15339 16952 15384 16980
rect 15378 16940 15384 16952
rect 15436 16940 15442 16992
rect 15841 16983 15899 16989
rect 15841 16949 15853 16983
rect 15887 16980 15899 16983
rect 16206 16980 16212 16992
rect 15887 16952 16212 16980
rect 15887 16949 15899 16952
rect 15841 16943 15899 16949
rect 16206 16940 16212 16952
rect 16264 16940 16270 16992
rect 16577 16983 16635 16989
rect 16577 16949 16589 16983
rect 16623 16980 16635 16983
rect 17328 16980 17356 17008
rect 16623 16952 17356 16980
rect 16623 16949 16635 16952
rect 16577 16943 16635 16949
rect 17402 16940 17408 16992
rect 17460 16980 17466 16992
rect 19518 16980 19524 16992
rect 17460 16952 19524 16980
rect 17460 16940 17466 16952
rect 19518 16940 19524 16952
rect 19576 16940 19582 16992
rect 19794 16980 19800 16992
rect 19755 16952 19800 16980
rect 19794 16940 19800 16952
rect 19852 16940 19858 16992
rect 21266 16980 21272 16992
rect 21227 16952 21272 16980
rect 21266 16940 21272 16952
rect 21324 16940 21330 16992
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 2038 16736 2044 16788
rect 2096 16776 2102 16788
rect 2133 16779 2191 16785
rect 2133 16776 2145 16779
rect 2096 16748 2145 16776
rect 2096 16736 2102 16748
rect 2133 16745 2145 16748
rect 2179 16745 2191 16779
rect 2133 16739 2191 16745
rect 2314 16736 2320 16788
rect 2372 16776 2378 16788
rect 3053 16779 3111 16785
rect 3053 16776 3065 16779
rect 2372 16748 3065 16776
rect 2372 16736 2378 16748
rect 3053 16745 3065 16748
rect 3099 16745 3111 16779
rect 5442 16776 5448 16788
rect 5403 16748 5448 16776
rect 3053 16739 3111 16745
rect 5442 16736 5448 16748
rect 5500 16736 5506 16788
rect 5813 16779 5871 16785
rect 5813 16745 5825 16779
rect 5859 16776 5871 16779
rect 6546 16776 6552 16788
rect 5859 16748 6552 16776
rect 5859 16745 5871 16748
rect 5813 16739 5871 16745
rect 6546 16736 6552 16748
rect 6604 16736 6610 16788
rect 6641 16779 6699 16785
rect 6641 16745 6653 16779
rect 6687 16776 6699 16779
rect 6917 16779 6975 16785
rect 6917 16776 6929 16779
rect 6687 16748 6929 16776
rect 6687 16745 6699 16748
rect 6641 16739 6699 16745
rect 6917 16745 6929 16748
rect 6963 16776 6975 16779
rect 8573 16779 8631 16785
rect 6963 16748 8248 16776
rect 6963 16745 6975 16748
rect 6917 16739 6975 16745
rect 1765 16711 1823 16717
rect 1765 16677 1777 16711
rect 1811 16708 1823 16711
rect 2958 16708 2964 16720
rect 1811 16680 2964 16708
rect 1811 16677 1823 16680
rect 1765 16671 1823 16677
rect 2958 16668 2964 16680
rect 3016 16668 3022 16720
rect 4709 16711 4767 16717
rect 4709 16708 4721 16711
rect 3160 16680 4721 16708
rect 1578 16640 1584 16652
rect 1539 16612 1584 16640
rect 1578 16600 1584 16612
rect 1636 16600 1642 16652
rect 2317 16643 2375 16649
rect 2317 16609 2329 16643
rect 2363 16640 2375 16643
rect 2777 16643 2835 16649
rect 2363 16612 2728 16640
rect 2363 16609 2375 16612
rect 2317 16603 2375 16609
rect 2700 16572 2728 16612
rect 2777 16609 2789 16643
rect 2823 16640 2835 16643
rect 3160 16640 3188 16680
rect 4709 16677 4721 16680
rect 4755 16708 4767 16711
rect 5626 16708 5632 16720
rect 4755 16680 5632 16708
rect 4755 16677 4767 16680
rect 4709 16671 4767 16677
rect 5626 16668 5632 16680
rect 5684 16668 5690 16720
rect 5902 16668 5908 16720
rect 5960 16708 5966 16720
rect 8113 16711 8171 16717
rect 8113 16708 8125 16711
rect 5960 16680 8125 16708
rect 5960 16668 5966 16680
rect 8113 16677 8125 16680
rect 8159 16677 8171 16711
rect 8220 16708 8248 16748
rect 8573 16745 8585 16779
rect 8619 16776 8631 16779
rect 10962 16776 10968 16788
rect 8619 16748 10968 16776
rect 8619 16745 8631 16748
rect 8573 16739 8631 16745
rect 10962 16736 10968 16748
rect 11020 16736 11026 16788
rect 11974 16776 11980 16788
rect 11935 16748 11980 16776
rect 11974 16736 11980 16748
rect 12032 16736 12038 16788
rect 14001 16779 14059 16785
rect 14001 16745 14013 16779
rect 14047 16776 14059 16779
rect 14642 16776 14648 16788
rect 14047 16748 14648 16776
rect 14047 16745 14059 16748
rect 14001 16739 14059 16745
rect 14642 16736 14648 16748
rect 14700 16736 14706 16788
rect 14829 16779 14887 16785
rect 14829 16745 14841 16779
rect 14875 16776 14887 16779
rect 15378 16776 15384 16788
rect 14875 16748 15384 16776
rect 14875 16745 14887 16748
rect 14829 16739 14887 16745
rect 15378 16736 15384 16748
rect 15436 16736 15442 16788
rect 16206 16776 16212 16788
rect 16167 16748 16212 16776
rect 16206 16736 16212 16748
rect 16264 16736 16270 16788
rect 16577 16779 16635 16785
rect 16577 16745 16589 16779
rect 16623 16776 16635 16779
rect 16758 16776 16764 16788
rect 16623 16748 16764 16776
rect 16623 16745 16635 16748
rect 16577 16739 16635 16745
rect 16758 16736 16764 16748
rect 16816 16736 16822 16788
rect 17218 16776 17224 16788
rect 17179 16748 17224 16776
rect 17218 16736 17224 16748
rect 17276 16736 17282 16788
rect 19245 16779 19303 16785
rect 19245 16745 19257 16779
rect 19291 16776 19303 16779
rect 20254 16776 20260 16788
rect 19291 16748 20260 16776
rect 19291 16745 19303 16748
rect 19245 16739 19303 16745
rect 20254 16736 20260 16748
rect 20312 16736 20318 16788
rect 20346 16736 20352 16788
rect 20404 16776 20410 16788
rect 20809 16779 20867 16785
rect 20404 16748 20449 16776
rect 20404 16736 20410 16748
rect 20809 16745 20821 16779
rect 20855 16776 20867 16779
rect 21174 16776 21180 16788
rect 20855 16748 21180 16776
rect 20855 16745 20867 16748
rect 20809 16739 20867 16745
rect 21174 16736 21180 16748
rect 21232 16736 21238 16788
rect 9122 16708 9128 16720
rect 8220 16680 9128 16708
rect 8113 16671 8171 16677
rect 9122 16668 9128 16680
rect 9180 16668 9186 16720
rect 9214 16668 9220 16720
rect 9272 16708 9278 16720
rect 10870 16708 10876 16720
rect 9272 16680 10876 16708
rect 9272 16668 9278 16680
rect 10870 16668 10876 16680
rect 10928 16708 10934 16720
rect 11241 16711 11299 16717
rect 11241 16708 11253 16711
rect 10928 16680 11253 16708
rect 10928 16668 10934 16680
rect 11241 16677 11253 16680
rect 11287 16677 11299 16711
rect 11241 16671 11299 16677
rect 11333 16711 11391 16717
rect 11333 16677 11345 16711
rect 11379 16708 11391 16711
rect 12345 16711 12403 16717
rect 11379 16680 12204 16708
rect 11379 16677 11391 16680
rect 11333 16671 11391 16677
rect 2823 16612 3188 16640
rect 3237 16643 3295 16649
rect 2823 16609 2835 16612
rect 2777 16603 2835 16609
rect 3237 16609 3249 16643
rect 3283 16640 3295 16643
rect 4154 16640 4160 16652
rect 3283 16612 4160 16640
rect 3283 16609 3295 16612
rect 3237 16603 3295 16609
rect 4154 16600 4160 16612
rect 4212 16600 4218 16652
rect 4341 16643 4399 16649
rect 4341 16609 4353 16643
rect 4387 16640 4399 16643
rect 6641 16643 6699 16649
rect 6641 16640 6653 16643
rect 4387 16612 6653 16640
rect 4387 16609 4399 16612
rect 4341 16603 4399 16609
rect 3510 16572 3516 16584
rect 2700 16544 3516 16572
rect 3510 16532 3516 16544
rect 3568 16532 3574 16584
rect 3602 16532 3608 16584
rect 3660 16572 3666 16584
rect 4356 16572 4384 16603
rect 5920 16581 5948 16612
rect 6641 16609 6653 16612
rect 6687 16609 6699 16643
rect 6641 16603 6699 16609
rect 8205 16643 8263 16649
rect 8205 16609 8217 16643
rect 8251 16640 8263 16643
rect 8386 16640 8392 16652
rect 8251 16612 8392 16640
rect 8251 16609 8263 16612
rect 8205 16603 8263 16609
rect 8386 16600 8392 16612
rect 8444 16640 8450 16652
rect 9306 16640 9312 16652
rect 8444 16612 9312 16640
rect 8444 16600 8450 16612
rect 9306 16600 9312 16612
rect 9364 16600 9370 16652
rect 10410 16600 10416 16652
rect 10468 16640 10474 16652
rect 10689 16643 10747 16649
rect 10689 16640 10701 16643
rect 10468 16612 10701 16640
rect 10468 16600 10474 16612
rect 10689 16609 10701 16612
rect 10735 16640 10747 16643
rect 11348 16640 11376 16671
rect 10735 16612 11376 16640
rect 12176 16640 12204 16680
rect 12345 16677 12357 16711
rect 12391 16708 12403 16711
rect 12710 16708 12716 16720
rect 12391 16680 12716 16708
rect 12391 16677 12403 16680
rect 12345 16671 12403 16677
rect 12710 16668 12716 16680
rect 12768 16668 12774 16720
rect 12820 16680 13768 16708
rect 12820 16640 12848 16680
rect 12176 16612 12848 16640
rect 10735 16609 10747 16612
rect 10689 16603 10747 16609
rect 12986 16600 12992 16652
rect 13044 16640 13050 16652
rect 13541 16643 13599 16649
rect 13541 16640 13553 16643
rect 13044 16612 13553 16640
rect 13044 16600 13050 16612
rect 13541 16609 13553 16612
rect 13587 16609 13599 16643
rect 13541 16603 13599 16609
rect 13633 16643 13691 16649
rect 13633 16609 13645 16643
rect 13679 16609 13691 16643
rect 13740 16640 13768 16680
rect 13906 16668 13912 16720
rect 13964 16708 13970 16720
rect 14921 16711 14979 16717
rect 14921 16708 14933 16711
rect 13964 16680 14933 16708
rect 13964 16668 13970 16680
rect 14921 16677 14933 16680
rect 14967 16677 14979 16711
rect 14921 16671 14979 16677
rect 15028 16680 19564 16708
rect 15028 16640 15056 16680
rect 16114 16640 16120 16652
rect 13740 16612 15056 16640
rect 15304 16612 16120 16640
rect 13633 16603 13691 16609
rect 3660 16544 4384 16572
rect 5905 16575 5963 16581
rect 3660 16532 3666 16544
rect 5905 16541 5917 16575
rect 5951 16541 5963 16575
rect 5905 16535 5963 16541
rect 5994 16532 6000 16584
rect 6052 16572 6058 16584
rect 8021 16575 8079 16581
rect 6052 16544 6097 16572
rect 6052 16532 6058 16544
rect 8021 16541 8033 16575
rect 8067 16572 8079 16575
rect 9398 16572 9404 16584
rect 8067 16544 9404 16572
rect 8067 16541 8079 16544
rect 8021 16535 8079 16541
rect 9398 16532 9404 16544
rect 9456 16572 9462 16584
rect 11149 16575 11207 16581
rect 11149 16572 11161 16575
rect 9456 16544 11161 16572
rect 9456 16532 9462 16544
rect 11149 16541 11161 16544
rect 11195 16572 11207 16575
rect 11422 16572 11428 16584
rect 11195 16544 11428 16572
rect 11195 16541 11207 16544
rect 11149 16535 11207 16541
rect 11422 16532 11428 16544
rect 11480 16532 11486 16584
rect 12437 16575 12495 16581
rect 12437 16572 12449 16575
rect 11716 16544 12449 16572
rect 2590 16504 2596 16516
rect 2551 16476 2596 16504
rect 2590 16464 2596 16476
rect 2648 16464 2654 16516
rect 11716 16513 11744 16544
rect 12437 16541 12449 16544
rect 12483 16541 12495 16575
rect 12437 16535 12495 16541
rect 12529 16575 12587 16581
rect 12529 16541 12541 16575
rect 12575 16541 12587 16575
rect 13354 16572 13360 16584
rect 13315 16544 13360 16572
rect 12529 16535 12587 16541
rect 11701 16507 11759 16513
rect 11701 16473 11713 16507
rect 11747 16473 11759 16507
rect 11701 16467 11759 16473
rect 12158 16464 12164 16516
rect 12216 16504 12222 16516
rect 12544 16504 12572 16535
rect 13354 16532 13360 16544
rect 13412 16532 13418 16584
rect 13648 16572 13676 16603
rect 13556 16544 13676 16572
rect 12216 16476 12572 16504
rect 12216 16464 12222 16476
rect 13078 16464 13084 16516
rect 13136 16504 13142 16516
rect 13556 16504 13584 16544
rect 14550 16532 14556 16584
rect 14608 16572 14614 16584
rect 14645 16575 14703 16581
rect 14645 16572 14657 16575
rect 14608 16544 14657 16572
rect 14608 16532 14614 16544
rect 14645 16541 14657 16544
rect 14691 16541 14703 16575
rect 14645 16535 14703 16541
rect 15304 16513 15332 16612
rect 16114 16600 16120 16612
rect 16172 16600 16178 16652
rect 16669 16643 16727 16649
rect 16669 16609 16681 16643
rect 16715 16640 16727 16643
rect 17402 16640 17408 16652
rect 16715 16612 17408 16640
rect 16715 16609 16727 16612
rect 16669 16603 16727 16609
rect 17402 16600 17408 16612
rect 17460 16600 17466 16652
rect 17589 16643 17647 16649
rect 17589 16609 17601 16643
rect 17635 16640 17647 16643
rect 17862 16640 17868 16652
rect 17635 16612 17868 16640
rect 17635 16609 17647 16612
rect 17589 16603 17647 16609
rect 17862 16600 17868 16612
rect 17920 16600 17926 16652
rect 18874 16600 18880 16652
rect 18932 16640 18938 16652
rect 19061 16643 19119 16649
rect 19061 16640 19073 16643
rect 18932 16612 19073 16640
rect 18932 16600 18938 16612
rect 19061 16609 19073 16612
rect 19107 16609 19119 16643
rect 19536 16640 19564 16680
rect 19978 16668 19984 16720
rect 20036 16708 20042 16720
rect 20036 16680 20668 16708
rect 20036 16668 20042 16680
rect 19794 16640 19800 16652
rect 19536 16612 19800 16640
rect 19061 16603 19119 16609
rect 19794 16600 19800 16612
rect 19852 16640 19858 16652
rect 20640 16649 20668 16680
rect 20165 16643 20223 16649
rect 20165 16640 20177 16643
rect 19852 16612 20177 16640
rect 19852 16600 19858 16612
rect 20165 16609 20177 16612
rect 20211 16609 20223 16643
rect 20165 16603 20223 16609
rect 20625 16643 20683 16649
rect 20625 16609 20637 16643
rect 20671 16609 20683 16643
rect 21177 16643 21235 16649
rect 21177 16640 21189 16643
rect 20625 16603 20683 16609
rect 20732 16612 21189 16640
rect 16761 16575 16819 16581
rect 16761 16572 16773 16575
rect 15396 16544 16773 16572
rect 13136 16476 13584 16504
rect 15289 16507 15347 16513
rect 13136 16464 13142 16476
rect 15289 16473 15301 16507
rect 15335 16473 15347 16507
rect 15289 16467 15347 16473
rect 2774 16396 2780 16448
rect 2832 16436 2838 16448
rect 3881 16439 3939 16445
rect 3881 16436 3893 16439
rect 2832 16408 3893 16436
rect 2832 16396 2838 16408
rect 3881 16405 3893 16408
rect 3927 16436 3939 16439
rect 5258 16436 5264 16448
rect 3927 16408 5264 16436
rect 3927 16405 3939 16408
rect 3881 16399 3939 16405
rect 5258 16396 5264 16408
rect 5316 16396 5322 16448
rect 13998 16396 14004 16448
rect 14056 16436 14062 16448
rect 15396 16436 15424 16544
rect 16761 16541 16773 16544
rect 16807 16541 16819 16575
rect 16761 16535 16819 16541
rect 16776 16504 16804 16535
rect 17310 16532 17316 16584
rect 17368 16572 17374 16584
rect 17681 16575 17739 16581
rect 17681 16572 17693 16575
rect 17368 16544 17693 16572
rect 17368 16532 17374 16544
rect 17681 16541 17693 16544
rect 17727 16541 17739 16575
rect 17681 16535 17739 16541
rect 17773 16575 17831 16581
rect 17773 16541 17785 16575
rect 17819 16541 17831 16575
rect 17773 16535 17831 16541
rect 17788 16504 17816 16535
rect 19886 16532 19892 16584
rect 19944 16572 19950 16584
rect 20732 16572 20760 16612
rect 21177 16609 21189 16612
rect 21223 16609 21235 16643
rect 21358 16640 21364 16652
rect 21319 16612 21364 16640
rect 21177 16603 21235 16609
rect 21358 16600 21364 16612
rect 21416 16600 21422 16652
rect 19944 16544 20760 16572
rect 19944 16532 19950 16544
rect 16776 16476 17816 16504
rect 14056 16408 15424 16436
rect 14056 16396 14062 16408
rect 15470 16396 15476 16448
rect 15528 16436 15534 16448
rect 18598 16436 18604 16448
rect 15528 16408 18604 16436
rect 15528 16396 15534 16408
rect 18598 16396 18604 16408
rect 18656 16396 18662 16448
rect 19610 16396 19616 16448
rect 19668 16436 19674 16448
rect 19797 16439 19855 16445
rect 19797 16436 19809 16439
rect 19668 16408 19809 16436
rect 19668 16396 19674 16408
rect 19797 16405 19809 16408
rect 19843 16405 19855 16439
rect 19797 16399 19855 16405
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 2958 16192 2964 16244
rect 3016 16232 3022 16244
rect 3053 16235 3111 16241
rect 3053 16232 3065 16235
rect 3016 16204 3065 16232
rect 3016 16192 3022 16204
rect 3053 16201 3065 16204
rect 3099 16201 3111 16235
rect 3510 16232 3516 16244
rect 3471 16204 3516 16232
rect 3053 16195 3111 16201
rect 3510 16192 3516 16204
rect 3568 16192 3574 16244
rect 5721 16235 5779 16241
rect 3988 16204 5672 16232
rect 3988 16173 4016 16204
rect 3973 16167 4031 16173
rect 3973 16164 3985 16167
rect 2332 16136 3985 16164
rect 1578 16096 1584 16108
rect 1539 16068 1584 16096
rect 1578 16056 1584 16068
rect 1636 16056 1642 16108
rect 2332 16037 2360 16136
rect 3973 16133 3985 16136
rect 4019 16133 4031 16167
rect 5644 16164 5672 16204
rect 5721 16201 5733 16235
rect 5767 16232 5779 16235
rect 5994 16232 6000 16244
rect 5767 16204 6000 16232
rect 5767 16201 5779 16204
rect 5721 16195 5779 16201
rect 5994 16192 6000 16204
rect 6052 16192 6058 16244
rect 7650 16192 7656 16244
rect 7708 16232 7714 16244
rect 7929 16235 7987 16241
rect 7929 16232 7941 16235
rect 7708 16204 7941 16232
rect 7708 16192 7714 16204
rect 7929 16201 7941 16204
rect 7975 16201 7987 16235
rect 7929 16195 7987 16201
rect 8573 16235 8631 16241
rect 8573 16201 8585 16235
rect 8619 16232 8631 16235
rect 9582 16232 9588 16244
rect 8619 16204 9588 16232
rect 8619 16201 8631 16204
rect 8573 16195 8631 16201
rect 7282 16164 7288 16176
rect 5644 16136 7288 16164
rect 3973 16127 4031 16133
rect 7282 16124 7288 16136
rect 7340 16124 7346 16176
rect 7377 16099 7435 16105
rect 3712 16068 4476 16096
rect 2317 16031 2375 16037
rect 2317 15997 2329 16031
rect 2363 15997 2375 16031
rect 2774 16028 2780 16040
rect 2735 16000 2780 16028
rect 2317 15991 2375 15997
rect 2774 15988 2780 16000
rect 2832 15988 2838 16040
rect 3237 16031 3295 16037
rect 3237 15997 3249 16031
rect 3283 16028 3295 16031
rect 3602 16028 3608 16040
rect 3283 16000 3608 16028
rect 3283 15997 3295 16000
rect 3237 15991 3295 15997
rect 3602 15988 3608 16000
rect 3660 15988 3666 16040
rect 3712 16037 3740 16068
rect 3697 16031 3755 16037
rect 3697 15997 3709 16031
rect 3743 15997 3755 16031
rect 4338 16028 4344 16040
rect 4299 16000 4344 16028
rect 3697 15991 3755 15997
rect 4338 15988 4344 16000
rect 4396 15988 4402 16040
rect 4448 16028 4476 16068
rect 7377 16065 7389 16099
rect 7423 16096 7435 16099
rect 8588 16096 8616 16195
rect 9582 16192 9588 16204
rect 9640 16192 9646 16244
rect 13078 16192 13084 16244
rect 13136 16232 13142 16244
rect 19610 16232 19616 16244
rect 13136 16204 19616 16232
rect 13136 16192 13142 16204
rect 19610 16192 19616 16204
rect 19668 16192 19674 16244
rect 19886 16232 19892 16244
rect 19847 16204 19892 16232
rect 19886 16192 19892 16204
rect 19944 16192 19950 16244
rect 19429 16167 19487 16173
rect 19429 16133 19441 16167
rect 19475 16164 19487 16167
rect 20622 16164 20628 16176
rect 19475 16136 20628 16164
rect 19475 16133 19487 16136
rect 19429 16127 19487 16133
rect 20622 16124 20628 16136
rect 20680 16124 20686 16176
rect 7423 16068 8616 16096
rect 7423 16065 7435 16068
rect 7377 16059 7435 16065
rect 11054 16056 11060 16108
rect 11112 16096 11118 16108
rect 17034 16096 17040 16108
rect 11112 16068 17040 16096
rect 11112 16056 11118 16068
rect 17034 16056 17040 16068
rect 17092 16056 17098 16108
rect 18598 16056 18604 16108
rect 18656 16096 18662 16108
rect 18656 16068 19748 16096
rect 18656 16056 18662 16068
rect 5718 16028 5724 16040
rect 4448 16000 5724 16028
rect 5718 15988 5724 16000
rect 5776 15988 5782 16040
rect 6270 15988 6276 16040
rect 6328 16028 6334 16040
rect 6825 16031 6883 16037
rect 6825 16028 6837 16031
rect 6328 16000 6837 16028
rect 6328 15988 6334 16000
rect 6825 15997 6837 16000
rect 6871 16028 6883 16031
rect 7469 16031 7527 16037
rect 7469 16028 7481 16031
rect 6871 16000 7481 16028
rect 6871 15997 6883 16000
rect 6825 15991 6883 15997
rect 7469 15997 7481 16000
rect 7515 15997 7527 16031
rect 9953 16031 10011 16037
rect 9953 16028 9965 16031
rect 7469 15991 7527 15997
rect 9508 16000 9965 16028
rect 9508 15972 9536 16000
rect 9953 15997 9965 16000
rect 9999 15997 10011 16031
rect 9953 15991 10011 15997
rect 15286 15988 15292 16040
rect 15344 16028 15350 16040
rect 19720 16037 19748 16068
rect 19245 16031 19303 16037
rect 19245 16028 19257 16031
rect 15344 16000 19257 16028
rect 15344 15988 15350 16000
rect 19245 15997 19257 16000
rect 19291 15997 19303 16031
rect 19245 15991 19303 15997
rect 19705 16031 19763 16037
rect 19705 15997 19717 16031
rect 19751 15997 19763 16031
rect 19705 15991 19763 15997
rect 20165 16031 20223 16037
rect 20165 15997 20177 16031
rect 20211 15997 20223 16031
rect 20165 15991 20223 15997
rect 1765 15963 1823 15969
rect 1765 15929 1777 15963
rect 1811 15960 1823 15963
rect 1811 15932 2636 15960
rect 1811 15929 1823 15932
rect 1765 15923 1823 15929
rect 2133 15895 2191 15901
rect 2133 15861 2145 15895
rect 2179 15892 2191 15895
rect 2314 15892 2320 15904
rect 2179 15864 2320 15892
rect 2179 15861 2191 15864
rect 2133 15855 2191 15861
rect 2314 15852 2320 15864
rect 2372 15852 2378 15904
rect 2608 15901 2636 15932
rect 3786 15920 3792 15972
rect 3844 15960 3850 15972
rect 3844 15932 4108 15960
rect 3844 15920 3850 15932
rect 2593 15895 2651 15901
rect 2593 15861 2605 15895
rect 2639 15861 2651 15895
rect 4080 15892 4108 15932
rect 4246 15920 4252 15972
rect 4304 15960 4310 15972
rect 4586 15963 4644 15969
rect 4586 15960 4598 15963
rect 4304 15932 4598 15960
rect 4304 15920 4310 15932
rect 4586 15929 4598 15932
rect 4632 15929 4644 15963
rect 4586 15923 4644 15929
rect 6549 15963 6607 15969
rect 6549 15929 6561 15963
rect 6595 15960 6607 15963
rect 7561 15963 7619 15969
rect 7561 15960 7573 15963
rect 6595 15932 7573 15960
rect 6595 15929 6607 15932
rect 6549 15923 6607 15929
rect 7561 15929 7573 15932
rect 7607 15929 7619 15963
rect 7561 15923 7619 15929
rect 6564 15892 6592 15923
rect 9490 15920 9496 15972
rect 9548 15920 9554 15972
rect 9708 15963 9766 15969
rect 9708 15929 9720 15963
rect 9754 15960 9766 15963
rect 9858 15960 9864 15972
rect 9754 15932 9864 15960
rect 9754 15929 9766 15932
rect 9708 15923 9766 15929
rect 9858 15920 9864 15932
rect 9916 15920 9922 15972
rect 20180 15960 20208 15991
rect 20254 15988 20260 16040
rect 20312 16028 20318 16040
rect 20625 16031 20683 16037
rect 20625 16028 20637 16031
rect 20312 16000 20637 16028
rect 20312 15988 20318 16000
rect 20625 15997 20637 16000
rect 20671 15997 20683 16031
rect 20625 15991 20683 15997
rect 21177 15963 21235 15969
rect 21177 15960 21189 15963
rect 18892 15932 20208 15960
rect 20824 15932 21189 15960
rect 4080 15864 6592 15892
rect 2593 15855 2651 15861
rect 11054 15852 11060 15904
rect 11112 15892 11118 15904
rect 11701 15895 11759 15901
rect 11701 15892 11713 15895
rect 11112 15864 11713 15892
rect 11112 15852 11118 15864
rect 11701 15861 11713 15864
rect 11747 15892 11759 15895
rect 12250 15892 12256 15904
rect 11747 15864 12256 15892
rect 11747 15861 11759 15864
rect 11701 15855 11759 15861
rect 12250 15852 12256 15864
rect 12308 15852 12314 15904
rect 13078 15892 13084 15904
rect 13039 15864 13084 15892
rect 13078 15852 13084 15864
rect 13136 15852 13142 15904
rect 16758 15852 16764 15904
rect 16816 15892 16822 15904
rect 17037 15895 17095 15901
rect 17037 15892 17049 15895
rect 16816 15864 17049 15892
rect 16816 15852 16822 15864
rect 17037 15861 17049 15864
rect 17083 15861 17095 15895
rect 17037 15855 17095 15861
rect 17310 15852 17316 15904
rect 17368 15892 17374 15904
rect 17405 15895 17463 15901
rect 17405 15892 17417 15895
rect 17368 15864 17417 15892
rect 17368 15852 17374 15864
rect 17405 15861 17417 15864
rect 17451 15861 17463 15895
rect 18598 15892 18604 15904
rect 18559 15864 18604 15892
rect 17405 15855 17463 15861
rect 18598 15852 18604 15864
rect 18656 15852 18662 15904
rect 18690 15852 18696 15904
rect 18748 15892 18754 15904
rect 18892 15901 18920 15932
rect 18877 15895 18935 15901
rect 18877 15892 18889 15895
rect 18748 15864 18889 15892
rect 18748 15852 18754 15864
rect 18877 15861 18889 15864
rect 18923 15861 18935 15895
rect 20346 15892 20352 15904
rect 20307 15864 20352 15892
rect 18877 15855 18935 15861
rect 20346 15852 20352 15864
rect 20404 15852 20410 15904
rect 20824 15901 20852 15932
rect 21177 15929 21189 15932
rect 21223 15929 21235 15963
rect 21177 15923 21235 15929
rect 21361 15963 21419 15969
rect 21361 15929 21373 15963
rect 21407 15960 21419 15963
rect 22005 15963 22063 15969
rect 22005 15960 22017 15963
rect 21407 15932 22017 15960
rect 21407 15929 21419 15932
rect 21361 15923 21419 15929
rect 22005 15929 22017 15932
rect 22051 15929 22063 15963
rect 22005 15923 22063 15929
rect 20809 15895 20867 15901
rect 20809 15861 20821 15895
rect 20855 15861 20867 15895
rect 20809 15855 20867 15861
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 4065 15691 4123 15697
rect 4065 15657 4077 15691
rect 4111 15688 4123 15691
rect 4246 15688 4252 15700
rect 4111 15660 4252 15688
rect 4111 15657 4123 15660
rect 4065 15651 4123 15657
rect 1765 15623 1823 15629
rect 1765 15589 1777 15623
rect 1811 15620 1823 15623
rect 1854 15620 1860 15632
rect 1811 15592 1860 15620
rect 1811 15589 1823 15592
rect 1765 15583 1823 15589
rect 1854 15580 1860 15592
rect 1912 15580 1918 15632
rect 2130 15620 2136 15632
rect 2091 15592 2136 15620
rect 2130 15580 2136 15592
rect 2188 15580 2194 15632
rect 2314 15620 2320 15632
rect 2275 15592 2320 15620
rect 2314 15580 2320 15592
rect 2372 15580 2378 15632
rect 4080 15620 4108 15651
rect 4246 15648 4252 15660
rect 4304 15648 4310 15700
rect 15286 15688 15292 15700
rect 15247 15660 15292 15688
rect 15286 15648 15292 15660
rect 15344 15648 15350 15700
rect 20257 15691 20315 15697
rect 20257 15657 20269 15691
rect 20303 15688 20315 15691
rect 20303 15660 21220 15688
rect 20303 15657 20315 15660
rect 20257 15651 20315 15657
rect 2884 15592 4108 15620
rect 2884 15493 2912 15592
rect 4338 15580 4344 15632
rect 4396 15620 4402 15632
rect 5350 15620 5356 15632
rect 4396 15592 5356 15620
rect 4396 15580 4402 15592
rect 5350 15580 5356 15592
rect 5408 15620 5414 15632
rect 12342 15620 12348 15632
rect 12400 15629 12406 15632
rect 5408 15592 5488 15620
rect 12312 15592 12348 15620
rect 5408 15580 5414 15592
rect 3050 15552 3056 15564
rect 3011 15524 3056 15552
rect 3050 15512 3056 15524
rect 3108 15512 3114 15564
rect 5166 15512 5172 15564
rect 5224 15561 5230 15564
rect 5224 15552 5236 15561
rect 5224 15524 5269 15552
rect 5224 15515 5236 15524
rect 5224 15512 5230 15515
rect 5460 15496 5488 15592
rect 12342 15580 12348 15592
rect 12400 15583 12412 15629
rect 15832 15623 15890 15629
rect 15832 15589 15844 15623
rect 15878 15620 15890 15623
rect 15930 15620 15936 15632
rect 15878 15592 15936 15620
rect 15878 15589 15890 15592
rect 15832 15583 15890 15589
rect 12400 15580 12406 15583
rect 15930 15580 15936 15592
rect 15988 15580 15994 15632
rect 20346 15580 20352 15632
rect 20404 15620 20410 15632
rect 21192 15629 21220 15660
rect 20625 15623 20683 15629
rect 20625 15620 20637 15623
rect 20404 15592 20637 15620
rect 20404 15580 20410 15592
rect 20625 15589 20637 15592
rect 20671 15589 20683 15623
rect 20625 15583 20683 15589
rect 21177 15623 21235 15629
rect 21177 15589 21189 15623
rect 21223 15589 21235 15623
rect 21177 15583 21235 15589
rect 7282 15512 7288 15564
rect 7340 15552 7346 15564
rect 7662 15555 7720 15561
rect 7662 15552 7674 15555
rect 7340 15524 7674 15552
rect 7340 15512 7346 15524
rect 7662 15521 7674 15524
rect 7708 15521 7720 15555
rect 7662 15515 7720 15521
rect 8478 15512 8484 15564
rect 8536 15552 8542 15564
rect 9309 15555 9367 15561
rect 9309 15552 9321 15555
rect 8536 15524 9321 15552
rect 8536 15512 8542 15524
rect 9309 15521 9321 15524
rect 9355 15521 9367 15555
rect 12618 15552 12624 15564
rect 12579 15524 12624 15552
rect 9309 15515 9367 15521
rect 12618 15512 12624 15524
rect 12676 15512 12682 15564
rect 14918 15552 14924 15564
rect 14879 15524 14924 15552
rect 14918 15512 14924 15524
rect 14976 15512 14982 15564
rect 17954 15561 17960 15564
rect 17948 15515 17960 15561
rect 18012 15552 18018 15564
rect 18012 15524 18048 15552
rect 17954 15512 17960 15515
rect 18012 15512 18018 15524
rect 19610 15512 19616 15564
rect 19668 15552 19674 15564
rect 20073 15555 20131 15561
rect 20073 15552 20085 15555
rect 19668 15524 20085 15552
rect 19668 15512 19674 15524
rect 20073 15521 20085 15524
rect 20119 15521 20131 15555
rect 20806 15552 20812 15564
rect 20767 15524 20812 15552
rect 20073 15515 20131 15521
rect 20806 15512 20812 15524
rect 20864 15512 20870 15564
rect 2869 15487 2927 15493
rect 2869 15453 2881 15487
rect 2915 15453 2927 15487
rect 2869 15447 2927 15453
rect 2961 15487 3019 15493
rect 2961 15453 2973 15487
rect 3007 15484 3019 15487
rect 4062 15484 4068 15496
rect 3007 15456 4068 15484
rect 3007 15453 3019 15456
rect 2961 15447 3019 15453
rect 4062 15444 4068 15456
rect 4120 15444 4126 15496
rect 5442 15484 5448 15496
rect 5403 15456 5448 15484
rect 5442 15444 5448 15456
rect 5500 15444 5506 15496
rect 7929 15487 7987 15493
rect 7929 15453 7941 15487
rect 7975 15484 7987 15487
rect 8386 15484 8392 15496
rect 7975 15456 8392 15484
rect 7975 15453 7987 15456
rect 7929 15447 7987 15453
rect 8386 15444 8392 15456
rect 8444 15444 8450 15496
rect 14550 15444 14556 15496
rect 14608 15484 14614 15496
rect 14645 15487 14703 15493
rect 14645 15484 14657 15487
rect 14608 15456 14657 15484
rect 14608 15444 14614 15456
rect 14645 15453 14657 15456
rect 14691 15453 14703 15487
rect 14645 15447 14703 15453
rect 14734 15444 14740 15496
rect 14792 15484 14798 15496
rect 14829 15487 14887 15493
rect 14829 15484 14841 15487
rect 14792 15456 14841 15484
rect 14792 15444 14798 15456
rect 14829 15453 14841 15456
rect 14875 15453 14887 15487
rect 15562 15484 15568 15496
rect 15523 15456 15568 15484
rect 14829 15447 14887 15453
rect 15562 15444 15568 15456
rect 15620 15444 15626 15496
rect 17126 15444 17132 15496
rect 17184 15484 17190 15496
rect 17681 15487 17739 15493
rect 17681 15484 17693 15487
rect 17184 15456 17693 15484
rect 17184 15444 17190 15456
rect 17681 15453 17693 15456
rect 17727 15453 17739 15487
rect 17681 15447 17739 15453
rect 1670 15348 1676 15360
rect 1631 15320 1676 15348
rect 1670 15308 1676 15320
rect 1728 15308 1734 15360
rect 3421 15351 3479 15357
rect 3421 15317 3433 15351
rect 3467 15348 3479 15351
rect 4246 15348 4252 15360
rect 3467 15320 4252 15348
rect 3467 15317 3479 15320
rect 3421 15311 3479 15317
rect 4246 15308 4252 15320
rect 4304 15308 4310 15360
rect 6546 15348 6552 15360
rect 6507 15320 6552 15348
rect 6546 15308 6552 15320
rect 6604 15308 6610 15360
rect 9490 15348 9496 15360
rect 9451 15320 9496 15348
rect 9490 15308 9496 15320
rect 9548 15308 9554 15360
rect 11241 15351 11299 15357
rect 11241 15317 11253 15351
rect 11287 15348 11299 15351
rect 11882 15348 11888 15360
rect 11287 15320 11888 15348
rect 11287 15317 11299 15320
rect 11241 15311 11299 15317
rect 11882 15308 11888 15320
rect 11940 15308 11946 15360
rect 16945 15351 17003 15357
rect 16945 15317 16957 15351
rect 16991 15348 17003 15351
rect 17586 15348 17592 15360
rect 16991 15320 17592 15348
rect 16991 15317 17003 15320
rect 16945 15311 17003 15317
rect 17586 15308 17592 15320
rect 17644 15308 17650 15360
rect 19058 15348 19064 15360
rect 19019 15320 19064 15348
rect 19058 15308 19064 15320
rect 19116 15308 19122 15360
rect 19334 15308 19340 15360
rect 19392 15348 19398 15360
rect 19610 15348 19616 15360
rect 19392 15320 19616 15348
rect 19392 15308 19398 15320
rect 19610 15308 19616 15320
rect 19668 15308 19674 15360
rect 21266 15348 21272 15360
rect 21227 15320 21272 15348
rect 21266 15308 21272 15320
rect 21324 15308 21330 15360
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 22002 15212 22008 15224
rect 1104 15184 21896 15206
rect 21963 15184 22008 15212
rect 22002 15172 22008 15184
rect 22060 15172 22066 15224
rect 4154 15144 4160 15156
rect 4115 15116 4160 15144
rect 4154 15104 4160 15116
rect 4212 15104 4218 15156
rect 7098 15104 7104 15156
rect 7156 15144 7162 15156
rect 8202 15144 8208 15156
rect 7156 15116 8208 15144
rect 7156 15104 7162 15116
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 9858 15104 9864 15156
rect 9916 15144 9922 15156
rect 9953 15147 10011 15153
rect 9953 15144 9965 15147
rect 9916 15116 9965 15144
rect 9916 15104 9922 15116
rect 9953 15113 9965 15116
rect 9999 15113 10011 15147
rect 9953 15107 10011 15113
rect 12250 15104 12256 15156
rect 12308 15144 12314 15156
rect 14737 15147 14795 15153
rect 12308 15116 14688 15144
rect 12308 15104 12314 15116
rect 9674 15036 9680 15088
rect 9732 15076 9738 15088
rect 14660 15076 14688 15116
rect 14737 15113 14749 15147
rect 14783 15144 14795 15147
rect 14918 15144 14924 15156
rect 14783 15116 14924 15144
rect 14783 15113 14795 15116
rect 14737 15107 14795 15113
rect 14918 15104 14924 15116
rect 14976 15104 14982 15156
rect 19702 15144 19708 15156
rect 18432 15116 19708 15144
rect 18432 15076 18460 15116
rect 19702 15104 19708 15116
rect 19760 15104 19766 15156
rect 9732 15048 9777 15076
rect 14660 15048 18460 15076
rect 18509 15079 18567 15085
rect 9732 15036 9738 15048
rect 18509 15045 18521 15079
rect 18555 15045 18567 15079
rect 18509 15039 18567 15045
rect 3789 15011 3847 15017
rect 3789 14977 3801 15011
rect 3835 15008 3847 15011
rect 4338 15008 4344 15020
rect 3835 14980 4344 15008
rect 3835 14977 3847 14980
rect 3789 14971 3847 14977
rect 4338 14968 4344 14980
rect 4396 14968 4402 15020
rect 12618 14968 12624 15020
rect 12676 15008 12682 15020
rect 13081 15011 13139 15017
rect 13081 15008 13093 15011
rect 12676 14980 13093 15008
rect 12676 14968 12682 14980
rect 13081 14977 13093 14980
rect 13127 14977 13139 15011
rect 15289 15011 15347 15017
rect 15289 15008 15301 15011
rect 13081 14971 13139 14977
rect 14108 14980 15301 15008
rect 6546 14900 6552 14952
rect 6604 14940 6610 14952
rect 8021 14943 8079 14949
rect 6604 14912 7880 14940
rect 6604 14900 6610 14912
rect 1765 14875 1823 14881
rect 1765 14841 1777 14875
rect 1811 14872 1823 14875
rect 2590 14872 2596 14884
rect 1811 14844 2596 14872
rect 1811 14841 1823 14844
rect 1765 14835 1823 14841
rect 2590 14832 2596 14844
rect 2648 14832 2654 14884
rect 3544 14875 3602 14881
rect 3544 14841 3556 14875
rect 3590 14872 3602 14875
rect 3694 14872 3700 14884
rect 3590 14844 3700 14872
rect 3590 14841 3602 14844
rect 3544 14835 3602 14841
rect 3694 14832 3700 14844
rect 3752 14832 3758 14884
rect 7558 14832 7564 14884
rect 7616 14872 7622 14884
rect 7754 14875 7812 14881
rect 7754 14872 7766 14875
rect 7616 14844 7766 14872
rect 7616 14832 7622 14844
rect 7754 14841 7766 14844
rect 7800 14841 7812 14875
rect 7852 14872 7880 14912
rect 8021 14909 8033 14943
rect 8067 14940 8079 14943
rect 8297 14943 8355 14949
rect 8297 14940 8309 14943
rect 8067 14912 8309 14940
rect 8067 14909 8079 14912
rect 8021 14903 8079 14909
rect 8297 14909 8309 14912
rect 8343 14940 8355 14943
rect 8386 14940 8392 14952
rect 8343 14912 8392 14940
rect 8343 14909 8355 14912
rect 8297 14903 8355 14909
rect 8386 14900 8392 14912
rect 8444 14940 8450 14952
rect 9490 14940 9496 14952
rect 8444 14912 9496 14940
rect 8444 14900 8450 14912
rect 9490 14900 9496 14912
rect 9548 14900 9554 14952
rect 11238 14900 11244 14952
rect 11296 14940 11302 14952
rect 11333 14943 11391 14949
rect 11333 14940 11345 14943
rect 11296 14912 11345 14940
rect 11296 14900 11302 14912
rect 11333 14909 11345 14912
rect 11379 14909 11391 14943
rect 11333 14903 11391 14909
rect 8542 14875 8600 14881
rect 8542 14872 8554 14875
rect 7852 14844 8554 14872
rect 7754 14835 7812 14841
rect 8542 14841 8554 14844
rect 8588 14841 8600 14875
rect 8542 14835 8600 14841
rect 10686 14832 10692 14884
rect 10744 14872 10750 14884
rect 11066 14875 11124 14881
rect 11066 14872 11078 14875
rect 10744 14844 11078 14872
rect 10744 14832 10750 14844
rect 11066 14841 11078 14844
rect 11112 14841 11124 14875
rect 13096 14872 13124 14971
rect 13170 14900 13176 14952
rect 13228 14940 13234 14952
rect 13348 14943 13406 14949
rect 13348 14940 13360 14943
rect 13228 14912 13360 14940
rect 13228 14900 13234 14912
rect 13348 14909 13360 14912
rect 13394 14940 13406 14943
rect 14108 14940 14136 14980
rect 15289 14977 15301 14980
rect 15335 14977 15347 15011
rect 17954 15008 17960 15020
rect 17915 14980 17960 15008
rect 15289 14971 15347 14977
rect 17954 14968 17960 14980
rect 18012 14968 18018 15020
rect 13394 14912 14136 14940
rect 18524 14940 18552 15039
rect 19058 15036 19064 15088
rect 19116 15076 19122 15088
rect 19116 15048 20392 15076
rect 19116 15036 19122 15048
rect 19242 14968 19248 15020
rect 19300 15008 19306 15020
rect 20364 15017 20392 15048
rect 19337 15011 19395 15017
rect 19337 15008 19349 15011
rect 19300 14980 19349 15008
rect 19300 14968 19306 14980
rect 19337 14977 19349 14980
rect 19383 14977 19395 15011
rect 19337 14971 19395 14977
rect 20349 15011 20407 15017
rect 20349 14977 20361 15011
rect 20395 14977 20407 15011
rect 20349 14971 20407 14977
rect 20165 14943 20223 14949
rect 20165 14940 20177 14943
rect 18524 14912 20177 14940
rect 13394 14909 13406 14912
rect 13348 14903 13406 14909
rect 20165 14909 20177 14912
rect 20211 14909 20223 14943
rect 20165 14903 20223 14909
rect 13630 14872 13636 14884
rect 13096 14844 13636 14872
rect 11066 14835 11124 14841
rect 13630 14832 13636 14844
rect 13688 14832 13694 14884
rect 15105 14875 15163 14881
rect 15105 14841 15117 14875
rect 15151 14872 15163 14875
rect 15286 14872 15292 14884
rect 15151 14844 15292 14872
rect 15151 14841 15163 14844
rect 15105 14835 15163 14841
rect 15286 14832 15292 14844
rect 15344 14832 15350 14884
rect 18141 14875 18199 14881
rect 18141 14841 18153 14875
rect 18187 14872 18199 14875
rect 18187 14844 18828 14872
rect 18187 14841 18199 14844
rect 18141 14835 18199 14841
rect 1670 14804 1676 14816
rect 1631 14776 1676 14804
rect 1670 14764 1676 14776
rect 1728 14764 1734 14816
rect 2409 14807 2467 14813
rect 2409 14773 2421 14807
rect 2455 14804 2467 14807
rect 2498 14804 2504 14816
rect 2455 14776 2504 14804
rect 2455 14773 2467 14776
rect 2409 14767 2467 14773
rect 2498 14764 2504 14776
rect 2556 14764 2562 14816
rect 6454 14764 6460 14816
rect 6512 14804 6518 14816
rect 6641 14807 6699 14813
rect 6641 14804 6653 14807
rect 6512 14776 6653 14804
rect 6512 14764 6518 14776
rect 6641 14773 6653 14776
rect 6687 14773 6699 14807
rect 6641 14767 6699 14773
rect 14461 14807 14519 14813
rect 14461 14773 14473 14807
rect 14507 14804 14519 14807
rect 14550 14804 14556 14816
rect 14507 14776 14556 14804
rect 14507 14773 14519 14776
rect 14461 14767 14519 14773
rect 14550 14764 14556 14776
rect 14608 14764 14614 14816
rect 14642 14764 14648 14816
rect 14700 14804 14706 14816
rect 15197 14807 15255 14813
rect 15197 14804 15209 14807
rect 14700 14776 15209 14804
rect 14700 14764 14706 14776
rect 15197 14773 15209 14776
rect 15243 14773 15255 14807
rect 15197 14767 15255 14773
rect 15378 14764 15384 14816
rect 15436 14804 15442 14816
rect 15749 14807 15807 14813
rect 15749 14804 15761 14807
rect 15436 14776 15761 14804
rect 15436 14764 15442 14776
rect 15749 14773 15761 14776
rect 15795 14773 15807 14807
rect 15749 14767 15807 14773
rect 16574 14764 16580 14816
rect 16632 14804 16638 14816
rect 18800 14813 18828 14844
rect 20346 14832 20352 14884
rect 20404 14872 20410 14884
rect 21177 14875 21235 14881
rect 21177 14872 21189 14875
rect 20404 14844 21189 14872
rect 20404 14832 20410 14844
rect 21177 14841 21189 14844
rect 21223 14841 21235 14875
rect 21358 14872 21364 14884
rect 21319 14844 21364 14872
rect 21177 14835 21235 14841
rect 21358 14832 21364 14844
rect 21416 14832 21422 14884
rect 18049 14807 18107 14813
rect 18049 14804 18061 14807
rect 16632 14776 18061 14804
rect 16632 14764 16638 14776
rect 18049 14773 18061 14776
rect 18095 14773 18107 14807
rect 18049 14767 18107 14773
rect 18785 14807 18843 14813
rect 18785 14773 18797 14807
rect 18831 14773 18843 14807
rect 19150 14804 19156 14816
rect 19111 14776 19156 14804
rect 18785 14767 18843 14773
rect 19150 14764 19156 14776
rect 19208 14764 19214 14816
rect 19245 14807 19303 14813
rect 19245 14773 19257 14807
rect 19291 14804 19303 14807
rect 19702 14804 19708 14816
rect 19291 14776 19708 14804
rect 19291 14773 19303 14776
rect 19245 14767 19303 14773
rect 19702 14764 19708 14776
rect 19760 14764 19766 14816
rect 19794 14764 19800 14816
rect 19852 14804 19858 14816
rect 19852 14776 19897 14804
rect 19852 14764 19858 14776
rect 19978 14764 19984 14816
rect 20036 14804 20042 14816
rect 20257 14807 20315 14813
rect 20257 14804 20269 14807
rect 20036 14776 20269 14804
rect 20036 14764 20042 14776
rect 20257 14773 20269 14776
rect 20303 14773 20315 14807
rect 20257 14767 20315 14773
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 3050 14560 3056 14612
rect 3108 14600 3114 14612
rect 3145 14603 3203 14609
rect 3145 14600 3157 14603
rect 3108 14572 3157 14600
rect 3108 14560 3114 14572
rect 3145 14569 3157 14572
rect 3191 14569 3203 14603
rect 3145 14563 3203 14569
rect 3234 14560 3240 14612
rect 3292 14600 3298 14612
rect 3513 14603 3571 14609
rect 3513 14600 3525 14603
rect 3292 14572 3525 14600
rect 3292 14560 3298 14572
rect 3513 14569 3525 14572
rect 3559 14600 3571 14603
rect 3786 14600 3792 14612
rect 3559 14572 3792 14600
rect 3559 14569 3571 14572
rect 3513 14563 3571 14569
rect 3786 14560 3792 14572
rect 3844 14560 3850 14612
rect 4062 14600 4068 14612
rect 4023 14572 4068 14600
rect 4062 14560 4068 14572
rect 4120 14560 4126 14612
rect 5718 14600 5724 14612
rect 5679 14572 5724 14600
rect 5718 14560 5724 14572
rect 5776 14560 5782 14612
rect 6181 14603 6239 14609
rect 6181 14569 6193 14603
rect 6227 14600 6239 14603
rect 6733 14603 6791 14609
rect 6733 14600 6745 14603
rect 6227 14572 6745 14600
rect 6227 14569 6239 14572
rect 6181 14563 6239 14569
rect 6733 14569 6745 14572
rect 6779 14569 6791 14603
rect 6733 14563 6791 14569
rect 7745 14603 7803 14609
rect 7745 14569 7757 14603
rect 7791 14569 7803 14603
rect 7745 14563 7803 14569
rect 5442 14492 5448 14544
rect 5500 14532 5506 14544
rect 7760 14532 7788 14563
rect 8202 14560 8208 14612
rect 8260 14600 8266 14612
rect 8297 14603 8355 14609
rect 8297 14600 8309 14603
rect 8260 14572 8309 14600
rect 8260 14560 8266 14572
rect 8297 14569 8309 14572
rect 8343 14600 8355 14603
rect 8343 14572 9812 14600
rect 8343 14569 8355 14572
rect 8297 14563 8355 14569
rect 5500 14504 7788 14532
rect 5500 14492 5506 14504
rect 9674 14492 9680 14544
rect 9732 14532 9738 14544
rect 9784 14532 9812 14572
rect 9858 14560 9864 14612
rect 9916 14600 9922 14612
rect 10686 14600 10692 14612
rect 9916 14572 10692 14600
rect 9916 14560 9922 14572
rect 10686 14560 10692 14572
rect 10744 14560 10750 14612
rect 12066 14600 12072 14612
rect 11716 14572 12072 14600
rect 11716 14532 11744 14572
rect 12066 14560 12072 14572
rect 12124 14560 12130 14612
rect 13170 14600 13176 14612
rect 13131 14572 13176 14600
rect 13170 14560 13176 14572
rect 13228 14560 13234 14612
rect 13630 14600 13636 14612
rect 13591 14572 13636 14600
rect 13630 14560 13636 14572
rect 13688 14560 13694 14612
rect 15286 14600 15292 14612
rect 15247 14572 15292 14600
rect 15286 14560 15292 14572
rect 15344 14560 15350 14612
rect 17954 14560 17960 14612
rect 18012 14600 18018 14612
rect 18601 14603 18659 14609
rect 18601 14600 18613 14603
rect 18012 14572 18613 14600
rect 18012 14560 18018 14572
rect 18601 14569 18613 14572
rect 18647 14569 18659 14603
rect 18601 14563 18659 14569
rect 19150 14560 19156 14612
rect 19208 14600 19214 14612
rect 19245 14603 19303 14609
rect 19245 14600 19257 14603
rect 19208 14572 19257 14600
rect 19208 14560 19214 14572
rect 19245 14569 19257 14572
rect 19291 14569 19303 14603
rect 19245 14563 19303 14569
rect 19702 14560 19708 14612
rect 19760 14600 19766 14612
rect 19797 14603 19855 14609
rect 19797 14600 19809 14603
rect 19760 14572 19809 14600
rect 19760 14560 19766 14572
rect 19797 14569 19809 14572
rect 19843 14569 19855 14603
rect 19797 14563 19855 14569
rect 12618 14532 12624 14544
rect 9732 14492 9751 14532
rect 9784 14504 11744 14532
rect 11808 14504 12624 14532
rect 1762 14464 1768 14476
rect 1723 14436 1768 14464
rect 1762 14424 1768 14436
rect 1820 14424 1826 14476
rect 2777 14467 2835 14473
rect 2777 14433 2789 14467
rect 2823 14464 2835 14467
rect 2958 14464 2964 14476
rect 2823 14436 2964 14464
rect 2823 14433 2835 14436
rect 2777 14427 2835 14433
rect 2958 14424 2964 14436
rect 3016 14424 3022 14476
rect 4338 14424 4344 14476
rect 4396 14464 4402 14476
rect 4433 14467 4491 14473
rect 4433 14464 4445 14467
rect 4396 14436 4445 14464
rect 4396 14424 4402 14436
rect 4433 14433 4445 14436
rect 4479 14433 4491 14467
rect 6086 14464 6092 14476
rect 6047 14436 6092 14464
rect 4433 14427 4491 14433
rect 6086 14424 6092 14436
rect 6144 14424 6150 14476
rect 7098 14464 7104 14476
rect 7059 14436 7104 14464
rect 7098 14424 7104 14436
rect 7156 14424 7162 14476
rect 7929 14467 7987 14473
rect 7929 14433 7941 14467
rect 7975 14464 7987 14467
rect 8478 14464 8484 14476
rect 7975 14436 8484 14464
rect 7975 14433 7987 14436
rect 7929 14427 7987 14433
rect 8478 14424 8484 14436
rect 8536 14424 8542 14476
rect 9576 14467 9634 14473
rect 9576 14433 9588 14467
rect 9622 14464 9634 14467
rect 9723 14464 9751 14492
rect 9950 14464 9956 14476
rect 9622 14436 9956 14464
rect 9622 14433 9634 14436
rect 9576 14427 9634 14433
rect 9950 14424 9956 14436
rect 10008 14424 10014 14476
rect 11808 14473 11836 14504
rect 12618 14492 12624 14504
rect 12676 14492 12682 14544
rect 14921 14535 14979 14541
rect 14921 14501 14933 14535
rect 14967 14532 14979 14535
rect 15378 14532 15384 14544
rect 14967 14504 15384 14532
rect 14967 14501 14979 14504
rect 14921 14495 14979 14501
rect 15378 14492 15384 14504
rect 15436 14492 15442 14544
rect 15838 14541 15844 14544
rect 15832 14495 15844 14541
rect 15896 14532 15902 14544
rect 19886 14532 19892 14544
rect 15896 14504 19892 14532
rect 15838 14492 15844 14495
rect 15896 14492 15902 14504
rect 19886 14492 19892 14504
rect 19944 14532 19950 14544
rect 19944 14504 20392 14532
rect 19944 14492 19950 14504
rect 11793 14467 11851 14473
rect 11793 14433 11805 14467
rect 11839 14433 11851 14467
rect 11793 14427 11851 14433
rect 11882 14424 11888 14476
rect 11940 14464 11946 14476
rect 12049 14467 12107 14473
rect 12049 14464 12061 14467
rect 11940 14436 12061 14464
rect 11940 14424 11946 14436
rect 12049 14433 12061 14436
rect 12095 14433 12107 14467
rect 13814 14464 13820 14476
rect 13775 14436 13820 14464
rect 12049 14427 12107 14433
rect 13814 14424 13820 14436
rect 13872 14424 13878 14476
rect 14826 14464 14832 14476
rect 14739 14436 14832 14464
rect 14826 14424 14832 14436
rect 14884 14464 14890 14476
rect 15470 14464 15476 14476
rect 14884 14436 15476 14464
rect 14884 14424 14890 14436
rect 15470 14424 15476 14436
rect 15528 14424 15534 14476
rect 17477 14467 17535 14473
rect 17477 14464 17489 14467
rect 16960 14436 17489 14464
rect 2498 14396 2504 14408
rect 2459 14368 2504 14396
rect 2498 14356 2504 14368
rect 2556 14356 2562 14408
rect 2685 14399 2743 14405
rect 2685 14365 2697 14399
rect 2731 14396 2743 14399
rect 3970 14396 3976 14408
rect 2731 14368 3976 14396
rect 2731 14365 2743 14368
rect 2685 14359 2743 14365
rect 3970 14356 3976 14368
rect 4028 14356 4034 14408
rect 4154 14356 4160 14408
rect 4212 14396 4218 14408
rect 4525 14399 4583 14405
rect 4525 14396 4537 14399
rect 4212 14368 4537 14396
rect 4212 14356 4218 14368
rect 4525 14365 4537 14368
rect 4571 14365 4583 14399
rect 4525 14359 4583 14365
rect 4617 14399 4675 14405
rect 4617 14365 4629 14399
rect 4663 14396 4675 14399
rect 5166 14396 5172 14408
rect 4663 14368 5172 14396
rect 4663 14365 4675 14368
rect 4617 14359 4675 14365
rect 2516 14328 2544 14356
rect 4632 14328 4660 14359
rect 5166 14356 5172 14368
rect 5224 14356 5230 14408
rect 6365 14399 6423 14405
rect 6365 14365 6377 14399
rect 6411 14396 6423 14399
rect 6546 14396 6552 14408
rect 6411 14368 6552 14396
rect 6411 14365 6423 14368
rect 6365 14359 6423 14365
rect 6546 14356 6552 14368
rect 6604 14356 6610 14408
rect 7190 14396 7196 14408
rect 7151 14368 7196 14396
rect 7190 14356 7196 14368
rect 7248 14356 7254 14408
rect 7282 14356 7288 14408
rect 7340 14396 7346 14408
rect 9309 14399 9367 14405
rect 7340 14368 7433 14396
rect 7340 14356 7346 14368
rect 9309 14365 9321 14399
rect 9355 14365 9367 14399
rect 14645 14399 14703 14405
rect 14645 14396 14657 14399
rect 9309 14359 9367 14365
rect 13556 14368 14657 14396
rect 2516 14300 4660 14328
rect 6454 14288 6460 14340
rect 6512 14328 6518 14340
rect 7300 14328 7328 14356
rect 6512 14300 7328 14328
rect 6512 14288 6518 14300
rect 1670 14260 1676 14272
rect 1631 14232 1676 14260
rect 1670 14220 1676 14232
rect 1728 14220 1734 14272
rect 9324 14260 9352 14359
rect 9490 14260 9496 14272
rect 9324 14232 9496 14260
rect 9490 14220 9496 14232
rect 9548 14260 9554 14272
rect 11146 14260 11152 14272
rect 9548 14232 11152 14260
rect 9548 14220 9554 14232
rect 11146 14220 11152 14232
rect 11204 14220 11210 14272
rect 11974 14220 11980 14272
rect 12032 14260 12038 14272
rect 13556 14260 13584 14368
rect 14645 14365 14657 14368
rect 14691 14365 14703 14399
rect 15562 14396 15568 14408
rect 15523 14368 15568 14396
rect 14645 14359 14703 14365
rect 14660 14328 14688 14359
rect 15562 14356 15568 14368
rect 15620 14356 15626 14408
rect 15378 14328 15384 14340
rect 14660 14300 15384 14328
rect 15378 14288 15384 14300
rect 15436 14288 15442 14340
rect 16960 14272 16988 14436
rect 17477 14433 17489 14436
rect 17523 14433 17535 14467
rect 17477 14427 17535 14433
rect 19610 14424 19616 14476
rect 19668 14464 19674 14476
rect 19705 14467 19763 14473
rect 19705 14464 19717 14467
rect 19668 14436 19717 14464
rect 19668 14424 19674 14436
rect 19705 14433 19717 14436
rect 19751 14464 19763 14467
rect 20165 14467 20223 14473
rect 20165 14464 20177 14467
rect 19751 14436 20177 14464
rect 19751 14433 19763 14436
rect 19705 14427 19763 14433
rect 20165 14433 20177 14436
rect 20211 14433 20223 14467
rect 20165 14427 20223 14433
rect 17126 14356 17132 14408
rect 17184 14396 17190 14408
rect 17221 14399 17279 14405
rect 17221 14396 17233 14399
rect 17184 14368 17233 14396
rect 17184 14356 17190 14368
rect 17221 14365 17233 14368
rect 17267 14365 17279 14399
rect 17221 14359 17279 14365
rect 18598 14356 18604 14408
rect 18656 14396 18662 14408
rect 20364 14405 20392 14504
rect 20806 14424 20812 14476
rect 20864 14464 20870 14476
rect 21177 14467 21235 14473
rect 21177 14464 21189 14467
rect 20864 14436 21189 14464
rect 20864 14424 20870 14436
rect 21177 14433 21189 14436
rect 21223 14433 21235 14467
rect 21177 14427 21235 14433
rect 20257 14399 20315 14405
rect 20257 14396 20269 14399
rect 18656 14368 20269 14396
rect 18656 14356 18662 14368
rect 20257 14365 20269 14368
rect 20303 14365 20315 14399
rect 20257 14359 20315 14365
rect 20349 14399 20407 14405
rect 20349 14365 20361 14399
rect 20395 14365 20407 14399
rect 20349 14359 20407 14365
rect 21361 14331 21419 14337
rect 21361 14297 21373 14331
rect 21407 14328 21419 14331
rect 21450 14328 21456 14340
rect 21407 14300 21456 14328
rect 21407 14297 21419 14300
rect 21361 14291 21419 14297
rect 21450 14288 21456 14300
rect 21508 14288 21514 14340
rect 16942 14260 16948 14272
rect 12032 14232 13584 14260
rect 16903 14232 16948 14260
rect 12032 14220 12038 14232
rect 16942 14220 16948 14232
rect 17000 14220 17006 14272
rect 17402 14220 17408 14272
rect 17460 14260 17466 14272
rect 19705 14263 19763 14269
rect 19705 14260 19717 14263
rect 17460 14232 19717 14260
rect 17460 14220 17466 14232
rect 19705 14229 19717 14232
rect 19751 14229 19763 14263
rect 19705 14223 19763 14229
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 2958 14056 2964 14068
rect 2919 14028 2964 14056
rect 2958 14016 2964 14028
rect 3016 14016 3022 14068
rect 4154 14056 4160 14068
rect 4115 14028 4160 14056
rect 4154 14016 4160 14028
rect 4212 14016 4218 14068
rect 7101 14059 7159 14065
rect 7101 14025 7113 14059
rect 7147 14056 7159 14059
rect 7190 14056 7196 14068
rect 7147 14028 7196 14056
rect 7147 14025 7159 14028
rect 7101 14019 7159 14025
rect 7190 14016 7196 14028
rect 7248 14016 7254 14068
rect 8294 14056 8300 14068
rect 8255 14028 8300 14056
rect 8294 14016 8300 14028
rect 8352 14016 8358 14068
rect 10502 14016 10508 14068
rect 10560 14056 10566 14068
rect 10686 14056 10692 14068
rect 10560 14028 10692 14056
rect 10560 14016 10566 14028
rect 10686 14016 10692 14028
rect 10744 14016 10750 14068
rect 14369 14059 14427 14065
rect 14369 14025 14381 14059
rect 14415 14056 14427 14059
rect 14734 14056 14740 14068
rect 14415 14028 14740 14056
rect 14415 14025 14427 14028
rect 14369 14019 14427 14025
rect 14734 14016 14740 14028
rect 14792 14016 14798 14068
rect 18601 14059 18659 14065
rect 18601 14025 18613 14059
rect 18647 14056 18659 14059
rect 19978 14056 19984 14068
rect 18647 14028 19984 14056
rect 18647 14025 18659 14028
rect 18601 14019 18659 14025
rect 19978 14016 19984 14028
rect 20036 14016 20042 14068
rect 20346 14056 20352 14068
rect 20307 14028 20352 14056
rect 20346 14016 20352 14028
rect 20404 14016 20410 14068
rect 20806 14056 20812 14068
rect 20767 14028 20812 14056
rect 20806 14016 20812 14028
rect 20864 14016 20870 14068
rect 1762 13948 1768 14000
rect 1820 13988 1826 14000
rect 3697 13991 3755 13997
rect 3697 13988 3709 13991
rect 1820 13960 3709 13988
rect 1820 13948 1826 13960
rect 3697 13957 3709 13960
rect 3743 13957 3755 13991
rect 9309 13991 9367 13997
rect 9309 13988 9321 13991
rect 3697 13951 3755 13957
rect 8772 13960 9321 13988
rect 2409 13923 2467 13929
rect 2409 13889 2421 13923
rect 2455 13920 2467 13923
rect 4709 13923 4767 13929
rect 4709 13920 4721 13923
rect 2455 13892 4721 13920
rect 2455 13889 2467 13892
rect 2409 13883 2467 13889
rect 3712 13864 3740 13892
rect 4709 13889 4721 13892
rect 4755 13889 4767 13923
rect 4709 13883 4767 13889
rect 5166 13880 5172 13932
rect 5224 13920 5230 13932
rect 5721 13923 5779 13929
rect 5721 13920 5733 13923
rect 5224 13892 5733 13920
rect 5224 13880 5230 13892
rect 5721 13889 5733 13892
rect 5767 13889 5779 13923
rect 5721 13883 5779 13889
rect 7558 13880 7564 13932
rect 7616 13920 7622 13932
rect 8772 13929 8800 13960
rect 9309 13957 9321 13960
rect 9355 13957 9367 13991
rect 9309 13951 9367 13957
rect 12621 13991 12679 13997
rect 12621 13957 12633 13991
rect 12667 13988 12679 13991
rect 14642 13988 14648 14000
rect 12667 13960 14648 13988
rect 12667 13957 12679 13960
rect 12621 13951 12679 13957
rect 14642 13948 14648 13960
rect 14700 13948 14706 14000
rect 18877 13991 18935 13997
rect 18877 13988 18889 13991
rect 18156 13960 18889 13988
rect 7653 13923 7711 13929
rect 7653 13920 7665 13923
rect 7616 13892 7665 13920
rect 7616 13880 7622 13892
rect 7653 13889 7665 13892
rect 7699 13889 7711 13923
rect 7653 13883 7711 13889
rect 8757 13923 8815 13929
rect 8757 13889 8769 13923
rect 8803 13889 8815 13923
rect 8757 13883 8815 13889
rect 8941 13923 8999 13929
rect 8941 13889 8953 13923
rect 8987 13920 8999 13923
rect 9766 13920 9772 13932
rect 8987 13892 9772 13920
rect 8987 13889 8999 13892
rect 8941 13883 8999 13889
rect 9766 13880 9772 13892
rect 9824 13880 9830 13932
rect 9858 13880 9864 13932
rect 9916 13920 9922 13932
rect 9916 13892 9961 13920
rect 9916 13880 9922 13892
rect 11882 13880 11888 13932
rect 11940 13920 11946 13932
rect 11977 13923 12035 13929
rect 11977 13920 11989 13923
rect 11940 13892 11989 13920
rect 11940 13880 11946 13892
rect 11977 13889 11989 13892
rect 12023 13889 12035 13923
rect 11977 13883 12035 13889
rect 13170 13880 13176 13932
rect 13228 13920 13234 13932
rect 13725 13923 13783 13929
rect 13725 13920 13737 13923
rect 13228 13892 13737 13920
rect 13228 13880 13234 13892
rect 13725 13889 13737 13892
rect 13771 13889 13783 13923
rect 13725 13883 13783 13889
rect 14737 13923 14795 13929
rect 14737 13889 14749 13923
rect 14783 13920 14795 13923
rect 14826 13920 14832 13932
rect 14783 13892 14832 13920
rect 14783 13889 14795 13892
rect 14737 13883 14795 13889
rect 14826 13880 14832 13892
rect 14884 13880 14890 13932
rect 17954 13920 17960 13932
rect 17915 13892 17960 13920
rect 17954 13880 17960 13892
rect 18012 13880 18018 13932
rect 18156 13929 18184 13960
rect 18877 13957 18889 13960
rect 18923 13957 18935 13991
rect 18877 13951 18935 13957
rect 18141 13923 18199 13929
rect 18141 13889 18153 13923
rect 18187 13889 18199 13923
rect 19242 13920 19248 13932
rect 18141 13883 18199 13889
rect 18892 13892 19248 13920
rect 18892 13864 18920 13892
rect 19242 13880 19248 13892
rect 19300 13920 19306 13932
rect 19429 13923 19487 13929
rect 19429 13920 19441 13923
rect 19300 13892 19441 13920
rect 19300 13880 19306 13892
rect 19429 13889 19441 13892
rect 19475 13889 19487 13923
rect 19429 13883 19487 13889
rect 1578 13852 1584 13864
rect 1539 13824 1584 13852
rect 1578 13812 1584 13824
rect 1636 13812 1642 13864
rect 3694 13812 3700 13864
rect 3752 13812 3758 13864
rect 3878 13852 3884 13864
rect 3839 13824 3884 13852
rect 3878 13812 3884 13824
rect 3936 13812 3942 13864
rect 5074 13812 5080 13864
rect 5132 13852 5138 13864
rect 5629 13855 5687 13861
rect 5132 13824 5304 13852
rect 5132 13812 5138 13824
rect 1762 13784 1768 13796
rect 1723 13756 1768 13784
rect 1762 13744 1768 13756
rect 1820 13744 1826 13796
rect 4525 13787 4583 13793
rect 4525 13753 4537 13787
rect 4571 13784 4583 13787
rect 5276 13784 5304 13824
rect 5629 13821 5641 13855
rect 5675 13852 5687 13855
rect 7742 13852 7748 13864
rect 5675 13824 7748 13852
rect 5675 13821 5687 13824
rect 5629 13815 5687 13821
rect 7742 13812 7748 13824
rect 7800 13812 7806 13864
rect 8202 13852 8208 13864
rect 7852 13824 8208 13852
rect 5350 13784 5356 13796
rect 4571 13756 5212 13784
rect 5276 13756 5356 13784
rect 4571 13753 4583 13756
rect 4525 13747 4583 13753
rect 2498 13716 2504 13728
rect 2459 13688 2504 13716
rect 2498 13676 2504 13688
rect 2556 13676 2562 13728
rect 2593 13719 2651 13725
rect 2593 13685 2605 13719
rect 2639 13716 2651 13719
rect 3237 13719 3295 13725
rect 3237 13716 3249 13719
rect 2639 13688 3249 13716
rect 2639 13685 2651 13688
rect 2593 13679 2651 13685
rect 3237 13685 3249 13688
rect 3283 13685 3295 13719
rect 3237 13679 3295 13685
rect 4614 13676 4620 13728
rect 4672 13716 4678 13728
rect 5184 13725 5212 13756
rect 5350 13744 5356 13756
rect 5408 13744 5414 13796
rect 7561 13787 7619 13793
rect 7561 13753 7573 13787
rect 7607 13784 7619 13787
rect 7852 13784 7880 13824
rect 8202 13812 8208 13824
rect 8260 13812 8266 13864
rect 11333 13855 11391 13861
rect 11333 13821 11345 13855
rect 11379 13852 11391 13855
rect 11790 13852 11796 13864
rect 11379 13824 11796 13852
rect 11379 13821 11391 13824
rect 11333 13815 11391 13821
rect 11790 13812 11796 13824
rect 11848 13852 11854 13864
rect 12250 13852 12256 13864
rect 11848 13824 12256 13852
rect 11848 13812 11854 13824
rect 12250 13812 12256 13824
rect 12308 13812 12314 13864
rect 13814 13812 13820 13864
rect 13872 13852 13878 13864
rect 16209 13855 16267 13861
rect 16209 13852 16221 13855
rect 13872 13824 16221 13852
rect 13872 13812 13878 13824
rect 16209 13821 16221 13824
rect 16255 13821 16267 13855
rect 16209 13815 16267 13821
rect 16850 13812 16856 13864
rect 16908 13852 16914 13864
rect 17497 13855 17555 13861
rect 17497 13852 17509 13855
rect 16908 13824 17509 13852
rect 16908 13812 16914 13824
rect 17497 13821 17509 13824
rect 17543 13852 17555 13855
rect 18598 13852 18604 13864
rect 17543 13824 18604 13852
rect 17543 13821 17555 13824
rect 17497 13815 17555 13821
rect 18598 13812 18604 13824
rect 18656 13812 18662 13864
rect 18874 13812 18880 13864
rect 18932 13812 18938 13864
rect 20162 13852 20168 13864
rect 20123 13824 20168 13852
rect 20162 13812 20168 13824
rect 20220 13812 20226 13864
rect 20622 13852 20628 13864
rect 20583 13824 20628 13852
rect 20622 13812 20628 13824
rect 20680 13812 20686 13864
rect 21174 13852 21180 13864
rect 21135 13824 21180 13852
rect 21174 13812 21180 13824
rect 21232 13812 21238 13864
rect 21358 13852 21364 13864
rect 21319 13824 21364 13852
rect 21358 13812 21364 13824
rect 21416 13812 21422 13864
rect 7607 13756 7880 13784
rect 8220 13756 9996 13784
rect 7607 13753 7619 13756
rect 7561 13747 7619 13753
rect 5169 13719 5227 13725
rect 4672 13688 4717 13716
rect 4672 13676 4678 13688
rect 5169 13685 5181 13719
rect 5215 13685 5227 13719
rect 5534 13716 5540 13728
rect 5495 13688 5540 13716
rect 5169 13679 5227 13685
rect 5534 13676 5540 13688
rect 5592 13676 5598 13728
rect 7469 13719 7527 13725
rect 7469 13685 7481 13719
rect 7515 13716 7527 13719
rect 7650 13716 7656 13728
rect 7515 13688 7656 13716
rect 7515 13685 7527 13688
rect 7469 13679 7527 13685
rect 7650 13676 7656 13688
rect 7708 13716 7714 13728
rect 8220 13716 8248 13756
rect 7708 13688 8248 13716
rect 8665 13719 8723 13725
rect 7708 13676 7714 13688
rect 8665 13685 8677 13719
rect 8711 13716 8723 13719
rect 9030 13716 9036 13728
rect 8711 13688 9036 13716
rect 8711 13685 8723 13688
rect 8665 13679 8723 13685
rect 9030 13676 9036 13688
rect 9088 13676 9094 13728
rect 9674 13716 9680 13728
rect 9635 13688 9680 13716
rect 9674 13676 9680 13688
rect 9732 13676 9738 13728
rect 9766 13676 9772 13728
rect 9824 13716 9830 13728
rect 9968 13716 9996 13756
rect 10042 13744 10048 13796
rect 10100 13784 10106 13796
rect 10100 13756 10640 13784
rect 10100 13744 10106 13756
rect 10502 13716 10508 13728
rect 9824 13688 9869 13716
rect 9968 13688 10508 13716
rect 9824 13676 9830 13688
rect 10502 13676 10508 13688
rect 10560 13676 10566 13728
rect 10612 13716 10640 13756
rect 11698 13744 11704 13796
rect 11756 13784 11762 13796
rect 14001 13787 14059 13793
rect 14001 13784 14013 13787
rect 11756 13756 14013 13784
rect 11756 13744 11762 13756
rect 14001 13753 14013 13756
rect 14047 13753 14059 13787
rect 14001 13747 14059 13753
rect 15746 13744 15752 13796
rect 15804 13784 15810 13796
rect 18782 13784 18788 13796
rect 15804 13756 18788 13784
rect 15804 13744 15810 13756
rect 18782 13744 18788 13756
rect 18840 13744 18846 13796
rect 19245 13787 19303 13793
rect 19245 13753 19257 13787
rect 19291 13784 19303 13787
rect 19794 13784 19800 13796
rect 19291 13756 19800 13784
rect 19291 13753 19303 13756
rect 19245 13747 19303 13753
rect 19794 13744 19800 13756
rect 19852 13744 19858 13796
rect 12161 13719 12219 13725
rect 12161 13716 12173 13719
rect 10612 13688 12173 13716
rect 12161 13685 12173 13688
rect 12207 13685 12219 13719
rect 13906 13716 13912 13728
rect 13867 13688 13912 13716
rect 12161 13679 12219 13685
rect 13906 13676 13912 13688
rect 13964 13676 13970 13728
rect 14458 13676 14464 13728
rect 14516 13716 14522 13728
rect 15562 13716 15568 13728
rect 14516 13688 15568 13716
rect 14516 13676 14522 13688
rect 15562 13676 15568 13688
rect 15620 13716 15626 13728
rect 16393 13719 16451 13725
rect 16393 13716 16405 13719
rect 15620 13688 16405 13716
rect 15620 13676 15626 13688
rect 16393 13685 16405 13688
rect 16439 13716 16451 13719
rect 17126 13716 17132 13728
rect 16439 13688 17132 13716
rect 16439 13685 16451 13688
rect 16393 13679 16451 13685
rect 17126 13676 17132 13688
rect 17184 13676 17190 13728
rect 18230 13716 18236 13728
rect 18191 13688 18236 13716
rect 18230 13676 18236 13688
rect 18288 13676 18294 13728
rect 19334 13676 19340 13728
rect 19392 13716 19398 13728
rect 19392 13688 19437 13716
rect 19392 13676 19398 13688
rect 19518 13676 19524 13728
rect 19576 13716 19582 13728
rect 20254 13716 20260 13728
rect 19576 13688 20260 13716
rect 19576 13676 19582 13688
rect 20254 13676 20260 13688
rect 20312 13676 20318 13728
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 2409 13515 2467 13521
rect 2409 13481 2421 13515
rect 2455 13512 2467 13515
rect 2498 13512 2504 13524
rect 2455 13484 2504 13512
rect 2455 13481 2467 13484
rect 2409 13475 2467 13481
rect 2498 13472 2504 13484
rect 2556 13472 2562 13524
rect 2869 13515 2927 13521
rect 2869 13481 2881 13515
rect 2915 13512 2927 13515
rect 3234 13512 3240 13524
rect 2915 13484 3240 13512
rect 2915 13481 2927 13484
rect 2869 13475 2927 13481
rect 3234 13472 3240 13484
rect 3292 13512 3298 13524
rect 3510 13512 3516 13524
rect 3292 13484 3516 13512
rect 3292 13472 3298 13484
rect 3510 13472 3516 13484
rect 3568 13472 3574 13524
rect 3878 13472 3884 13524
rect 3936 13512 3942 13524
rect 4065 13515 4123 13521
rect 4065 13512 4077 13515
rect 3936 13484 4077 13512
rect 3936 13472 3942 13484
rect 4065 13481 4077 13484
rect 4111 13481 4123 13515
rect 4065 13475 4123 13481
rect 4614 13472 4620 13524
rect 4672 13512 4678 13524
rect 4801 13515 4859 13521
rect 4801 13512 4813 13515
rect 4672 13484 4813 13512
rect 4672 13472 4678 13484
rect 4801 13481 4813 13484
rect 4847 13481 4859 13515
rect 5258 13512 5264 13524
rect 5219 13484 5264 13512
rect 4801 13475 4859 13481
rect 5258 13472 5264 13484
rect 5316 13472 5322 13524
rect 5813 13515 5871 13521
rect 5813 13481 5825 13515
rect 5859 13512 5871 13515
rect 6086 13512 6092 13524
rect 5859 13484 6092 13512
rect 5859 13481 5871 13484
rect 5813 13475 5871 13481
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 6181 13515 6239 13521
rect 6181 13481 6193 13515
rect 6227 13512 6239 13515
rect 6825 13515 6883 13521
rect 6825 13512 6837 13515
rect 6227 13484 6837 13512
rect 6227 13481 6239 13484
rect 6181 13475 6239 13481
rect 6825 13481 6837 13484
rect 6871 13481 6883 13515
rect 6825 13475 6883 13481
rect 7650 13472 7656 13524
rect 7708 13512 7714 13524
rect 7929 13515 7987 13521
rect 7929 13512 7941 13515
rect 7708 13484 7941 13512
rect 7708 13472 7714 13484
rect 7929 13481 7941 13484
rect 7975 13481 7987 13515
rect 7929 13475 7987 13481
rect 8478 13472 8484 13524
rect 8536 13512 8542 13524
rect 8757 13515 8815 13521
rect 8757 13512 8769 13515
rect 8536 13484 8769 13512
rect 8536 13472 8542 13484
rect 8757 13481 8769 13484
rect 8803 13481 8815 13515
rect 8757 13475 8815 13481
rect 9677 13515 9735 13521
rect 9677 13481 9689 13515
rect 9723 13512 9735 13515
rect 9766 13512 9772 13524
rect 9723 13484 9772 13512
rect 9723 13481 9735 13484
rect 9677 13475 9735 13481
rect 9766 13472 9772 13484
rect 9824 13472 9830 13524
rect 11698 13512 11704 13524
rect 11659 13484 11704 13512
rect 11698 13472 11704 13484
rect 11756 13472 11762 13524
rect 13906 13472 13912 13524
rect 13964 13512 13970 13524
rect 14829 13515 14887 13521
rect 14829 13512 14841 13515
rect 13964 13484 14841 13512
rect 13964 13472 13970 13484
rect 14829 13481 14841 13484
rect 14875 13481 14887 13515
rect 16574 13512 16580 13524
rect 16535 13484 16580 13512
rect 14829 13475 14887 13481
rect 16574 13472 16580 13484
rect 16632 13472 16638 13524
rect 17494 13472 17500 13524
rect 17552 13512 17558 13524
rect 19245 13515 19303 13521
rect 17552 13484 19196 13512
rect 17552 13472 17558 13484
rect 2777 13447 2835 13453
rect 2777 13413 2789 13447
rect 2823 13444 2835 13447
rect 4154 13444 4160 13456
rect 2823 13416 4160 13444
rect 2823 13413 2835 13416
rect 2777 13407 2835 13413
rect 4154 13404 4160 13416
rect 4212 13444 4218 13456
rect 5074 13444 5080 13456
rect 4212 13416 5080 13444
rect 4212 13404 4218 13416
rect 5074 13404 5080 13416
rect 5132 13404 5138 13456
rect 5169 13447 5227 13453
rect 5169 13413 5181 13447
rect 5215 13444 5227 13447
rect 5350 13444 5356 13456
rect 5215 13416 5356 13444
rect 5215 13413 5227 13416
rect 5169 13407 5227 13413
rect 5350 13404 5356 13416
rect 5408 13444 5414 13456
rect 5408 13416 7696 13444
rect 5408 13404 5414 13416
rect 1765 13379 1823 13385
rect 1765 13345 1777 13379
rect 1811 13376 1823 13379
rect 2130 13376 2136 13388
rect 1811 13348 2136 13376
rect 1811 13345 1823 13348
rect 1765 13339 1823 13345
rect 2130 13336 2136 13348
rect 2188 13336 2194 13388
rect 4246 13376 4252 13388
rect 4207 13348 4252 13376
rect 4246 13336 4252 13348
rect 4304 13336 4310 13388
rect 6273 13379 6331 13385
rect 6273 13345 6285 13379
rect 6319 13376 6331 13379
rect 7006 13376 7012 13388
rect 6319 13348 7012 13376
rect 6319 13345 6331 13348
rect 6273 13339 6331 13345
rect 7006 13336 7012 13348
rect 7064 13336 7070 13388
rect 7190 13376 7196 13388
rect 7151 13348 7196 13376
rect 7190 13336 7196 13348
rect 7248 13336 7254 13388
rect 3053 13311 3111 13317
rect 3053 13277 3065 13311
rect 3099 13277 3111 13311
rect 3053 13271 3111 13277
rect 5353 13311 5411 13317
rect 5353 13277 5365 13311
rect 5399 13277 5411 13311
rect 6454 13308 6460 13320
rect 6415 13280 6460 13308
rect 5353 13271 5411 13277
rect 1578 13240 1584 13252
rect 1539 13212 1584 13240
rect 1578 13200 1584 13212
rect 1636 13200 1642 13252
rect 3068 13240 3096 13271
rect 4154 13240 4160 13252
rect 3068 13212 4160 13240
rect 4154 13200 4160 13212
rect 4212 13240 4218 13252
rect 5166 13240 5172 13252
rect 4212 13212 5172 13240
rect 4212 13200 4218 13212
rect 5166 13200 5172 13212
rect 5224 13240 5230 13252
rect 5368 13240 5396 13271
rect 6454 13268 6460 13280
rect 6512 13268 6518 13320
rect 7282 13308 7288 13320
rect 7243 13280 7288 13308
rect 7282 13268 7288 13280
rect 7340 13268 7346 13320
rect 7469 13311 7527 13317
rect 7469 13277 7481 13311
rect 7515 13308 7527 13311
rect 7558 13308 7564 13320
rect 7515 13280 7564 13308
rect 7515 13277 7527 13280
rect 7469 13271 7527 13277
rect 7558 13268 7564 13280
rect 7616 13268 7622 13320
rect 7668 13308 7696 13416
rect 7742 13404 7748 13456
rect 7800 13444 7806 13456
rect 10226 13444 10232 13456
rect 7800 13416 10232 13444
rect 7800 13404 7806 13416
rect 10226 13404 10232 13416
rect 10284 13404 10290 13456
rect 10962 13404 10968 13456
rect 11020 13444 11026 13456
rect 11241 13447 11299 13453
rect 11241 13444 11253 13447
rect 11020 13416 11253 13444
rect 11020 13404 11026 13416
rect 11241 13413 11253 13416
rect 11287 13413 11299 13447
rect 16942 13444 16948 13456
rect 11241 13407 11299 13413
rect 16040 13416 16948 13444
rect 8570 13376 8576 13388
rect 8531 13348 8576 13376
rect 8570 13336 8576 13348
rect 8628 13336 8634 13388
rect 9766 13336 9772 13388
rect 9824 13376 9830 13388
rect 10045 13379 10103 13385
rect 10045 13376 10057 13379
rect 9824 13348 10057 13376
rect 9824 13336 9830 13348
rect 10045 13345 10057 13348
rect 10091 13345 10103 13379
rect 10045 13339 10103 13345
rect 10137 13379 10195 13385
rect 10137 13345 10149 13379
rect 10183 13376 10195 13379
rect 10686 13376 10692 13388
rect 10183 13348 10692 13376
rect 10183 13345 10195 13348
rect 10137 13339 10195 13345
rect 10686 13336 10692 13348
rect 10744 13336 10750 13388
rect 11333 13379 11391 13385
rect 11333 13376 11345 13379
rect 10980 13348 11345 13376
rect 10226 13308 10232 13320
rect 7668 13280 10232 13308
rect 10226 13268 10232 13280
rect 10284 13268 10290 13320
rect 10321 13311 10379 13317
rect 10321 13277 10333 13311
rect 10367 13277 10379 13311
rect 10321 13271 10379 13277
rect 5224 13212 5396 13240
rect 5224 13200 5230 13212
rect 9950 13200 9956 13252
rect 10008 13240 10014 13252
rect 10336 13240 10364 13271
rect 10980 13240 11008 13348
rect 11333 13345 11345 13348
rect 11379 13345 11391 13379
rect 11333 13339 11391 13345
rect 12437 13379 12495 13385
rect 12437 13345 12449 13379
rect 12483 13376 12495 13379
rect 12802 13376 12808 13388
rect 12483 13348 12808 13376
rect 12483 13345 12495 13348
rect 12437 13339 12495 13345
rect 12802 13336 12808 13348
rect 12860 13336 12866 13388
rect 15194 13376 15200 13388
rect 15155 13348 15200 13376
rect 15194 13336 15200 13348
rect 15252 13336 15258 13388
rect 11149 13311 11207 13317
rect 11149 13277 11161 13311
rect 11195 13277 11207 13311
rect 11149 13271 11207 13277
rect 12253 13311 12311 13317
rect 12253 13277 12265 13311
rect 12299 13277 12311 13311
rect 12253 13271 12311 13277
rect 12345 13311 12403 13317
rect 12345 13277 12357 13311
rect 12391 13308 12403 13311
rect 12618 13308 12624 13320
rect 12391 13280 12624 13308
rect 12391 13277 12403 13280
rect 12345 13271 12403 13277
rect 10008 13212 10364 13240
rect 10428 13212 11008 13240
rect 11164 13240 11192 13271
rect 11882 13240 11888 13252
rect 11164 13212 11888 13240
rect 10008 13200 10014 13212
rect 3418 13172 3424 13184
rect 3379 13144 3424 13172
rect 3418 13132 3424 13144
rect 3476 13132 3482 13184
rect 5534 13132 5540 13184
rect 5592 13172 5598 13184
rect 7466 13172 7472 13184
rect 5592 13144 7472 13172
rect 5592 13132 5598 13144
rect 7466 13132 7472 13144
rect 7524 13172 7530 13184
rect 10428 13172 10456 13212
rect 11882 13200 11888 13212
rect 11940 13200 11946 13252
rect 12268 13240 12296 13271
rect 12618 13268 12624 13280
rect 12676 13268 12682 13320
rect 15289 13311 15347 13317
rect 15289 13277 15301 13311
rect 15335 13277 15347 13311
rect 15289 13271 15347 13277
rect 12434 13240 12440 13252
rect 12268 13212 12440 13240
rect 12434 13200 12440 13212
rect 12492 13200 12498 13252
rect 15304 13240 15332 13271
rect 15378 13268 15384 13320
rect 15436 13308 15442 13320
rect 16040 13317 16068 13416
rect 16942 13404 16948 13416
rect 17000 13444 17006 13456
rect 18874 13444 18880 13456
rect 17000 13416 18880 13444
rect 17000 13404 17006 13416
rect 18874 13404 18880 13416
rect 18932 13404 18938 13456
rect 16206 13376 16212 13388
rect 16167 13348 16212 13376
rect 16206 13336 16212 13348
rect 16264 13336 16270 13388
rect 16298 13336 16304 13388
rect 16356 13376 16362 13388
rect 16758 13376 16764 13388
rect 16356 13348 16764 13376
rect 16356 13336 16362 13348
rect 16758 13336 16764 13348
rect 16816 13376 16822 13388
rect 17497 13379 17555 13385
rect 17497 13376 17509 13379
rect 16816 13348 17509 13376
rect 16816 13336 16822 13348
rect 17497 13345 17509 13348
rect 17543 13345 17555 13379
rect 17497 13339 17555 13345
rect 18601 13379 18659 13385
rect 18601 13345 18613 13379
rect 18647 13345 18659 13379
rect 19058 13376 19064 13388
rect 19019 13348 19064 13376
rect 18601 13339 18659 13345
rect 16025 13311 16083 13317
rect 15436 13280 15481 13308
rect 15436 13268 15442 13280
rect 16025 13277 16037 13311
rect 16071 13277 16083 13311
rect 16025 13271 16083 13277
rect 16117 13311 16175 13317
rect 16117 13277 16129 13311
rect 16163 13308 16175 13311
rect 16390 13308 16396 13320
rect 16163 13280 16396 13308
rect 16163 13277 16175 13280
rect 16117 13271 16175 13277
rect 16390 13268 16396 13280
rect 16448 13268 16454 13320
rect 16942 13268 16948 13320
rect 17000 13308 17006 13320
rect 17218 13308 17224 13320
rect 17000 13280 17224 13308
rect 17000 13268 17006 13280
rect 17218 13268 17224 13280
rect 17276 13268 17282 13320
rect 18616 13308 18644 13339
rect 19058 13336 19064 13348
rect 19116 13336 19122 13388
rect 19168 13376 19196 13484
rect 19245 13481 19257 13515
rect 19291 13481 19303 13515
rect 19245 13475 19303 13481
rect 19260 13444 19288 13475
rect 19334 13472 19340 13524
rect 19392 13512 19398 13524
rect 19797 13515 19855 13521
rect 19797 13512 19809 13515
rect 19392 13484 19809 13512
rect 19392 13472 19398 13484
rect 19797 13481 19809 13484
rect 19843 13481 19855 13515
rect 20254 13512 20260 13524
rect 20215 13484 20260 13512
rect 19797 13475 19855 13481
rect 20254 13472 20260 13484
rect 20312 13472 20318 13524
rect 20622 13444 20628 13456
rect 19260 13416 20628 13444
rect 20622 13404 20628 13416
rect 20680 13404 20686 13456
rect 20165 13379 20223 13385
rect 20165 13376 20177 13379
rect 19168 13348 20177 13376
rect 20165 13345 20177 13348
rect 20211 13345 20223 13379
rect 21269 13379 21327 13385
rect 21269 13376 21281 13379
rect 20165 13339 20223 13345
rect 20272 13348 21281 13376
rect 19702 13308 19708 13320
rect 18616 13280 19708 13308
rect 19702 13268 19708 13280
rect 19760 13268 19766 13320
rect 17494 13240 17500 13252
rect 12728 13212 14412 13240
rect 15304 13212 17500 13240
rect 7524 13144 10456 13172
rect 7524 13132 7530 13144
rect 10502 13132 10508 13184
rect 10560 13172 10566 13184
rect 12728 13172 12756 13212
rect 10560 13144 12756 13172
rect 12805 13175 12863 13181
rect 10560 13132 10566 13144
rect 12805 13141 12817 13175
rect 12851 13172 12863 13175
rect 14274 13172 14280 13184
rect 12851 13144 14280 13172
rect 12851 13141 12863 13144
rect 12805 13135 12863 13141
rect 14274 13132 14280 13144
rect 14332 13132 14338 13184
rect 14384 13172 14412 13212
rect 17494 13200 17500 13212
rect 17552 13200 17558 13252
rect 17957 13243 18015 13249
rect 17957 13209 17969 13243
rect 18003 13240 18015 13243
rect 18785 13243 18843 13249
rect 18003 13212 18736 13240
rect 18003 13209 18015 13212
rect 17957 13203 18015 13209
rect 16574 13172 16580 13184
rect 14384 13144 16580 13172
rect 16574 13132 16580 13144
rect 16632 13132 16638 13184
rect 18325 13175 18383 13181
rect 18325 13141 18337 13175
rect 18371 13172 18383 13175
rect 18598 13172 18604 13184
rect 18371 13144 18604 13172
rect 18371 13141 18383 13144
rect 18325 13135 18383 13141
rect 18598 13132 18604 13144
rect 18656 13132 18662 13184
rect 18708 13172 18736 13212
rect 18785 13209 18797 13243
rect 18831 13240 18843 13243
rect 20162 13240 20168 13252
rect 18831 13212 20168 13240
rect 18831 13209 18843 13212
rect 18785 13203 18843 13209
rect 20162 13200 20168 13212
rect 20220 13200 20226 13252
rect 20272 13172 20300 13348
rect 21269 13345 21281 13348
rect 21315 13376 21327 13379
rect 22005 13379 22063 13385
rect 22005 13376 22017 13379
rect 21315 13348 22017 13376
rect 21315 13345 21327 13348
rect 21269 13339 21327 13345
rect 22005 13345 22017 13348
rect 22051 13345 22063 13379
rect 22005 13339 22063 13345
rect 20441 13311 20499 13317
rect 20441 13277 20453 13311
rect 20487 13277 20499 13311
rect 20441 13271 20499 13277
rect 20346 13200 20352 13252
rect 20404 13240 20410 13252
rect 20456 13240 20484 13271
rect 21082 13240 21088 13252
rect 20404 13212 20484 13240
rect 21043 13212 21088 13240
rect 20404 13200 20410 13212
rect 21082 13200 21088 13212
rect 21140 13200 21146 13252
rect 18708 13144 20300 13172
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 1762 12928 1768 12980
rect 1820 12968 1826 12980
rect 2133 12971 2191 12977
rect 2133 12968 2145 12971
rect 1820 12940 2145 12968
rect 1820 12928 1826 12940
rect 2133 12937 2145 12940
rect 2179 12937 2191 12971
rect 2590 12968 2596 12980
rect 2551 12940 2596 12968
rect 2133 12931 2191 12937
rect 2590 12928 2596 12940
rect 2648 12928 2654 12980
rect 4338 12968 4344 12980
rect 4299 12940 4344 12968
rect 4338 12928 4344 12940
rect 4396 12928 4402 12980
rect 5258 12928 5264 12980
rect 5316 12968 5322 12980
rect 5997 12971 6055 12977
rect 5997 12968 6009 12971
rect 5316 12940 6009 12968
rect 5316 12928 5322 12940
rect 5997 12937 6009 12940
rect 6043 12937 6055 12971
rect 5997 12931 6055 12937
rect 7098 12928 7104 12980
rect 7156 12968 7162 12980
rect 7377 12971 7435 12977
rect 7377 12968 7389 12971
rect 7156 12940 7389 12968
rect 7156 12928 7162 12940
rect 7377 12937 7389 12940
rect 7423 12937 7435 12971
rect 9030 12968 9036 12980
rect 8991 12940 9036 12968
rect 7377 12931 7435 12937
rect 9030 12928 9036 12940
rect 9088 12928 9094 12980
rect 9766 12928 9772 12980
rect 9824 12968 9830 12980
rect 10134 12968 10140 12980
rect 9824 12940 10140 12968
rect 9824 12928 9830 12940
rect 10134 12928 10140 12940
rect 10192 12968 10198 12980
rect 10597 12971 10655 12977
rect 10597 12968 10609 12971
rect 10192 12940 10609 12968
rect 10192 12928 10198 12940
rect 10597 12937 10609 12940
rect 10643 12968 10655 12971
rect 10643 12940 13768 12968
rect 10643 12937 10655 12940
rect 10597 12931 10655 12937
rect 1581 12903 1639 12909
rect 1581 12869 1593 12903
rect 1627 12900 1639 12903
rect 10502 12900 10508 12912
rect 1627 12872 10508 12900
rect 1627 12869 1639 12872
rect 1581 12863 1639 12869
rect 10502 12860 10508 12872
rect 10560 12860 10566 12912
rect 13740 12900 13768 12940
rect 13814 12928 13820 12980
rect 13872 12968 13878 12980
rect 14737 12971 14795 12977
rect 14737 12968 14749 12971
rect 13872 12940 14749 12968
rect 13872 12928 13878 12940
rect 14737 12937 14749 12940
rect 14783 12937 14795 12971
rect 14737 12931 14795 12937
rect 15381 12971 15439 12977
rect 15381 12937 15393 12971
rect 15427 12968 15439 12971
rect 15654 12968 15660 12980
rect 15427 12940 15660 12968
rect 15427 12937 15439 12940
rect 15381 12931 15439 12937
rect 15654 12928 15660 12940
rect 15712 12928 15718 12980
rect 16390 12968 16396 12980
rect 16351 12940 16396 12968
rect 16390 12928 16396 12940
rect 16448 12928 16454 12980
rect 18138 12928 18144 12980
rect 18196 12968 18202 12980
rect 18325 12971 18383 12977
rect 18325 12968 18337 12971
rect 18196 12940 18337 12968
rect 18196 12928 18202 12940
rect 18325 12937 18337 12940
rect 18371 12937 18383 12971
rect 18325 12931 18383 12937
rect 16022 12900 16028 12912
rect 13740 12872 16028 12900
rect 16022 12860 16028 12872
rect 16080 12860 16086 12912
rect 18049 12903 18107 12909
rect 18049 12869 18061 12903
rect 18095 12900 18107 12903
rect 20898 12900 20904 12912
rect 18095 12872 20904 12900
rect 18095 12869 18107 12872
rect 18049 12863 18107 12869
rect 20898 12860 20904 12872
rect 20956 12860 20962 12912
rect 20990 12860 20996 12912
rect 21048 12900 21054 12912
rect 21085 12903 21143 12909
rect 21085 12900 21097 12903
rect 21048 12872 21097 12900
rect 21048 12860 21054 12872
rect 21085 12869 21097 12872
rect 21131 12869 21143 12903
rect 21085 12863 21143 12869
rect 3418 12832 3424 12844
rect 1412 12804 3424 12832
rect 1412 12776 1440 12804
rect 3418 12792 3424 12804
rect 3476 12792 3482 12844
rect 3694 12832 3700 12844
rect 3655 12804 3700 12832
rect 3694 12792 3700 12804
rect 3752 12792 3758 12844
rect 5166 12832 5172 12844
rect 5127 12804 5172 12832
rect 5166 12792 5172 12804
rect 5224 12832 5230 12844
rect 5442 12832 5448 12844
rect 5224 12804 5448 12832
rect 5224 12792 5230 12804
rect 5442 12792 5448 12804
rect 5500 12792 5506 12844
rect 7558 12792 7564 12844
rect 7616 12832 7622 12844
rect 7929 12835 7987 12841
rect 7929 12832 7941 12835
rect 7616 12804 7941 12832
rect 7616 12792 7622 12804
rect 7929 12801 7941 12804
rect 7975 12801 7987 12835
rect 7929 12795 7987 12801
rect 8297 12835 8355 12841
rect 8297 12801 8309 12835
rect 8343 12832 8355 12835
rect 8481 12835 8539 12841
rect 8481 12832 8493 12835
rect 8343 12804 8493 12832
rect 8343 12801 8355 12804
rect 8297 12795 8355 12801
rect 8481 12801 8493 12804
rect 8527 12832 8539 12835
rect 9030 12832 9036 12844
rect 8527 12804 9036 12832
rect 8527 12801 8539 12804
rect 8481 12795 8539 12801
rect 9030 12792 9036 12804
rect 9088 12792 9094 12844
rect 9677 12835 9735 12841
rect 9677 12801 9689 12835
rect 9723 12832 9735 12835
rect 9858 12832 9864 12844
rect 9723 12804 9864 12832
rect 9723 12801 9735 12804
rect 9677 12795 9735 12801
rect 9858 12792 9864 12804
rect 9916 12792 9922 12844
rect 10686 12792 10692 12844
rect 10744 12832 10750 12844
rect 12710 12832 12716 12844
rect 10744 12804 12716 12832
rect 10744 12792 10750 12804
rect 12710 12792 12716 12804
rect 12768 12792 12774 12844
rect 15838 12832 15844 12844
rect 15799 12804 15844 12832
rect 15838 12792 15844 12804
rect 15896 12792 15902 12844
rect 17589 12835 17647 12841
rect 17589 12801 17601 12835
rect 17635 12832 17647 12835
rect 17635 12804 18828 12832
rect 17635 12801 17647 12804
rect 17589 12795 17647 12801
rect 1394 12764 1400 12776
rect 1355 12736 1400 12764
rect 1394 12724 1400 12736
rect 1452 12724 1458 12776
rect 2317 12767 2375 12773
rect 2317 12733 2329 12767
rect 2363 12733 2375 12767
rect 2317 12727 2375 12733
rect 2777 12767 2835 12773
rect 2777 12733 2789 12767
rect 2823 12764 2835 12767
rect 4430 12764 4436 12776
rect 2823 12736 4436 12764
rect 2823 12733 2835 12736
rect 2777 12727 2835 12733
rect 2332 12696 2360 12727
rect 4430 12724 4436 12736
rect 4488 12724 4494 12776
rect 5350 12724 5356 12776
rect 5408 12764 5414 12776
rect 5629 12767 5687 12773
rect 5629 12764 5641 12767
rect 5408 12736 5641 12764
rect 5408 12724 5414 12736
rect 5629 12733 5641 12736
rect 5675 12733 5687 12767
rect 5629 12727 5687 12733
rect 7837 12767 7895 12773
rect 7837 12733 7849 12767
rect 7883 12764 7895 12767
rect 8202 12764 8208 12776
rect 7883 12736 8208 12764
rect 7883 12733 7895 12736
rect 7837 12727 7895 12733
rect 8202 12724 8208 12736
rect 8260 12764 8266 12776
rect 8260 12736 10640 12764
rect 8260 12724 8266 12736
rect 2958 12696 2964 12708
rect 2332 12668 2964 12696
rect 2958 12656 2964 12668
rect 3016 12656 3022 12708
rect 3881 12699 3939 12705
rect 3881 12665 3893 12699
rect 3927 12696 3939 12699
rect 5077 12699 5135 12705
rect 3927 12668 4660 12696
rect 3927 12665 3939 12668
rect 3881 12659 3939 12665
rect 3050 12628 3056 12640
rect 3011 12600 3056 12628
rect 3050 12588 3056 12600
rect 3108 12588 3114 12640
rect 3973 12631 4031 12637
rect 3973 12597 3985 12631
rect 4019 12628 4031 12631
rect 4522 12628 4528 12640
rect 4019 12600 4528 12628
rect 4019 12597 4031 12600
rect 3973 12591 4031 12597
rect 4522 12588 4528 12600
rect 4580 12588 4586 12640
rect 4632 12637 4660 12668
rect 5077 12665 5089 12699
rect 5123 12696 5135 12699
rect 7098 12696 7104 12708
rect 5123 12668 7104 12696
rect 5123 12665 5135 12668
rect 5077 12659 5135 12665
rect 7098 12656 7104 12668
rect 7156 12656 7162 12708
rect 7745 12699 7803 12705
rect 7745 12665 7757 12699
rect 7791 12696 7803 12699
rect 8297 12699 8355 12705
rect 8297 12696 8309 12699
rect 7791 12668 8309 12696
rect 7791 12665 7803 12668
rect 7745 12659 7803 12665
rect 8297 12665 8309 12668
rect 8343 12665 8355 12699
rect 8297 12659 8355 12665
rect 8386 12656 8392 12708
rect 8444 12696 8450 12708
rect 10042 12696 10048 12708
rect 8444 12668 10048 12696
rect 8444 12656 8450 12668
rect 10042 12656 10048 12668
rect 10100 12656 10106 12708
rect 4617 12631 4675 12637
rect 4617 12597 4629 12631
rect 4663 12597 4675 12631
rect 4982 12628 4988 12640
rect 4943 12600 4988 12628
rect 4617 12591 4675 12597
rect 4982 12588 4988 12600
rect 5040 12588 5046 12640
rect 9398 12628 9404 12640
rect 9359 12600 9404 12628
rect 9398 12588 9404 12600
rect 9456 12588 9462 12640
rect 9490 12588 9496 12640
rect 9548 12628 9554 12640
rect 10612 12628 10640 12736
rect 12526 12724 12532 12776
rect 12584 12764 12590 12776
rect 12805 12767 12863 12773
rect 12805 12764 12817 12767
rect 12584 12736 12817 12764
rect 12584 12724 12590 12736
rect 12805 12733 12817 12736
rect 12851 12764 12863 12767
rect 13354 12764 13360 12776
rect 12851 12736 13360 12764
rect 12851 12733 12863 12736
rect 12805 12727 12863 12733
rect 13354 12724 13360 12736
rect 13412 12724 13418 12776
rect 14553 12767 14611 12773
rect 14553 12733 14565 12767
rect 14599 12764 14611 12767
rect 15194 12764 15200 12776
rect 14599 12736 15200 12764
rect 14599 12733 14611 12736
rect 14553 12727 14611 12733
rect 15194 12724 15200 12736
rect 15252 12724 15258 12776
rect 15286 12724 15292 12776
rect 15344 12764 15350 12776
rect 17221 12767 17279 12773
rect 15344 12736 17172 12764
rect 15344 12724 15350 12736
rect 12434 12656 12440 12708
rect 12492 12696 12498 12708
rect 13050 12699 13108 12705
rect 13050 12696 13062 12699
rect 12492 12668 13062 12696
rect 12492 12656 12498 12668
rect 13050 12665 13062 12668
rect 13096 12696 13108 12699
rect 13262 12696 13268 12708
rect 13096 12668 13268 12696
rect 13096 12665 13108 12668
rect 13050 12659 13108 12665
rect 13262 12656 13268 12668
rect 13320 12656 13326 12708
rect 16025 12699 16083 12705
rect 16025 12696 16037 12699
rect 14016 12668 16037 12696
rect 14016 12628 14044 12668
rect 16025 12665 16037 12668
rect 16071 12665 16083 12699
rect 17144 12696 17172 12736
rect 17221 12733 17233 12767
rect 17267 12764 17279 12767
rect 17865 12767 17923 12773
rect 17865 12764 17877 12767
rect 17267 12736 17877 12764
rect 17267 12733 17279 12736
rect 17221 12727 17279 12733
rect 17865 12733 17877 12736
rect 17911 12764 17923 12767
rect 17954 12764 17960 12776
rect 17911 12736 17960 12764
rect 17911 12733 17923 12736
rect 17865 12727 17923 12733
rect 17954 12724 17960 12736
rect 18012 12724 18018 12776
rect 18800 12764 18828 12804
rect 18874 12792 18880 12844
rect 18932 12832 18938 12844
rect 19886 12832 19892 12844
rect 18932 12804 18977 12832
rect 19847 12804 19892 12832
rect 18932 12792 18938 12804
rect 19886 12792 19892 12804
rect 19944 12832 19950 12844
rect 20346 12832 20352 12844
rect 19944 12804 20352 12832
rect 19944 12792 19950 12804
rect 20346 12792 20352 12804
rect 20404 12792 20410 12844
rect 20622 12764 20628 12776
rect 18800 12736 20628 12764
rect 20622 12724 20628 12736
rect 20680 12724 20686 12776
rect 18414 12696 18420 12708
rect 17144 12668 18420 12696
rect 16025 12659 16083 12665
rect 18414 12656 18420 12668
rect 18472 12656 18478 12708
rect 18693 12699 18751 12705
rect 18693 12665 18705 12699
rect 18739 12696 18751 12699
rect 19426 12696 19432 12708
rect 18739 12668 19432 12696
rect 18739 12665 18751 12668
rect 18693 12659 18751 12665
rect 19426 12656 19432 12668
rect 19484 12656 19490 12708
rect 19518 12656 19524 12708
rect 19576 12696 19582 12708
rect 19797 12699 19855 12705
rect 19797 12696 19809 12699
rect 19576 12668 19809 12696
rect 19576 12656 19582 12668
rect 19797 12665 19809 12668
rect 19843 12665 19855 12699
rect 21266 12696 21272 12708
rect 21227 12668 21272 12696
rect 19797 12659 19855 12665
rect 21266 12656 21272 12668
rect 21324 12656 21330 12708
rect 14182 12628 14188 12640
rect 9548 12600 9593 12628
rect 10612 12600 14044 12628
rect 14143 12600 14188 12628
rect 9548 12588 9554 12600
rect 14182 12588 14188 12600
rect 14240 12588 14246 12640
rect 15654 12588 15660 12640
rect 15712 12628 15718 12640
rect 15933 12631 15991 12637
rect 15933 12628 15945 12631
rect 15712 12600 15945 12628
rect 15712 12588 15718 12600
rect 15933 12597 15945 12600
rect 15979 12628 15991 12631
rect 16390 12628 16396 12640
rect 15979 12600 16396 12628
rect 15979 12597 15991 12600
rect 15933 12591 15991 12597
rect 16390 12588 16396 12600
rect 16448 12588 16454 12640
rect 18785 12631 18843 12637
rect 18785 12597 18797 12631
rect 18831 12628 18843 12631
rect 19337 12631 19395 12637
rect 19337 12628 19349 12631
rect 18831 12600 19349 12628
rect 18831 12597 18843 12600
rect 18785 12591 18843 12597
rect 19337 12597 19349 12600
rect 19383 12597 19395 12631
rect 19702 12628 19708 12640
rect 19663 12600 19708 12628
rect 19337 12591 19395 12597
rect 19702 12588 19708 12600
rect 19760 12588 19766 12640
rect 20714 12628 20720 12640
rect 20675 12600 20720 12628
rect 20714 12588 20720 12600
rect 20772 12588 20778 12640
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 22002 12492 22008 12504
rect 1104 12464 21896 12486
rect 21963 12464 22008 12492
rect 22002 12452 22008 12464
rect 22060 12452 22066 12504
rect 2682 12424 2688 12436
rect 2643 12396 2688 12424
rect 2682 12384 2688 12396
rect 2740 12384 2746 12436
rect 2777 12427 2835 12433
rect 2777 12393 2789 12427
rect 2823 12424 2835 12427
rect 2866 12424 2872 12436
rect 2823 12396 2872 12424
rect 2823 12393 2835 12396
rect 2777 12387 2835 12393
rect 2866 12384 2872 12396
rect 2924 12384 2930 12436
rect 3510 12384 3516 12436
rect 3568 12424 3574 12436
rect 4798 12424 4804 12436
rect 3568 12396 4804 12424
rect 3568 12384 3574 12396
rect 4798 12384 4804 12396
rect 4856 12384 4862 12436
rect 5721 12427 5779 12433
rect 5721 12424 5733 12427
rect 4908 12396 5733 12424
rect 1670 12356 1676 12368
rect 1631 12328 1676 12356
rect 1670 12316 1676 12328
rect 1728 12356 1734 12368
rect 3050 12356 3056 12368
rect 1728 12328 3056 12356
rect 1728 12316 1734 12328
rect 3050 12316 3056 12328
rect 3108 12316 3114 12368
rect 3237 12359 3295 12365
rect 3237 12325 3249 12359
rect 3283 12356 3295 12359
rect 4154 12356 4160 12368
rect 3283 12328 4160 12356
rect 3283 12325 3295 12328
rect 3237 12319 3295 12325
rect 4154 12316 4160 12328
rect 4212 12316 4218 12368
rect 4908 12356 4936 12396
rect 5721 12393 5733 12396
rect 5767 12424 5779 12427
rect 6270 12424 6276 12436
rect 5767 12396 6276 12424
rect 5767 12393 5779 12396
rect 5721 12387 5779 12393
rect 6270 12384 6276 12396
rect 6328 12384 6334 12436
rect 7006 12384 7012 12436
rect 7064 12424 7070 12436
rect 7193 12427 7251 12433
rect 7193 12424 7205 12427
rect 7064 12396 7205 12424
rect 7064 12384 7070 12396
rect 7193 12393 7205 12396
rect 7239 12393 7251 12427
rect 7193 12387 7251 12393
rect 9401 12427 9459 12433
rect 9401 12393 9413 12427
rect 9447 12424 9459 12427
rect 9490 12424 9496 12436
rect 9447 12396 9496 12424
rect 9447 12393 9459 12396
rect 9401 12387 9459 12393
rect 9490 12384 9496 12396
rect 9548 12384 9554 12436
rect 9861 12427 9919 12433
rect 9861 12393 9873 12427
rect 9907 12424 9919 12427
rect 12158 12424 12164 12436
rect 9907 12396 12164 12424
rect 9907 12393 9919 12396
rect 9861 12387 9919 12393
rect 12158 12384 12164 12396
rect 12216 12384 12222 12436
rect 12434 12384 12440 12436
rect 12492 12424 12498 12436
rect 15470 12424 15476 12436
rect 12492 12396 12537 12424
rect 14108 12396 15476 12424
rect 12492 12384 12498 12396
rect 14108 12356 14136 12396
rect 15470 12384 15476 12396
rect 15528 12384 15534 12436
rect 15838 12384 15844 12436
rect 15896 12424 15902 12436
rect 15933 12427 15991 12433
rect 15933 12424 15945 12427
rect 15896 12396 15945 12424
rect 15896 12384 15902 12396
rect 15933 12393 15945 12396
rect 15979 12393 15991 12427
rect 15933 12387 15991 12393
rect 17126 12384 17132 12436
rect 17184 12424 17190 12436
rect 17957 12427 18015 12433
rect 17957 12424 17969 12427
rect 17184 12396 17969 12424
rect 17184 12384 17190 12396
rect 17957 12393 17969 12396
rect 18003 12393 18015 12427
rect 18414 12424 18420 12436
rect 18375 12396 18420 12424
rect 17957 12387 18015 12393
rect 18414 12384 18420 12396
rect 18472 12384 18478 12436
rect 18506 12384 18512 12436
rect 18564 12424 18570 12436
rect 18966 12424 18972 12436
rect 18564 12396 18972 12424
rect 18564 12384 18570 12396
rect 18966 12384 18972 12396
rect 19024 12384 19030 12436
rect 19794 12424 19800 12436
rect 19755 12396 19800 12424
rect 19794 12384 19800 12396
rect 19852 12384 19858 12436
rect 20162 12424 20168 12436
rect 20123 12396 20168 12424
rect 20162 12384 20168 12396
rect 20220 12384 20226 12436
rect 4264 12328 4936 12356
rect 5000 12328 14136 12356
rect 1854 12248 1860 12300
rect 1912 12288 1918 12300
rect 1912 12260 2774 12288
rect 1912 12248 1918 12260
rect 2590 12220 2596 12232
rect 2551 12192 2596 12220
rect 2590 12180 2596 12192
rect 2648 12180 2654 12232
rect 2746 12220 2774 12260
rect 3510 12248 3516 12300
rect 3568 12288 3574 12300
rect 4264 12288 4292 12328
rect 3568 12260 4292 12288
rect 4341 12291 4399 12297
rect 3568 12248 3574 12260
rect 4341 12257 4353 12291
rect 4387 12288 4399 12291
rect 4430 12288 4436 12300
rect 4387 12260 4436 12288
rect 4387 12257 4399 12260
rect 4341 12251 4399 12257
rect 4430 12248 4436 12260
rect 4488 12248 4494 12300
rect 5000 12220 5028 12328
rect 14182 12316 14188 12368
rect 14240 12356 14246 12368
rect 14798 12359 14856 12365
rect 14798 12356 14810 12359
rect 14240 12328 14810 12356
rect 14240 12316 14246 12328
rect 14798 12325 14810 12328
rect 14844 12325 14856 12359
rect 14798 12319 14856 12325
rect 14918 12316 14924 12368
rect 14976 12356 14982 12368
rect 15746 12356 15752 12368
rect 14976 12328 15752 12356
rect 14976 12316 14982 12328
rect 15746 12316 15752 12328
rect 15804 12316 15810 12368
rect 17586 12316 17592 12368
rect 17644 12365 17650 12368
rect 17644 12356 17656 12365
rect 18230 12356 18236 12368
rect 17644 12328 18236 12356
rect 17644 12319 17656 12328
rect 17644 12316 17650 12319
rect 18230 12316 18236 12328
rect 18288 12316 18294 12368
rect 19245 12359 19303 12365
rect 19245 12325 19257 12359
rect 19291 12356 19303 12359
rect 19291 12328 21312 12356
rect 19291 12325 19303 12328
rect 19245 12319 19303 12325
rect 5077 12291 5135 12297
rect 5077 12257 5089 12291
rect 5123 12257 5135 12291
rect 5077 12251 5135 12257
rect 5169 12291 5227 12297
rect 5169 12257 5181 12291
rect 5215 12288 5227 12291
rect 5994 12288 6000 12300
rect 5215 12260 6000 12288
rect 5215 12257 5227 12260
rect 5169 12251 5227 12257
rect 2746 12192 5028 12220
rect 2608 12152 2636 12180
rect 3145 12155 3203 12161
rect 2608 12124 2774 12152
rect 1762 12084 1768 12096
rect 1723 12056 1768 12084
rect 1762 12044 1768 12056
rect 1820 12044 1826 12096
rect 2746 12084 2774 12124
rect 3145 12121 3157 12155
rect 3191 12152 3203 12155
rect 4338 12152 4344 12164
rect 3191 12124 4344 12152
rect 3191 12121 3203 12124
rect 3145 12115 3203 12121
rect 4338 12112 4344 12124
rect 4396 12112 4402 12164
rect 4614 12112 4620 12164
rect 4672 12152 4678 12164
rect 4709 12155 4767 12161
rect 4709 12152 4721 12155
rect 4672 12124 4721 12152
rect 4672 12112 4678 12124
rect 4709 12121 4721 12124
rect 4755 12121 4767 12155
rect 4709 12115 4767 12121
rect 4798 12112 4804 12164
rect 4856 12152 4862 12164
rect 5092 12152 5120 12251
rect 5994 12248 6000 12260
rect 6052 12288 6058 12300
rect 7561 12291 7619 12297
rect 7561 12288 7573 12291
rect 6052 12260 7573 12288
rect 6052 12248 6058 12260
rect 7561 12257 7573 12260
rect 7607 12257 7619 12291
rect 7561 12251 7619 12257
rect 7653 12291 7711 12297
rect 7653 12257 7665 12291
rect 7699 12288 7711 12291
rect 8754 12288 8760 12300
rect 7699 12260 8760 12288
rect 7699 12257 7711 12260
rect 7653 12251 7711 12257
rect 8754 12248 8760 12260
rect 8812 12248 8818 12300
rect 9769 12291 9827 12297
rect 9769 12257 9781 12291
rect 9815 12257 9827 12291
rect 9769 12251 9827 12257
rect 11057 12291 11115 12297
rect 11057 12257 11069 12291
rect 11103 12288 11115 12291
rect 11146 12288 11152 12300
rect 11103 12260 11152 12288
rect 11103 12257 11115 12260
rect 11057 12251 11115 12257
rect 5258 12180 5264 12232
rect 5316 12220 5322 12232
rect 7742 12220 7748 12232
rect 5316 12192 5361 12220
rect 7703 12192 7748 12220
rect 5316 12180 5322 12192
rect 7742 12180 7748 12192
rect 7800 12180 7806 12232
rect 9784 12220 9812 12251
rect 11146 12248 11152 12260
rect 11204 12248 11210 12300
rect 11324 12291 11382 12297
rect 11324 12257 11336 12291
rect 11370 12288 11382 12291
rect 11698 12288 11704 12300
rect 11370 12260 11704 12288
rect 11370 12257 11382 12260
rect 11324 12251 11382 12257
rect 11698 12248 11704 12260
rect 11756 12248 11762 12300
rect 11790 12248 11796 12300
rect 11848 12288 11854 12300
rect 13541 12291 13599 12297
rect 13541 12288 13553 12291
rect 11848 12260 13553 12288
rect 11848 12248 11854 12260
rect 13541 12257 13553 12260
rect 13587 12257 13599 12291
rect 18138 12288 18144 12300
rect 13541 12251 13599 12257
rect 14476 12260 18144 12288
rect 9950 12220 9956 12232
rect 7852 12192 9812 12220
rect 9911 12192 9956 12220
rect 7852 12152 7880 12192
rect 9950 12180 9956 12192
rect 10008 12180 10014 12232
rect 12894 12220 12900 12232
rect 12855 12192 12900 12220
rect 12894 12180 12900 12192
rect 12952 12180 12958 12232
rect 13262 12220 13268 12232
rect 13223 12192 13268 12220
rect 13262 12180 13268 12192
rect 13320 12180 13326 12232
rect 13449 12223 13507 12229
rect 13449 12189 13461 12223
rect 13495 12220 13507 12223
rect 14476 12220 14504 12260
rect 18138 12248 18144 12260
rect 18196 12248 18202 12300
rect 18509 12291 18567 12297
rect 18509 12257 18521 12291
rect 18555 12288 18567 12291
rect 18690 12288 18696 12300
rect 18555 12260 18696 12288
rect 18555 12257 18567 12260
rect 18509 12251 18567 12257
rect 18690 12248 18696 12260
rect 18748 12248 18754 12300
rect 18782 12248 18788 12300
rect 18840 12288 18846 12300
rect 20257 12291 20315 12297
rect 20257 12288 20269 12291
rect 18840 12260 20269 12288
rect 18840 12248 18846 12260
rect 20257 12257 20269 12260
rect 20303 12288 20315 12291
rect 20806 12288 20812 12300
rect 20303 12260 20812 12288
rect 20303 12257 20315 12260
rect 20257 12251 20315 12257
rect 20806 12248 20812 12260
rect 20864 12248 20870 12300
rect 21284 12297 21312 12328
rect 21269 12291 21327 12297
rect 21269 12257 21281 12291
rect 21315 12288 21327 12291
rect 22005 12291 22063 12297
rect 22005 12288 22017 12291
rect 21315 12260 22017 12288
rect 21315 12257 21327 12260
rect 21269 12251 21327 12257
rect 22005 12257 22017 12260
rect 22051 12257 22063 12291
rect 22005 12251 22063 12257
rect 13495 12192 14504 12220
rect 14553 12223 14611 12229
rect 13495 12189 13507 12192
rect 13449 12183 13507 12189
rect 14553 12189 14565 12223
rect 14599 12189 14611 12223
rect 14553 12183 14611 12189
rect 17865 12223 17923 12229
rect 17865 12189 17877 12223
rect 17911 12189 17923 12223
rect 18230 12220 18236 12232
rect 18191 12192 18236 12220
rect 17865 12183 17923 12189
rect 4856 12124 7880 12152
rect 4856 12112 4862 12124
rect 8754 12112 8760 12164
rect 8812 12152 8818 12164
rect 8812 12124 9720 12152
rect 8812 12112 8818 12124
rect 3237 12087 3295 12093
rect 3237 12084 3249 12087
rect 2746 12056 3249 12084
rect 3237 12053 3249 12056
rect 3283 12053 3295 12087
rect 3418 12084 3424 12096
rect 3379 12056 3424 12084
rect 3237 12047 3295 12053
rect 3418 12044 3424 12056
rect 3476 12044 3482 12096
rect 3973 12087 4031 12093
rect 3973 12053 3985 12087
rect 4019 12084 4031 12087
rect 4062 12084 4068 12096
rect 4019 12056 4068 12084
rect 4019 12053 4031 12056
rect 3973 12047 4031 12053
rect 4062 12044 4068 12056
rect 4120 12044 4126 12096
rect 7006 12044 7012 12096
rect 7064 12084 7070 12096
rect 7282 12084 7288 12096
rect 7064 12056 7288 12084
rect 7064 12044 7070 12056
rect 7282 12044 7288 12056
rect 7340 12044 7346 12096
rect 9692 12084 9720 12124
rect 13170 12112 13176 12164
rect 13228 12152 13234 12164
rect 13228 12124 14412 12152
rect 13228 12112 13234 12124
rect 11974 12084 11980 12096
rect 9692 12056 11980 12084
rect 11974 12044 11980 12056
rect 12032 12044 12038 12096
rect 13909 12087 13967 12093
rect 13909 12053 13921 12087
rect 13955 12084 13967 12087
rect 14182 12084 14188 12096
rect 13955 12056 14188 12084
rect 13955 12053 13967 12056
rect 13909 12047 13967 12053
rect 14182 12044 14188 12056
rect 14240 12044 14246 12096
rect 14384 12084 14412 12124
rect 14458 12112 14464 12164
rect 14516 12152 14522 12164
rect 14568 12152 14596 12183
rect 17880 12152 17908 12183
rect 18230 12180 18236 12192
rect 18288 12180 18294 12232
rect 19150 12180 19156 12232
rect 19208 12220 19214 12232
rect 20162 12220 20168 12232
rect 19208 12192 20168 12220
rect 19208 12180 19214 12192
rect 20162 12180 20168 12192
rect 20220 12180 20226 12232
rect 20346 12180 20352 12232
rect 20404 12220 20410 12232
rect 20404 12192 20449 12220
rect 20404 12180 20410 12192
rect 17957 12155 18015 12161
rect 17957 12152 17969 12155
rect 14516 12124 14596 12152
rect 17867 12124 17969 12152
rect 14516 12112 14522 12124
rect 17957 12121 17969 12124
rect 18003 12152 18015 12155
rect 20070 12152 20076 12164
rect 18003 12124 20076 12152
rect 18003 12121 18015 12124
rect 17957 12115 18015 12121
rect 20070 12112 20076 12124
rect 20128 12112 20134 12164
rect 14918 12084 14924 12096
rect 14384 12056 14924 12084
rect 14918 12044 14924 12056
rect 14976 12044 14982 12096
rect 15286 12044 15292 12096
rect 15344 12084 15350 12096
rect 15838 12084 15844 12096
rect 15344 12056 15844 12084
rect 15344 12044 15350 12056
rect 15838 12044 15844 12056
rect 15896 12044 15902 12096
rect 16485 12087 16543 12093
rect 16485 12053 16497 12087
rect 16531 12084 16543 12087
rect 17678 12084 17684 12096
rect 16531 12056 17684 12084
rect 16531 12053 16543 12056
rect 16485 12047 16543 12053
rect 17678 12044 17684 12056
rect 17736 12044 17742 12096
rect 18782 12044 18788 12096
rect 18840 12084 18846 12096
rect 18877 12087 18935 12093
rect 18877 12084 18889 12087
rect 18840 12056 18889 12084
rect 18840 12044 18846 12056
rect 18877 12053 18889 12056
rect 18923 12053 18935 12087
rect 18877 12047 18935 12053
rect 18966 12044 18972 12096
rect 19024 12084 19030 12096
rect 21177 12087 21235 12093
rect 21177 12084 21189 12087
rect 19024 12056 21189 12084
rect 19024 12044 19030 12056
rect 21177 12053 21189 12056
rect 21223 12053 21235 12087
rect 21177 12047 21235 12053
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 1104 11920 21896 11942
rect 1762 11840 1768 11892
rect 1820 11880 1826 11892
rect 3694 11880 3700 11892
rect 1820 11852 3556 11880
rect 3607 11852 3700 11880
rect 1820 11840 1826 11852
rect 1854 11812 1860 11824
rect 1815 11784 1860 11812
rect 1854 11772 1860 11784
rect 1912 11772 1918 11824
rect 1670 11676 1676 11688
rect 1631 11648 1676 11676
rect 1670 11636 1676 11648
rect 1728 11636 1734 11688
rect 2038 11636 2044 11688
rect 2096 11676 2102 11688
rect 2317 11679 2375 11685
rect 2317 11676 2329 11679
rect 2096 11648 2329 11676
rect 2096 11636 2102 11648
rect 2317 11645 2329 11648
rect 2363 11645 2375 11679
rect 3418 11676 3424 11688
rect 2317 11639 2375 11645
rect 2424 11648 3424 11676
rect 1688 11608 1716 11636
rect 2424 11608 2452 11648
rect 3418 11636 3424 11648
rect 3476 11636 3482 11688
rect 2590 11617 2596 11620
rect 2584 11608 2596 11617
rect 1688 11580 2452 11608
rect 2551 11580 2596 11608
rect 2584 11571 2596 11580
rect 2590 11568 2596 11571
rect 2648 11568 2654 11620
rect 3528 11608 3556 11852
rect 3694 11840 3700 11852
rect 3752 11840 3758 11892
rect 3970 11880 3976 11892
rect 3931 11852 3976 11880
rect 3970 11840 3976 11852
rect 4028 11840 4034 11892
rect 4246 11840 4252 11892
rect 4304 11880 4310 11892
rect 7006 11880 7012 11892
rect 4304 11852 7012 11880
rect 4304 11840 4310 11852
rect 7006 11840 7012 11852
rect 7064 11840 7070 11892
rect 7282 11840 7288 11892
rect 7340 11880 7346 11892
rect 7834 11880 7840 11892
rect 7340 11852 7840 11880
rect 7340 11840 7346 11852
rect 7834 11840 7840 11852
rect 7892 11840 7898 11892
rect 9217 11883 9275 11889
rect 9217 11849 9229 11883
rect 9263 11880 9275 11883
rect 9398 11880 9404 11892
rect 9263 11852 9404 11880
rect 9263 11849 9275 11852
rect 9217 11843 9275 11849
rect 9398 11840 9404 11852
rect 9456 11840 9462 11892
rect 9493 11883 9551 11889
rect 9493 11849 9505 11883
rect 9539 11880 9551 11883
rect 9674 11880 9680 11892
rect 9539 11852 9680 11880
rect 9539 11849 9551 11852
rect 9493 11843 9551 11849
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 11241 11883 11299 11889
rect 11241 11849 11253 11883
rect 11287 11880 11299 11883
rect 11790 11880 11796 11892
rect 11287 11852 11796 11880
rect 11287 11849 11299 11852
rect 11241 11843 11299 11849
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 12618 11880 12624 11892
rect 12579 11852 12624 11880
rect 12618 11840 12624 11852
rect 12676 11840 12682 11892
rect 12802 11840 12808 11892
rect 12860 11880 12866 11892
rect 12897 11883 12955 11889
rect 12897 11880 12909 11883
rect 12860 11852 12909 11880
rect 12860 11840 12866 11852
rect 12897 11849 12909 11852
rect 12943 11849 12955 11883
rect 12897 11843 12955 11849
rect 13924 11852 15424 11880
rect 3712 11812 3740 11840
rect 3712 11784 4568 11812
rect 4540 11753 4568 11784
rect 4890 11772 4896 11824
rect 4948 11812 4954 11824
rect 7742 11812 7748 11824
rect 4948 11784 7748 11812
rect 4948 11772 4954 11784
rect 7742 11772 7748 11784
rect 7800 11772 7806 11824
rect 7926 11772 7932 11824
rect 7984 11812 7990 11824
rect 13924 11812 13952 11852
rect 14090 11812 14096 11824
rect 7984 11784 13952 11812
rect 14016 11784 14096 11812
rect 7984 11772 7990 11784
rect 4525 11747 4583 11753
rect 4525 11713 4537 11747
rect 4571 11713 4583 11747
rect 4525 11707 4583 11713
rect 5077 11747 5135 11753
rect 5077 11713 5089 11747
rect 5123 11744 5135 11747
rect 5166 11744 5172 11756
rect 5123 11716 5172 11744
rect 5123 11713 5135 11716
rect 5077 11707 5135 11713
rect 5166 11704 5172 11716
rect 5224 11704 5230 11756
rect 5810 11704 5816 11756
rect 5868 11744 5874 11756
rect 7650 11744 7656 11756
rect 5868 11716 7656 11744
rect 5868 11704 5874 11716
rect 7650 11704 7656 11716
rect 7708 11704 7714 11756
rect 8665 11747 8723 11753
rect 8665 11713 8677 11747
rect 8711 11744 8723 11747
rect 9950 11744 9956 11756
rect 8711 11716 9956 11744
rect 8711 11713 8723 11716
rect 8665 11707 8723 11713
rect 9950 11704 9956 11716
rect 10008 11744 10014 11756
rect 10045 11747 10103 11753
rect 10045 11744 10057 11747
rect 10008 11716 10057 11744
rect 10008 11704 10014 11716
rect 10045 11713 10057 11716
rect 10091 11713 10103 11747
rect 10045 11707 10103 11713
rect 10689 11747 10747 11753
rect 10689 11713 10701 11747
rect 10735 11744 10747 11747
rect 11698 11744 11704 11756
rect 10735 11716 11704 11744
rect 10735 11713 10747 11716
rect 10689 11707 10747 11713
rect 11698 11704 11704 11716
rect 11756 11744 11762 11756
rect 14016 11753 14044 11784
rect 14090 11772 14096 11784
rect 14148 11772 14154 11824
rect 14645 11815 14703 11821
rect 14645 11781 14657 11815
rect 14691 11812 14703 11815
rect 14691 11784 15148 11812
rect 14691 11781 14703 11784
rect 14645 11775 14703 11781
rect 11977 11747 12035 11753
rect 11977 11744 11989 11747
rect 11756 11716 11989 11744
rect 11756 11704 11762 11716
rect 11977 11713 11989 11716
rect 12023 11744 12035 11747
rect 13541 11747 13599 11753
rect 13541 11744 13553 11747
rect 12023 11716 13553 11744
rect 12023 11713 12035 11716
rect 11977 11707 12035 11713
rect 13541 11713 13553 11716
rect 13587 11744 13599 11747
rect 14001 11747 14059 11753
rect 13587 11716 13952 11744
rect 13587 11713 13599 11716
rect 13541 11707 13599 11713
rect 4154 11636 4160 11688
rect 4212 11676 4218 11688
rect 8757 11679 8815 11685
rect 8757 11676 8769 11679
rect 4212 11648 8769 11676
rect 4212 11636 4218 11648
rect 8757 11645 8769 11648
rect 8803 11645 8815 11679
rect 8757 11639 8815 11645
rect 9858 11636 9864 11688
rect 9916 11676 9922 11688
rect 10873 11679 10931 11685
rect 10873 11676 10885 11679
rect 9916 11648 10885 11676
rect 9916 11636 9922 11648
rect 10873 11645 10885 11648
rect 10919 11645 10931 11679
rect 10873 11639 10931 11645
rect 12894 11636 12900 11688
rect 12952 11676 12958 11688
rect 13265 11679 13323 11685
rect 13265 11676 13277 11679
rect 12952 11648 13277 11676
rect 12952 11636 12958 11648
rect 13265 11645 13277 11648
rect 13311 11645 13323 11679
rect 13265 11639 13323 11645
rect 13814 11608 13820 11620
rect 3528 11580 13820 11608
rect 13814 11568 13820 11580
rect 13872 11568 13878 11620
rect 13924 11608 13952 11716
rect 14001 11713 14013 11747
rect 14047 11713 14059 11747
rect 14182 11744 14188 11756
rect 14143 11716 14188 11744
rect 14001 11707 14059 11713
rect 14182 11704 14188 11716
rect 14240 11704 14246 11756
rect 14274 11676 14280 11688
rect 14235 11648 14280 11676
rect 14274 11636 14280 11648
rect 14332 11636 14338 11688
rect 15120 11676 15148 11784
rect 15286 11744 15292 11756
rect 15247 11716 15292 11744
rect 15286 11704 15292 11716
rect 15344 11704 15350 11756
rect 15396 11744 15424 11852
rect 16022 11840 16028 11892
rect 16080 11880 16086 11892
rect 16117 11883 16175 11889
rect 16117 11880 16129 11883
rect 16080 11852 16129 11880
rect 16080 11840 16086 11852
rect 16117 11849 16129 11852
rect 16163 11849 16175 11883
rect 16117 11843 16175 11849
rect 18138 11840 18144 11892
rect 18196 11880 18202 11892
rect 18417 11883 18475 11889
rect 18417 11880 18429 11883
rect 18196 11852 18429 11880
rect 18196 11840 18202 11852
rect 18417 11849 18429 11852
rect 18463 11849 18475 11883
rect 18417 11843 18475 11849
rect 18782 11840 18788 11892
rect 18840 11880 18846 11892
rect 19245 11883 19303 11889
rect 19245 11880 19257 11883
rect 18840 11852 19257 11880
rect 18840 11840 18846 11852
rect 19245 11849 19257 11852
rect 19291 11849 19303 11883
rect 19426 11880 19432 11892
rect 19387 11852 19432 11880
rect 19245 11843 19303 11849
rect 19426 11840 19432 11852
rect 19484 11840 19490 11892
rect 15841 11815 15899 11821
rect 15841 11781 15853 11815
rect 15887 11812 15899 11815
rect 16206 11812 16212 11824
rect 15887 11784 16212 11812
rect 15887 11781 15899 11784
rect 15841 11775 15899 11781
rect 16206 11772 16212 11784
rect 16264 11772 16270 11824
rect 19058 11812 19064 11824
rect 16960 11784 19064 11812
rect 16850 11744 16856 11756
rect 15396 11716 16856 11744
rect 16850 11704 16856 11716
rect 16908 11704 16914 11756
rect 16960 11676 16988 11784
rect 19058 11772 19064 11784
rect 19116 11772 19122 11824
rect 17034 11704 17040 11756
rect 17092 11744 17098 11756
rect 17586 11744 17592 11756
rect 17092 11716 17137 11744
rect 17547 11716 17592 11744
rect 17092 11704 17098 11716
rect 17586 11704 17592 11716
rect 17644 11704 17650 11756
rect 17678 11704 17684 11756
rect 17736 11744 17742 11756
rect 18969 11747 19027 11753
rect 18969 11744 18981 11747
rect 17736 11716 18981 11744
rect 17736 11704 17742 11716
rect 18969 11713 18981 11716
rect 19015 11713 19027 11747
rect 18969 11707 19027 11713
rect 20073 11747 20131 11753
rect 20073 11713 20085 11747
rect 20119 11744 20131 11747
rect 20346 11744 20352 11756
rect 20119 11716 20352 11744
rect 20119 11713 20131 11716
rect 20073 11707 20131 11713
rect 20346 11704 20352 11716
rect 20404 11704 20410 11756
rect 20714 11704 20720 11756
rect 20772 11744 20778 11756
rect 20993 11747 21051 11753
rect 20993 11744 21005 11747
rect 20772 11716 21005 11744
rect 20772 11704 20778 11716
rect 20993 11713 21005 11716
rect 21039 11713 21051 11747
rect 20993 11707 21051 11713
rect 21085 11747 21143 11753
rect 21085 11713 21097 11747
rect 21131 11713 21143 11747
rect 21085 11707 21143 11713
rect 15120 11648 16988 11676
rect 17696 11608 17724 11704
rect 17773 11679 17831 11685
rect 17773 11645 17785 11679
rect 17819 11676 17831 11679
rect 17862 11676 17868 11688
rect 17819 11648 17868 11676
rect 17819 11645 17831 11648
rect 17773 11639 17831 11645
rect 17862 11636 17868 11648
rect 17920 11636 17926 11688
rect 19889 11679 19947 11685
rect 19889 11676 19901 11679
rect 18064 11648 19901 11676
rect 18064 11608 18092 11648
rect 19889 11645 19901 11648
rect 19935 11645 19947 11679
rect 20898 11676 20904 11688
rect 20859 11648 20904 11676
rect 19889 11639 19947 11645
rect 20898 11636 20904 11648
rect 20956 11636 20962 11688
rect 13924 11580 17724 11608
rect 17788 11580 18092 11608
rect 18785 11611 18843 11617
rect 17788 11552 17816 11580
rect 18785 11577 18797 11611
rect 18831 11608 18843 11611
rect 19245 11611 19303 11617
rect 19245 11608 19257 11611
rect 18831 11580 19257 11608
rect 18831 11577 18843 11580
rect 18785 11571 18843 11577
rect 19245 11577 19257 11580
rect 19291 11577 19303 11611
rect 19245 11571 19303 11577
rect 20346 11568 20352 11620
rect 20404 11608 20410 11620
rect 21100 11608 21128 11707
rect 20404 11580 21128 11608
rect 20404 11568 20410 11580
rect 2682 11500 2688 11552
rect 2740 11540 2746 11552
rect 3510 11540 3516 11552
rect 2740 11512 3516 11540
rect 2740 11500 2746 11512
rect 3510 11500 3516 11512
rect 3568 11500 3574 11552
rect 4338 11540 4344 11552
rect 4299 11512 4344 11540
rect 4338 11500 4344 11512
rect 4396 11500 4402 11552
rect 4430 11500 4436 11552
rect 4488 11540 4494 11552
rect 4488 11512 4533 11540
rect 4488 11500 4494 11512
rect 5074 11500 5080 11552
rect 5132 11540 5138 11552
rect 5442 11540 5448 11552
rect 5132 11512 5448 11540
rect 5132 11500 5138 11512
rect 5442 11500 5448 11512
rect 5500 11500 5506 11552
rect 7190 11500 7196 11552
rect 7248 11540 7254 11552
rect 7285 11543 7343 11549
rect 7285 11540 7297 11543
rect 7248 11512 7297 11540
rect 7248 11500 7254 11512
rect 7285 11509 7297 11512
rect 7331 11509 7343 11543
rect 8846 11540 8852 11552
rect 8807 11512 8852 11540
rect 7285 11503 7343 11509
rect 8846 11500 8852 11512
rect 8904 11500 8910 11552
rect 9858 11540 9864 11552
rect 9819 11512 9864 11540
rect 9858 11500 9864 11512
rect 9916 11500 9922 11552
rect 9953 11543 10011 11549
rect 9953 11509 9965 11543
rect 9999 11540 10011 11543
rect 10410 11540 10416 11552
rect 9999 11512 10416 11540
rect 9999 11509 10011 11512
rect 9953 11503 10011 11509
rect 10410 11500 10416 11512
rect 10468 11540 10474 11552
rect 10781 11543 10839 11549
rect 10781 11540 10793 11543
rect 10468 11512 10793 11540
rect 10468 11500 10474 11512
rect 10781 11509 10793 11512
rect 10827 11509 10839 11543
rect 12158 11540 12164 11552
rect 12119 11512 12164 11540
rect 10781 11503 10839 11509
rect 12158 11500 12164 11512
rect 12216 11500 12222 11552
rect 12250 11500 12256 11552
rect 12308 11540 12314 11552
rect 12308 11512 12353 11540
rect 12308 11500 12314 11512
rect 13170 11500 13176 11552
rect 13228 11540 13234 11552
rect 13357 11543 13415 11549
rect 13357 11540 13369 11543
rect 13228 11512 13369 11540
rect 13228 11500 13234 11512
rect 13357 11509 13369 11512
rect 13403 11509 13415 11543
rect 15378 11540 15384 11552
rect 15339 11512 15384 11540
rect 13357 11503 13415 11509
rect 15378 11500 15384 11512
rect 15436 11500 15442 11552
rect 15470 11500 15476 11552
rect 15528 11540 15534 11552
rect 16574 11540 16580 11552
rect 15528 11512 15573 11540
rect 16535 11512 16580 11540
rect 15528 11500 15534 11512
rect 16574 11500 16580 11512
rect 16632 11500 16638 11552
rect 17586 11500 17592 11552
rect 17644 11540 17650 11552
rect 17681 11543 17739 11549
rect 17681 11540 17693 11543
rect 17644 11512 17693 11540
rect 17644 11500 17650 11512
rect 17681 11509 17693 11512
rect 17727 11509 17739 11543
rect 17681 11503 17739 11509
rect 17770 11500 17776 11552
rect 17828 11500 17834 11552
rect 18141 11543 18199 11549
rect 18141 11509 18153 11543
rect 18187 11540 18199 11543
rect 18877 11543 18935 11549
rect 18877 11540 18889 11543
rect 18187 11512 18889 11540
rect 18187 11509 18199 11512
rect 18141 11503 18199 11509
rect 18877 11509 18889 11512
rect 18923 11509 18935 11543
rect 18877 11503 18935 11509
rect 19058 11500 19064 11552
rect 19116 11540 19122 11552
rect 19797 11543 19855 11549
rect 19797 11540 19809 11543
rect 19116 11512 19809 11540
rect 19116 11500 19122 11512
rect 19797 11509 19809 11512
rect 19843 11509 19855 11543
rect 19797 11503 19855 11509
rect 20254 11500 20260 11552
rect 20312 11540 20318 11552
rect 20533 11543 20591 11549
rect 20533 11540 20545 11543
rect 20312 11512 20545 11540
rect 20312 11500 20318 11512
rect 20533 11509 20545 11512
rect 20579 11509 20591 11543
rect 20533 11503 20591 11509
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 3145 11339 3203 11345
rect 3145 11305 3157 11339
rect 3191 11336 3203 11339
rect 4338 11336 4344 11348
rect 3191 11308 4344 11336
rect 3191 11305 3203 11308
rect 3145 11299 3203 11305
rect 4338 11296 4344 11308
rect 4396 11296 4402 11348
rect 4433 11339 4491 11345
rect 4433 11305 4445 11339
rect 4479 11336 4491 11339
rect 5258 11336 5264 11348
rect 4479 11308 5264 11336
rect 4479 11305 4491 11308
rect 4433 11299 4491 11305
rect 5258 11296 5264 11308
rect 5316 11296 5322 11348
rect 6270 11336 6276 11348
rect 6231 11308 6276 11336
rect 6270 11296 6276 11308
rect 6328 11296 6334 11348
rect 6457 11339 6515 11345
rect 6457 11305 6469 11339
rect 6503 11336 6515 11339
rect 6503 11308 8340 11336
rect 6503 11305 6515 11308
rect 6457 11299 6515 11305
rect 1670 11268 1676 11280
rect 1631 11240 1676 11268
rect 1670 11228 1676 11240
rect 1728 11268 1734 11280
rect 3421 11271 3479 11277
rect 3421 11268 3433 11271
rect 1728 11240 3433 11268
rect 1728 11228 1734 11240
rect 3421 11237 3433 11240
rect 3467 11237 3479 11271
rect 3421 11231 3479 11237
rect 3878 11228 3884 11280
rect 3936 11268 3942 11280
rect 3936 11240 5856 11268
rect 3936 11228 3942 11240
rect 2777 11203 2835 11209
rect 2777 11169 2789 11203
rect 2823 11200 2835 11203
rect 4154 11200 4160 11212
rect 2823 11172 4160 11200
rect 2823 11169 2835 11172
rect 2777 11163 2835 11169
rect 4154 11160 4160 11172
rect 4212 11160 4218 11212
rect 5557 11203 5615 11209
rect 5557 11169 5569 11203
rect 5603 11200 5615 11203
rect 5718 11200 5724 11212
rect 5603 11172 5724 11200
rect 5603 11169 5615 11172
rect 5557 11163 5615 11169
rect 5718 11160 5724 11172
rect 5776 11160 5782 11212
rect 5828 11209 5856 11240
rect 5813 11203 5871 11209
rect 5813 11169 5825 11203
rect 5859 11169 5871 11203
rect 6288 11200 6316 11296
rect 7006 11268 7012 11280
rect 6967 11240 7012 11268
rect 7006 11228 7012 11240
rect 7064 11228 7070 11280
rect 7742 11228 7748 11280
rect 7800 11228 7806 11280
rect 8021 11271 8079 11277
rect 8021 11237 8033 11271
rect 8067 11268 8079 11271
rect 8202 11268 8208 11280
rect 8067 11240 8208 11268
rect 8067 11237 8079 11240
rect 8021 11231 8079 11237
rect 8202 11228 8208 11240
rect 8260 11228 8266 11280
rect 8312 11268 8340 11308
rect 8846 11296 8852 11348
rect 8904 11336 8910 11348
rect 9401 11339 9459 11345
rect 9401 11336 9413 11339
rect 8904 11308 9413 11336
rect 8904 11296 8910 11308
rect 9401 11305 9413 11308
rect 9447 11305 9459 11339
rect 9401 11299 9459 11305
rect 11238 11296 11244 11348
rect 11296 11336 11302 11348
rect 12250 11336 12256 11348
rect 11296 11308 12256 11336
rect 11296 11296 11302 11308
rect 12250 11296 12256 11308
rect 12308 11336 12314 11348
rect 13909 11339 13967 11345
rect 12308 11308 13860 11336
rect 12308 11296 12314 11308
rect 10870 11268 10876 11280
rect 8312 11240 10876 11268
rect 10870 11228 10876 11240
rect 10928 11228 10934 11280
rect 13832 11268 13860 11308
rect 13909 11305 13921 11339
rect 13955 11336 13967 11339
rect 15194 11336 15200 11348
rect 13955 11308 15200 11336
rect 13955 11305 13967 11308
rect 13909 11299 13967 11305
rect 15194 11296 15200 11308
rect 15252 11336 15258 11348
rect 15838 11336 15844 11348
rect 15252 11308 15844 11336
rect 15252 11296 15258 11308
rect 15838 11296 15844 11308
rect 15896 11296 15902 11348
rect 15930 11296 15936 11348
rect 15988 11336 15994 11348
rect 16945 11339 17003 11345
rect 16945 11336 16957 11339
rect 15988 11308 16957 11336
rect 15988 11296 15994 11308
rect 16945 11305 16957 11308
rect 16991 11336 17003 11339
rect 18046 11336 18052 11348
rect 16991 11308 18052 11336
rect 16991 11305 17003 11308
rect 16945 11299 17003 11305
rect 18046 11296 18052 11308
rect 18104 11336 18110 11348
rect 20622 11336 20628 11348
rect 18104 11308 20628 11336
rect 18104 11296 18110 11308
rect 20622 11296 20628 11308
rect 20680 11296 20686 11348
rect 18874 11268 18880 11280
rect 12406 11240 13768 11268
rect 13832 11240 18880 11268
rect 6917 11203 6975 11209
rect 6917 11200 6929 11203
rect 6288 11172 6929 11200
rect 5813 11163 5871 11169
rect 6917 11169 6929 11172
rect 6963 11169 6975 11203
rect 7760 11200 7788 11228
rect 8113 11203 8171 11209
rect 8113 11200 8125 11203
rect 7760 11172 8125 11200
rect 6917 11163 6975 11169
rect 8113 11169 8125 11172
rect 8159 11169 8171 11203
rect 8113 11163 8171 11169
rect 10045 11203 10103 11209
rect 10045 11169 10057 11203
rect 10091 11200 10103 11203
rect 11701 11203 11759 11209
rect 11701 11200 11713 11203
rect 10091 11172 11713 11200
rect 10091 11169 10103 11172
rect 10045 11163 10103 11169
rect 11701 11169 11713 11172
rect 11747 11200 11759 11203
rect 12406 11200 12434 11240
rect 13446 11200 13452 11212
rect 11747 11172 12434 11200
rect 13407 11172 13452 11200
rect 11747 11169 11759 11172
rect 11701 11163 11759 11169
rect 13446 11160 13452 11172
rect 13504 11160 13510 11212
rect 13740 11209 13768 11240
rect 18874 11228 18880 11240
rect 18932 11228 18938 11280
rect 20248 11271 20306 11277
rect 20248 11237 20260 11271
rect 20294 11268 20306 11271
rect 20346 11268 20352 11280
rect 20294 11240 20352 11268
rect 20294 11237 20306 11240
rect 20248 11231 20306 11237
rect 20346 11228 20352 11240
rect 20404 11228 20410 11280
rect 13725 11203 13783 11209
rect 13725 11169 13737 11203
rect 13771 11169 13783 11203
rect 17954 11200 17960 11212
rect 17915 11172 17960 11200
rect 13725 11163 13783 11169
rect 17954 11160 17960 11172
rect 18012 11160 18018 11212
rect 18785 11203 18843 11209
rect 18785 11169 18797 11203
rect 18831 11200 18843 11203
rect 19058 11200 19064 11212
rect 18831 11172 19064 11200
rect 18831 11169 18843 11172
rect 18785 11163 18843 11169
rect 19058 11160 19064 11172
rect 19116 11160 19122 11212
rect 19981 11203 20039 11209
rect 19981 11169 19993 11203
rect 20027 11200 20039 11203
rect 20070 11200 20076 11212
rect 20027 11172 20076 11200
rect 20027 11169 20039 11172
rect 19981 11163 20039 11169
rect 20070 11160 20076 11172
rect 20128 11160 20134 11212
rect 2590 11132 2596 11144
rect 2551 11104 2596 11132
rect 2590 11092 2596 11104
rect 2648 11092 2654 11144
rect 2685 11135 2743 11141
rect 2685 11101 2697 11135
rect 2731 11132 2743 11135
rect 4246 11132 4252 11144
rect 2731 11104 4252 11132
rect 2731 11101 2743 11104
rect 2685 11095 2743 11101
rect 4246 11092 4252 11104
rect 4304 11092 4310 11144
rect 6825 11135 6883 11141
rect 6825 11101 6837 11135
rect 6871 11101 6883 11135
rect 6825 11095 6883 11101
rect 8205 11135 8263 11141
rect 8205 11101 8217 11135
rect 8251 11101 8263 11135
rect 8205 11095 8263 11101
rect 1857 11067 1915 11073
rect 1857 11033 1869 11067
rect 1903 11064 1915 11067
rect 6840 11064 6868 11095
rect 8018 11064 8024 11076
rect 1903 11036 4936 11064
rect 6840 11036 8024 11064
rect 1903 11033 1915 11036
rect 1857 11027 1915 11033
rect 3786 10956 3792 11008
rect 3844 10996 3850 11008
rect 3881 10999 3939 11005
rect 3881 10996 3893 10999
rect 3844 10968 3893 10996
rect 3844 10956 3850 10968
rect 3881 10965 3893 10968
rect 3927 10965 3939 10999
rect 4908 10996 4936 11036
rect 8018 11024 8024 11036
rect 8076 11064 8082 11076
rect 8220 11064 8248 11095
rect 8846 11092 8852 11144
rect 8904 11132 8910 11144
rect 9030 11132 9036 11144
rect 8904 11104 9036 11132
rect 8904 11092 8910 11104
rect 9030 11092 9036 11104
rect 9088 11132 9094 11144
rect 9088 11104 10180 11132
rect 9088 11092 9094 11104
rect 8076 11036 8248 11064
rect 8076 11024 8082 11036
rect 8570 11024 8576 11076
rect 8628 11064 8634 11076
rect 9861 11067 9919 11073
rect 9861 11064 9873 11067
rect 8628 11036 9873 11064
rect 8628 11024 8634 11036
rect 9861 11033 9873 11036
rect 9907 11033 9919 11067
rect 10152 11064 10180 11104
rect 11238 11092 11244 11144
rect 11296 11132 11302 11144
rect 11333 11135 11391 11141
rect 11333 11132 11345 11135
rect 11296 11104 11345 11132
rect 11296 11092 11302 11104
rect 11333 11101 11345 11104
rect 11379 11101 11391 11135
rect 11333 11095 11391 11101
rect 11974 11092 11980 11144
rect 12032 11132 12038 11144
rect 15470 11132 15476 11144
rect 12032 11104 15476 11132
rect 12032 11092 12038 11104
rect 15470 11092 15476 11104
rect 15528 11092 15534 11144
rect 16022 11132 16028 11144
rect 15580 11104 16028 11132
rect 14921 11067 14979 11073
rect 14921 11064 14933 11067
rect 10152 11036 14933 11064
rect 9861 11027 9919 11033
rect 14921 11033 14933 11036
rect 14967 11064 14979 11067
rect 15378 11064 15384 11076
rect 14967 11036 15384 11064
rect 14967 11033 14979 11036
rect 14921 11027 14979 11033
rect 15378 11024 15384 11036
rect 15436 11024 15442 11076
rect 15580 11064 15608 11104
rect 16022 11092 16028 11104
rect 16080 11132 16086 11144
rect 16485 11135 16543 11141
rect 16485 11132 16497 11135
rect 16080 11104 16497 11132
rect 16080 11092 16086 11104
rect 16485 11101 16497 11104
rect 16531 11132 16543 11135
rect 18046 11132 18052 11144
rect 16531 11104 17908 11132
rect 18007 11104 18052 11132
rect 16531 11101 16543 11104
rect 16485 11095 16543 11101
rect 15488 11036 15608 11064
rect 15657 11067 15715 11073
rect 6457 10999 6515 11005
rect 6457 10996 6469 10999
rect 4908 10968 6469 10996
rect 3881 10959 3939 10965
rect 6457 10965 6469 10968
rect 6503 10965 6515 10999
rect 6457 10959 6515 10965
rect 7098 10956 7104 11008
rect 7156 10996 7162 11008
rect 7377 10999 7435 11005
rect 7377 10996 7389 10999
rect 7156 10968 7389 10996
rect 7156 10956 7162 10968
rect 7377 10965 7389 10968
rect 7423 10965 7435 10999
rect 7650 10996 7656 11008
rect 7611 10968 7656 10996
rect 7377 10959 7435 10965
rect 7650 10956 7656 10968
rect 7708 10956 7714 11008
rect 10134 10956 10140 11008
rect 10192 10996 10198 11008
rect 15488 10996 15516 11036
rect 15657 11033 15669 11067
rect 15703 11064 15715 11067
rect 16206 11064 16212 11076
rect 15703 11036 16212 11064
rect 15703 11033 15715 11036
rect 15657 11027 15715 11033
rect 16206 11024 16212 11036
rect 16264 11024 16270 11076
rect 16758 11024 16764 11076
rect 16816 11064 16822 11076
rect 17589 11067 17647 11073
rect 17589 11064 17601 11067
rect 16816 11036 17601 11064
rect 16816 11024 16822 11036
rect 17589 11033 17601 11036
rect 17635 11033 17647 11067
rect 17880 11064 17908 11104
rect 18046 11092 18052 11104
rect 18104 11092 18110 11144
rect 18233 11135 18291 11141
rect 18233 11101 18245 11135
rect 18279 11132 18291 11135
rect 19150 11132 19156 11144
rect 18279 11104 19156 11132
rect 18279 11101 18291 11104
rect 18233 11095 18291 11101
rect 19150 11092 19156 11104
rect 19208 11092 19214 11144
rect 19886 11132 19892 11144
rect 19260 11104 19892 11132
rect 18966 11064 18972 11076
rect 17880 11036 18972 11064
rect 17589 11027 17647 11033
rect 18966 11024 18972 11036
rect 19024 11024 19030 11076
rect 19260 11073 19288 11104
rect 19886 11092 19892 11104
rect 19944 11092 19950 11144
rect 19245 11067 19303 11073
rect 19245 11033 19257 11067
rect 19291 11033 19303 11067
rect 19702 11064 19708 11076
rect 19663 11036 19708 11064
rect 19245 11027 19303 11033
rect 19702 11024 19708 11036
rect 19760 11024 19766 11076
rect 22002 11064 22008 11076
rect 21963 11036 22008 11064
rect 22002 11024 22008 11036
rect 22060 11024 22066 11076
rect 10192 10968 15516 10996
rect 16025 10999 16083 11005
rect 10192 10956 10198 10968
rect 16025 10965 16037 10999
rect 16071 10996 16083 10999
rect 16114 10996 16120 11008
rect 16071 10968 16120 10996
rect 16071 10965 16083 10968
rect 16025 10959 16083 10965
rect 16114 10956 16120 10968
rect 16172 10956 16178 11008
rect 17218 10996 17224 11008
rect 17179 10968 17224 10996
rect 17218 10956 17224 10968
rect 17276 10956 17282 11008
rect 21358 10996 21364 11008
rect 21319 10968 21364 10996
rect 21358 10956 21364 10968
rect 21416 10956 21422 11008
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 2130 10792 2136 10804
rect 2091 10764 2136 10792
rect 2130 10752 2136 10764
rect 2188 10752 2194 10804
rect 2958 10752 2964 10804
rect 3016 10792 3022 10804
rect 3053 10795 3111 10801
rect 3053 10792 3065 10795
rect 3016 10764 3065 10792
rect 3016 10752 3022 10764
rect 3053 10761 3065 10764
rect 3099 10761 3111 10795
rect 3053 10755 3111 10761
rect 4890 10752 4896 10804
rect 4948 10792 4954 10804
rect 5166 10792 5172 10804
rect 4948 10764 5172 10792
rect 4948 10752 4954 10764
rect 5166 10752 5172 10764
rect 5224 10752 5230 10804
rect 5261 10795 5319 10801
rect 5261 10761 5273 10795
rect 5307 10792 5319 10795
rect 5718 10792 5724 10804
rect 5307 10764 5724 10792
rect 5307 10761 5319 10764
rect 5261 10755 5319 10761
rect 5718 10752 5724 10764
rect 5776 10752 5782 10804
rect 6086 10752 6092 10804
rect 6144 10792 6150 10804
rect 6549 10795 6607 10801
rect 6549 10792 6561 10795
rect 6144 10764 6561 10792
rect 6144 10752 6150 10764
rect 6549 10761 6561 10764
rect 6595 10792 6607 10795
rect 10226 10792 10232 10804
rect 6595 10764 10232 10792
rect 6595 10761 6607 10764
rect 6549 10755 6607 10761
rect 10226 10752 10232 10764
rect 10284 10752 10290 10804
rect 15562 10752 15568 10804
rect 15620 10792 15626 10804
rect 16485 10795 16543 10801
rect 16485 10792 16497 10795
rect 15620 10764 16497 10792
rect 15620 10752 15626 10764
rect 16485 10761 16497 10764
rect 16531 10792 16543 10795
rect 16666 10792 16672 10804
rect 16531 10764 16672 10792
rect 16531 10761 16543 10764
rect 16485 10755 16543 10761
rect 16666 10752 16672 10764
rect 16724 10752 16730 10804
rect 18046 10752 18052 10804
rect 18104 10792 18110 10804
rect 18141 10795 18199 10801
rect 18141 10792 18153 10795
rect 18104 10764 18153 10792
rect 18104 10752 18110 10764
rect 18141 10761 18153 10764
rect 18187 10761 18199 10795
rect 18141 10755 18199 10761
rect 20346 10752 20352 10804
rect 20404 10792 20410 10804
rect 20625 10795 20683 10801
rect 20625 10792 20637 10795
rect 20404 10764 20637 10792
rect 20404 10752 20410 10764
rect 20625 10761 20637 10764
rect 20671 10761 20683 10795
rect 20625 10755 20683 10761
rect 1857 10727 1915 10733
rect 1857 10693 1869 10727
rect 1903 10724 1915 10727
rect 1903 10696 3924 10724
rect 1903 10693 1915 10696
rect 1857 10687 1915 10693
rect 3513 10659 3571 10665
rect 3513 10656 3525 10659
rect 1688 10628 3525 10656
rect 1688 10532 1716 10628
rect 3513 10625 3525 10628
rect 3559 10625 3571 10659
rect 3896 10656 3924 10696
rect 8404 10696 12434 10724
rect 5629 10659 5687 10665
rect 3896 10628 4016 10656
rect 3513 10619 3571 10625
rect 2317 10591 2375 10597
rect 2317 10557 2329 10591
rect 2363 10588 2375 10591
rect 2777 10591 2835 10597
rect 2363 10560 2636 10588
rect 2363 10557 2375 10560
rect 2317 10551 2375 10557
rect 1670 10520 1676 10532
rect 1631 10492 1676 10520
rect 1670 10480 1676 10492
rect 1728 10480 1734 10532
rect 2608 10461 2636 10560
rect 2777 10557 2789 10591
rect 2823 10588 2835 10591
rect 3050 10588 3056 10600
rect 2823 10560 3056 10588
rect 2823 10557 2835 10560
rect 2777 10551 2835 10557
rect 3050 10548 3056 10560
rect 3108 10548 3114 10600
rect 3237 10591 3295 10597
rect 3237 10557 3249 10591
rect 3283 10588 3295 10591
rect 3602 10588 3608 10600
rect 3283 10560 3608 10588
rect 3283 10557 3295 10560
rect 3237 10551 3295 10557
rect 3602 10548 3608 10560
rect 3660 10548 3666 10600
rect 3878 10588 3884 10600
rect 3839 10560 3884 10588
rect 3878 10548 3884 10560
rect 3936 10548 3942 10600
rect 3988 10588 4016 10628
rect 5629 10625 5641 10659
rect 5675 10656 5687 10659
rect 6270 10656 6276 10668
rect 5675 10628 6276 10656
rect 5675 10625 5687 10628
rect 5629 10619 5687 10625
rect 6270 10616 6276 10628
rect 6328 10616 6334 10668
rect 8404 10656 8432 10696
rect 8754 10656 8760 10668
rect 8312 10628 8432 10656
rect 8496 10628 8760 10656
rect 8312 10600 8340 10628
rect 3988 10560 8248 10588
rect 4148 10523 4206 10529
rect 4148 10489 4160 10523
rect 4194 10520 4206 10523
rect 6546 10520 6552 10532
rect 4194 10492 6552 10520
rect 4194 10489 4206 10492
rect 4148 10483 4206 10489
rect 6546 10480 6552 10492
rect 6604 10520 6610 10532
rect 6604 10492 7052 10520
rect 6604 10480 6610 10492
rect 2593 10455 2651 10461
rect 2593 10421 2605 10455
rect 2639 10421 2651 10455
rect 2593 10415 2651 10421
rect 5997 10455 6055 10461
rect 5997 10421 6009 10455
rect 6043 10452 6055 10455
rect 6178 10452 6184 10464
rect 6043 10424 6184 10452
rect 6043 10421 6055 10424
rect 5997 10415 6055 10421
rect 6178 10412 6184 10424
rect 6236 10452 6242 10464
rect 6914 10452 6920 10464
rect 6236 10424 6920 10452
rect 6236 10412 6242 10424
rect 6914 10412 6920 10424
rect 6972 10412 6978 10464
rect 7024 10461 7052 10492
rect 7558 10480 7564 10532
rect 7616 10520 7622 10532
rect 8018 10520 8024 10532
rect 7616 10492 8024 10520
rect 7616 10480 7622 10492
rect 8018 10480 8024 10492
rect 8076 10520 8082 10532
rect 8122 10523 8180 10529
rect 8122 10520 8134 10523
rect 8076 10492 8134 10520
rect 8076 10480 8082 10492
rect 8122 10489 8134 10492
rect 8168 10489 8180 10523
rect 8220 10520 8248 10560
rect 8294 10548 8300 10600
rect 8352 10548 8358 10600
rect 8389 10591 8447 10597
rect 8389 10557 8401 10591
rect 8435 10588 8447 10591
rect 8496 10588 8524 10628
rect 8754 10616 8760 10628
rect 8812 10616 8818 10668
rect 9674 10656 9680 10668
rect 9635 10628 9680 10656
rect 9674 10616 9680 10628
rect 9732 10616 9738 10668
rect 9766 10616 9772 10668
rect 9824 10656 9830 10668
rect 10686 10656 10692 10668
rect 9824 10628 10692 10656
rect 9824 10616 9830 10628
rect 10686 10616 10692 10628
rect 10744 10656 10750 10668
rect 10962 10656 10968 10668
rect 10744 10628 10968 10656
rect 10744 10616 10750 10628
rect 10962 10616 10968 10628
rect 11020 10656 11026 10668
rect 11057 10659 11115 10665
rect 11057 10656 11069 10659
rect 11020 10628 11069 10656
rect 11020 10616 11026 10628
rect 11057 10625 11069 10628
rect 11103 10625 11115 10659
rect 12406 10656 12434 10696
rect 15470 10684 15476 10736
rect 15528 10724 15534 10736
rect 16114 10724 16120 10736
rect 15528 10696 16120 10724
rect 15528 10684 15534 10696
rect 16114 10684 16120 10696
rect 16172 10724 16178 10736
rect 16172 10696 18184 10724
rect 16172 10684 16178 10696
rect 12805 10659 12863 10665
rect 12805 10656 12817 10659
rect 12406 10628 12817 10656
rect 11057 10619 11115 10625
rect 12805 10625 12817 10628
rect 12851 10656 12863 10659
rect 13170 10656 13176 10668
rect 12851 10628 13176 10656
rect 12851 10625 12863 10628
rect 12805 10619 12863 10625
rect 13170 10616 13176 10628
rect 13228 10616 13234 10668
rect 13354 10616 13360 10668
rect 13412 10656 13418 10668
rect 14461 10659 14519 10665
rect 14461 10656 14473 10659
rect 13412 10628 14473 10656
rect 13412 10616 13418 10628
rect 14461 10625 14473 10628
rect 14507 10625 14519 10659
rect 14461 10619 14519 10625
rect 17589 10659 17647 10665
rect 17589 10625 17601 10659
rect 17635 10656 17647 10659
rect 18046 10656 18052 10668
rect 17635 10628 18052 10656
rect 17635 10625 17647 10628
rect 17589 10619 17647 10625
rect 18046 10616 18052 10628
rect 18104 10616 18110 10668
rect 18156 10656 18184 10696
rect 18156 10628 19380 10656
rect 14274 10588 14280 10600
rect 8435 10560 8524 10588
rect 8588 10560 14280 10588
rect 8435 10557 8447 10560
rect 8389 10551 8447 10557
rect 8588 10520 8616 10560
rect 14274 10548 14280 10560
rect 14332 10548 14338 10600
rect 14550 10548 14556 10600
rect 14608 10588 14614 10600
rect 14717 10591 14775 10597
rect 14717 10588 14729 10591
rect 14608 10560 14729 10588
rect 14608 10548 14614 10560
rect 14717 10557 14729 10560
rect 14763 10557 14775 10591
rect 14717 10551 14775 10557
rect 16574 10548 16580 10600
rect 16632 10588 16638 10600
rect 17681 10591 17739 10597
rect 17681 10588 17693 10591
rect 16632 10560 17693 10588
rect 16632 10548 16638 10560
rect 17681 10557 17693 10560
rect 17727 10557 17739 10591
rect 19245 10591 19303 10597
rect 19245 10588 19257 10591
rect 17681 10551 17739 10557
rect 17972 10560 19257 10588
rect 8220 10492 8616 10520
rect 9861 10523 9919 10529
rect 8122 10483 8180 10489
rect 9861 10489 9873 10523
rect 9907 10520 9919 10523
rect 10505 10523 10563 10529
rect 10505 10520 10517 10523
rect 9907 10492 10517 10520
rect 9907 10489 9919 10492
rect 9861 10483 9919 10489
rect 10505 10489 10517 10492
rect 10551 10489 10563 10523
rect 10505 10483 10563 10489
rect 10870 10480 10876 10532
rect 10928 10520 10934 10532
rect 17218 10520 17224 10532
rect 10928 10492 17224 10520
rect 10928 10480 10934 10492
rect 17218 10480 17224 10492
rect 17276 10520 17282 10532
rect 17773 10523 17831 10529
rect 17773 10520 17785 10523
rect 17276 10492 17785 10520
rect 17276 10480 17282 10492
rect 17773 10489 17785 10492
rect 17819 10489 17831 10523
rect 17773 10483 17831 10489
rect 7009 10455 7067 10461
rect 7009 10421 7021 10455
rect 7055 10421 7067 10455
rect 7009 10415 7067 10421
rect 7190 10412 7196 10464
rect 7248 10452 7254 10464
rect 7374 10452 7380 10464
rect 7248 10424 7380 10452
rect 7248 10412 7254 10424
rect 7374 10412 7380 10424
rect 7432 10452 7438 10464
rect 8662 10452 8668 10464
rect 7432 10424 8668 10452
rect 7432 10412 7438 10424
rect 8662 10412 8668 10424
rect 8720 10412 8726 10464
rect 9030 10452 9036 10464
rect 8991 10424 9036 10452
rect 9030 10412 9036 10424
rect 9088 10412 9094 10464
rect 9214 10412 9220 10464
rect 9272 10452 9278 10464
rect 9769 10455 9827 10461
rect 9769 10452 9781 10455
rect 9272 10424 9781 10452
rect 9272 10412 9278 10424
rect 9769 10421 9781 10424
rect 9815 10421 9827 10455
rect 10226 10452 10232 10464
rect 10187 10424 10232 10452
rect 9769 10415 9827 10421
rect 10226 10412 10232 10424
rect 10284 10412 10290 10464
rect 12710 10412 12716 10464
rect 12768 10452 12774 10464
rect 13630 10452 13636 10464
rect 12768 10424 13636 10452
rect 12768 10412 12774 10424
rect 13630 10412 13636 10424
rect 13688 10412 13694 10464
rect 15378 10412 15384 10464
rect 15436 10452 15442 10464
rect 15841 10455 15899 10461
rect 15841 10452 15853 10455
rect 15436 10424 15853 10452
rect 15436 10412 15442 10424
rect 15841 10421 15853 10424
rect 15887 10421 15899 10455
rect 15841 10415 15899 10421
rect 16942 10412 16948 10464
rect 17000 10452 17006 10464
rect 17037 10455 17095 10461
rect 17037 10452 17049 10455
rect 17000 10424 17049 10452
rect 17000 10412 17006 10424
rect 17037 10421 17049 10424
rect 17083 10421 17095 10455
rect 17037 10415 17095 10421
rect 17126 10412 17132 10464
rect 17184 10452 17190 10464
rect 17972 10452 18000 10560
rect 19245 10557 19257 10560
rect 19291 10557 19303 10591
rect 19352 10588 19380 10628
rect 21085 10591 21143 10597
rect 21085 10588 21097 10591
rect 19352 10560 21097 10588
rect 19245 10551 19303 10557
rect 21085 10557 21097 10560
rect 21131 10557 21143 10591
rect 21085 10551 21143 10557
rect 19150 10480 19156 10532
rect 19208 10520 19214 10532
rect 19490 10523 19548 10529
rect 19490 10520 19502 10523
rect 19208 10492 19502 10520
rect 19208 10480 19214 10492
rect 19490 10489 19502 10492
rect 19536 10489 19548 10523
rect 19490 10483 19548 10489
rect 19702 10480 19708 10532
rect 19760 10520 19766 10532
rect 21266 10520 21272 10532
rect 19760 10492 21272 10520
rect 19760 10480 19766 10492
rect 21266 10480 21272 10492
rect 21324 10480 21330 10532
rect 18414 10452 18420 10464
rect 17184 10424 18000 10452
rect 18375 10424 18420 10452
rect 17184 10412 17190 10424
rect 18414 10412 18420 10424
rect 18472 10412 18478 10464
rect 18782 10412 18788 10464
rect 18840 10452 18846 10464
rect 18877 10455 18935 10461
rect 18877 10452 18889 10455
rect 18840 10424 18889 10452
rect 18840 10412 18846 10424
rect 18877 10421 18889 10424
rect 18923 10421 18935 10455
rect 18877 10415 18935 10421
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 3050 10248 3056 10260
rect 3011 10220 3056 10248
rect 3050 10208 3056 10220
rect 3108 10208 3114 10260
rect 3602 10208 3608 10260
rect 3660 10248 3666 10260
rect 4893 10251 4951 10257
rect 4893 10248 4905 10251
rect 3660 10220 4905 10248
rect 3660 10208 3666 10220
rect 4893 10217 4905 10220
rect 4939 10217 4951 10251
rect 4893 10211 4951 10217
rect 5353 10251 5411 10257
rect 5353 10217 5365 10251
rect 5399 10248 5411 10251
rect 5905 10251 5963 10257
rect 5905 10248 5917 10251
rect 5399 10220 5917 10248
rect 5399 10217 5411 10220
rect 5353 10211 5411 10217
rect 5905 10217 5917 10220
rect 5951 10217 5963 10251
rect 5905 10211 5963 10217
rect 6917 10251 6975 10257
rect 6917 10217 6929 10251
rect 6963 10217 6975 10251
rect 6917 10211 6975 10217
rect 3881 10183 3939 10189
rect 3881 10180 3893 10183
rect 1688 10152 3893 10180
rect 1688 10124 1716 10152
rect 3881 10149 3893 10152
rect 3927 10149 3939 10183
rect 3881 10143 3939 10149
rect 5261 10183 5319 10189
rect 5261 10149 5273 10183
rect 5307 10180 5319 10183
rect 6932 10180 6960 10211
rect 7006 10208 7012 10260
rect 7064 10248 7070 10260
rect 8113 10251 8171 10257
rect 7064 10220 7788 10248
rect 7064 10208 7070 10220
rect 5307 10152 6960 10180
rect 5307 10149 5319 10152
rect 5261 10143 5319 10149
rect 7098 10140 7104 10192
rect 7156 10180 7162 10192
rect 7377 10183 7435 10189
rect 7377 10180 7389 10183
rect 7156 10152 7389 10180
rect 7156 10140 7162 10152
rect 7377 10149 7389 10152
rect 7423 10149 7435 10183
rect 7650 10180 7656 10192
rect 7377 10143 7435 10149
rect 7484 10152 7656 10180
rect 1670 10112 1676 10124
rect 1631 10084 1676 10112
rect 1670 10072 1676 10084
rect 1728 10072 1734 10124
rect 2498 10072 2504 10124
rect 2556 10112 2562 10124
rect 2685 10115 2743 10121
rect 2685 10112 2697 10115
rect 2556 10084 2697 10112
rect 2556 10072 2562 10084
rect 2685 10081 2697 10084
rect 2731 10081 2743 10115
rect 3326 10112 3332 10124
rect 3287 10084 3332 10112
rect 2685 10075 2743 10081
rect 3326 10072 3332 10084
rect 3384 10112 3390 10124
rect 4249 10115 4307 10121
rect 4249 10112 4261 10115
rect 3384 10084 4261 10112
rect 3384 10072 3390 10084
rect 4249 10081 4261 10084
rect 4295 10081 4307 10115
rect 4249 10075 4307 10081
rect 6273 10115 6331 10121
rect 6273 10081 6285 10115
rect 6319 10112 6331 10115
rect 7006 10112 7012 10124
rect 6319 10084 7012 10112
rect 6319 10081 6331 10084
rect 6273 10075 6331 10081
rect 7006 10072 7012 10084
rect 7064 10072 7070 10124
rect 7285 10115 7343 10121
rect 7285 10081 7297 10115
rect 7331 10112 7343 10115
rect 7484 10112 7512 10152
rect 7650 10140 7656 10152
rect 7708 10140 7714 10192
rect 7760 10180 7788 10220
rect 8113 10217 8125 10251
rect 8159 10248 8171 10251
rect 8202 10248 8208 10260
rect 8159 10220 8208 10248
rect 8159 10217 8171 10220
rect 8113 10211 8171 10217
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 8662 10208 8668 10260
rect 8720 10248 8726 10260
rect 9125 10251 9183 10257
rect 9125 10248 9137 10251
rect 8720 10220 9137 10248
rect 8720 10208 8726 10220
rect 9125 10217 9137 10220
rect 9171 10217 9183 10251
rect 10870 10248 10876 10260
rect 9125 10211 9183 10217
rect 9232 10220 10876 10248
rect 9232 10180 9260 10220
rect 10870 10208 10876 10220
rect 10928 10208 10934 10260
rect 10962 10208 10968 10260
rect 11020 10248 11026 10260
rect 11333 10251 11391 10257
rect 11333 10248 11345 10251
rect 11020 10220 11345 10248
rect 11020 10208 11026 10220
rect 11333 10217 11345 10220
rect 11379 10217 11391 10251
rect 11333 10211 11391 10217
rect 11698 10208 11704 10260
rect 11756 10248 11762 10260
rect 11793 10251 11851 10257
rect 11793 10248 11805 10251
rect 11756 10220 11805 10248
rect 11756 10208 11762 10220
rect 11793 10217 11805 10220
rect 11839 10248 11851 10251
rect 12066 10248 12072 10260
rect 11839 10220 12072 10248
rect 11839 10217 11851 10220
rect 11793 10211 11851 10217
rect 12066 10208 12072 10220
rect 12124 10208 12130 10260
rect 13814 10208 13820 10260
rect 13872 10248 13878 10260
rect 14553 10251 14611 10257
rect 14553 10248 14565 10251
rect 13872 10220 14565 10248
rect 13872 10208 13878 10220
rect 14553 10217 14565 10220
rect 14599 10248 14611 10251
rect 15289 10251 15347 10257
rect 15289 10248 15301 10251
rect 14599 10220 15301 10248
rect 14599 10217 14611 10220
rect 14553 10211 14611 10217
rect 15289 10217 15301 10220
rect 15335 10248 15347 10251
rect 15930 10248 15936 10260
rect 15335 10220 15936 10248
rect 15335 10217 15347 10220
rect 15289 10211 15347 10217
rect 15930 10208 15936 10220
rect 15988 10208 15994 10260
rect 16666 10208 16672 10260
rect 16724 10248 16730 10260
rect 17037 10251 17095 10257
rect 17037 10248 17049 10251
rect 16724 10220 17049 10248
rect 16724 10208 16730 10220
rect 17037 10217 17049 10220
rect 17083 10217 17095 10251
rect 17037 10211 17095 10217
rect 17129 10251 17187 10257
rect 17129 10217 17141 10251
rect 17175 10248 17187 10251
rect 18414 10248 18420 10260
rect 17175 10220 18420 10248
rect 17175 10217 17187 10220
rect 17129 10211 17187 10217
rect 18414 10208 18420 10220
rect 18472 10208 18478 10260
rect 19150 10248 19156 10260
rect 19111 10220 19156 10248
rect 19150 10208 19156 10220
rect 19208 10208 19214 10260
rect 20622 10248 20628 10260
rect 20583 10220 20628 10248
rect 20622 10208 20628 10220
rect 20680 10208 20686 10260
rect 7760 10152 9260 10180
rect 9674 10140 9680 10192
rect 9732 10180 9738 10192
rect 9922 10183 9980 10189
rect 9922 10180 9934 10183
rect 9732 10152 9934 10180
rect 9732 10140 9738 10152
rect 9922 10149 9934 10152
rect 9968 10180 9980 10183
rect 10134 10180 10140 10192
rect 9968 10152 10140 10180
rect 9968 10149 9980 10152
rect 9922 10143 9980 10149
rect 10134 10140 10140 10152
rect 10192 10140 10198 10192
rect 14001 10183 14059 10189
rect 14001 10180 14013 10183
rect 10980 10152 14013 10180
rect 7331 10084 7512 10112
rect 7331 10081 7343 10084
rect 7285 10075 7343 10081
rect 8202 10072 8208 10124
rect 8260 10112 8266 10124
rect 8386 10112 8392 10124
rect 8260 10084 8392 10112
rect 8260 10072 8266 10084
rect 8386 10072 8392 10084
rect 8444 10072 8450 10124
rect 8570 10112 8576 10124
rect 8531 10084 8576 10112
rect 8570 10072 8576 10084
rect 8628 10072 8634 10124
rect 9766 10072 9772 10124
rect 9824 10112 9830 10124
rect 10778 10112 10784 10124
rect 9824 10084 10784 10112
rect 9824 10072 9830 10084
rect 10778 10072 10784 10084
rect 10836 10112 10842 10124
rect 10980 10112 11008 10152
rect 14001 10149 14013 10152
rect 14047 10180 14059 10183
rect 21082 10180 21088 10192
rect 14047 10152 21088 10180
rect 14047 10149 14059 10152
rect 14001 10143 14059 10149
rect 21082 10140 21088 10152
rect 21140 10140 21146 10192
rect 10836 10084 11008 10112
rect 12253 10115 12311 10121
rect 10836 10072 10842 10084
rect 12253 10081 12265 10115
rect 12299 10112 12311 10115
rect 12342 10112 12348 10124
rect 12299 10084 12348 10112
rect 12299 10081 12311 10084
rect 12253 10075 12311 10081
rect 12342 10072 12348 10084
rect 12400 10072 12406 10124
rect 12526 10121 12532 10124
rect 12520 10112 12532 10121
rect 12487 10084 12532 10112
rect 12520 10075 12532 10084
rect 12584 10112 12590 10124
rect 15194 10112 15200 10124
rect 12584 10084 14504 10112
rect 15155 10084 15200 10112
rect 12526 10072 12532 10075
rect 12584 10072 12590 10084
rect 2409 10047 2467 10053
rect 2409 10013 2421 10047
rect 2455 10013 2467 10047
rect 2409 10007 2467 10013
rect 2593 10047 2651 10053
rect 2593 10013 2605 10047
rect 2639 10044 2651 10047
rect 2774 10044 2780 10056
rect 2639 10016 2780 10044
rect 2639 10013 2651 10016
rect 2593 10007 2651 10013
rect 2424 9976 2452 10007
rect 2774 10004 2780 10016
rect 2832 10004 2838 10056
rect 5445 10047 5503 10053
rect 5445 10013 5457 10047
rect 5491 10044 5503 10047
rect 5718 10044 5724 10056
rect 5491 10016 5724 10044
rect 5491 10013 5503 10016
rect 5445 10007 5503 10013
rect 5718 10004 5724 10016
rect 5776 10004 5782 10056
rect 6362 10044 6368 10056
rect 6323 10016 6368 10044
rect 6362 10004 6368 10016
rect 6420 10004 6426 10056
rect 6546 10044 6552 10056
rect 6507 10016 6552 10044
rect 6546 10004 6552 10016
rect 6604 10044 6610 10056
rect 7469 10047 7527 10053
rect 7469 10044 7481 10047
rect 6604 10016 7481 10044
rect 6604 10004 6610 10016
rect 7469 10013 7481 10016
rect 7515 10013 7527 10047
rect 7469 10007 7527 10013
rect 8754 10004 8760 10056
rect 8812 10044 8818 10056
rect 9677 10047 9735 10053
rect 9677 10044 9689 10047
rect 8812 10016 9689 10044
rect 8812 10004 8818 10016
rect 9677 10013 9689 10016
rect 9723 10013 9735 10047
rect 14476 10044 14504 10084
rect 15194 10072 15200 10084
rect 15252 10072 15258 10124
rect 15838 10112 15844 10124
rect 15799 10084 15844 10112
rect 15838 10072 15844 10084
rect 15896 10072 15902 10124
rect 18046 10121 18052 10124
rect 18040 10112 18052 10121
rect 16960 10084 18052 10112
rect 15378 10044 15384 10056
rect 14476 10016 15384 10044
rect 9677 10007 9735 10013
rect 15378 10004 15384 10016
rect 15436 10044 15442 10056
rect 16960 10053 16988 10084
rect 18040 10075 18052 10084
rect 18046 10072 18052 10075
rect 18104 10072 18110 10124
rect 20533 10115 20591 10121
rect 20533 10081 20545 10115
rect 20579 10112 20591 10115
rect 21177 10115 21235 10121
rect 21177 10112 21189 10115
rect 20579 10084 21189 10112
rect 20579 10081 20591 10084
rect 20533 10075 20591 10081
rect 21177 10081 21189 10084
rect 21223 10081 21235 10115
rect 21177 10075 21235 10081
rect 16945 10047 17003 10053
rect 15436 10016 16344 10044
rect 15436 10004 15442 10016
rect 3418 9976 3424 9988
rect 2424 9948 3424 9976
rect 3418 9936 3424 9948
rect 3476 9936 3482 9988
rect 3513 9979 3571 9985
rect 3513 9945 3525 9979
rect 3559 9976 3571 9979
rect 9214 9976 9220 9988
rect 3559 9948 9220 9976
rect 3559 9945 3571 9948
rect 3513 9939 3571 9945
rect 9214 9936 9220 9948
rect 9272 9936 9278 9988
rect 11054 9976 11060 9988
rect 10967 9948 11060 9976
rect 11054 9936 11060 9948
rect 11112 9976 11118 9988
rect 12066 9976 12072 9988
rect 11112 9948 12072 9976
rect 11112 9936 11118 9948
rect 12066 9936 12072 9948
rect 12124 9936 12130 9988
rect 16316 9920 16344 10016
rect 16945 10013 16957 10047
rect 16991 10013 17003 10047
rect 16945 10007 17003 10013
rect 17126 10004 17132 10056
rect 17184 10044 17190 10056
rect 17773 10047 17831 10053
rect 17773 10044 17785 10047
rect 17184 10016 17785 10044
rect 17184 10004 17190 10016
rect 17773 10013 17785 10016
rect 17819 10013 17831 10047
rect 20806 10044 20812 10056
rect 20719 10016 20812 10044
rect 17773 10007 17831 10013
rect 20806 10004 20812 10016
rect 20864 10044 20870 10056
rect 21358 10044 21364 10056
rect 20864 10016 21364 10044
rect 20864 10004 20870 10016
rect 21358 10004 21364 10016
rect 21416 10004 21422 10056
rect 16482 9976 16488 9988
rect 16395 9948 16488 9976
rect 16482 9936 16488 9948
rect 16540 9976 16546 9988
rect 17678 9976 17684 9988
rect 16540 9948 17684 9976
rect 16540 9936 16546 9948
rect 17678 9936 17684 9948
rect 17736 9936 17742 9988
rect 1765 9911 1823 9917
rect 1765 9877 1777 9911
rect 1811 9908 1823 9911
rect 8294 9908 8300 9920
rect 1811 9880 8300 9908
rect 1811 9877 1823 9880
rect 1765 9871 1823 9877
rect 8294 9868 8300 9880
rect 8352 9868 8358 9920
rect 8386 9868 8392 9920
rect 8444 9908 8450 9920
rect 13633 9911 13691 9917
rect 8444 9880 8489 9908
rect 8444 9868 8450 9880
rect 13633 9877 13645 9911
rect 13679 9908 13691 9911
rect 13722 9908 13728 9920
rect 13679 9880 13728 9908
rect 13679 9877 13691 9880
rect 13633 9871 13691 9877
rect 13722 9868 13728 9880
rect 13780 9868 13786 9920
rect 13814 9868 13820 9920
rect 13872 9908 13878 9920
rect 14829 9911 14887 9917
rect 14829 9908 14841 9911
rect 13872 9880 14841 9908
rect 13872 9868 13878 9880
rect 14829 9877 14841 9880
rect 14875 9877 14887 9911
rect 14829 9871 14887 9877
rect 16025 9911 16083 9917
rect 16025 9877 16037 9911
rect 16071 9908 16083 9911
rect 16114 9908 16120 9920
rect 16071 9880 16120 9908
rect 16071 9877 16083 9880
rect 16025 9871 16083 9877
rect 16114 9868 16120 9880
rect 16172 9868 16178 9920
rect 16298 9868 16304 9920
rect 16356 9868 16362 9920
rect 17497 9911 17555 9917
rect 17497 9877 17509 9911
rect 17543 9908 17555 9911
rect 17954 9908 17960 9920
rect 17543 9880 17960 9908
rect 17543 9877 17555 9880
rect 17497 9871 17555 9877
rect 17954 9868 17960 9880
rect 18012 9868 18018 9920
rect 19518 9868 19524 9920
rect 19576 9908 19582 9920
rect 19613 9911 19671 9917
rect 19613 9908 19625 9911
rect 19576 9880 19625 9908
rect 19576 9868 19582 9880
rect 19613 9877 19625 9880
rect 19659 9877 19671 9911
rect 20162 9908 20168 9920
rect 20123 9880 20168 9908
rect 19613 9871 19671 9877
rect 20162 9868 20168 9880
rect 20220 9868 20226 9920
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 2038 9664 2044 9716
rect 2096 9704 2102 9716
rect 3878 9704 3884 9716
rect 2096 9676 3884 9704
rect 2096 9664 2102 9676
rect 3878 9664 3884 9676
rect 3936 9664 3942 9716
rect 7006 9664 7012 9716
rect 7064 9704 7070 9716
rect 7064 9676 7696 9704
rect 7064 9664 7070 9676
rect 3418 9636 3424 9648
rect 3379 9608 3424 9636
rect 3418 9596 3424 9608
rect 3476 9596 3482 9648
rect 7668 9636 7696 9676
rect 10244 9676 11100 9704
rect 7745 9639 7803 9645
rect 7745 9636 7757 9639
rect 7668 9608 7757 9636
rect 7745 9605 7757 9608
rect 7791 9605 7803 9639
rect 7745 9599 7803 9605
rect 7834 9596 7840 9648
rect 7892 9636 7898 9648
rect 9125 9639 9183 9645
rect 9125 9636 9137 9639
rect 7892 9608 9137 9636
rect 7892 9596 7898 9608
rect 9125 9605 9137 9608
rect 9171 9636 9183 9639
rect 10244 9636 10272 9676
rect 9171 9608 10272 9636
rect 9171 9605 9183 9608
rect 9125 9599 9183 9605
rect 10318 9596 10324 9648
rect 10376 9636 10382 9648
rect 10962 9636 10968 9648
rect 10376 9608 10968 9636
rect 10376 9596 10382 9608
rect 10962 9596 10968 9608
rect 11020 9596 11026 9648
rect 11072 9636 11100 9676
rect 11698 9664 11704 9716
rect 11756 9704 11762 9716
rect 11756 9676 12848 9704
rect 11756 9664 11762 9676
rect 11790 9636 11796 9648
rect 11072 9608 11796 9636
rect 11790 9596 11796 9608
rect 11848 9596 11854 9648
rect 12820 9636 12848 9676
rect 14274 9664 14280 9716
rect 14332 9704 14338 9716
rect 14642 9704 14648 9716
rect 14332 9676 14648 9704
rect 14332 9664 14338 9676
rect 14642 9664 14648 9676
rect 14700 9704 14706 9716
rect 17310 9704 17316 9716
rect 14700 9676 17316 9704
rect 14700 9664 14706 9676
rect 17310 9664 17316 9676
rect 17368 9664 17374 9716
rect 18046 9664 18052 9716
rect 18104 9704 18110 9716
rect 18509 9707 18567 9713
rect 18509 9704 18521 9707
rect 18104 9676 18521 9704
rect 18104 9664 18110 9676
rect 18509 9673 18521 9676
rect 18555 9673 18567 9707
rect 18509 9667 18567 9673
rect 13449 9639 13507 9645
rect 13449 9636 13461 9639
rect 12820 9608 13461 9636
rect 13449 9605 13461 9608
rect 13495 9605 13507 9639
rect 13449 9599 13507 9605
rect 19337 9639 19395 9645
rect 19337 9605 19349 9639
rect 19383 9636 19395 9639
rect 19426 9636 19432 9648
rect 19383 9608 19432 9636
rect 19383 9605 19395 9608
rect 19337 9599 19395 9605
rect 19426 9596 19432 9608
rect 19484 9596 19490 9648
rect 21082 9636 21088 9648
rect 21043 9608 21088 9636
rect 21082 9596 21088 9608
rect 21140 9596 21146 9648
rect 1596 9540 2176 9568
rect 1596 9512 1624 9540
rect 1578 9500 1584 9512
rect 1539 9472 1584 9500
rect 1578 9460 1584 9472
rect 1636 9460 1642 9512
rect 2038 9500 2044 9512
rect 1999 9472 2044 9500
rect 2038 9460 2044 9472
rect 2096 9460 2102 9512
rect 2148 9500 2176 9540
rect 7098 9528 7104 9580
rect 7156 9568 7162 9580
rect 7193 9571 7251 9577
rect 7193 9568 7205 9571
rect 7156 9540 7205 9568
rect 7156 9528 7162 9540
rect 7193 9537 7205 9540
rect 7239 9537 7251 9571
rect 7374 9568 7380 9580
rect 7335 9540 7380 9568
rect 7193 9531 7251 9537
rect 7374 9528 7380 9540
rect 7432 9528 7438 9580
rect 7558 9528 7564 9580
rect 7616 9568 7622 9580
rect 8297 9571 8355 9577
rect 8297 9568 8309 9571
rect 7616 9540 8309 9568
rect 7616 9528 7622 9540
rect 8297 9537 8309 9540
rect 8343 9537 8355 9571
rect 8297 9531 8355 9537
rect 9582 9528 9588 9580
rect 9640 9568 9646 9580
rect 10137 9571 10195 9577
rect 9640 9528 9674 9568
rect 10137 9537 10149 9571
rect 10183 9568 10195 9571
rect 11054 9568 11060 9580
rect 10183 9540 11060 9568
rect 10183 9537 10195 9540
rect 10137 9531 10195 9537
rect 11054 9528 11060 9540
rect 11112 9528 11118 9580
rect 15194 9568 15200 9580
rect 15155 9540 15200 9568
rect 15194 9528 15200 9540
rect 15252 9528 15258 9580
rect 16206 9568 16212 9580
rect 16167 9540 16212 9568
rect 16206 9528 16212 9540
rect 16264 9528 16270 9580
rect 16298 9528 16304 9580
rect 16356 9568 16362 9580
rect 17126 9568 17132 9580
rect 16356 9540 16401 9568
rect 17087 9540 17132 9568
rect 16356 9528 16362 9540
rect 17126 9528 17132 9540
rect 17184 9528 17190 9580
rect 20254 9568 20260 9580
rect 19352 9540 19656 9568
rect 20215 9540 20260 9568
rect 3697 9503 3755 9509
rect 3697 9500 3709 9503
rect 2148 9472 3709 9500
rect 3697 9469 3709 9472
rect 3743 9469 3755 9503
rect 3697 9463 3755 9469
rect 3970 9460 3976 9512
rect 4028 9500 4034 9512
rect 4433 9503 4491 9509
rect 4433 9500 4445 9503
rect 4028 9472 4445 9500
rect 4028 9460 4034 9472
rect 4433 9469 4445 9472
rect 4479 9469 4491 9503
rect 4433 9463 4491 9469
rect 6089 9503 6147 9509
rect 6089 9469 6101 9503
rect 6135 9500 6147 9503
rect 8386 9500 8392 9512
rect 6135 9472 8392 9500
rect 6135 9469 6147 9472
rect 6089 9463 6147 9469
rect 8386 9460 8392 9472
rect 8444 9460 8450 9512
rect 9646 9500 9674 9528
rect 10318 9500 10324 9512
rect 9646 9472 10088 9500
rect 10279 9472 10324 9500
rect 1854 9392 1860 9444
rect 1912 9432 1918 9444
rect 2286 9435 2344 9441
rect 2286 9432 2298 9435
rect 1912 9404 2298 9432
rect 1912 9392 1918 9404
rect 2286 9401 2298 9404
rect 2332 9401 2344 9435
rect 2286 9395 2344 9401
rect 2682 9392 2688 9444
rect 2740 9432 2746 9444
rect 2740 9404 4292 9432
rect 2740 9392 2746 9404
rect 1670 9364 1676 9376
rect 1631 9336 1676 9364
rect 1670 9324 1676 9336
rect 1728 9324 1734 9376
rect 3142 9324 3148 9376
rect 3200 9364 3206 9376
rect 4065 9367 4123 9373
rect 4065 9364 4077 9367
rect 3200 9336 4077 9364
rect 3200 9324 3206 9336
rect 4065 9333 4077 9336
rect 4111 9333 4123 9367
rect 4264 9364 4292 9404
rect 4338 9392 4344 9444
rect 4396 9432 4402 9444
rect 4801 9435 4859 9441
rect 4801 9432 4813 9435
rect 4396 9404 4813 9432
rect 4396 9392 4402 9404
rect 4801 9401 4813 9404
rect 4847 9401 4859 9435
rect 4801 9395 4859 9401
rect 7101 9435 7159 9441
rect 7101 9401 7113 9435
rect 7147 9432 7159 9435
rect 7650 9432 7656 9444
rect 7147 9404 7656 9432
rect 7147 9401 7159 9404
rect 7101 9395 7159 9401
rect 7650 9392 7656 9404
rect 7708 9392 7714 9444
rect 8205 9435 8263 9441
rect 8205 9401 8217 9435
rect 8251 9432 8263 9435
rect 9950 9432 9956 9444
rect 8251 9404 9956 9432
rect 8251 9401 8263 9404
rect 8205 9395 8263 9401
rect 9950 9392 9956 9404
rect 10008 9392 10014 9444
rect 4890 9364 4896 9376
rect 4264 9336 4896 9364
rect 4065 9327 4123 9333
rect 4890 9324 4896 9336
rect 4948 9324 4954 9376
rect 5074 9324 5080 9376
rect 5132 9364 5138 9376
rect 5169 9367 5227 9373
rect 5169 9364 5181 9367
rect 5132 9336 5181 9364
rect 5132 9324 5138 9336
rect 5169 9333 5181 9336
rect 5215 9333 5227 9367
rect 5169 9327 5227 9333
rect 5350 9324 5356 9376
rect 5408 9364 5414 9376
rect 5537 9367 5595 9373
rect 5537 9364 5549 9367
rect 5408 9336 5549 9364
rect 5408 9324 5414 9336
rect 5537 9333 5549 9336
rect 5583 9333 5595 9367
rect 5537 9327 5595 9333
rect 5810 9324 5816 9376
rect 5868 9364 5874 9376
rect 5905 9367 5963 9373
rect 5905 9364 5917 9367
rect 5868 9336 5917 9364
rect 5868 9324 5874 9336
rect 5905 9333 5917 9336
rect 5951 9333 5963 9367
rect 5905 9327 5963 9333
rect 6733 9367 6791 9373
rect 6733 9333 6745 9367
rect 6779 9364 6791 9367
rect 7006 9364 7012 9376
rect 6779 9336 7012 9364
rect 6779 9333 6791 9336
rect 6733 9327 6791 9333
rect 7006 9324 7012 9336
rect 7064 9324 7070 9376
rect 8113 9367 8171 9373
rect 8113 9333 8125 9367
rect 8159 9364 8171 9367
rect 8294 9364 8300 9376
rect 8159 9336 8300 9364
rect 8159 9333 8171 9336
rect 8113 9327 8171 9333
rect 8294 9324 8300 9336
rect 8352 9324 8358 9376
rect 8570 9324 8576 9376
rect 8628 9364 8634 9376
rect 8757 9367 8815 9373
rect 8757 9364 8769 9367
rect 8628 9336 8769 9364
rect 8628 9324 8634 9336
rect 8757 9333 8769 9336
rect 8803 9333 8815 9367
rect 8757 9327 8815 9333
rect 9677 9367 9735 9373
rect 9677 9333 9689 9367
rect 9723 9364 9735 9367
rect 9766 9364 9772 9376
rect 9723 9336 9772 9364
rect 9723 9333 9735 9336
rect 9677 9327 9735 9333
rect 9766 9324 9772 9336
rect 9824 9324 9830 9376
rect 10060 9364 10088 9472
rect 10318 9460 10324 9472
rect 10376 9460 10382 9512
rect 11885 9503 11943 9509
rect 11885 9469 11897 9503
rect 11931 9500 11943 9503
rect 13541 9503 13599 9509
rect 13541 9500 13553 9503
rect 11931 9472 13553 9500
rect 11931 9469 11943 9472
rect 11885 9463 11943 9469
rect 12268 9444 12296 9472
rect 13541 9469 13553 9472
rect 13587 9469 13599 9503
rect 13541 9463 13599 9469
rect 16942 9460 16948 9512
rect 17000 9500 17006 9512
rect 19352 9500 19380 9540
rect 19518 9500 19524 9512
rect 17000 9472 19380 9500
rect 19479 9472 19524 9500
rect 17000 9460 17006 9472
rect 19518 9460 19524 9472
rect 19576 9460 19582 9512
rect 19628 9500 19656 9540
rect 20254 9528 20260 9540
rect 20312 9528 20318 9580
rect 20441 9571 20499 9577
rect 20441 9537 20453 9571
rect 20487 9568 20499 9571
rect 20806 9568 20812 9580
rect 20487 9540 20812 9568
rect 20487 9537 20499 9540
rect 20441 9531 20499 9537
rect 20806 9528 20812 9540
rect 20864 9528 20870 9580
rect 20165 9503 20223 9509
rect 20165 9500 20177 9503
rect 19628 9472 20177 9500
rect 20165 9469 20177 9472
rect 20211 9469 20223 9503
rect 20165 9463 20223 9469
rect 12066 9392 12072 9444
rect 12124 9441 12130 9444
rect 12124 9435 12188 9441
rect 12124 9401 12142 9435
rect 12176 9401 12188 9435
rect 12124 9395 12188 9401
rect 12124 9392 12130 9395
rect 12250 9392 12256 9444
rect 12308 9392 12314 9444
rect 13722 9392 13728 9444
rect 13780 9441 13786 9444
rect 17402 9441 17408 9444
rect 13780 9435 13844 9441
rect 13780 9401 13798 9435
rect 13832 9401 13844 9435
rect 17396 9432 17408 9441
rect 13780 9395 13844 9401
rect 14660 9404 16896 9432
rect 17363 9404 17408 9432
rect 13780 9392 13786 9395
rect 10229 9367 10287 9373
rect 10229 9364 10241 9367
rect 10060 9336 10241 9364
rect 10229 9333 10241 9336
rect 10275 9333 10287 9367
rect 10686 9364 10692 9376
rect 10647 9336 10692 9364
rect 10229 9327 10287 9333
rect 10686 9324 10692 9336
rect 10744 9324 10750 9376
rect 11057 9367 11115 9373
rect 11057 9333 11069 9367
rect 11103 9364 11115 9367
rect 11330 9364 11336 9376
rect 11103 9336 11336 9364
rect 11103 9333 11115 9336
rect 11057 9327 11115 9333
rect 11330 9324 11336 9336
rect 11388 9364 11394 9376
rect 11882 9364 11888 9376
rect 11388 9336 11888 9364
rect 11388 9324 11394 9336
rect 11882 9324 11888 9336
rect 11940 9324 11946 9376
rect 13262 9364 13268 9376
rect 13223 9336 13268 9364
rect 13262 9324 13268 9336
rect 13320 9324 13326 9376
rect 13449 9367 13507 9373
rect 13449 9333 13461 9367
rect 13495 9364 13507 9367
rect 14660 9364 14688 9404
rect 13495 9336 14688 9364
rect 13495 9333 13507 9336
rect 13449 9327 13507 9333
rect 14734 9324 14740 9376
rect 14792 9364 14798 9376
rect 14921 9367 14979 9373
rect 14921 9364 14933 9367
rect 14792 9336 14933 9364
rect 14792 9324 14798 9336
rect 14921 9333 14933 9336
rect 14967 9333 14979 9367
rect 14921 9327 14979 9333
rect 15194 9324 15200 9376
rect 15252 9364 15258 9376
rect 15749 9367 15807 9373
rect 15749 9364 15761 9367
rect 15252 9336 15761 9364
rect 15252 9324 15258 9336
rect 15749 9333 15761 9336
rect 15795 9333 15807 9367
rect 16114 9364 16120 9376
rect 16075 9336 16120 9364
rect 15749 9327 15807 9333
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 16868 9364 16896 9404
rect 17396 9395 17408 9404
rect 17402 9392 17408 9395
rect 17460 9392 17466 9444
rect 19061 9435 19119 9441
rect 19061 9401 19073 9435
rect 19107 9432 19119 9435
rect 21266 9432 21272 9444
rect 19107 9404 21272 9432
rect 19107 9401 19119 9404
rect 19061 9395 19119 9401
rect 21266 9392 21272 9404
rect 21324 9392 21330 9444
rect 19610 9364 19616 9376
rect 16868 9336 19616 9364
rect 19610 9324 19616 9336
rect 19668 9324 19674 9376
rect 19794 9364 19800 9376
rect 19755 9336 19800 9364
rect 19794 9324 19800 9336
rect 19852 9324 19858 9376
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 2498 9160 2504 9172
rect 2459 9132 2504 9160
rect 2498 9120 2504 9132
rect 2556 9120 2562 9172
rect 2774 9120 2780 9172
rect 2832 9160 2838 9172
rect 3694 9160 3700 9172
rect 2832 9132 2877 9160
rect 2976 9132 3700 9160
rect 2832 9120 2838 9132
rect 1946 9052 1952 9104
rect 2004 9092 2010 9104
rect 2976 9092 3004 9132
rect 3694 9120 3700 9132
rect 3752 9120 3758 9172
rect 5445 9163 5503 9169
rect 5445 9129 5457 9163
rect 5491 9160 5503 9163
rect 5491 9132 5948 9160
rect 5491 9129 5503 9132
rect 5445 9123 5503 9129
rect 2004 9064 3004 9092
rect 2004 9052 2010 9064
rect 3418 9052 3424 9104
rect 3476 9092 3482 9104
rect 4310 9095 4368 9101
rect 4310 9092 4322 9095
rect 3476 9064 4322 9092
rect 3476 9052 3482 9064
rect 4310 9061 4322 9064
rect 4356 9061 4368 9095
rect 4310 9055 4368 9061
rect 2130 9024 2136 9036
rect 2091 8996 2136 9024
rect 2130 8984 2136 8996
rect 2188 8984 2194 9036
rect 3145 9027 3203 9033
rect 3145 8993 3157 9027
rect 3191 9024 3203 9027
rect 3602 9024 3608 9036
rect 3191 8996 3608 9024
rect 3191 8993 3203 8996
rect 3145 8987 3203 8993
rect 3602 8984 3608 8996
rect 3660 8984 3666 9036
rect 5721 9027 5779 9033
rect 5721 9024 5733 9027
rect 4080 8996 5733 9024
rect 1854 8956 1860 8968
rect 1815 8928 1860 8956
rect 1854 8916 1860 8928
rect 1912 8916 1918 8968
rect 2038 8956 2044 8968
rect 1999 8928 2044 8956
rect 2038 8916 2044 8928
rect 2096 8916 2102 8968
rect 2958 8916 2964 8968
rect 3016 8956 3022 8968
rect 3237 8959 3295 8965
rect 3237 8956 3249 8959
rect 3016 8928 3249 8956
rect 3016 8916 3022 8928
rect 3237 8925 3249 8928
rect 3283 8925 3295 8959
rect 3237 8919 3295 8925
rect 3329 8959 3387 8965
rect 3329 8925 3341 8959
rect 3375 8925 3387 8959
rect 3329 8919 3387 8925
rect 1872 8888 1900 8916
rect 3344 8888 3372 8919
rect 3418 8916 3424 8968
rect 3476 8956 3482 8968
rect 3878 8956 3884 8968
rect 3476 8928 3884 8956
rect 3476 8916 3482 8928
rect 3878 8916 3884 8928
rect 3936 8956 3942 8968
rect 4080 8965 4108 8996
rect 5721 8993 5733 8996
rect 5767 9024 5779 9027
rect 5810 9024 5816 9036
rect 5767 8996 5816 9024
rect 5767 8993 5779 8996
rect 5721 8987 5779 8993
rect 5810 8984 5816 8996
rect 5868 8984 5874 9036
rect 5920 9024 5948 9132
rect 5994 9120 6000 9172
rect 6052 9120 6058 9172
rect 7101 9163 7159 9169
rect 7101 9129 7113 9163
rect 7147 9160 7159 9163
rect 7558 9160 7564 9172
rect 7147 9132 7564 9160
rect 7147 9129 7159 9132
rect 7101 9123 7159 9129
rect 7558 9120 7564 9132
rect 7616 9120 7622 9172
rect 7742 9160 7748 9172
rect 7703 9132 7748 9160
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 9582 9120 9588 9172
rect 9640 9160 9646 9172
rect 10321 9163 10379 9169
rect 10321 9160 10333 9163
rect 9640 9132 10333 9160
rect 9640 9120 9646 9132
rect 10321 9129 10333 9132
rect 10367 9129 10379 9163
rect 10321 9123 10379 9129
rect 10870 9120 10876 9172
rect 10928 9160 10934 9172
rect 11609 9163 11667 9169
rect 11609 9160 11621 9163
rect 10928 9132 11621 9160
rect 10928 9120 10934 9132
rect 11609 9129 11621 9132
rect 11655 9129 11667 9163
rect 11609 9123 11667 9129
rect 12069 9163 12127 9169
rect 12069 9129 12081 9163
rect 12115 9160 12127 9163
rect 13541 9163 13599 9169
rect 13541 9160 13553 9163
rect 12115 9132 13553 9160
rect 12115 9129 12127 9132
rect 12069 9123 12127 9129
rect 13541 9129 13553 9132
rect 13587 9129 13599 9163
rect 13541 9123 13599 9129
rect 13633 9163 13691 9169
rect 13633 9129 13645 9163
rect 13679 9160 13691 9163
rect 13814 9160 13820 9172
rect 13679 9132 13820 9160
rect 13679 9129 13691 9132
rect 13633 9123 13691 9129
rect 13814 9120 13820 9132
rect 13872 9120 13878 9172
rect 14001 9163 14059 9169
rect 14001 9129 14013 9163
rect 14047 9160 14059 9163
rect 14185 9163 14243 9169
rect 14185 9160 14197 9163
rect 14047 9132 14197 9160
rect 14047 9129 14059 9132
rect 14001 9123 14059 9129
rect 14185 9129 14197 9132
rect 14231 9129 14243 9163
rect 14185 9123 14243 9129
rect 14829 9163 14887 9169
rect 14829 9129 14841 9163
rect 14875 9160 14887 9163
rect 15194 9160 15200 9172
rect 14875 9132 15200 9160
rect 14875 9129 14887 9132
rect 14829 9123 14887 9129
rect 15194 9120 15200 9132
rect 15252 9120 15258 9172
rect 15289 9163 15347 9169
rect 15289 9129 15301 9163
rect 15335 9160 15347 9163
rect 15841 9163 15899 9169
rect 15841 9160 15853 9163
rect 15335 9132 15853 9160
rect 15335 9129 15347 9132
rect 15289 9123 15347 9129
rect 15841 9129 15853 9132
rect 15887 9129 15899 9163
rect 15841 9123 15899 9129
rect 16301 9163 16359 9169
rect 16301 9129 16313 9163
rect 16347 9160 16359 9163
rect 18969 9163 19027 9169
rect 16347 9132 18736 9160
rect 16347 9129 16359 9132
rect 16301 9123 16359 9129
rect 6012 9092 6040 9120
rect 8294 9092 8300 9104
rect 6012 9064 8300 9092
rect 8294 9052 8300 9064
rect 8352 9052 8358 9104
rect 14921 9095 14979 9101
rect 14921 9092 14933 9095
rect 8496 9064 14933 9092
rect 8496 9036 8524 9064
rect 14921 9061 14933 9064
rect 14967 9061 14979 9095
rect 14921 9055 14979 9061
rect 16114 9052 16120 9104
rect 16172 9092 16178 9104
rect 17770 9092 17776 9104
rect 16172 9064 17776 9092
rect 16172 9052 16178 9064
rect 17770 9052 17776 9064
rect 17828 9052 17834 9104
rect 5988 9027 6046 9033
rect 5988 9024 6000 9027
rect 5920 8996 6000 9024
rect 5988 8993 6000 8996
rect 6034 9024 6046 9027
rect 7374 9024 7380 9036
rect 6034 8996 7380 9024
rect 6034 8993 6046 8996
rect 5988 8987 6046 8993
rect 7374 8984 7380 8996
rect 7432 9024 7438 9036
rect 7432 8996 7972 9024
rect 7432 8984 7438 8996
rect 4065 8959 4123 8965
rect 4065 8956 4077 8959
rect 3936 8928 4077 8956
rect 3936 8916 3942 8928
rect 4065 8925 4077 8928
rect 4111 8925 4123 8959
rect 4065 8919 4123 8925
rect 7190 8916 7196 8968
rect 7248 8956 7254 8968
rect 7944 8965 7972 8996
rect 8478 8984 8484 9036
rect 8536 8984 8542 9036
rect 9674 9024 9680 9036
rect 8680 8996 9680 9024
rect 7837 8959 7895 8965
rect 7837 8956 7849 8959
rect 7248 8928 7849 8956
rect 7248 8916 7254 8928
rect 7837 8925 7849 8928
rect 7883 8925 7895 8959
rect 7837 8919 7895 8925
rect 7929 8959 7987 8965
rect 7929 8925 7941 8959
rect 7975 8925 7987 8959
rect 7929 8919 7987 8925
rect 8680 8897 8708 8996
rect 9674 8984 9680 8996
rect 9732 9024 9738 9036
rect 10689 9027 10747 9033
rect 10689 9024 10701 9027
rect 9732 8996 9825 9024
rect 9968 8996 10701 9024
rect 9732 8984 9738 8996
rect 9398 8956 9404 8968
rect 9359 8928 9404 8956
rect 9398 8916 9404 8928
rect 9456 8916 9462 8968
rect 9585 8959 9643 8965
rect 9585 8925 9597 8959
rect 9631 8925 9643 8959
rect 9585 8919 9643 8925
rect 8665 8891 8723 8897
rect 8665 8888 8677 8891
rect 1872 8860 3372 8888
rect 6647 8860 8677 8888
rect 1394 8820 1400 8832
rect 1355 8792 1400 8820
rect 1394 8780 1400 8792
rect 1452 8780 1458 8832
rect 2498 8780 2504 8832
rect 2556 8820 2562 8832
rect 3786 8820 3792 8832
rect 2556 8792 3792 8820
rect 2556 8780 2562 8792
rect 3786 8780 3792 8792
rect 3844 8820 3850 8832
rect 6647 8820 6675 8860
rect 8665 8857 8677 8860
rect 8711 8857 8723 8891
rect 8665 8851 8723 8857
rect 7374 8820 7380 8832
rect 3844 8792 6675 8820
rect 7335 8792 7380 8820
rect 3844 8780 3850 8792
rect 7374 8780 7380 8792
rect 7432 8780 7438 8832
rect 9600 8820 9628 8919
rect 9674 8848 9680 8900
rect 9732 8888 9738 8900
rect 9968 8888 9996 8996
rect 10689 8993 10701 8996
rect 10735 9024 10747 9027
rect 11330 9024 11336 9036
rect 10735 8996 11336 9024
rect 10735 8993 10747 8996
rect 10689 8987 10747 8993
rect 11330 8984 11336 8996
rect 11388 8984 11394 9036
rect 11701 9027 11759 9033
rect 11701 8993 11713 9027
rect 11747 9024 11759 9027
rect 12434 9024 12440 9036
rect 11747 8996 12440 9024
rect 11747 8993 11759 8996
rect 11701 8987 11759 8993
rect 12434 8984 12440 8996
rect 12492 9024 12498 9036
rect 14185 9027 14243 9033
rect 12492 8996 13584 9024
rect 12492 8984 12498 8996
rect 10781 8959 10839 8965
rect 10781 8956 10793 8959
rect 10060 8928 10793 8956
rect 10060 8897 10088 8928
rect 10781 8925 10793 8928
rect 10827 8925 10839 8959
rect 10781 8919 10839 8925
rect 10873 8959 10931 8965
rect 10873 8925 10885 8959
rect 10919 8925 10931 8959
rect 10873 8919 10931 8925
rect 9732 8860 9996 8888
rect 10045 8891 10103 8897
rect 9732 8848 9738 8860
rect 10045 8857 10057 8891
rect 10091 8857 10103 8891
rect 10045 8851 10103 8857
rect 10134 8848 10140 8900
rect 10192 8888 10198 8900
rect 10888 8888 10916 8919
rect 11238 8916 11244 8968
rect 11296 8956 11302 8968
rect 11425 8959 11483 8965
rect 11425 8956 11437 8959
rect 11296 8928 11437 8956
rect 11296 8916 11302 8928
rect 11425 8925 11437 8928
rect 11471 8956 11483 8959
rect 12526 8956 12532 8968
rect 11471 8928 12532 8956
rect 11471 8925 11483 8928
rect 11425 8919 11483 8925
rect 12526 8916 12532 8928
rect 12584 8916 12590 8968
rect 13449 8959 13507 8965
rect 13449 8925 13461 8959
rect 13495 8925 13507 8959
rect 13449 8919 13507 8925
rect 10192 8860 10916 8888
rect 10192 8848 10198 8860
rect 10962 8848 10968 8900
rect 11020 8888 11026 8900
rect 11020 8860 12848 8888
rect 11020 8848 11026 8860
rect 12820 8832 12848 8860
rect 11698 8820 11704 8832
rect 9600 8792 11704 8820
rect 11698 8780 11704 8792
rect 11756 8780 11762 8832
rect 12802 8820 12808 8832
rect 12763 8792 12808 8820
rect 12802 8780 12808 8792
rect 12860 8780 12866 8832
rect 13464 8820 13492 8919
rect 13556 8888 13584 8996
rect 14185 8993 14197 9027
rect 14231 9024 14243 9027
rect 15933 9027 15991 9033
rect 15933 9024 15945 9027
rect 14231 8996 15945 9024
rect 14231 8993 14243 8996
rect 14185 8987 14243 8993
rect 15933 8993 15945 8996
rect 15979 8993 15991 9027
rect 15933 8987 15991 8993
rect 16206 8984 16212 9036
rect 16264 9024 16270 9036
rect 16577 9027 16635 9033
rect 16577 9024 16589 9027
rect 16264 8996 16589 9024
rect 16264 8984 16270 8996
rect 16577 8993 16589 8996
rect 16623 8993 16635 9027
rect 18598 9024 18604 9036
rect 16577 8987 16635 8993
rect 16684 8996 18604 9024
rect 14093 8959 14151 8965
rect 14093 8925 14105 8959
rect 14139 8956 14151 8959
rect 14645 8959 14703 8965
rect 14645 8956 14657 8959
rect 14139 8928 14657 8956
rect 14139 8925 14151 8928
rect 14093 8919 14151 8925
rect 14645 8925 14657 8928
rect 14691 8925 14703 8959
rect 14645 8919 14703 8925
rect 14734 8916 14740 8968
rect 14792 8956 14798 8968
rect 15657 8959 15715 8965
rect 15657 8956 15669 8959
rect 14792 8928 15669 8956
rect 14792 8916 14798 8928
rect 15657 8925 15669 8928
rect 15703 8925 15715 8959
rect 15657 8919 15715 8925
rect 16684 8888 16712 8996
rect 18598 8984 18604 8996
rect 18656 8984 18662 9036
rect 18708 9024 18736 9132
rect 18969 9129 18981 9163
rect 19015 9160 19027 9163
rect 19794 9160 19800 9172
rect 19015 9132 19800 9160
rect 19015 9129 19027 9132
rect 18969 9123 19027 9129
rect 19794 9120 19800 9132
rect 19852 9120 19858 9172
rect 18877 9095 18935 9101
rect 18877 9061 18889 9095
rect 18923 9092 18935 9095
rect 20162 9092 20168 9104
rect 18923 9064 20168 9092
rect 18923 9061 18935 9064
rect 18877 9055 18935 9061
rect 20162 9052 20168 9064
rect 20220 9052 20226 9104
rect 20806 9052 20812 9104
rect 20864 9092 20870 9104
rect 20910 9095 20968 9101
rect 20910 9092 20922 9095
rect 20864 9064 20922 9092
rect 20864 9052 20870 9064
rect 20910 9061 20922 9064
rect 20956 9061 20968 9095
rect 20910 9055 20968 9061
rect 19334 9024 19340 9036
rect 18708 8996 19340 9024
rect 19334 8984 19340 8996
rect 19392 8984 19398 9036
rect 17497 8959 17555 8965
rect 17497 8925 17509 8959
rect 17543 8956 17555 8959
rect 18874 8956 18880 8968
rect 17543 8928 18880 8956
rect 17543 8925 17555 8928
rect 17497 8919 17555 8925
rect 18874 8916 18880 8928
rect 18932 8916 18938 8968
rect 19153 8959 19211 8965
rect 19153 8925 19165 8959
rect 19199 8925 19211 8959
rect 21174 8956 21180 8968
rect 21135 8928 21180 8956
rect 19153 8919 19211 8925
rect 13556 8860 16712 8888
rect 17129 8891 17187 8897
rect 17129 8857 17141 8891
rect 17175 8888 17187 8891
rect 17175 8860 19012 8888
rect 17175 8857 17187 8860
rect 17129 8851 17187 8857
rect 13722 8820 13728 8832
rect 13464 8792 13728 8820
rect 13722 8780 13728 8792
rect 13780 8820 13786 8832
rect 14093 8823 14151 8829
rect 14093 8820 14105 8823
rect 13780 8792 14105 8820
rect 13780 8780 13786 8792
rect 14093 8789 14105 8792
rect 14139 8789 14151 8823
rect 14093 8783 14151 8789
rect 16761 8823 16819 8829
rect 16761 8789 16773 8823
rect 16807 8820 16819 8823
rect 17218 8820 17224 8832
rect 16807 8792 17224 8820
rect 16807 8789 16819 8792
rect 16761 8783 16819 8789
rect 17218 8780 17224 8792
rect 17276 8780 17282 8832
rect 17865 8823 17923 8829
rect 17865 8789 17877 8823
rect 17911 8820 17923 8823
rect 17954 8820 17960 8832
rect 17911 8792 17960 8820
rect 17911 8789 17923 8792
rect 17865 8783 17923 8789
rect 17954 8780 17960 8792
rect 18012 8780 18018 8832
rect 18138 8820 18144 8832
rect 18099 8792 18144 8820
rect 18138 8780 18144 8792
rect 18196 8780 18202 8832
rect 18509 8823 18567 8829
rect 18509 8789 18521 8823
rect 18555 8820 18567 8823
rect 18598 8820 18604 8832
rect 18555 8792 18604 8820
rect 18555 8789 18567 8792
rect 18509 8783 18567 8789
rect 18598 8780 18604 8792
rect 18656 8780 18662 8832
rect 18984 8820 19012 8860
rect 19058 8848 19064 8900
rect 19116 8888 19122 8900
rect 19168 8888 19196 8919
rect 21174 8916 21180 8928
rect 21232 8916 21238 8968
rect 19797 8891 19855 8897
rect 19797 8888 19809 8891
rect 19116 8860 19809 8888
rect 19116 8848 19122 8860
rect 19797 8857 19809 8860
rect 19843 8857 19855 8891
rect 19797 8851 19855 8857
rect 19242 8820 19248 8832
rect 18984 8792 19248 8820
rect 19242 8780 19248 8792
rect 19300 8780 19306 8832
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 1670 8576 1676 8628
rect 1728 8616 1734 8628
rect 1728 8588 3556 8616
rect 1728 8576 1734 8588
rect 1854 8548 1860 8560
rect 1815 8520 1860 8548
rect 1854 8508 1860 8520
rect 1912 8508 1918 8560
rect 3237 8415 3295 8421
rect 3237 8381 3249 8415
rect 3283 8381 3295 8415
rect 3237 8375 3295 8381
rect 3050 8353 3056 8356
rect 2992 8347 3056 8353
rect 2992 8313 3004 8347
rect 3038 8313 3056 8347
rect 2992 8307 3056 8313
rect 3050 8304 3056 8307
rect 3108 8304 3114 8356
rect 1578 8276 1584 8288
rect 1539 8248 1584 8276
rect 1578 8236 1584 8248
rect 1636 8236 1642 8288
rect 3252 8276 3280 8375
rect 3528 8344 3556 8588
rect 3602 8576 3608 8628
rect 3660 8616 3666 8628
rect 3881 8619 3939 8625
rect 3881 8616 3893 8619
rect 3660 8588 3893 8616
rect 3660 8576 3666 8588
rect 3881 8585 3893 8588
rect 3927 8585 3939 8619
rect 3881 8579 3939 8585
rect 6362 8576 6368 8628
rect 6420 8616 6426 8628
rect 6641 8619 6699 8625
rect 6641 8616 6653 8619
rect 6420 8588 6653 8616
rect 6420 8576 6426 8588
rect 6641 8585 6653 8588
rect 6687 8585 6699 8619
rect 11238 8616 11244 8628
rect 6641 8579 6699 8585
rect 8005 8588 11244 8616
rect 4062 8508 4068 8560
rect 4120 8548 4126 8560
rect 5353 8551 5411 8557
rect 5353 8548 5365 8551
rect 4120 8520 5365 8548
rect 4120 8508 4126 8520
rect 4525 8483 4583 8489
rect 4525 8449 4537 8483
rect 4571 8480 4583 8483
rect 4614 8480 4620 8492
rect 4571 8452 4620 8480
rect 4571 8449 4583 8452
rect 4525 8443 4583 8449
rect 4614 8440 4620 8452
rect 4672 8440 4678 8492
rect 4982 8440 4988 8492
rect 5040 8440 5046 8492
rect 3602 8372 3608 8424
rect 3660 8412 3666 8424
rect 4341 8415 4399 8421
rect 3660 8384 3705 8412
rect 3660 8372 3666 8384
rect 4341 8381 4353 8415
rect 4387 8412 4399 8415
rect 5000 8412 5028 8440
rect 5092 8421 5120 8520
rect 5353 8517 5365 8520
rect 5399 8517 5411 8551
rect 7374 8548 7380 8560
rect 5353 8511 5411 8517
rect 7116 8520 7380 8548
rect 5442 8440 5448 8492
rect 5500 8480 5506 8492
rect 6730 8480 6736 8492
rect 5500 8452 6736 8480
rect 5500 8440 5506 8452
rect 6730 8440 6736 8452
rect 6788 8440 6794 8492
rect 7116 8489 7144 8520
rect 7374 8508 7380 8520
rect 7432 8508 7438 8560
rect 8005 8548 8033 8588
rect 11238 8576 11244 8588
rect 11296 8576 11302 8628
rect 12434 8616 12440 8628
rect 12395 8588 12440 8616
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 12802 8576 12808 8628
rect 12860 8616 12866 8628
rect 21177 8619 21235 8625
rect 21177 8616 21189 8619
rect 12860 8588 21189 8616
rect 12860 8576 12866 8588
rect 21177 8585 21189 8588
rect 21223 8585 21235 8619
rect 21177 8579 21235 8585
rect 8478 8548 8484 8560
rect 7944 8520 8033 8548
rect 8439 8520 8484 8548
rect 7101 8483 7159 8489
rect 7101 8449 7113 8483
rect 7147 8449 7159 8483
rect 7101 8443 7159 8449
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8480 7343 8483
rect 7558 8480 7564 8492
rect 7331 8452 7564 8480
rect 7331 8449 7343 8452
rect 7285 8443 7343 8449
rect 7558 8440 7564 8452
rect 7616 8440 7622 8492
rect 7944 8489 7972 8520
rect 8478 8508 8484 8520
rect 8536 8508 8542 8560
rect 10134 8548 10140 8560
rect 10095 8520 10140 8548
rect 10134 8508 10140 8520
rect 10192 8508 10198 8560
rect 11698 8548 11704 8560
rect 10796 8520 11704 8548
rect 7929 8483 7987 8489
rect 7929 8449 7941 8483
rect 7975 8449 7987 8483
rect 7929 8443 7987 8449
rect 8018 8440 8024 8492
rect 8076 8480 8082 8492
rect 10318 8480 10324 8492
rect 8076 8452 8121 8480
rect 9784 8452 10324 8480
rect 8076 8440 8082 8452
rect 4387 8384 5028 8412
rect 5077 8415 5135 8421
rect 4387 8381 4399 8384
rect 4341 8375 4399 8381
rect 5077 8381 5089 8415
rect 5123 8381 5135 8415
rect 5718 8412 5724 8424
rect 5679 8384 5724 8412
rect 5077 8375 5135 8381
rect 5718 8372 5724 8384
rect 5776 8372 5782 8424
rect 7006 8412 7012 8424
rect 6967 8384 7012 8412
rect 7006 8372 7012 8384
rect 7064 8372 7070 8424
rect 7650 8372 7656 8424
rect 7708 8412 7714 8424
rect 8113 8415 8171 8421
rect 8113 8412 8125 8415
rect 7708 8384 8125 8412
rect 7708 8372 7714 8384
rect 8113 8381 8125 8384
rect 8159 8381 8171 8415
rect 8754 8412 8760 8424
rect 8715 8384 8760 8412
rect 8113 8375 8171 8381
rect 8754 8372 8760 8384
rect 8812 8372 8818 8424
rect 9024 8415 9082 8421
rect 9024 8381 9036 8415
rect 9070 8412 9082 8415
rect 9398 8412 9404 8424
rect 9070 8384 9404 8412
rect 9070 8381 9082 8384
rect 9024 8375 9082 8381
rect 9398 8372 9404 8384
rect 9456 8372 9462 8424
rect 9490 8372 9496 8424
rect 9548 8412 9554 8424
rect 9784 8412 9812 8452
rect 10318 8440 10324 8452
rect 10376 8440 10382 8492
rect 10796 8489 10824 8520
rect 11698 8508 11704 8520
rect 11756 8548 11762 8560
rect 12713 8551 12771 8557
rect 12713 8548 12725 8551
rect 11756 8520 12725 8548
rect 11756 8508 11762 8520
rect 12713 8517 12725 8520
rect 12759 8548 12771 8551
rect 12894 8548 12900 8560
rect 12759 8520 12900 8548
rect 12759 8517 12771 8520
rect 12713 8511 12771 8517
rect 12894 8508 12900 8520
rect 12952 8508 12958 8560
rect 14553 8551 14611 8557
rect 14553 8517 14565 8551
rect 14599 8548 14611 8551
rect 14642 8548 14648 8560
rect 14599 8520 14648 8548
rect 14599 8517 14611 8520
rect 14553 8511 14611 8517
rect 14642 8508 14648 8520
rect 14700 8508 14706 8560
rect 16577 8551 16635 8557
rect 16577 8517 16589 8551
rect 16623 8548 16635 8551
rect 17402 8548 17408 8560
rect 16623 8520 17408 8548
rect 16623 8517 16635 8520
rect 16577 8511 16635 8517
rect 17402 8508 17408 8520
rect 17460 8548 17466 8560
rect 17460 8520 17724 8548
rect 17460 8508 17466 8520
rect 10781 8483 10839 8489
rect 10781 8449 10793 8483
rect 10827 8449 10839 8483
rect 10781 8443 10839 8449
rect 14274 8440 14280 8492
rect 14332 8480 14338 8492
rect 17696 8489 17724 8520
rect 18046 8508 18052 8560
rect 18104 8548 18110 8560
rect 18325 8551 18383 8557
rect 18325 8548 18337 8551
rect 18104 8520 18337 8548
rect 18104 8508 18110 8520
rect 18325 8517 18337 8520
rect 18371 8548 18383 8551
rect 18690 8548 18696 8560
rect 18371 8520 18696 8548
rect 18371 8517 18383 8520
rect 18325 8511 18383 8517
rect 18690 8508 18696 8520
rect 18748 8508 18754 8560
rect 17681 8483 17739 8489
rect 14332 8452 15332 8480
rect 14332 8440 14338 8452
rect 9548 8384 9812 8412
rect 9876 8384 12940 8412
rect 9548 8372 9554 8384
rect 3528 8316 9536 8344
rect 3418 8276 3424 8288
rect 3252 8248 3424 8276
rect 3418 8236 3424 8248
rect 3476 8276 3482 8288
rect 3786 8276 3792 8288
rect 3476 8248 3792 8276
rect 3476 8236 3482 8248
rect 3786 8236 3792 8248
rect 3844 8236 3850 8288
rect 3878 8236 3884 8288
rect 3936 8276 3942 8288
rect 4249 8279 4307 8285
rect 4249 8276 4261 8279
rect 3936 8248 4261 8276
rect 3936 8236 3942 8248
rect 4249 8245 4261 8248
rect 4295 8276 4307 8279
rect 4522 8276 4528 8288
rect 4295 8248 4528 8276
rect 4295 8245 4307 8248
rect 4249 8239 4307 8245
rect 4522 8236 4528 8248
rect 4580 8236 4586 8288
rect 4890 8276 4896 8288
rect 4851 8248 4896 8276
rect 4890 8236 4896 8248
rect 4948 8236 4954 8288
rect 4982 8236 4988 8288
rect 5040 8276 5046 8288
rect 9214 8276 9220 8288
rect 5040 8248 9220 8276
rect 5040 8236 5046 8248
rect 9214 8236 9220 8248
rect 9272 8236 9278 8288
rect 9508 8276 9536 8316
rect 9876 8276 9904 8384
rect 10502 8304 10508 8356
rect 10560 8344 10566 8356
rect 10873 8347 10931 8353
rect 10873 8344 10885 8347
rect 10560 8316 10885 8344
rect 10560 8304 10566 8316
rect 10873 8313 10885 8316
rect 10919 8313 10931 8347
rect 10873 8307 10931 8313
rect 10965 8347 11023 8353
rect 10965 8313 10977 8347
rect 11011 8344 11023 8347
rect 11885 8347 11943 8353
rect 11885 8344 11897 8347
rect 11011 8316 11897 8344
rect 11011 8313 11023 8316
rect 10965 8307 11023 8313
rect 11885 8313 11897 8316
rect 11931 8313 11943 8347
rect 12912 8344 12940 8384
rect 13262 8372 13268 8424
rect 13320 8412 13326 8424
rect 13826 8415 13884 8421
rect 13826 8412 13838 8415
rect 13320 8384 13838 8412
rect 13320 8372 13326 8384
rect 13826 8381 13838 8384
rect 13872 8381 13884 8415
rect 13826 8375 13884 8381
rect 14093 8415 14151 8421
rect 14093 8381 14105 8415
rect 14139 8381 14151 8415
rect 14093 8375 14151 8381
rect 13998 8344 14004 8356
rect 11885 8307 11943 8313
rect 12544 8316 12848 8344
rect 12912 8316 14004 8344
rect 9508 8248 9904 8276
rect 11333 8279 11391 8285
rect 11333 8245 11345 8279
rect 11379 8276 11391 8279
rect 11790 8276 11796 8288
rect 11379 8248 11796 8276
rect 11379 8245 11391 8248
rect 11333 8239 11391 8245
rect 11790 8236 11796 8248
rect 11848 8236 11854 8288
rect 12066 8236 12072 8288
rect 12124 8276 12130 8288
rect 12544 8276 12572 8316
rect 12124 8248 12572 8276
rect 12820 8276 12848 8316
rect 13998 8304 14004 8316
rect 14056 8304 14062 8356
rect 14108 8344 14136 8375
rect 14458 8372 14464 8424
rect 14516 8412 14522 8424
rect 15197 8415 15255 8421
rect 15197 8412 15209 8415
rect 14516 8384 15209 8412
rect 14516 8372 14522 8384
rect 15197 8381 15209 8384
rect 15243 8381 15255 8415
rect 15304 8412 15332 8452
rect 17681 8449 17693 8483
rect 17727 8449 17739 8483
rect 17681 8443 17739 8449
rect 18230 8440 18236 8492
rect 18288 8480 18294 8492
rect 18785 8483 18843 8489
rect 18785 8480 18797 8483
rect 18288 8452 18797 8480
rect 18288 8440 18294 8452
rect 18785 8449 18797 8452
rect 18831 8449 18843 8483
rect 18785 8443 18843 8449
rect 15304 8384 16712 8412
rect 15197 8375 15255 8381
rect 14550 8344 14556 8356
rect 14108 8316 14556 8344
rect 14550 8304 14556 8316
rect 14608 8304 14614 8356
rect 14829 8347 14887 8353
rect 14829 8313 14841 8347
rect 14875 8313 14887 8347
rect 14829 8307 14887 8313
rect 15464 8347 15522 8353
rect 15464 8313 15476 8347
rect 15510 8344 15522 8347
rect 16574 8344 16580 8356
rect 15510 8316 16580 8344
rect 15510 8313 15522 8316
rect 15464 8307 15522 8313
rect 14642 8276 14648 8288
rect 12820 8248 14648 8276
rect 12124 8236 12130 8248
rect 14642 8236 14648 8248
rect 14700 8276 14706 8288
rect 14844 8276 14872 8307
rect 16574 8304 16580 8316
rect 16632 8304 16638 8356
rect 16684 8344 16712 8384
rect 16942 8372 16948 8424
rect 17000 8412 17006 8424
rect 17589 8415 17647 8421
rect 17589 8412 17601 8415
rect 17000 8384 17601 8412
rect 17000 8372 17006 8384
rect 17589 8381 17601 8384
rect 17635 8381 17647 8415
rect 17589 8375 17647 8381
rect 18509 8415 18567 8421
rect 18509 8381 18521 8415
rect 18555 8412 18567 8415
rect 18690 8412 18696 8424
rect 18555 8384 18696 8412
rect 18555 8381 18567 8384
rect 18509 8375 18567 8381
rect 18690 8372 18696 8384
rect 18748 8372 18754 8424
rect 19058 8421 19064 8424
rect 19052 8412 19064 8421
rect 19019 8384 19064 8412
rect 19052 8375 19064 8384
rect 19058 8372 19064 8375
rect 19116 8372 19122 8424
rect 20533 8415 20591 8421
rect 20533 8412 20545 8415
rect 19168 8384 20545 8412
rect 19168 8344 19196 8384
rect 20533 8381 20545 8384
rect 20579 8381 20591 8415
rect 21266 8412 21272 8424
rect 21227 8384 21272 8412
rect 20533 8375 20591 8381
rect 21266 8372 21272 8384
rect 21324 8372 21330 8424
rect 16684 8316 19196 8344
rect 19242 8304 19248 8356
rect 19300 8344 19306 8356
rect 20714 8344 20720 8356
rect 19300 8316 20720 8344
rect 19300 8304 19306 8316
rect 20714 8304 20720 8316
rect 20772 8304 20778 8356
rect 17126 8276 17132 8288
rect 14700 8248 14872 8276
rect 17087 8248 17132 8276
rect 14700 8236 14706 8248
rect 17126 8236 17132 8248
rect 17184 8236 17190 8288
rect 17310 8236 17316 8288
rect 17368 8276 17374 8288
rect 17497 8279 17555 8285
rect 17497 8276 17509 8279
rect 17368 8248 17509 8276
rect 17368 8236 17374 8248
rect 17497 8245 17509 8248
rect 17543 8245 17555 8279
rect 20162 8276 20168 8288
rect 20123 8248 20168 8276
rect 17497 8239 17555 8245
rect 20162 8236 20168 8248
rect 20220 8236 20226 8288
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 2038 8032 2044 8084
rect 2096 8072 2102 8084
rect 2409 8075 2467 8081
rect 2409 8072 2421 8075
rect 2096 8044 2421 8072
rect 2096 8032 2102 8044
rect 2409 8041 2421 8044
rect 2455 8041 2467 8075
rect 2409 8035 2467 8041
rect 2777 8075 2835 8081
rect 2777 8041 2789 8075
rect 2823 8072 2835 8075
rect 4249 8075 4307 8081
rect 2823 8044 4016 8072
rect 2823 8041 2835 8044
rect 2777 8035 2835 8041
rect 1486 7964 1492 8016
rect 1544 8004 1550 8016
rect 1673 8007 1731 8013
rect 1673 8004 1685 8007
rect 1544 7976 1685 8004
rect 1544 7964 1550 7976
rect 1673 7973 1685 7976
rect 1719 8004 1731 8007
rect 3421 8007 3479 8013
rect 3421 8004 3433 8007
rect 1719 7976 3433 8004
rect 1719 7973 1731 7976
rect 1673 7967 1731 7973
rect 3421 7973 3433 7976
rect 3467 7973 3479 8007
rect 3421 7967 3479 7973
rect 2866 7896 2872 7948
rect 2924 7936 2930 7948
rect 3234 7936 3240 7948
rect 2924 7908 3240 7936
rect 2924 7896 2930 7908
rect 3234 7896 3240 7908
rect 3292 7896 3298 7948
rect 3988 7936 4016 8044
rect 4249 8041 4261 8075
rect 4295 8072 4307 8075
rect 8478 8072 8484 8084
rect 4295 8044 8484 8072
rect 4295 8041 4307 8044
rect 4249 8035 4307 8041
rect 8478 8032 8484 8044
rect 8536 8032 8542 8084
rect 9490 8032 9496 8084
rect 9548 8072 9554 8084
rect 10321 8075 10379 8081
rect 10321 8072 10333 8075
rect 9548 8044 10333 8072
rect 9548 8032 9554 8044
rect 10321 8041 10333 8044
rect 10367 8072 10379 8075
rect 12066 8072 12072 8084
rect 10367 8044 12072 8072
rect 10367 8041 10379 8044
rect 10321 8035 10379 8041
rect 12066 8032 12072 8044
rect 12124 8032 12130 8084
rect 14642 8032 14648 8084
rect 14700 8072 14706 8084
rect 16577 8075 16635 8081
rect 16577 8072 16589 8075
rect 14700 8044 16589 8072
rect 14700 8032 14706 8044
rect 16577 8041 16589 8044
rect 16623 8041 16635 8075
rect 16942 8072 16948 8084
rect 16903 8044 16948 8072
rect 16577 8035 16635 8041
rect 16942 8032 16948 8044
rect 17000 8032 17006 8084
rect 17310 8072 17316 8084
rect 17271 8044 17316 8072
rect 17310 8032 17316 8044
rect 17368 8032 17374 8084
rect 17678 8032 17684 8084
rect 17736 8072 17742 8084
rect 17773 8075 17831 8081
rect 17773 8072 17785 8075
rect 17736 8044 17785 8072
rect 17736 8032 17742 8044
rect 17773 8041 17785 8044
rect 17819 8041 17831 8075
rect 17773 8035 17831 8041
rect 18138 8032 18144 8084
rect 18196 8072 18202 8084
rect 18196 8044 21312 8072
rect 18196 8032 18202 8044
rect 4062 7964 4068 8016
rect 4120 8004 4126 8016
rect 4157 8007 4215 8013
rect 4157 8004 4169 8007
rect 4120 7976 4169 8004
rect 4120 7964 4126 7976
rect 4157 7973 4169 7976
rect 4203 8004 4215 8007
rect 6457 8007 6515 8013
rect 6457 8004 6469 8007
rect 4203 7976 6469 8004
rect 4203 7973 4215 7976
rect 4157 7967 4215 7973
rect 6457 7973 6469 7976
rect 6503 7973 6515 8007
rect 6457 7967 6515 7973
rect 6546 7964 6552 8016
rect 6604 8004 6610 8016
rect 9125 8007 9183 8013
rect 9125 8004 9137 8007
rect 6604 7976 9137 8004
rect 6604 7964 6610 7976
rect 9125 7973 9137 7976
rect 9171 7973 9183 8007
rect 9125 7967 9183 7973
rect 11698 7964 11704 8016
rect 11756 8004 11762 8016
rect 11802 8007 11860 8013
rect 11802 8004 11814 8007
rect 11756 7976 11814 8004
rect 11756 7964 11762 7976
rect 11802 7973 11814 7976
rect 11848 7973 11860 8007
rect 11802 7967 11860 7973
rect 13265 8007 13323 8013
rect 13265 7973 13277 8007
rect 13311 8004 13323 8007
rect 13630 8004 13636 8016
rect 13311 7976 13636 8004
rect 13311 7973 13323 7976
rect 13265 7967 13323 7973
rect 13630 7964 13636 7976
rect 13688 8004 13694 8016
rect 14274 8004 14280 8016
rect 13688 7976 14280 8004
rect 13688 7964 13694 7976
rect 14274 7964 14280 7976
rect 14332 7964 14338 8016
rect 14826 8013 14832 8016
rect 14820 7967 14832 8013
rect 14884 8004 14890 8016
rect 16485 8007 16543 8013
rect 14884 7976 14920 8004
rect 14826 7964 14832 7967
rect 14884 7964 14890 7976
rect 16485 7973 16497 8007
rect 16531 8004 16543 8007
rect 17034 8004 17040 8016
rect 16531 7976 17040 8004
rect 16531 7973 16543 7976
rect 16485 7967 16543 7973
rect 17034 7964 17040 7976
rect 17092 7964 17098 8016
rect 17862 8004 17868 8016
rect 17604 7976 17868 8004
rect 3988 7908 4200 7936
rect 4172 7880 4200 7908
rect 4982 7896 4988 7948
rect 5040 7936 5046 7948
rect 5445 7939 5503 7945
rect 5445 7936 5457 7939
rect 5040 7908 5457 7936
rect 5040 7896 5046 7908
rect 5445 7905 5457 7908
rect 5491 7905 5503 7939
rect 5445 7899 5503 7905
rect 5810 7896 5816 7948
rect 5868 7936 5874 7948
rect 7929 7939 7987 7945
rect 7929 7936 7941 7939
rect 5868 7908 7941 7936
rect 5868 7896 5874 7908
rect 7929 7905 7941 7908
rect 7975 7905 7987 7939
rect 7929 7899 7987 7905
rect 8386 7896 8392 7948
rect 8444 7936 8450 7948
rect 8481 7939 8539 7945
rect 8481 7936 8493 7939
rect 8444 7908 8493 7936
rect 8444 7896 8450 7908
rect 8481 7905 8493 7908
rect 8527 7905 8539 7939
rect 8481 7899 8539 7905
rect 9214 7896 9220 7948
rect 9272 7936 9278 7948
rect 12342 7936 12348 7948
rect 9272 7908 12348 7936
rect 9272 7896 9278 7908
rect 12342 7896 12348 7908
rect 12400 7896 12406 7948
rect 12529 7939 12587 7945
rect 12529 7905 12541 7939
rect 12575 7936 12587 7939
rect 12621 7939 12679 7945
rect 12621 7936 12633 7939
rect 12575 7908 12633 7936
rect 12575 7905 12587 7908
rect 12529 7899 12587 7905
rect 12621 7905 12633 7908
rect 12667 7936 12679 7939
rect 13173 7939 13231 7945
rect 13173 7936 13185 7939
rect 12667 7908 13185 7936
rect 12667 7905 12679 7908
rect 12621 7899 12679 7905
rect 13173 7905 13185 7908
rect 13219 7936 13231 7939
rect 13538 7936 13544 7948
rect 13219 7908 13544 7936
rect 13219 7905 13231 7908
rect 13173 7899 13231 7905
rect 13538 7896 13544 7908
rect 13596 7896 13602 7948
rect 14001 7939 14059 7945
rect 14001 7905 14013 7939
rect 14047 7936 14059 7939
rect 16206 7936 16212 7948
rect 14047 7908 16212 7936
rect 14047 7905 14059 7908
rect 14001 7899 14059 7905
rect 16206 7896 16212 7908
rect 16264 7896 16270 7948
rect 16574 7896 16580 7948
rect 16632 7936 16638 7948
rect 17604 7936 17632 7976
rect 17862 7964 17868 7976
rect 17920 7964 17926 8016
rect 17954 7964 17960 8016
rect 18012 8004 18018 8016
rect 18012 7976 18460 8004
rect 18012 7964 18018 7976
rect 16632 7908 17632 7936
rect 17681 7939 17739 7945
rect 16632 7896 16638 7908
rect 17681 7905 17693 7939
rect 17727 7936 17739 7939
rect 18325 7939 18383 7945
rect 18325 7936 18337 7939
rect 17727 7908 18337 7936
rect 17727 7905 17739 7908
rect 17681 7899 17739 7905
rect 18325 7905 18337 7908
rect 18371 7905 18383 7939
rect 18432 7936 18460 7976
rect 18874 7964 18880 8016
rect 18932 8004 18938 8016
rect 20714 8004 20720 8016
rect 18932 7976 20720 8004
rect 18932 7964 18938 7976
rect 20714 7964 20720 7976
rect 20772 7964 20778 8016
rect 19061 7939 19119 7945
rect 19061 7936 19073 7939
rect 18432 7908 19073 7936
rect 18325 7899 18383 7905
rect 19061 7905 19073 7908
rect 19107 7936 19119 7939
rect 19150 7936 19156 7948
rect 19107 7908 19156 7936
rect 19107 7905 19119 7908
rect 19061 7899 19119 7905
rect 19150 7896 19156 7908
rect 19208 7896 19214 7948
rect 19797 7939 19855 7945
rect 19797 7905 19809 7939
rect 19843 7936 19855 7939
rect 20070 7936 20076 7948
rect 19843 7908 20076 7936
rect 19843 7905 19855 7908
rect 19797 7899 19855 7905
rect 20070 7896 20076 7908
rect 20128 7896 20134 7948
rect 21284 7945 21312 8044
rect 21269 7939 21327 7945
rect 21269 7905 21281 7939
rect 21315 7936 21327 7939
rect 22005 7939 22063 7945
rect 22005 7936 22017 7939
rect 21315 7908 22017 7936
rect 21315 7905 21327 7908
rect 21269 7899 21327 7905
rect 22005 7905 22017 7908
rect 22051 7905 22063 7939
rect 22005 7899 22063 7905
rect 3050 7868 3056 7880
rect 2963 7840 3056 7868
rect 3050 7828 3056 7840
rect 3108 7828 3114 7880
rect 4154 7828 4160 7880
rect 4212 7828 4218 7880
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7868 4675 7871
rect 4798 7868 4804 7880
rect 4663 7840 4804 7868
rect 4663 7837 4675 7840
rect 4617 7831 4675 7837
rect 4798 7828 4804 7840
rect 4856 7828 4862 7880
rect 5169 7871 5227 7877
rect 5169 7837 5181 7871
rect 5215 7837 5227 7871
rect 5169 7831 5227 7837
rect 1854 7800 1860 7812
rect 1815 7772 1860 7800
rect 1854 7760 1860 7772
rect 1912 7760 1918 7812
rect 3068 7800 3096 7828
rect 4522 7800 4528 7812
rect 3068 7772 4528 7800
rect 4522 7760 4528 7772
rect 4580 7760 4586 7812
rect 5184 7800 5212 7831
rect 5258 7828 5264 7880
rect 5316 7868 5322 7880
rect 5353 7871 5411 7877
rect 5353 7868 5365 7871
rect 5316 7840 5365 7868
rect 5316 7828 5322 7840
rect 5353 7837 5365 7840
rect 5399 7837 5411 7871
rect 5353 7831 5411 7837
rect 5626 7828 5632 7880
rect 5684 7868 5690 7880
rect 7561 7871 7619 7877
rect 7561 7868 7573 7871
rect 5684 7840 7573 7868
rect 5684 7828 5690 7840
rect 7561 7837 7573 7840
rect 7607 7837 7619 7871
rect 7561 7831 7619 7837
rect 7742 7828 7748 7880
rect 7800 7868 7806 7880
rect 9493 7871 9551 7877
rect 9493 7868 9505 7871
rect 7800 7840 9505 7868
rect 7800 7828 7806 7840
rect 9493 7837 9505 7840
rect 9539 7868 9551 7871
rect 12069 7871 12127 7877
rect 9539 7840 9996 7868
rect 9539 7837 9551 7840
rect 9493 7831 9551 7837
rect 5718 7800 5724 7812
rect 5184 7772 5724 7800
rect 5718 7760 5724 7772
rect 5776 7760 5782 7812
rect 5813 7803 5871 7809
rect 5813 7769 5825 7803
rect 5859 7800 5871 7803
rect 8294 7800 8300 7812
rect 5859 7772 8300 7800
rect 5859 7769 5871 7772
rect 5813 7763 5871 7769
rect 8294 7760 8300 7772
rect 8352 7760 8358 7812
rect 8386 7760 8392 7812
rect 8444 7800 8450 7812
rect 9674 7800 9680 7812
rect 8444 7772 9680 7800
rect 8444 7760 8450 7772
rect 9674 7760 9680 7772
rect 9732 7760 9738 7812
rect 9968 7809 9996 7840
rect 12069 7837 12081 7871
rect 12115 7868 12127 7871
rect 12250 7868 12256 7880
rect 12115 7840 12256 7868
rect 12115 7837 12127 7840
rect 12069 7831 12127 7837
rect 12250 7828 12256 7840
rect 12308 7868 12314 7880
rect 12308 7840 13308 7868
rect 12308 7828 12314 7840
rect 9953 7803 10011 7809
rect 9953 7769 9965 7803
rect 9999 7800 10011 7803
rect 9999 7772 11192 7800
rect 9999 7769 10011 7772
rect 9953 7763 10011 7769
rect 3326 7692 3332 7744
rect 3384 7732 3390 7744
rect 6089 7735 6147 7741
rect 6089 7732 6101 7735
rect 3384 7704 6101 7732
rect 3384 7692 3390 7704
rect 6089 7701 6101 7704
rect 6135 7701 6147 7735
rect 6914 7732 6920 7744
rect 6875 7704 6920 7732
rect 6089 7695 6147 7701
rect 6914 7692 6920 7704
rect 6972 7692 6978 7744
rect 7006 7692 7012 7744
rect 7064 7732 7070 7744
rect 7193 7735 7251 7741
rect 7193 7732 7205 7735
rect 7064 7704 7205 7732
rect 7064 7692 7070 7704
rect 7193 7701 7205 7704
rect 7239 7701 7251 7735
rect 7193 7695 7251 7701
rect 8665 7735 8723 7741
rect 8665 7701 8677 7735
rect 8711 7732 8723 7735
rect 8754 7732 8760 7744
rect 8711 7704 8760 7732
rect 8711 7701 8723 7704
rect 8665 7695 8723 7701
rect 8754 7692 8760 7704
rect 8812 7692 8818 7744
rect 10689 7735 10747 7741
rect 10689 7701 10701 7735
rect 10735 7732 10747 7735
rect 10778 7732 10784 7744
rect 10735 7704 10784 7732
rect 10735 7701 10747 7704
rect 10689 7695 10747 7701
rect 10778 7692 10784 7704
rect 10836 7692 10842 7744
rect 11164 7732 11192 7772
rect 13280 7744 13308 7840
rect 13354 7828 13360 7880
rect 13412 7868 13418 7880
rect 14550 7868 14556 7880
rect 13412 7840 13457 7868
rect 14511 7840 14556 7868
rect 13412 7828 13418 7840
rect 14550 7828 14556 7840
rect 14608 7828 14614 7880
rect 16393 7871 16451 7877
rect 16393 7837 16405 7871
rect 16439 7868 16451 7871
rect 16592 7868 16620 7896
rect 16439 7840 16620 7868
rect 16439 7837 16451 7840
rect 16393 7831 16451 7837
rect 17862 7828 17868 7880
rect 17920 7868 17926 7880
rect 17920 7840 17965 7868
rect 17920 7828 17926 7840
rect 19610 7828 19616 7880
rect 19668 7868 19674 7880
rect 20533 7871 20591 7877
rect 20533 7868 20545 7871
rect 19668 7840 20545 7868
rect 19668 7828 19674 7840
rect 20533 7837 20545 7840
rect 20579 7837 20591 7871
rect 20533 7831 20591 7837
rect 16574 7760 16580 7812
rect 16632 7800 16638 7812
rect 21085 7803 21143 7809
rect 21085 7800 21097 7803
rect 16632 7772 21097 7800
rect 16632 7760 16638 7772
rect 21085 7769 21097 7772
rect 21131 7769 21143 7803
rect 21085 7763 21143 7769
rect 12621 7735 12679 7741
rect 12621 7732 12633 7735
rect 11164 7704 12633 7732
rect 12621 7701 12633 7704
rect 12667 7701 12679 7735
rect 12802 7732 12808 7744
rect 12763 7704 12808 7732
rect 12621 7695 12679 7701
rect 12802 7692 12808 7704
rect 12860 7692 12866 7744
rect 13262 7692 13268 7744
rect 13320 7732 13326 7744
rect 13817 7735 13875 7741
rect 13817 7732 13829 7735
rect 13320 7704 13829 7732
rect 13320 7692 13326 7704
rect 13817 7701 13829 7704
rect 13863 7732 13875 7735
rect 14458 7732 14464 7744
rect 13863 7704 14464 7732
rect 13863 7701 13875 7704
rect 13817 7695 13875 7701
rect 14458 7692 14464 7704
rect 14516 7692 14522 7744
rect 15194 7692 15200 7744
rect 15252 7732 15258 7744
rect 15933 7735 15991 7741
rect 15933 7732 15945 7735
rect 15252 7704 15945 7732
rect 15252 7692 15258 7704
rect 15933 7701 15945 7704
rect 15979 7701 15991 7735
rect 15933 7695 15991 7701
rect 17034 7692 17040 7744
rect 17092 7732 17098 7744
rect 17218 7732 17224 7744
rect 17092 7704 17224 7732
rect 17092 7692 17098 7704
rect 17218 7692 17224 7704
rect 17276 7732 17282 7744
rect 18138 7732 18144 7744
rect 17276 7704 18144 7732
rect 17276 7692 17282 7704
rect 18138 7692 18144 7704
rect 18196 7692 18202 7744
rect 19242 7732 19248 7744
rect 19203 7704 19248 7732
rect 19242 7692 19248 7704
rect 19300 7692 19306 7744
rect 20254 7732 20260 7744
rect 20215 7704 20260 7732
rect 20254 7692 20260 7704
rect 20312 7692 20318 7744
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 2130 7488 2136 7540
rect 2188 7528 2194 7540
rect 2317 7531 2375 7537
rect 2317 7528 2329 7531
rect 2188 7500 2329 7528
rect 2188 7488 2194 7500
rect 2317 7497 2329 7500
rect 2363 7497 2375 7531
rect 2317 7491 2375 7497
rect 3513 7531 3571 7537
rect 3513 7497 3525 7531
rect 3559 7528 3571 7531
rect 3694 7528 3700 7540
rect 3559 7500 3700 7528
rect 3559 7497 3571 7500
rect 3513 7491 3571 7497
rect 3694 7488 3700 7500
rect 3752 7488 3758 7540
rect 5258 7528 5264 7540
rect 3804 7500 5120 7528
rect 5219 7500 5264 7528
rect 1857 7463 1915 7469
rect 1857 7429 1869 7463
rect 1903 7460 1915 7463
rect 1946 7460 1952 7472
rect 1903 7432 1952 7460
rect 1903 7429 1915 7432
rect 1857 7423 1915 7429
rect 1946 7420 1952 7432
rect 2004 7420 2010 7472
rect 3804 7460 3832 7500
rect 5092 7460 5120 7500
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 5442 7488 5448 7540
rect 5500 7528 5506 7540
rect 9125 7531 9183 7537
rect 5500 7500 8708 7528
rect 5500 7488 5506 7500
rect 6730 7460 6736 7472
rect 2792 7432 3832 7460
rect 4448 7432 4936 7460
rect 5092 7432 6736 7460
rect 2792 7401 2820 7432
rect 4448 7404 4476 7432
rect 2777 7395 2835 7401
rect 2777 7361 2789 7395
rect 2823 7361 2835 7395
rect 2777 7355 2835 7361
rect 2961 7395 3019 7401
rect 2961 7361 2973 7395
rect 3007 7392 3019 7395
rect 3050 7392 3056 7404
rect 3007 7364 3056 7392
rect 3007 7361 3019 7364
rect 2961 7355 3019 7361
rect 3050 7352 3056 7364
rect 3108 7352 3114 7404
rect 3694 7352 3700 7404
rect 3752 7392 3758 7404
rect 3878 7392 3884 7404
rect 3752 7364 3884 7392
rect 3752 7352 3758 7364
rect 3878 7352 3884 7364
rect 3936 7352 3942 7404
rect 4430 7392 4436 7404
rect 4391 7364 4436 7392
rect 4430 7352 4436 7364
rect 4488 7352 4494 7404
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7392 4583 7395
rect 4706 7392 4712 7404
rect 4571 7364 4712 7392
rect 4571 7361 4583 7364
rect 4525 7355 4583 7361
rect 4706 7352 4712 7364
rect 4764 7352 4770 7404
rect 4908 7392 4936 7432
rect 6730 7420 6736 7432
rect 6788 7420 6794 7472
rect 6822 7420 6828 7472
rect 6880 7460 6886 7472
rect 7742 7460 7748 7472
rect 6880 7432 7748 7460
rect 6880 7420 6886 7432
rect 7742 7420 7748 7432
rect 7800 7420 7806 7472
rect 8680 7460 8708 7500
rect 9125 7497 9137 7531
rect 9171 7528 9183 7531
rect 9398 7528 9404 7540
rect 9171 7500 9404 7528
rect 9171 7497 9183 7500
rect 9125 7491 9183 7497
rect 9398 7488 9404 7500
rect 9456 7488 9462 7540
rect 10870 7528 10876 7540
rect 10831 7500 10876 7528
rect 10870 7488 10876 7500
rect 10928 7488 10934 7540
rect 13998 7528 14004 7540
rect 12406 7500 13124 7528
rect 13959 7500 14004 7528
rect 9493 7463 9551 7469
rect 9493 7460 9505 7463
rect 8680 7432 9505 7460
rect 9493 7429 9505 7432
rect 9539 7429 9551 7463
rect 9493 7423 9551 7429
rect 9674 7420 9680 7472
rect 9732 7460 9738 7472
rect 9953 7463 10011 7469
rect 9953 7460 9965 7463
rect 9732 7432 9965 7460
rect 9732 7420 9738 7432
rect 9953 7429 9965 7432
rect 9999 7429 10011 7463
rect 9953 7423 10011 7429
rect 5534 7392 5540 7404
rect 4908 7364 5540 7392
rect 5534 7352 5540 7364
rect 5592 7392 5598 7404
rect 5813 7395 5871 7401
rect 5813 7392 5825 7395
rect 5592 7364 5825 7392
rect 5592 7352 5598 7364
rect 5813 7361 5825 7364
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 9030 7352 9036 7404
rect 9088 7392 9094 7404
rect 10321 7395 10379 7401
rect 10321 7392 10333 7395
rect 9088 7364 10333 7392
rect 9088 7352 9094 7364
rect 10321 7361 10333 7364
rect 10367 7361 10379 7395
rect 10321 7355 10379 7361
rect 1578 7284 1584 7336
rect 1636 7324 1642 7336
rect 2685 7327 2743 7333
rect 2685 7324 2697 7327
rect 1636 7296 2697 7324
rect 1636 7284 1642 7296
rect 2685 7293 2697 7296
rect 2731 7293 2743 7327
rect 2685 7287 2743 7293
rect 4617 7327 4675 7333
rect 4617 7293 4629 7327
rect 4663 7324 4675 7327
rect 4798 7324 4804 7336
rect 4663 7296 4804 7324
rect 4663 7293 4675 7296
rect 4617 7287 4675 7293
rect 4798 7284 4804 7296
rect 4856 7284 4862 7336
rect 5721 7327 5779 7333
rect 5721 7293 5733 7327
rect 5767 7324 5779 7327
rect 6178 7324 6184 7336
rect 5767 7296 6184 7324
rect 5767 7293 5779 7296
rect 5721 7287 5779 7293
rect 6178 7284 6184 7296
rect 6236 7284 6242 7336
rect 6362 7284 6368 7336
rect 6420 7324 6426 7336
rect 7745 7327 7803 7333
rect 7745 7324 7757 7327
rect 6420 7296 7757 7324
rect 6420 7284 6426 7296
rect 7745 7293 7757 7296
rect 7791 7324 7803 7327
rect 7791 7296 8524 7324
rect 7791 7293 7803 7296
rect 7745 7287 7803 7293
rect 1673 7259 1731 7265
rect 1673 7225 1685 7259
rect 1719 7225 1731 7259
rect 3418 7256 3424 7268
rect 3379 7228 3424 7256
rect 1673 7219 1731 7225
rect 1578 7148 1584 7200
rect 1636 7188 1642 7200
rect 1688 7188 1716 7219
rect 3418 7216 3424 7228
rect 3476 7216 3482 7268
rect 6825 7259 6883 7265
rect 6825 7256 6837 7259
rect 3528 7228 6837 7256
rect 3528 7188 3556 7228
rect 6825 7225 6837 7228
rect 6871 7225 6883 7259
rect 6825 7219 6883 7225
rect 7990 7259 8048 7265
rect 7990 7225 8002 7259
rect 8036 7225 8048 7259
rect 8496 7256 8524 7296
rect 9122 7284 9128 7336
rect 9180 7324 9186 7336
rect 11146 7324 11152 7336
rect 9180 7296 11152 7324
rect 9180 7284 9186 7296
rect 11146 7284 11152 7296
rect 11204 7324 11210 7336
rect 11241 7327 11299 7333
rect 11241 7324 11253 7327
rect 11204 7296 11253 7324
rect 11204 7284 11210 7296
rect 11241 7293 11253 7296
rect 11287 7324 11299 7327
rect 12406 7324 12434 7500
rect 12802 7392 12808 7404
rect 12763 7364 12808 7392
rect 12802 7352 12808 7364
rect 12860 7352 12866 7404
rect 12894 7352 12900 7404
rect 12952 7392 12958 7404
rect 12952 7364 12997 7392
rect 12952 7352 12958 7364
rect 11287 7296 12434 7324
rect 13096 7324 13124 7500
rect 13998 7488 14004 7500
rect 14056 7488 14062 7540
rect 14185 7531 14243 7537
rect 14185 7497 14197 7531
rect 14231 7528 14243 7531
rect 14369 7531 14427 7537
rect 14369 7528 14381 7531
rect 14231 7500 14381 7528
rect 14231 7497 14243 7500
rect 14185 7491 14243 7497
rect 14369 7497 14381 7500
rect 14415 7528 14427 7531
rect 16114 7528 16120 7540
rect 14415 7500 16120 7528
rect 14415 7497 14427 7500
rect 14369 7491 14427 7497
rect 16114 7488 16120 7500
rect 16172 7488 16178 7540
rect 16209 7531 16267 7537
rect 16209 7497 16221 7531
rect 16255 7528 16267 7531
rect 17494 7528 17500 7540
rect 16255 7500 17500 7528
rect 16255 7497 16267 7500
rect 16209 7491 16267 7497
rect 17494 7488 17500 7500
rect 17552 7488 17558 7540
rect 17862 7488 17868 7540
rect 17920 7528 17926 7540
rect 18509 7531 18567 7537
rect 18509 7528 18521 7531
rect 17920 7500 18521 7528
rect 17920 7488 17926 7500
rect 18509 7497 18521 7500
rect 18555 7497 18567 7531
rect 20438 7528 20444 7540
rect 18509 7491 18567 7497
rect 18616 7500 20444 7528
rect 13170 7420 13176 7472
rect 13228 7460 13234 7472
rect 13633 7463 13691 7469
rect 13633 7460 13645 7463
rect 13228 7432 13645 7460
rect 13228 7420 13234 7432
rect 13633 7429 13645 7432
rect 13679 7460 13691 7463
rect 16482 7460 16488 7472
rect 13679 7432 16488 7460
rect 13679 7429 13691 7432
rect 13633 7423 13691 7429
rect 16482 7420 16488 7432
rect 16540 7420 16546 7472
rect 18322 7420 18328 7472
rect 18380 7460 18386 7472
rect 18616 7460 18644 7500
rect 20438 7488 20444 7500
rect 20496 7488 20502 7540
rect 20809 7531 20867 7537
rect 20809 7497 20821 7531
rect 20855 7528 20867 7531
rect 21266 7528 21272 7540
rect 20855 7500 21272 7528
rect 20855 7497 20867 7500
rect 20809 7491 20867 7497
rect 21266 7488 21272 7500
rect 21324 7488 21330 7540
rect 18380 7432 18644 7460
rect 18380 7420 18386 7432
rect 18690 7420 18696 7472
rect 18748 7460 18754 7472
rect 21085 7463 21143 7469
rect 21085 7460 21097 7463
rect 18748 7432 21097 7460
rect 18748 7420 18754 7432
rect 21085 7429 21097 7432
rect 21131 7429 21143 7463
rect 21085 7423 21143 7429
rect 13538 7352 13544 7404
rect 13596 7392 13602 7404
rect 15105 7395 15163 7401
rect 15105 7392 15117 7395
rect 13596 7364 15117 7392
rect 13596 7352 13602 7364
rect 15105 7361 15117 7364
rect 15151 7392 15163 7395
rect 16301 7395 16359 7401
rect 16301 7392 16313 7395
rect 15151 7364 16313 7392
rect 15151 7361 15163 7364
rect 15105 7355 15163 7361
rect 16301 7361 16313 7364
rect 16347 7361 16359 7395
rect 16301 7355 16359 7361
rect 16577 7395 16635 7401
rect 16577 7361 16589 7395
rect 16623 7392 16635 7395
rect 16623 7364 17264 7392
rect 16623 7361 16635 7364
rect 16577 7355 16635 7361
rect 14185 7327 14243 7333
rect 14185 7324 14197 7327
rect 13096 7296 14197 7324
rect 11287 7293 11299 7296
rect 11241 7287 11299 7293
rect 14185 7293 14197 7296
rect 14231 7293 14243 7327
rect 14185 7287 14243 7293
rect 15473 7327 15531 7333
rect 15473 7293 15485 7327
rect 15519 7324 15531 7327
rect 16850 7324 16856 7336
rect 15519 7296 16856 7324
rect 15519 7293 15531 7296
rect 15473 7287 15531 7293
rect 16850 7284 16856 7296
rect 16908 7284 16914 7336
rect 17034 7284 17040 7336
rect 17092 7324 17098 7336
rect 17129 7327 17187 7333
rect 17129 7324 17141 7327
rect 17092 7296 17141 7324
rect 17092 7284 17098 7296
rect 17129 7293 17141 7296
rect 17175 7293 17187 7327
rect 17236 7324 17264 7364
rect 18892 7364 20116 7392
rect 18892 7324 18920 7364
rect 19058 7324 19064 7336
rect 17236 7296 18920 7324
rect 19019 7296 19064 7324
rect 17129 7287 17187 7293
rect 19058 7284 19064 7296
rect 19116 7284 19122 7336
rect 20088 7324 20116 7364
rect 20162 7352 20168 7404
rect 20220 7392 20226 7404
rect 20257 7395 20315 7401
rect 20257 7392 20269 7395
rect 20220 7364 20269 7392
rect 20220 7352 20226 7364
rect 20257 7361 20269 7364
rect 20303 7361 20315 7395
rect 20257 7355 20315 7361
rect 21266 7324 21272 7336
rect 20088 7296 21272 7324
rect 21266 7284 21272 7296
rect 21324 7284 21330 7336
rect 8754 7256 8760 7268
rect 8496 7228 8760 7256
rect 7990 7219 8048 7225
rect 3878 7188 3884 7200
rect 1636 7160 3556 7188
rect 3839 7160 3884 7188
rect 1636 7148 1642 7160
rect 3878 7148 3884 7160
rect 3936 7148 3942 7200
rect 4982 7188 4988 7200
rect 4943 7160 4988 7188
rect 4982 7148 4988 7160
rect 5040 7148 5046 7200
rect 5629 7191 5687 7197
rect 5629 7157 5641 7191
rect 5675 7188 5687 7191
rect 6086 7188 6092 7200
rect 5675 7160 6092 7188
rect 5675 7157 5687 7160
rect 5629 7151 5687 7157
rect 6086 7148 6092 7160
rect 6144 7148 6150 7200
rect 6454 7188 6460 7200
rect 6415 7160 6460 7188
rect 6454 7148 6460 7160
rect 6512 7148 6518 7200
rect 7285 7191 7343 7197
rect 7285 7157 7297 7191
rect 7331 7188 7343 7191
rect 7374 7188 7380 7200
rect 7331 7160 7380 7188
rect 7331 7157 7343 7160
rect 7285 7151 7343 7157
rect 7374 7148 7380 7160
rect 7432 7148 7438 7200
rect 7742 7148 7748 7200
rect 7800 7188 7806 7200
rect 8005 7188 8033 7219
rect 8754 7216 8760 7228
rect 8812 7256 8818 7268
rect 9582 7256 9588 7268
rect 8812 7228 9588 7256
rect 8812 7216 8818 7228
rect 9582 7216 9588 7228
rect 9640 7216 9646 7268
rect 9674 7216 9680 7268
rect 9732 7256 9738 7268
rect 10137 7259 10195 7265
rect 10137 7256 10149 7259
rect 9732 7228 10149 7256
rect 9732 7216 9738 7228
rect 10137 7225 10149 7228
rect 10183 7225 10195 7259
rect 10137 7219 10195 7225
rect 10321 7259 10379 7265
rect 10321 7225 10333 7259
rect 10367 7256 10379 7259
rect 16574 7256 16580 7268
rect 10367 7228 16580 7256
rect 10367 7225 10379 7228
rect 10321 7219 10379 7225
rect 16574 7216 16580 7228
rect 16632 7216 16638 7268
rect 16666 7216 16672 7268
rect 16724 7256 16730 7268
rect 17374 7259 17432 7265
rect 17374 7256 17386 7259
rect 16724 7228 17386 7256
rect 16724 7216 16730 7228
rect 17374 7225 17386 7228
rect 17420 7225 17432 7259
rect 17374 7219 17432 7225
rect 17512 7228 19840 7256
rect 7800 7160 8033 7188
rect 7800 7148 7806 7160
rect 9214 7148 9220 7200
rect 9272 7188 9278 7200
rect 9769 7191 9827 7197
rect 9769 7188 9781 7191
rect 9272 7160 9781 7188
rect 9272 7148 9278 7160
rect 9769 7157 9781 7160
rect 9815 7157 9827 7191
rect 9769 7151 9827 7157
rect 9953 7191 10011 7197
rect 9953 7157 9965 7191
rect 9999 7188 10011 7191
rect 10597 7191 10655 7197
rect 10597 7188 10609 7191
rect 9999 7160 10609 7188
rect 9999 7157 10011 7160
rect 9953 7151 10011 7157
rect 10597 7157 10609 7160
rect 10643 7188 10655 7191
rect 10870 7188 10876 7200
rect 10643 7160 10876 7188
rect 10643 7157 10655 7160
rect 10597 7151 10655 7157
rect 10870 7148 10876 7160
rect 10928 7148 10934 7200
rect 11054 7148 11060 7200
rect 11112 7188 11118 7200
rect 11701 7191 11759 7197
rect 11701 7188 11713 7191
rect 11112 7160 11713 7188
rect 11112 7148 11118 7160
rect 11701 7157 11713 7160
rect 11747 7157 11759 7191
rect 12342 7188 12348 7200
rect 12303 7160 12348 7188
rect 11701 7151 11759 7157
rect 12342 7148 12348 7160
rect 12400 7148 12406 7200
rect 12434 7148 12440 7200
rect 12492 7188 12498 7200
rect 12713 7191 12771 7197
rect 12713 7188 12725 7191
rect 12492 7160 12725 7188
rect 12492 7148 12498 7160
rect 12713 7157 12725 7160
rect 12759 7157 12771 7191
rect 14642 7188 14648 7200
rect 14603 7160 14648 7188
rect 12713 7151 12771 7157
rect 14642 7148 14648 7160
rect 14700 7148 14706 7200
rect 15841 7191 15899 7197
rect 15841 7157 15853 7191
rect 15887 7188 15899 7191
rect 16206 7188 16212 7200
rect 15887 7160 16212 7188
rect 15887 7157 15899 7160
rect 15841 7151 15899 7157
rect 16206 7148 16212 7160
rect 16264 7148 16270 7200
rect 16301 7191 16359 7197
rect 16301 7157 16313 7191
rect 16347 7188 16359 7191
rect 17512 7188 17540 7228
rect 18874 7188 18880 7200
rect 16347 7160 17540 7188
rect 18835 7160 18880 7188
rect 16347 7157 16359 7160
rect 16301 7151 16359 7157
rect 18874 7148 18880 7160
rect 18932 7148 18938 7200
rect 18966 7148 18972 7200
rect 19024 7188 19030 7200
rect 19337 7191 19395 7197
rect 19337 7188 19349 7191
rect 19024 7160 19349 7188
rect 19024 7148 19030 7160
rect 19337 7157 19349 7160
rect 19383 7157 19395 7191
rect 19702 7188 19708 7200
rect 19663 7160 19708 7188
rect 19337 7151 19395 7157
rect 19702 7148 19708 7160
rect 19760 7148 19766 7200
rect 19812 7188 19840 7228
rect 19886 7216 19892 7268
rect 19944 7256 19950 7268
rect 20165 7259 20223 7265
rect 20165 7256 20177 7259
rect 19944 7228 20177 7256
rect 19944 7216 19950 7228
rect 20165 7225 20177 7228
rect 20211 7225 20223 7259
rect 20165 7219 20223 7225
rect 20073 7191 20131 7197
rect 20073 7188 20085 7191
rect 19812 7160 20085 7188
rect 20073 7157 20085 7160
rect 20119 7157 20131 7191
rect 20073 7151 20131 7157
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 2774 6944 2780 6996
rect 2832 6984 2838 6996
rect 2832 6956 2877 6984
rect 2832 6944 2838 6956
rect 3326 6944 3332 6996
rect 3384 6984 3390 6996
rect 3384 6956 3648 6984
rect 3384 6944 3390 6956
rect 1949 6919 2007 6925
rect 1949 6885 1961 6919
rect 1995 6916 2007 6919
rect 3510 6916 3516 6928
rect 1995 6888 3516 6916
rect 1995 6885 2007 6888
rect 1949 6879 2007 6885
rect 3510 6876 3516 6888
rect 3568 6876 3574 6928
rect 2314 6808 2320 6860
rect 2372 6848 2378 6860
rect 2685 6851 2743 6857
rect 2685 6848 2697 6851
rect 2372 6820 2697 6848
rect 2372 6808 2378 6820
rect 2685 6817 2697 6820
rect 2731 6848 2743 6851
rect 3142 6848 3148 6860
rect 2731 6820 3148 6848
rect 2731 6817 2743 6820
rect 2685 6811 2743 6817
rect 3142 6808 3148 6820
rect 3200 6808 3206 6860
rect 3337 6851 3395 6857
rect 3337 6817 3349 6851
rect 3383 6848 3395 6851
rect 3620 6848 3648 6956
rect 3694 6944 3700 6996
rect 3752 6984 3758 6996
rect 4062 6984 4068 6996
rect 3752 6956 4068 6984
rect 3752 6944 3758 6956
rect 4062 6944 4068 6956
rect 4120 6944 4126 6996
rect 5718 6944 5724 6996
rect 5776 6984 5782 6996
rect 5813 6987 5871 6993
rect 5813 6984 5825 6987
rect 5776 6956 5825 6984
rect 5776 6944 5782 6956
rect 5813 6953 5825 6956
rect 5859 6953 5871 6987
rect 7742 6984 7748 6996
rect 7703 6956 7748 6984
rect 5813 6947 5871 6953
rect 7742 6944 7748 6956
rect 7800 6944 7806 6996
rect 8294 6944 8300 6996
rect 8352 6984 8358 6996
rect 8389 6987 8447 6993
rect 8389 6984 8401 6987
rect 8352 6956 8401 6984
rect 8352 6944 8358 6956
rect 8389 6953 8401 6956
rect 8435 6953 8447 6987
rect 8389 6947 8447 6953
rect 8478 6944 8484 6996
rect 8536 6984 8542 6996
rect 12342 6984 12348 6996
rect 8536 6956 9674 6984
rect 12303 6956 12348 6984
rect 8536 6944 8542 6956
rect 4430 6876 4436 6928
rect 4488 6916 4494 6928
rect 4678 6919 4736 6925
rect 4678 6916 4690 6919
rect 4488 6888 4690 6916
rect 4488 6876 4494 6888
rect 4678 6885 4690 6888
rect 4724 6885 4736 6919
rect 9646 6916 9674 6956
rect 12342 6944 12348 6956
rect 12400 6944 12406 6996
rect 16666 6984 16672 6996
rect 16627 6956 16672 6984
rect 16666 6944 16672 6956
rect 16724 6944 16730 6996
rect 17586 6984 17592 6996
rect 17547 6956 17592 6984
rect 17586 6944 17592 6956
rect 17644 6944 17650 6996
rect 18138 6984 18144 6996
rect 17972 6956 18144 6984
rect 12434 6916 12440 6928
rect 9646 6888 12440 6916
rect 4678 6879 4736 6885
rect 12434 6876 12440 6888
rect 12492 6876 12498 6928
rect 15488 6888 15976 6916
rect 6362 6848 6368 6860
rect 3383 6820 3648 6848
rect 6323 6820 6368 6848
rect 3383 6817 3395 6820
rect 3337 6811 3395 6817
rect 6362 6808 6368 6820
rect 6420 6808 6426 6860
rect 6638 6857 6644 6860
rect 6632 6848 6644 6857
rect 6599 6820 6644 6848
rect 6632 6811 6644 6820
rect 6638 6808 6644 6811
rect 6696 6808 6702 6860
rect 7558 6808 7564 6860
rect 7616 6848 7622 6860
rect 9493 6851 9551 6857
rect 9493 6848 9505 6851
rect 7616 6820 9505 6848
rect 7616 6808 7622 6820
rect 9493 6817 9505 6820
rect 9539 6817 9551 6851
rect 9493 6811 9551 6817
rect 9582 6808 9588 6860
rect 9640 6848 9646 6860
rect 10229 6851 10287 6857
rect 10229 6848 10241 6851
rect 9640 6820 10241 6848
rect 9640 6808 9646 6820
rect 10229 6817 10241 6820
rect 10275 6817 10287 6851
rect 10229 6811 10287 6817
rect 10496 6851 10554 6857
rect 10496 6817 10508 6851
rect 10542 6848 10554 6851
rect 10778 6848 10784 6860
rect 10542 6820 10784 6848
rect 10542 6817 10554 6820
rect 10496 6811 10554 6817
rect 10778 6808 10784 6820
rect 10836 6848 10842 6860
rect 10836 6820 11284 6848
rect 10836 6808 10842 6820
rect 2041 6783 2099 6789
rect 2041 6749 2053 6783
rect 2087 6749 2099 6783
rect 2041 6743 2099 6749
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6780 2283 6783
rect 3050 6780 3056 6792
rect 2271 6752 3056 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 2056 6712 2084 6743
rect 3050 6740 3056 6752
rect 3108 6740 3114 6792
rect 3786 6740 3792 6792
rect 3844 6780 3850 6792
rect 4433 6783 4491 6789
rect 4433 6780 4445 6783
rect 3844 6752 4445 6780
rect 3844 6740 3850 6752
rect 4433 6749 4445 6752
rect 4479 6749 4491 6783
rect 4433 6743 4491 6749
rect 7742 6740 7748 6792
rect 7800 6780 7806 6792
rect 8113 6783 8171 6789
rect 8113 6780 8125 6783
rect 7800 6752 8125 6780
rect 7800 6740 7806 6752
rect 8113 6749 8125 6752
rect 8159 6749 8171 6783
rect 8294 6780 8300 6792
rect 8255 6752 8300 6780
rect 8113 6743 8171 6749
rect 8294 6740 8300 6752
rect 8352 6740 8358 6792
rect 8386 6740 8392 6792
rect 8444 6780 8450 6792
rect 9030 6780 9036 6792
rect 8444 6752 9036 6780
rect 8444 6740 8450 6752
rect 9030 6740 9036 6752
rect 9088 6740 9094 6792
rect 9122 6740 9128 6792
rect 9180 6780 9186 6792
rect 9861 6783 9919 6789
rect 9861 6780 9873 6783
rect 9180 6752 9873 6780
rect 9180 6740 9186 6752
rect 9861 6749 9873 6752
rect 9907 6749 9919 6783
rect 11256 6780 11284 6820
rect 11790 6808 11796 6860
rect 11848 6848 11854 6860
rect 12253 6851 12311 6857
rect 12253 6848 12265 6851
rect 11848 6820 12265 6848
rect 11848 6808 11854 6820
rect 12253 6817 12265 6820
rect 12299 6817 12311 6851
rect 12253 6811 12311 6817
rect 14645 6851 14703 6857
rect 14645 6817 14657 6851
rect 14691 6848 14703 6851
rect 15488 6848 15516 6888
rect 14691 6820 15516 6848
rect 15556 6851 15614 6857
rect 14691 6817 14703 6820
rect 14645 6811 14703 6817
rect 15556 6817 15568 6851
rect 15602 6848 15614 6851
rect 15838 6848 15844 6860
rect 15602 6820 15844 6848
rect 15602 6817 15614 6820
rect 15556 6811 15614 6817
rect 15838 6808 15844 6820
rect 15896 6808 15902 6860
rect 15948 6848 15976 6888
rect 16206 6876 16212 6928
rect 16264 6916 16270 6928
rect 17972 6916 18000 6956
rect 18138 6944 18144 6956
rect 18196 6944 18202 6996
rect 19058 6944 19064 6996
rect 19116 6984 19122 6996
rect 19245 6987 19303 6993
rect 19245 6984 19257 6987
rect 19116 6956 19257 6984
rect 19116 6944 19122 6956
rect 19245 6953 19257 6956
rect 19291 6953 19303 6987
rect 19245 6947 19303 6953
rect 18966 6916 18972 6928
rect 16264 6888 18000 6916
rect 18064 6888 18972 6916
rect 16264 6876 16270 6888
rect 16482 6848 16488 6860
rect 15948 6820 16488 6848
rect 16482 6808 16488 6820
rect 16540 6808 16546 6860
rect 17586 6808 17592 6860
rect 17644 6848 17650 6860
rect 18064 6857 18092 6888
rect 18966 6876 18972 6888
rect 19024 6876 19030 6928
rect 20064 6919 20122 6925
rect 20064 6885 20076 6919
rect 20110 6916 20122 6919
rect 20162 6916 20168 6928
rect 20110 6888 20168 6916
rect 20110 6885 20122 6888
rect 20064 6879 20122 6885
rect 20162 6876 20168 6888
rect 20220 6876 20226 6928
rect 22002 6916 22008 6928
rect 21963 6888 22008 6916
rect 22002 6876 22008 6888
rect 22060 6876 22066 6928
rect 17773 6851 17831 6857
rect 17773 6848 17785 6851
rect 17644 6820 17785 6848
rect 17644 6808 17650 6820
rect 17773 6817 17785 6820
rect 17819 6817 17831 6851
rect 17773 6811 17831 6817
rect 18049 6851 18107 6857
rect 18049 6817 18061 6851
rect 18095 6817 18107 6851
rect 18049 6811 18107 6817
rect 18877 6851 18935 6857
rect 18877 6817 18889 6851
rect 18923 6848 18935 6851
rect 19150 6848 19156 6860
rect 18923 6820 19156 6848
rect 18923 6817 18935 6820
rect 18877 6811 18935 6817
rect 19150 6808 19156 6820
rect 19208 6808 19214 6860
rect 19797 6851 19855 6857
rect 19797 6817 19809 6851
rect 19843 6848 19855 6851
rect 21174 6848 21180 6860
rect 19843 6820 21180 6848
rect 19843 6817 19855 6820
rect 19797 6811 19855 6817
rect 21174 6808 21180 6820
rect 21232 6808 21238 6860
rect 12437 6783 12495 6789
rect 12437 6780 12449 6783
rect 11256 6752 12449 6780
rect 9861 6743 9919 6749
rect 12437 6749 12449 6752
rect 12483 6749 12495 6783
rect 12437 6743 12495 6749
rect 14550 6740 14556 6792
rect 14608 6780 14614 6792
rect 15102 6780 15108 6792
rect 14608 6752 15108 6780
rect 14608 6740 14614 6752
rect 15102 6740 15108 6752
rect 15160 6780 15166 6792
rect 15289 6783 15347 6789
rect 15289 6780 15301 6783
rect 15160 6752 15301 6780
rect 15160 6740 15166 6752
rect 15289 6749 15301 6752
rect 15335 6749 15347 6783
rect 15289 6743 15347 6749
rect 17221 6783 17279 6789
rect 17221 6749 17233 6783
rect 17267 6780 17279 6783
rect 17494 6780 17500 6792
rect 17267 6752 17500 6780
rect 17267 6749 17279 6752
rect 17221 6743 17279 6749
rect 17494 6740 17500 6752
rect 17552 6740 17558 6792
rect 18693 6783 18751 6789
rect 18693 6749 18705 6783
rect 18739 6749 18751 6783
rect 18693 6743 18751 6749
rect 18785 6783 18843 6789
rect 18785 6749 18797 6783
rect 18831 6780 18843 6783
rect 19702 6780 19708 6792
rect 18831 6752 19708 6780
rect 18831 6749 18843 6752
rect 18785 6743 18843 6749
rect 3145 6715 3203 6721
rect 3145 6712 3157 6715
rect 2056 6684 3157 6712
rect 3145 6681 3157 6684
rect 3191 6681 3203 6715
rect 3145 6675 3203 6681
rect 8757 6715 8815 6721
rect 8757 6681 8769 6715
rect 8803 6712 8815 6715
rect 12618 6712 12624 6724
rect 8803 6684 10272 6712
rect 8803 6681 8815 6684
rect 8757 6675 8815 6681
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 1854 6644 1860 6656
rect 1627 6616 1860 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 1854 6604 1860 6616
rect 1912 6604 1918 6656
rect 3694 6604 3700 6656
rect 3752 6644 3758 6656
rect 3881 6647 3939 6653
rect 3881 6644 3893 6647
rect 3752 6616 3893 6644
rect 3752 6604 3758 6616
rect 3881 6613 3893 6616
rect 3927 6613 3939 6647
rect 3881 6607 3939 6613
rect 4246 6604 4252 6656
rect 4304 6644 4310 6656
rect 4798 6644 4804 6656
rect 4304 6616 4804 6644
rect 4304 6604 4310 6616
rect 4798 6604 4804 6616
rect 4856 6604 4862 6656
rect 5718 6604 5724 6656
rect 5776 6644 5782 6656
rect 6638 6644 6644 6656
rect 5776 6616 6644 6644
rect 5776 6604 5782 6616
rect 6638 6604 6644 6616
rect 6696 6604 6702 6656
rect 7098 6604 7104 6656
rect 7156 6644 7162 6656
rect 9125 6647 9183 6653
rect 9125 6644 9137 6647
rect 7156 6616 9137 6644
rect 7156 6604 7162 6616
rect 9125 6613 9137 6616
rect 9171 6613 9183 6647
rect 10244 6644 10272 6684
rect 11164 6684 12624 6712
rect 11164 6644 11192 6684
rect 12618 6672 12624 6684
rect 12676 6672 12682 6724
rect 18708 6712 18736 6743
rect 19702 6740 19708 6752
rect 19760 6740 19766 6792
rect 18708 6684 19840 6712
rect 10244 6616 11192 6644
rect 11609 6647 11667 6653
rect 9125 6607 9183 6613
rect 11609 6613 11621 6647
rect 11655 6644 11667 6647
rect 11698 6644 11704 6656
rect 11655 6616 11704 6644
rect 11655 6613 11667 6616
rect 11609 6607 11667 6613
rect 11698 6604 11704 6616
rect 11756 6604 11762 6656
rect 11885 6647 11943 6653
rect 11885 6613 11897 6647
rect 11931 6644 11943 6647
rect 12158 6644 12164 6656
rect 11931 6616 12164 6644
rect 11931 6613 11943 6616
rect 11885 6607 11943 6613
rect 12158 6604 12164 6616
rect 12216 6604 12222 6656
rect 13170 6644 13176 6656
rect 13131 6616 13176 6644
rect 13170 6604 13176 6616
rect 13228 6604 13234 6656
rect 13630 6644 13636 6656
rect 13591 6616 13636 6644
rect 13630 6604 13636 6616
rect 13688 6604 13694 6656
rect 15013 6647 15071 6653
rect 15013 6613 15025 6647
rect 15059 6644 15071 6647
rect 15562 6644 15568 6656
rect 15059 6616 15568 6644
rect 15059 6613 15071 6616
rect 15013 6607 15071 6613
rect 15562 6604 15568 6616
rect 15620 6604 15626 6656
rect 18233 6647 18291 6653
rect 18233 6613 18245 6647
rect 18279 6644 18291 6647
rect 19058 6644 19064 6656
rect 18279 6616 19064 6644
rect 18279 6613 18291 6616
rect 18233 6607 18291 6613
rect 19058 6604 19064 6616
rect 19116 6604 19122 6656
rect 19812 6644 19840 6684
rect 21082 6644 21088 6656
rect 19812 6616 21088 6644
rect 21082 6604 21088 6616
rect 21140 6644 21146 6656
rect 21177 6647 21235 6653
rect 21177 6644 21189 6647
rect 21140 6616 21189 6644
rect 21140 6604 21146 6616
rect 21177 6613 21189 6616
rect 21223 6613 21235 6647
rect 21177 6607 21235 6613
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 3234 6400 3240 6452
rect 3292 6440 3298 6452
rect 3973 6443 4031 6449
rect 3973 6440 3985 6443
rect 3292 6412 3985 6440
rect 3292 6400 3298 6412
rect 3973 6409 3985 6412
rect 4019 6409 4031 6443
rect 3973 6403 4031 6409
rect 4154 6400 4160 6452
rect 4212 6440 4218 6452
rect 4893 6443 4951 6449
rect 4893 6440 4905 6443
rect 4212 6412 4905 6440
rect 4212 6400 4218 6412
rect 4893 6409 4905 6412
rect 4939 6409 4951 6443
rect 4893 6403 4951 6409
rect 6089 6443 6147 6449
rect 6089 6409 6101 6443
rect 6135 6440 6147 6443
rect 8294 6440 8300 6452
rect 6135 6412 8300 6440
rect 6135 6409 6147 6412
rect 6089 6403 6147 6409
rect 8294 6400 8300 6412
rect 8352 6400 8358 6452
rect 11517 6443 11575 6449
rect 11517 6440 11529 6443
rect 8404 6412 11529 6440
rect 4433 6375 4491 6381
rect 4433 6341 4445 6375
rect 4479 6372 4491 6375
rect 4798 6372 4804 6384
rect 4479 6344 4804 6372
rect 4479 6341 4491 6344
rect 4433 6335 4491 6341
rect 4798 6332 4804 6344
rect 4856 6332 4862 6384
rect 6362 6332 6368 6384
rect 6420 6372 6426 6384
rect 6420 6344 6684 6372
rect 6420 6332 6426 6344
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6304 1731 6307
rect 2314 6304 2320 6316
rect 1719 6276 2320 6304
rect 1719 6273 1731 6276
rect 1673 6267 1731 6273
rect 2314 6264 2320 6276
rect 2372 6264 2378 6316
rect 3050 6304 3056 6316
rect 3011 6276 3056 6304
rect 3050 6264 3056 6276
rect 3108 6264 3114 6316
rect 3510 6304 3516 6316
rect 3471 6276 3516 6304
rect 3510 6264 3516 6276
rect 3568 6264 3574 6316
rect 4246 6304 4252 6316
rect 4159 6276 4252 6304
rect 1854 6236 1860 6248
rect 1815 6208 1860 6236
rect 1854 6196 1860 6208
rect 1912 6196 1918 6248
rect 1946 6196 1952 6248
rect 2004 6236 2010 6248
rect 4172 6245 4200 6276
rect 4246 6264 4252 6276
rect 4304 6304 4310 6316
rect 5350 6304 5356 6316
rect 4304 6276 5356 6304
rect 4304 6264 4310 6276
rect 5350 6264 5356 6276
rect 5408 6264 5414 6316
rect 5537 6307 5595 6313
rect 5537 6273 5549 6307
rect 5583 6304 5595 6307
rect 5718 6304 5724 6316
rect 5583 6276 5724 6304
rect 5583 6273 5595 6276
rect 5537 6267 5595 6273
rect 5718 6264 5724 6276
rect 5776 6264 5782 6316
rect 2869 6239 2927 6245
rect 2869 6236 2881 6239
rect 2004 6208 2881 6236
rect 2004 6196 2010 6208
rect 2869 6205 2881 6208
rect 2915 6205 2927 6239
rect 2869 6199 2927 6205
rect 4157 6239 4215 6245
rect 4157 6205 4169 6239
rect 4203 6205 4215 6239
rect 4157 6199 4215 6205
rect 4617 6239 4675 6245
rect 4617 6205 4629 6239
rect 4663 6205 4675 6239
rect 4617 6199 4675 6205
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6236 4767 6239
rect 5077 6239 5135 6245
rect 5077 6236 5089 6239
rect 4755 6208 5089 6236
rect 4755 6205 4767 6208
rect 4709 6199 4767 6205
rect 5077 6205 5089 6208
rect 5123 6236 5135 6239
rect 6546 6236 6552 6248
rect 5123 6208 6552 6236
rect 5123 6205 5135 6208
rect 5077 6199 5135 6205
rect 1765 6171 1823 6177
rect 1765 6137 1777 6171
rect 1811 6168 1823 6171
rect 1811 6140 2544 6168
rect 1811 6137 1823 6140
rect 1765 6131 1823 6137
rect 2222 6100 2228 6112
rect 2183 6072 2228 6100
rect 2222 6060 2228 6072
rect 2280 6060 2286 6112
rect 2516 6109 2544 6140
rect 3510 6128 3516 6180
rect 3568 6168 3574 6180
rect 4632 6168 4660 6199
rect 6546 6196 6552 6208
rect 6604 6196 6610 6248
rect 6656 6236 6684 6344
rect 6730 6332 6736 6384
rect 6788 6372 6794 6384
rect 8404 6372 8432 6412
rect 11517 6409 11529 6412
rect 11563 6409 11575 6443
rect 11517 6403 11575 6409
rect 12894 6400 12900 6452
rect 12952 6440 12958 6452
rect 19981 6443 20039 6449
rect 19981 6440 19993 6443
rect 12952 6412 19993 6440
rect 12952 6400 12958 6412
rect 19981 6409 19993 6412
rect 20027 6409 20039 6443
rect 19981 6403 20039 6409
rect 6788 6344 8432 6372
rect 6788 6332 6794 6344
rect 10318 6332 10324 6384
rect 10376 6372 10382 6384
rect 10376 6344 15792 6372
rect 10376 6332 10382 6344
rect 7285 6307 7343 6313
rect 7285 6273 7297 6307
rect 7331 6304 7343 6307
rect 7742 6304 7748 6316
rect 7331 6276 7748 6304
rect 7331 6273 7343 6276
rect 7285 6267 7343 6273
rect 7742 6264 7748 6276
rect 7800 6264 7806 6316
rect 13354 6304 13360 6316
rect 13267 6276 13360 6304
rect 13354 6264 13360 6276
rect 13412 6304 13418 6316
rect 14737 6307 14795 6313
rect 14737 6304 14749 6307
rect 13412 6276 14749 6304
rect 13412 6264 13418 6276
rect 14737 6273 14749 6276
rect 14783 6273 14795 6307
rect 14737 6267 14795 6273
rect 6822 6236 6828 6248
rect 6656 6208 6828 6236
rect 6822 6196 6828 6208
rect 6880 6236 6886 6248
rect 7009 6239 7067 6245
rect 7009 6236 7021 6239
rect 6880 6208 7021 6236
rect 6880 6196 6886 6208
rect 7009 6205 7021 6208
rect 7055 6205 7067 6239
rect 7009 6199 7067 6205
rect 7101 6239 7159 6245
rect 7101 6205 7113 6239
rect 7147 6236 7159 6239
rect 8386 6236 8392 6248
rect 7147 6208 8392 6236
rect 7147 6205 7159 6208
rect 7101 6199 7159 6205
rect 8386 6196 8392 6208
rect 8444 6196 8450 6248
rect 9030 6196 9036 6248
rect 9088 6236 9094 6248
rect 9582 6236 9588 6248
rect 9088 6208 9588 6236
rect 9088 6196 9094 6208
rect 9582 6196 9588 6208
rect 9640 6236 9646 6248
rect 9677 6239 9735 6245
rect 9677 6236 9689 6239
rect 9640 6208 9689 6236
rect 9640 6196 9646 6208
rect 9677 6205 9689 6208
rect 9723 6205 9735 6239
rect 9677 6199 9735 6205
rect 9766 6196 9772 6248
rect 9824 6236 9830 6248
rect 13449 6239 13507 6245
rect 13449 6236 13461 6239
rect 9824 6208 13461 6236
rect 9824 6196 9830 6208
rect 13449 6205 13461 6208
rect 13495 6205 13507 6239
rect 13449 6199 13507 6205
rect 13998 6196 14004 6248
rect 14056 6236 14062 6248
rect 14645 6239 14703 6245
rect 14645 6236 14657 6239
rect 14056 6208 14657 6236
rect 14056 6196 14062 6208
rect 14645 6205 14657 6208
rect 14691 6205 14703 6239
rect 15764 6236 15792 6344
rect 15838 6332 15844 6384
rect 15896 6372 15902 6384
rect 17218 6372 17224 6384
rect 15896 6344 17224 6372
rect 15896 6332 15902 6344
rect 17218 6332 17224 6344
rect 17276 6372 17282 6384
rect 18325 6375 18383 6381
rect 17276 6344 17724 6372
rect 17276 6332 17282 6344
rect 16025 6307 16083 6313
rect 16025 6273 16037 6307
rect 16071 6304 16083 6307
rect 16666 6304 16672 6316
rect 16071 6276 16672 6304
rect 16071 6273 16083 6276
rect 16025 6267 16083 6273
rect 16666 6264 16672 6276
rect 16724 6264 16730 6316
rect 17402 6264 17408 6316
rect 17460 6304 17466 6316
rect 17696 6313 17724 6344
rect 18325 6341 18337 6375
rect 18371 6372 18383 6375
rect 18690 6372 18696 6384
rect 18371 6344 18696 6372
rect 18371 6341 18383 6344
rect 18325 6335 18383 6341
rect 18690 6332 18696 6344
rect 18748 6332 18754 6384
rect 18782 6332 18788 6384
rect 18840 6372 18846 6384
rect 19426 6372 19432 6384
rect 18840 6344 19432 6372
rect 18840 6332 18846 6344
rect 19426 6332 19432 6344
rect 19484 6332 19490 6384
rect 17589 6307 17647 6313
rect 17589 6304 17601 6307
rect 17460 6276 17601 6304
rect 17460 6264 17466 6276
rect 17589 6273 17601 6276
rect 17635 6273 17647 6307
rect 17589 6267 17647 6273
rect 17681 6307 17739 6313
rect 17681 6273 17693 6307
rect 17727 6273 17739 6307
rect 17681 6267 17739 6273
rect 18046 6264 18052 6316
rect 18104 6304 18110 6316
rect 18414 6304 18420 6316
rect 18104 6276 18420 6304
rect 18104 6264 18110 6276
rect 18414 6264 18420 6276
rect 18472 6264 18478 6316
rect 18506 6264 18512 6316
rect 18564 6304 18570 6316
rect 18564 6276 18828 6304
rect 18564 6264 18570 6276
rect 17310 6236 17316 6248
rect 15764 6208 17316 6236
rect 14645 6199 14703 6205
rect 17310 6196 17316 6208
rect 17368 6196 17374 6248
rect 17494 6236 17500 6248
rect 17455 6208 17500 6236
rect 17494 6196 17500 6208
rect 17552 6196 17558 6248
rect 18141 6239 18199 6245
rect 18141 6205 18153 6239
rect 18187 6236 18199 6239
rect 18598 6236 18604 6248
rect 18187 6208 18604 6236
rect 18187 6205 18199 6208
rect 18141 6199 18199 6205
rect 18598 6196 18604 6208
rect 18656 6196 18662 6248
rect 18800 6245 18828 6276
rect 19150 6264 19156 6316
rect 19208 6304 19214 6316
rect 19521 6307 19579 6313
rect 19521 6304 19533 6307
rect 19208 6276 19533 6304
rect 19208 6264 19214 6276
rect 19521 6273 19533 6276
rect 19567 6273 19579 6307
rect 19521 6267 19579 6273
rect 18785 6239 18843 6245
rect 18785 6205 18797 6239
rect 18831 6205 18843 6239
rect 18785 6199 18843 6205
rect 19245 6239 19303 6245
rect 19245 6205 19257 6239
rect 19291 6205 19303 6239
rect 19245 6199 19303 6205
rect 5166 6168 5172 6180
rect 3568 6140 4568 6168
rect 4632 6140 5172 6168
rect 3568 6128 3574 6140
rect 2501 6103 2559 6109
rect 2501 6069 2513 6103
rect 2547 6069 2559 6103
rect 2501 6063 2559 6069
rect 2961 6103 3019 6109
rect 2961 6069 2973 6103
rect 3007 6100 3019 6103
rect 4430 6100 4436 6112
rect 3007 6072 4436 6100
rect 3007 6069 3019 6072
rect 2961 6063 3019 6069
rect 4430 6060 4436 6072
rect 4488 6060 4494 6112
rect 4540 6100 4568 6140
rect 5166 6128 5172 6140
rect 5224 6168 5230 6180
rect 5442 6168 5448 6180
rect 5224 6140 5448 6168
rect 5224 6128 5230 6140
rect 5442 6128 5448 6140
rect 5500 6128 5506 6180
rect 5629 6171 5687 6177
rect 5629 6137 5641 6171
rect 5675 6168 5687 6171
rect 8662 6168 8668 6180
rect 5675 6140 6500 6168
rect 5675 6137 5687 6140
rect 5629 6131 5687 6137
rect 4709 6103 4767 6109
rect 4709 6100 4721 6103
rect 4540 6072 4721 6100
rect 4709 6069 4721 6072
rect 4755 6069 4767 6103
rect 5718 6100 5724 6112
rect 5679 6072 5724 6100
rect 4709 6063 4767 6069
rect 5718 6060 5724 6072
rect 5776 6060 5782 6112
rect 6472 6100 6500 6140
rect 8312 6140 8668 6168
rect 6641 6103 6699 6109
rect 6641 6100 6653 6103
rect 6472 6072 6653 6100
rect 6641 6069 6653 6072
rect 6687 6069 6699 6103
rect 6641 6063 6699 6069
rect 6822 6060 6828 6112
rect 6880 6100 6886 6112
rect 8312 6109 8340 6140
rect 8662 6128 8668 6140
rect 8720 6128 8726 6180
rect 9398 6128 9404 6180
rect 9456 6177 9462 6180
rect 9456 6168 9468 6177
rect 11517 6171 11575 6177
rect 9456 6140 9501 6168
rect 9456 6131 9468 6140
rect 11517 6137 11529 6171
rect 11563 6168 11575 6171
rect 13541 6171 13599 6177
rect 13541 6168 13553 6171
rect 11563 6140 13553 6168
rect 11563 6137 11575 6140
rect 11517 6131 11575 6137
rect 13541 6137 13553 6140
rect 13587 6137 13599 6171
rect 13541 6131 13599 6137
rect 16209 6171 16267 6177
rect 16209 6137 16221 6171
rect 16255 6168 16267 6171
rect 16255 6140 17172 6168
rect 16255 6137 16267 6140
rect 16209 6131 16267 6137
rect 9456 6128 9462 6131
rect 7653 6103 7711 6109
rect 7653 6100 7665 6103
rect 6880 6072 7665 6100
rect 6880 6060 6886 6072
rect 7653 6069 7665 6072
rect 7699 6069 7711 6103
rect 7653 6063 7711 6069
rect 8297 6103 8355 6109
rect 8297 6069 8309 6103
rect 8343 6069 8355 6103
rect 8297 6063 8355 6069
rect 8386 6060 8392 6112
rect 8444 6100 8450 6112
rect 9953 6103 10011 6109
rect 9953 6100 9965 6103
rect 8444 6072 9965 6100
rect 8444 6060 8450 6072
rect 9953 6069 9965 6072
rect 9999 6069 10011 6103
rect 10318 6100 10324 6112
rect 10279 6072 10324 6100
rect 9953 6063 10011 6069
rect 10318 6060 10324 6072
rect 10376 6060 10382 6112
rect 10778 6100 10784 6112
rect 10739 6072 10784 6100
rect 10778 6060 10784 6072
rect 10836 6060 10842 6112
rect 11238 6100 11244 6112
rect 11199 6072 11244 6100
rect 11238 6060 11244 6072
rect 11296 6060 11302 6112
rect 11790 6100 11796 6112
rect 11751 6072 11796 6100
rect 11790 6060 11796 6072
rect 11848 6060 11854 6112
rect 12250 6100 12256 6112
rect 12211 6072 12256 6100
rect 12250 6060 12256 6072
rect 12308 6060 12314 6112
rect 12710 6100 12716 6112
rect 12671 6072 12716 6100
rect 12710 6060 12716 6072
rect 12768 6060 12774 6112
rect 13906 6100 13912 6112
rect 13867 6072 13912 6100
rect 13906 6060 13912 6072
rect 13964 6060 13970 6112
rect 14182 6100 14188 6112
rect 14143 6072 14188 6100
rect 14182 6060 14188 6072
rect 14240 6060 14246 6112
rect 14550 6100 14556 6112
rect 14511 6072 14556 6100
rect 14550 6060 14556 6072
rect 14608 6060 14614 6112
rect 15565 6103 15623 6109
rect 15565 6069 15577 6103
rect 15611 6100 15623 6103
rect 15930 6100 15936 6112
rect 15611 6072 15936 6100
rect 15611 6069 15623 6072
rect 15565 6063 15623 6069
rect 15930 6060 15936 6072
rect 15988 6060 15994 6112
rect 16117 6103 16175 6109
rect 16117 6069 16129 6103
rect 16163 6100 16175 6103
rect 16298 6100 16304 6112
rect 16163 6072 16304 6100
rect 16163 6069 16175 6072
rect 16117 6063 16175 6069
rect 16298 6060 16304 6072
rect 16356 6060 16362 6112
rect 16574 6100 16580 6112
rect 16535 6072 16580 6100
rect 16574 6060 16580 6072
rect 16632 6060 16638 6112
rect 17144 6109 17172 6140
rect 17678 6128 17684 6180
rect 17736 6168 17742 6180
rect 19260 6168 19288 6199
rect 21082 6196 21088 6248
rect 21140 6245 21146 6248
rect 21140 6236 21152 6245
rect 21361 6239 21419 6245
rect 21140 6208 21185 6236
rect 21140 6199 21152 6208
rect 21361 6205 21373 6239
rect 21407 6205 21419 6239
rect 21361 6199 21419 6205
rect 21140 6196 21146 6199
rect 17736 6140 19288 6168
rect 17736 6128 17742 6140
rect 21174 6128 21180 6180
rect 21232 6168 21238 6180
rect 21376 6168 21404 6199
rect 21232 6140 21404 6168
rect 21232 6128 21238 6140
rect 17129 6103 17187 6109
rect 17129 6069 17141 6103
rect 17175 6069 17187 6103
rect 17129 6063 17187 6069
rect 18601 6103 18659 6109
rect 18601 6069 18613 6103
rect 18647 6100 18659 6103
rect 18782 6100 18788 6112
rect 18647 6072 18788 6100
rect 18647 6069 18659 6072
rect 18601 6063 18659 6069
rect 18782 6060 18788 6072
rect 18840 6060 18846 6112
rect 18966 6060 18972 6112
rect 19024 6100 19030 6112
rect 19061 6103 19119 6109
rect 19061 6100 19073 6103
rect 19024 6072 19073 6100
rect 19024 6060 19030 6072
rect 19061 6069 19073 6072
rect 19107 6069 19119 6103
rect 19061 6063 19119 6069
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 2774 5896 2780 5908
rect 2148 5868 2780 5896
rect 1670 5828 1676 5840
rect 1631 5800 1676 5828
rect 1670 5788 1676 5800
rect 1728 5788 1734 5840
rect 2148 5769 2176 5868
rect 2774 5856 2780 5868
rect 2832 5856 2838 5908
rect 3513 5899 3571 5905
rect 3513 5865 3525 5899
rect 3559 5865 3571 5899
rect 3513 5859 3571 5865
rect 5445 5899 5503 5905
rect 5445 5865 5457 5899
rect 5491 5896 5503 5899
rect 5534 5896 5540 5908
rect 5491 5868 5540 5896
rect 5491 5865 5503 5868
rect 5445 5859 5503 5865
rect 3528 5828 3556 5859
rect 5534 5856 5540 5868
rect 5592 5856 5598 5908
rect 5718 5856 5724 5908
rect 5776 5896 5782 5908
rect 6089 5899 6147 5905
rect 6089 5896 6101 5899
rect 5776 5868 6101 5896
rect 5776 5856 5782 5868
rect 6089 5865 6101 5868
rect 6135 5865 6147 5899
rect 6089 5859 6147 5865
rect 6549 5899 6607 5905
rect 6549 5865 6561 5899
rect 6595 5896 6607 5899
rect 7377 5899 7435 5905
rect 6595 5868 6868 5896
rect 6595 5865 6607 5868
rect 6549 5859 6607 5865
rect 3970 5828 3976 5840
rect 3528 5800 3976 5828
rect 3970 5788 3976 5800
rect 4028 5828 4034 5840
rect 4310 5831 4368 5837
rect 4310 5828 4322 5831
rect 4028 5800 4322 5828
rect 4028 5788 4034 5800
rect 4310 5797 4322 5800
rect 4356 5797 4368 5831
rect 5552 5828 5580 5856
rect 6840 5840 6868 5868
rect 7377 5865 7389 5899
rect 7423 5896 7435 5899
rect 7466 5896 7472 5908
rect 7423 5868 7472 5896
rect 7423 5865 7435 5868
rect 7377 5859 7435 5865
rect 7466 5856 7472 5868
rect 7524 5856 7530 5908
rect 8754 5896 8760 5908
rect 8715 5868 8760 5896
rect 8754 5856 8760 5868
rect 8812 5856 8818 5908
rect 9677 5899 9735 5905
rect 9677 5865 9689 5899
rect 9723 5896 9735 5899
rect 9766 5896 9772 5908
rect 9723 5868 9772 5896
rect 9723 5865 9735 5868
rect 9677 5859 9735 5865
rect 9766 5856 9772 5868
rect 9824 5856 9830 5908
rect 12894 5896 12900 5908
rect 9876 5868 12900 5896
rect 5552 5800 6684 5828
rect 4310 5791 4368 5797
rect 2406 5769 2412 5772
rect 2133 5763 2191 5769
rect 2133 5729 2145 5763
rect 2179 5729 2191 5763
rect 2400 5760 2412 5769
rect 2367 5732 2412 5760
rect 2133 5723 2191 5729
rect 2400 5723 2412 5732
rect 2406 5720 2412 5723
rect 2464 5720 2470 5772
rect 2774 5720 2780 5772
rect 2832 5760 2838 5772
rect 3786 5760 3792 5772
rect 2832 5732 3792 5760
rect 2832 5720 2838 5732
rect 3786 5720 3792 5732
rect 3844 5760 3850 5772
rect 4065 5763 4123 5769
rect 4065 5760 4077 5763
rect 3844 5732 4077 5760
rect 3844 5720 3850 5732
rect 4065 5729 4077 5732
rect 4111 5729 4123 5763
rect 4065 5723 4123 5729
rect 6457 5763 6515 5769
rect 6457 5729 6469 5763
rect 6503 5760 6515 5763
rect 6503 5732 6592 5760
rect 6503 5729 6515 5732
rect 6457 5723 6515 5729
rect 5534 5652 5540 5704
rect 5592 5692 5598 5704
rect 6178 5692 6184 5704
rect 5592 5664 6184 5692
rect 5592 5652 5598 5664
rect 6178 5652 6184 5664
rect 6236 5652 6242 5704
rect 6564 5624 6592 5732
rect 6656 5701 6684 5800
rect 6822 5788 6828 5840
rect 6880 5788 6886 5840
rect 9398 5828 9404 5840
rect 8312 5800 9404 5828
rect 7558 5760 7564 5772
rect 7519 5732 7564 5760
rect 7558 5720 7564 5732
rect 7616 5720 7622 5772
rect 8312 5760 8340 5800
rect 9398 5788 9404 5800
rect 9456 5828 9462 5840
rect 9876 5828 9904 5868
rect 12894 5856 12900 5868
rect 12952 5856 12958 5908
rect 14550 5896 14556 5908
rect 14511 5868 14556 5896
rect 14550 5856 14556 5868
rect 14608 5856 14614 5908
rect 15473 5899 15531 5905
rect 15473 5865 15485 5899
rect 15519 5896 15531 5899
rect 15519 5868 16160 5896
rect 15519 5865 15531 5868
rect 15473 5859 15531 5865
rect 10502 5828 10508 5840
rect 9456 5800 9904 5828
rect 10060 5800 10508 5828
rect 9456 5788 9462 5800
rect 8220 5732 8340 5760
rect 8389 5763 8447 5769
rect 6641 5695 6699 5701
rect 6641 5661 6653 5695
rect 6687 5692 6699 5695
rect 7742 5692 7748 5704
rect 6687 5664 7748 5692
rect 6687 5661 6699 5664
rect 6641 5655 6699 5661
rect 7742 5652 7748 5664
rect 7800 5652 7806 5704
rect 8220 5701 8248 5732
rect 8389 5729 8401 5763
rect 8435 5760 8447 5763
rect 9490 5760 9496 5772
rect 8435 5732 9496 5760
rect 8435 5729 8447 5732
rect 8389 5723 8447 5729
rect 9490 5720 9496 5732
rect 9548 5720 9554 5772
rect 8205 5695 8263 5701
rect 8205 5661 8217 5695
rect 8251 5661 8263 5695
rect 8205 5655 8263 5661
rect 8294 5652 8300 5704
rect 8352 5692 8358 5704
rect 9692 5692 9720 5800
rect 9769 5763 9827 5769
rect 9769 5729 9781 5763
rect 9815 5760 9827 5763
rect 10060 5760 10088 5800
rect 10502 5788 10508 5800
rect 10560 5788 10566 5840
rect 11548 5831 11606 5837
rect 11548 5797 11560 5831
rect 11594 5828 11606 5831
rect 11698 5828 11704 5840
rect 11594 5800 11704 5828
rect 11594 5797 11606 5800
rect 11548 5791 11606 5797
rect 11698 5788 11704 5800
rect 11756 5788 11762 5840
rect 16022 5828 16028 5840
rect 11808 5800 15700 5828
rect 15983 5800 16028 5828
rect 11808 5760 11836 5800
rect 9815 5732 10088 5760
rect 10152 5732 11836 5760
rect 12888 5763 12946 5769
rect 9815 5729 9827 5732
rect 9769 5723 9827 5729
rect 9861 5695 9919 5701
rect 9861 5692 9873 5695
rect 8352 5664 8397 5692
rect 8496 5664 9444 5692
rect 9692 5664 9873 5692
rect 8352 5652 8358 5664
rect 6730 5624 6736 5636
rect 5736 5596 6408 5624
rect 6564 5596 6736 5624
rect 1765 5559 1823 5565
rect 1765 5525 1777 5559
rect 1811 5556 1823 5559
rect 5736 5556 5764 5596
rect 1811 5528 5764 5556
rect 5813 5559 5871 5565
rect 1811 5525 1823 5528
rect 1765 5519 1823 5525
rect 5813 5525 5825 5559
rect 5859 5556 5871 5559
rect 6086 5556 6092 5568
rect 5859 5528 6092 5556
rect 5859 5525 5871 5528
rect 5813 5519 5871 5525
rect 6086 5516 6092 5528
rect 6144 5516 6150 5568
rect 6380 5556 6408 5596
rect 6730 5584 6736 5596
rect 6788 5624 6794 5636
rect 8496 5624 8524 5664
rect 6788 5596 8524 5624
rect 6788 5584 6794 5596
rect 8570 5584 8576 5636
rect 8628 5624 8634 5636
rect 9309 5627 9367 5633
rect 9309 5624 9321 5627
rect 8628 5596 9321 5624
rect 8628 5584 8634 5596
rect 9309 5593 9321 5596
rect 9355 5593 9367 5627
rect 9416 5624 9444 5664
rect 9861 5661 9873 5664
rect 9907 5661 9919 5695
rect 9861 5655 9919 5661
rect 10152 5624 10180 5732
rect 12888 5729 12900 5763
rect 12934 5760 12946 5763
rect 13354 5760 13360 5772
rect 12934 5732 13360 5760
rect 12934 5729 12946 5732
rect 12888 5723 12946 5729
rect 13354 5720 13360 5732
rect 13412 5720 13418 5772
rect 15289 5763 15347 5769
rect 15289 5729 15301 5763
rect 15335 5760 15347 5763
rect 15562 5760 15568 5772
rect 15335 5732 15568 5760
rect 15335 5729 15347 5732
rect 15289 5723 15347 5729
rect 15562 5720 15568 5732
rect 15620 5720 15626 5772
rect 15672 5760 15700 5800
rect 16022 5788 16028 5800
rect 16080 5788 16086 5840
rect 16132 5828 16160 5868
rect 16298 5856 16304 5908
rect 16356 5896 16362 5908
rect 16485 5899 16543 5905
rect 16485 5896 16497 5899
rect 16356 5868 16497 5896
rect 16356 5856 16362 5868
rect 16485 5865 16497 5868
rect 16531 5865 16543 5899
rect 16485 5859 16543 5865
rect 17310 5856 17316 5908
rect 17368 5896 17374 5908
rect 21177 5899 21235 5905
rect 21177 5896 21189 5899
rect 17368 5868 21189 5896
rect 17368 5856 17374 5868
rect 21177 5865 21189 5868
rect 21223 5865 21235 5899
rect 21177 5859 21235 5865
rect 17770 5828 17776 5840
rect 16132 5800 17776 5828
rect 17770 5788 17776 5800
rect 17828 5828 17834 5840
rect 18141 5831 18199 5837
rect 18141 5828 18153 5831
rect 17828 5800 18153 5828
rect 17828 5788 17834 5800
rect 18141 5797 18153 5800
rect 18187 5797 18199 5831
rect 18141 5791 18199 5797
rect 18233 5831 18291 5837
rect 18233 5797 18245 5831
rect 18279 5828 18291 5831
rect 18322 5828 18328 5840
rect 18279 5800 18328 5828
rect 18279 5797 18291 5800
rect 18233 5791 18291 5797
rect 18322 5788 18328 5800
rect 18380 5788 18386 5840
rect 20257 5831 20315 5837
rect 20257 5797 20269 5831
rect 20303 5828 20315 5831
rect 20438 5828 20444 5840
rect 20303 5800 20444 5828
rect 20303 5797 20315 5800
rect 20257 5791 20315 5797
rect 20438 5788 20444 5800
rect 20496 5788 20502 5840
rect 16117 5763 16175 5769
rect 16117 5760 16129 5763
rect 15672 5732 16129 5760
rect 16117 5729 16129 5732
rect 16163 5729 16175 5763
rect 16758 5760 16764 5772
rect 16719 5732 16764 5760
rect 16117 5723 16175 5729
rect 16758 5720 16764 5732
rect 16816 5720 16822 5772
rect 17126 5720 17132 5772
rect 17184 5760 17190 5772
rect 17221 5763 17279 5769
rect 17221 5760 17233 5763
rect 17184 5732 17233 5760
rect 17184 5720 17190 5732
rect 17221 5729 17233 5732
rect 17267 5729 17279 5763
rect 18506 5760 18512 5772
rect 17221 5723 17279 5729
rect 17696 5732 18512 5760
rect 11793 5695 11851 5701
rect 11793 5661 11805 5695
rect 11839 5661 11851 5695
rect 12066 5692 12072 5704
rect 12027 5664 12072 5692
rect 11793 5655 11851 5661
rect 11808 5624 11836 5655
rect 12066 5652 12072 5664
rect 12124 5652 12130 5704
rect 12621 5695 12679 5701
rect 12621 5661 12633 5695
rect 12667 5661 12679 5695
rect 15838 5692 15844 5704
rect 15799 5664 15844 5692
rect 12621 5655 12679 5661
rect 11882 5624 11888 5636
rect 9416 5596 10180 5624
rect 10244 5596 10916 5624
rect 11795 5596 11888 5624
rect 9309 5587 9367 5593
rect 6638 5556 6644 5568
rect 6380 5528 6644 5556
rect 6638 5516 6644 5528
rect 6696 5556 6702 5568
rect 10244 5556 10272 5596
rect 10410 5556 10416 5568
rect 6696 5528 10272 5556
rect 10371 5528 10416 5556
rect 6696 5516 6702 5528
rect 10410 5516 10416 5528
rect 10468 5516 10474 5568
rect 10888 5556 10916 5596
rect 11882 5584 11888 5596
rect 11940 5624 11946 5636
rect 12636 5624 12664 5655
rect 15838 5652 15844 5664
rect 15896 5652 15902 5704
rect 17696 5692 17724 5732
rect 18506 5720 18512 5732
rect 18564 5720 18570 5772
rect 19058 5760 19064 5772
rect 19019 5732 19064 5760
rect 19058 5720 19064 5732
rect 19116 5720 19122 5772
rect 20162 5760 20168 5772
rect 20123 5732 20168 5760
rect 20162 5720 20168 5732
rect 20220 5720 20226 5772
rect 20622 5720 20628 5772
rect 20680 5760 20686 5772
rect 21269 5763 21327 5769
rect 21269 5760 21281 5763
rect 20680 5732 21281 5760
rect 20680 5720 20686 5732
rect 21269 5729 21281 5732
rect 21315 5729 21327 5763
rect 21269 5723 21327 5729
rect 16868 5664 17724 5692
rect 11940 5596 12664 5624
rect 11940 5584 11946 5596
rect 11054 5556 11060 5568
rect 10888 5528 11060 5556
rect 11054 5516 11060 5528
rect 11112 5516 11118 5568
rect 12636 5556 12664 5596
rect 14642 5584 14648 5636
rect 14700 5624 14706 5636
rect 16868 5624 16896 5664
rect 17770 5652 17776 5704
rect 17828 5692 17834 5704
rect 17957 5695 18015 5701
rect 17957 5692 17969 5695
rect 17828 5664 17969 5692
rect 17828 5652 17834 5664
rect 17957 5661 17969 5664
rect 18003 5661 18015 5695
rect 17957 5655 18015 5661
rect 20346 5652 20352 5704
rect 20404 5692 20410 5704
rect 20404 5664 20449 5692
rect 20404 5652 20410 5664
rect 14700 5596 16896 5624
rect 16945 5627 17003 5633
rect 14700 5584 14706 5596
rect 16945 5593 16957 5627
rect 16991 5624 17003 5627
rect 18046 5624 18052 5636
rect 16991 5596 18052 5624
rect 16991 5593 17003 5596
rect 16945 5587 17003 5593
rect 18046 5584 18052 5596
rect 18104 5584 18110 5636
rect 13262 5556 13268 5568
rect 12636 5528 13268 5556
rect 13262 5516 13268 5528
rect 13320 5516 13326 5568
rect 14001 5559 14059 5565
rect 14001 5525 14013 5559
rect 14047 5556 14059 5559
rect 14090 5556 14096 5568
rect 14047 5528 14096 5556
rect 14047 5525 14059 5528
rect 14001 5519 14059 5525
rect 14090 5516 14096 5528
rect 14148 5516 14154 5568
rect 17405 5559 17463 5565
rect 17405 5525 17417 5559
rect 17451 5556 17463 5559
rect 17954 5556 17960 5568
rect 17451 5528 17960 5556
rect 17451 5525 17463 5528
rect 17405 5519 17463 5525
rect 17954 5516 17960 5528
rect 18012 5516 18018 5568
rect 18598 5556 18604 5568
rect 18559 5528 18604 5556
rect 18598 5516 18604 5528
rect 18656 5516 18662 5568
rect 19058 5516 19064 5568
rect 19116 5556 19122 5568
rect 19245 5559 19303 5565
rect 19245 5556 19257 5559
rect 19116 5528 19257 5556
rect 19116 5516 19122 5528
rect 19245 5525 19257 5528
rect 19291 5525 19303 5559
rect 19794 5556 19800 5568
rect 19755 5528 19800 5556
rect 19245 5519 19303 5525
rect 19794 5516 19800 5528
rect 19852 5516 19858 5568
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 2958 5312 2964 5364
rect 3016 5352 3022 5364
rect 7469 5355 7527 5361
rect 7469 5352 7481 5355
rect 3016 5324 7481 5352
rect 3016 5312 3022 5324
rect 7469 5321 7481 5324
rect 7515 5321 7527 5355
rect 7469 5315 7527 5321
rect 7650 5312 7656 5364
rect 7708 5352 7714 5364
rect 7745 5355 7803 5361
rect 7745 5352 7757 5355
rect 7708 5324 7757 5352
rect 7708 5312 7714 5324
rect 7745 5321 7757 5324
rect 7791 5321 7803 5355
rect 9125 5355 9183 5361
rect 7745 5315 7803 5321
rect 8312 5324 8708 5352
rect 8312 5296 8340 5324
rect 4154 5244 4160 5296
rect 4212 5284 4218 5296
rect 4433 5287 4491 5293
rect 4433 5284 4445 5287
rect 4212 5256 4445 5284
rect 4212 5244 4218 5256
rect 4433 5253 4445 5256
rect 4479 5253 4491 5287
rect 5718 5284 5724 5296
rect 5679 5256 5724 5284
rect 4433 5247 4491 5253
rect 5718 5244 5724 5256
rect 5776 5244 5782 5296
rect 6178 5244 6184 5296
rect 6236 5284 6242 5296
rect 6362 5284 6368 5296
rect 6236 5256 6368 5284
rect 6236 5244 6242 5256
rect 6362 5244 6368 5256
rect 6420 5244 6426 5296
rect 7285 5287 7343 5293
rect 7285 5253 7297 5287
rect 7331 5284 7343 5287
rect 8294 5284 8300 5296
rect 7331 5256 8300 5284
rect 7331 5253 7343 5256
rect 7285 5247 7343 5253
rect 8294 5244 8300 5256
rect 8352 5244 8358 5296
rect 8680 5284 8708 5324
rect 9125 5321 9137 5355
rect 9171 5352 9183 5355
rect 9306 5352 9312 5364
rect 9171 5324 9312 5352
rect 9171 5321 9183 5324
rect 9125 5315 9183 5321
rect 9306 5312 9312 5324
rect 9364 5312 9370 5364
rect 10410 5312 10416 5364
rect 10468 5352 10474 5364
rect 13265 5355 13323 5361
rect 10468 5324 11192 5352
rect 10468 5312 10474 5324
rect 10321 5287 10379 5293
rect 8680 5256 10272 5284
rect 2866 5216 2872 5228
rect 2827 5188 2872 5216
rect 2866 5176 2872 5188
rect 2924 5176 2930 5228
rect 3050 5216 3056 5228
rect 3011 5188 3056 5216
rect 3050 5176 3056 5188
rect 3108 5176 3114 5228
rect 3970 5216 3976 5228
rect 3931 5188 3976 5216
rect 3970 5176 3976 5188
rect 4028 5176 4034 5228
rect 8570 5216 8576 5228
rect 5092 5188 5672 5216
rect 8531 5188 8576 5216
rect 1394 5148 1400 5160
rect 1355 5120 1400 5148
rect 1394 5108 1400 5120
rect 1452 5108 1458 5160
rect 1854 5148 1860 5160
rect 1815 5120 1860 5148
rect 1854 5108 1860 5120
rect 1912 5108 1918 5160
rect 2498 5108 2504 5160
rect 2556 5108 2562 5160
rect 2682 5108 2688 5160
rect 2740 5148 2746 5160
rect 2740 5120 4016 5148
rect 2740 5108 2746 5120
rect 2130 5040 2136 5092
rect 2188 5080 2194 5092
rect 2516 5080 2544 5108
rect 2777 5083 2835 5089
rect 2777 5080 2789 5083
rect 2188 5052 2789 5080
rect 2188 5040 2194 5052
rect 2777 5049 2789 5052
rect 2823 5049 2835 5083
rect 2777 5043 2835 5049
rect 2958 5040 2964 5092
rect 3016 5080 3022 5092
rect 3881 5083 3939 5089
rect 3881 5080 3893 5083
rect 3016 5052 3893 5080
rect 3016 5040 3022 5052
rect 3881 5049 3893 5052
rect 3927 5049 3939 5083
rect 3988 5080 4016 5120
rect 4154 5108 4160 5160
rect 4212 5148 4218 5160
rect 4338 5148 4344 5160
rect 4212 5120 4344 5148
rect 4212 5108 4218 5120
rect 4338 5108 4344 5120
rect 4396 5148 4402 5160
rect 5092 5157 5120 5188
rect 4617 5151 4675 5157
rect 4617 5148 4629 5151
rect 4396 5120 4629 5148
rect 4396 5108 4402 5120
rect 4617 5117 4629 5120
rect 4663 5117 4675 5151
rect 4617 5111 4675 5117
rect 5077 5151 5135 5157
rect 5077 5117 5089 5151
rect 5123 5117 5135 5151
rect 5077 5111 5135 5117
rect 5442 5108 5448 5160
rect 5500 5148 5506 5160
rect 5537 5151 5595 5157
rect 5537 5148 5549 5151
rect 5500 5120 5549 5148
rect 5500 5108 5506 5120
rect 5537 5117 5549 5120
rect 5583 5117 5595 5151
rect 5644 5148 5672 5188
rect 8570 5176 8576 5188
rect 8628 5176 8634 5228
rect 8757 5219 8815 5225
rect 8757 5185 8769 5219
rect 8803 5216 8815 5219
rect 9769 5219 9827 5225
rect 8803 5188 8892 5216
rect 8803 5185 8815 5188
rect 8757 5179 8815 5185
rect 5810 5148 5816 5160
rect 5644 5120 5816 5148
rect 5537 5111 5595 5117
rect 5810 5108 5816 5120
rect 5868 5108 5874 5160
rect 7098 5148 7104 5160
rect 7059 5120 7104 5148
rect 7098 5108 7104 5120
rect 7156 5108 7162 5160
rect 7466 5108 7472 5160
rect 7524 5148 7530 5160
rect 7561 5151 7619 5157
rect 7561 5148 7573 5151
rect 7524 5120 7573 5148
rect 7524 5108 7530 5120
rect 7561 5117 7573 5120
rect 7607 5148 7619 5151
rect 8386 5148 8392 5160
rect 7607 5120 8392 5148
rect 7607 5117 7619 5120
rect 7561 5111 7619 5117
rect 8386 5108 8392 5120
rect 8444 5108 8450 5160
rect 5997 5083 6055 5089
rect 5997 5080 6009 5083
rect 3988 5052 6009 5080
rect 3881 5043 3939 5049
rect 5997 5049 6009 5052
rect 6043 5049 6055 5083
rect 5997 5043 6055 5049
rect 8662 5040 8668 5092
rect 8720 5080 8726 5092
rect 8864 5080 8892 5188
rect 9769 5185 9781 5219
rect 9815 5185 9827 5219
rect 10244 5216 10272 5256
rect 10321 5253 10333 5287
rect 10367 5284 10379 5287
rect 11054 5284 11060 5296
rect 10367 5256 11060 5284
rect 10367 5253 10379 5256
rect 10321 5247 10379 5253
rect 11054 5244 11060 5256
rect 11112 5244 11118 5296
rect 10244 5188 10916 5216
rect 9769 5179 9827 5185
rect 9122 5108 9128 5160
rect 9180 5148 9186 5160
rect 9309 5151 9367 5157
rect 9309 5148 9321 5151
rect 9180 5120 9321 5148
rect 9180 5108 9186 5120
rect 9309 5117 9321 5120
rect 9355 5117 9367 5151
rect 9784 5148 9812 5179
rect 10410 5148 10416 5160
rect 9784 5120 10416 5148
rect 9309 5111 9367 5117
rect 10410 5108 10416 5120
rect 10468 5108 10474 5160
rect 10505 5151 10563 5157
rect 10505 5117 10517 5151
rect 10551 5148 10563 5151
rect 10551 5120 10732 5148
rect 10551 5117 10563 5120
rect 10505 5111 10563 5117
rect 8720 5052 8892 5080
rect 9861 5083 9919 5089
rect 8720 5040 8726 5052
rect 9861 5049 9873 5083
rect 9907 5080 9919 5083
rect 9907 5052 10640 5080
rect 9907 5049 9919 5052
rect 9861 5043 9919 5049
rect 1578 5012 1584 5024
rect 1539 4984 1584 5012
rect 1578 4972 1584 4984
rect 1636 4972 1642 5024
rect 2038 5012 2044 5024
rect 1999 4984 2044 5012
rect 2038 4972 2044 4984
rect 2096 4972 2102 5024
rect 2409 5015 2467 5021
rect 2409 4981 2421 5015
rect 2455 5012 2467 5015
rect 2498 5012 2504 5024
rect 2455 4984 2504 5012
rect 2455 4981 2467 4984
rect 2409 4975 2467 4981
rect 2498 4972 2504 4984
rect 2556 4972 2562 5024
rect 3326 4972 3332 5024
rect 3384 5012 3390 5024
rect 3421 5015 3479 5021
rect 3421 5012 3433 5015
rect 3384 4984 3433 5012
rect 3384 4972 3390 4984
rect 3421 4981 3433 4984
rect 3467 4981 3479 5015
rect 3786 5012 3792 5024
rect 3747 4984 3792 5012
rect 3421 4975 3479 4981
rect 3786 4972 3792 4984
rect 3844 4972 3850 5024
rect 5258 5012 5264 5024
rect 5219 4984 5264 5012
rect 5258 4972 5264 4984
rect 5316 4972 5322 5024
rect 6825 5015 6883 5021
rect 6825 4981 6837 5015
rect 6871 5012 6883 5015
rect 7190 5012 7196 5024
rect 6871 4984 7196 5012
rect 6871 4981 6883 4984
rect 6825 4975 6883 4981
rect 7190 4972 7196 4984
rect 7248 4972 7254 5024
rect 7469 5015 7527 5021
rect 7469 4981 7481 5015
rect 7515 5012 7527 5015
rect 8113 5015 8171 5021
rect 8113 5012 8125 5015
rect 7515 4984 8125 5012
rect 7515 4981 7527 4984
rect 7469 4975 7527 4981
rect 8113 4981 8125 4984
rect 8159 4981 8171 5015
rect 8113 4975 8171 4981
rect 8481 5015 8539 5021
rect 8481 4981 8493 5015
rect 8527 5012 8539 5015
rect 8754 5012 8760 5024
rect 8527 4984 8760 5012
rect 8527 4981 8539 4984
rect 8481 4975 8539 4981
rect 8754 4972 8760 4984
rect 8812 4972 8818 5024
rect 9950 5012 9956 5024
rect 9911 4984 9956 5012
rect 9950 4972 9956 4984
rect 10008 4972 10014 5024
rect 10410 4972 10416 5024
rect 10468 5012 10474 5024
rect 10612 5021 10640 5052
rect 10505 5015 10563 5021
rect 10505 5012 10517 5015
rect 10468 4984 10517 5012
rect 10468 4972 10474 4984
rect 10505 4981 10517 4984
rect 10551 4981 10563 5015
rect 10505 4975 10563 4981
rect 10597 5015 10655 5021
rect 10597 4981 10609 5015
rect 10643 4981 10655 5015
rect 10704 5012 10732 5120
rect 10888 5080 10916 5188
rect 10962 5108 10968 5160
rect 11020 5148 11026 5160
rect 11057 5151 11115 5157
rect 11057 5148 11069 5151
rect 11020 5120 11069 5148
rect 11020 5108 11026 5120
rect 11057 5117 11069 5120
rect 11103 5117 11115 5151
rect 11164 5148 11192 5324
rect 13265 5321 13277 5355
rect 13311 5352 13323 5355
rect 13354 5352 13360 5364
rect 13311 5324 13360 5352
rect 13311 5321 13323 5324
rect 13265 5315 13323 5321
rect 13354 5312 13360 5324
rect 13412 5312 13418 5364
rect 16117 5355 16175 5361
rect 16117 5321 16129 5355
rect 16163 5352 16175 5355
rect 17678 5352 17684 5364
rect 16163 5324 17684 5352
rect 16163 5321 16175 5324
rect 16117 5315 16175 5321
rect 17678 5312 17684 5324
rect 17736 5312 17742 5364
rect 21174 5352 21180 5364
rect 19168 5324 21180 5352
rect 15838 5244 15844 5296
rect 15896 5284 15902 5296
rect 16669 5287 16727 5293
rect 16669 5284 16681 5287
rect 15896 5256 16681 5284
rect 15896 5244 15902 5256
rect 16669 5253 16681 5256
rect 16715 5253 16727 5287
rect 16669 5247 16727 5253
rect 11241 5219 11299 5225
rect 11241 5185 11253 5219
rect 11287 5216 11299 5219
rect 11698 5216 11704 5228
rect 11287 5188 11704 5216
rect 11287 5185 11299 5188
rect 11241 5179 11299 5185
rect 11698 5176 11704 5188
rect 11756 5176 11762 5228
rect 11882 5216 11888 5228
rect 11843 5188 11888 5216
rect 11882 5176 11888 5188
rect 11940 5176 11946 5228
rect 13906 5176 13912 5228
rect 13964 5216 13970 5228
rect 14001 5219 14059 5225
rect 14001 5216 14013 5219
rect 13964 5188 14013 5216
rect 13964 5176 13970 5188
rect 14001 5185 14013 5188
rect 14047 5185 14059 5219
rect 14001 5179 14059 5185
rect 14090 5176 14096 5228
rect 14148 5216 14154 5228
rect 14829 5219 14887 5225
rect 14148 5188 14193 5216
rect 14148 5176 14154 5188
rect 14829 5185 14841 5219
rect 14875 5216 14887 5219
rect 15194 5216 15200 5228
rect 14875 5188 15200 5216
rect 14875 5185 14887 5188
rect 14829 5179 14887 5185
rect 15194 5176 15200 5188
rect 15252 5216 15258 5228
rect 19168 5225 19196 5324
rect 21174 5312 21180 5324
rect 21232 5312 21238 5364
rect 19153 5219 19211 5225
rect 15252 5188 17632 5216
rect 15252 5176 15258 5188
rect 12141 5151 12199 5157
rect 12141 5148 12153 5151
rect 11164 5120 12153 5148
rect 11057 5111 11115 5117
rect 12141 5117 12153 5120
rect 12187 5117 12199 5151
rect 14921 5151 14979 5157
rect 14921 5148 14933 5151
rect 12141 5111 12199 5117
rect 12268 5120 14933 5148
rect 12268 5080 12296 5120
rect 14921 5117 14933 5120
rect 14967 5117 14979 5151
rect 14921 5111 14979 5117
rect 15933 5151 15991 5157
rect 15933 5117 15945 5151
rect 15979 5117 15991 5151
rect 15933 5111 15991 5117
rect 16393 5151 16451 5157
rect 16393 5117 16405 5151
rect 16439 5148 16451 5151
rect 16574 5148 16580 5160
rect 16439 5120 16580 5148
rect 16439 5117 16451 5120
rect 16393 5111 16451 5117
rect 10888 5052 12296 5080
rect 13909 5083 13967 5089
rect 13909 5049 13921 5083
rect 13955 5080 13967 5083
rect 14182 5080 14188 5092
rect 13955 5052 14188 5080
rect 13955 5049 13967 5052
rect 13909 5043 13967 5049
rect 14182 5040 14188 5052
rect 14240 5040 14246 5092
rect 15948 5080 15976 5111
rect 16574 5108 16580 5120
rect 16632 5108 16638 5160
rect 16669 5151 16727 5157
rect 16669 5117 16681 5151
rect 16715 5148 16727 5151
rect 17034 5148 17040 5160
rect 16715 5120 17040 5148
rect 16715 5117 16727 5120
rect 16669 5111 16727 5117
rect 17034 5108 17040 5120
rect 17092 5148 17098 5160
rect 17497 5151 17555 5157
rect 17497 5148 17509 5151
rect 17092 5120 17509 5148
rect 17092 5108 17098 5120
rect 17497 5117 17509 5120
rect 17543 5117 17555 5151
rect 17604 5148 17632 5188
rect 19153 5185 19165 5219
rect 19199 5185 19211 5219
rect 19153 5179 19211 5185
rect 17770 5157 17776 5160
rect 17753 5151 17776 5157
rect 17753 5148 17765 5151
rect 17604 5120 17765 5148
rect 17497 5111 17555 5117
rect 17753 5117 17765 5120
rect 17828 5148 17834 5160
rect 17828 5120 17901 5148
rect 17753 5111 17776 5117
rect 17512 5080 17540 5111
rect 17770 5108 17776 5111
rect 17828 5108 17834 5120
rect 18138 5108 18144 5160
rect 18196 5148 18202 5160
rect 18506 5148 18512 5160
rect 18196 5120 18512 5148
rect 18196 5108 18202 5120
rect 18506 5108 18512 5120
rect 18564 5108 18570 5160
rect 19168 5080 19196 5179
rect 20162 5176 20168 5228
rect 20220 5216 20226 5228
rect 20809 5219 20867 5225
rect 20809 5216 20821 5219
rect 20220 5188 20821 5216
rect 20220 5176 20226 5188
rect 20809 5185 20821 5188
rect 20855 5185 20867 5219
rect 20809 5179 20867 5185
rect 19420 5151 19478 5157
rect 19420 5148 19432 5151
rect 15948 5052 17080 5080
rect 17512 5052 19196 5080
rect 19260 5120 19432 5148
rect 10965 5015 11023 5021
rect 10965 5012 10977 5015
rect 10704 4984 10977 5012
rect 10597 4975 10655 4981
rect 10965 4981 10977 4984
rect 11011 4981 11023 5015
rect 10965 4975 11023 4981
rect 13541 5015 13599 5021
rect 13541 4981 13553 5015
rect 13587 5012 13599 5015
rect 13814 5012 13820 5024
rect 13587 4984 13820 5012
rect 13587 4981 13599 4984
rect 13541 4975 13599 4981
rect 13814 4972 13820 4984
rect 13872 4972 13878 5024
rect 13998 4972 14004 5024
rect 14056 5012 14062 5024
rect 15013 5015 15071 5021
rect 15013 5012 15025 5015
rect 14056 4984 15025 5012
rect 14056 4972 14062 4984
rect 15013 4981 15025 4984
rect 15059 4981 15071 5015
rect 15378 5012 15384 5024
rect 15339 4984 15384 5012
rect 15013 4975 15071 4981
rect 15378 4972 15384 4984
rect 15436 4972 15442 5024
rect 16574 5012 16580 5024
rect 16535 4984 16580 5012
rect 16574 4972 16580 4984
rect 16632 4972 16638 5024
rect 17052 5021 17080 5052
rect 17037 5015 17095 5021
rect 17037 4981 17049 5015
rect 17083 5012 17095 5015
rect 17862 5012 17868 5024
rect 17083 4984 17868 5012
rect 17083 4981 17095 4984
rect 17037 4975 17095 4981
rect 17862 4972 17868 4984
rect 17920 4972 17926 5024
rect 18138 4972 18144 5024
rect 18196 5012 18202 5024
rect 18877 5015 18935 5021
rect 18877 5012 18889 5015
rect 18196 4984 18889 5012
rect 18196 4972 18202 4984
rect 18877 4981 18889 4984
rect 18923 5012 18935 5015
rect 19260 5012 19288 5120
rect 19420 5117 19432 5120
rect 19466 5148 19478 5151
rect 20346 5148 20352 5160
rect 19466 5120 20352 5148
rect 19466 5117 19478 5120
rect 19420 5111 19478 5117
rect 20346 5108 20352 5120
rect 20404 5108 20410 5160
rect 20530 5012 20536 5024
rect 18923 4984 19288 5012
rect 20491 4984 20536 5012
rect 18923 4981 18935 4984
rect 18877 4975 18935 4981
rect 20530 4972 20536 4984
rect 20588 4972 20594 5024
rect 21358 5012 21364 5024
rect 21319 4984 21364 5012
rect 21358 4972 21364 4984
rect 21416 4972 21422 5024
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 2498 4808 2504 4820
rect 2459 4780 2504 4808
rect 2498 4768 2504 4780
rect 2556 4768 2562 4820
rect 2958 4808 2964 4820
rect 2919 4780 2964 4808
rect 2958 4768 2964 4780
rect 3016 4768 3022 4820
rect 3421 4811 3479 4817
rect 3421 4777 3433 4811
rect 3467 4808 3479 4811
rect 5169 4811 5227 4817
rect 5169 4808 5181 4811
rect 3467 4780 5181 4808
rect 3467 4777 3479 4780
rect 3421 4771 3479 4777
rect 5169 4777 5181 4780
rect 5215 4777 5227 4811
rect 5169 4771 5227 4777
rect 5350 4768 5356 4820
rect 5408 4808 5414 4820
rect 5994 4808 6000 4820
rect 5408 4780 6000 4808
rect 5408 4768 5414 4780
rect 5994 4768 6000 4780
rect 6052 4768 6058 4820
rect 6273 4811 6331 4817
rect 6273 4777 6285 4811
rect 6319 4808 6331 4811
rect 6454 4808 6460 4820
rect 6319 4780 6460 4808
rect 6319 4777 6331 4780
rect 6273 4771 6331 4777
rect 6454 4768 6460 4780
rect 6512 4768 6518 4820
rect 6546 4768 6552 4820
rect 6604 4808 6610 4820
rect 8205 4811 8263 4817
rect 8205 4808 8217 4811
rect 6604 4780 8217 4808
rect 6604 4768 6610 4780
rect 8205 4777 8217 4780
rect 8251 4808 8263 4811
rect 8251 4780 8432 4808
rect 8251 4777 8263 4780
rect 8205 4771 8263 4777
rect 1673 4743 1731 4749
rect 1673 4709 1685 4743
rect 1719 4740 1731 4743
rect 1762 4740 1768 4752
rect 1719 4712 1768 4740
rect 1719 4709 1731 4712
rect 1673 4703 1731 4709
rect 1762 4700 1768 4712
rect 1820 4700 1826 4752
rect 2406 4700 2412 4752
rect 2464 4740 2470 4752
rect 6178 4740 6184 4752
rect 2464 4712 6184 4740
rect 2464 4700 2470 4712
rect 6178 4700 6184 4712
rect 6236 4700 6242 4752
rect 7190 4700 7196 4752
rect 7248 4740 7254 4752
rect 8294 4740 8300 4752
rect 7248 4712 7293 4740
rect 8255 4712 8300 4740
rect 7248 4700 7254 4712
rect 8294 4700 8300 4712
rect 8352 4700 8358 4752
rect 8404 4740 8432 4780
rect 9398 4768 9404 4820
rect 9456 4808 9462 4820
rect 9769 4811 9827 4817
rect 9769 4808 9781 4811
rect 9456 4780 9781 4808
rect 9456 4768 9462 4780
rect 9769 4777 9781 4780
rect 9815 4777 9827 4811
rect 9769 4771 9827 4777
rect 9950 4768 9956 4820
rect 10008 4808 10014 4820
rect 10965 4811 11023 4817
rect 10965 4808 10977 4811
rect 10008 4780 10977 4808
rect 10008 4768 10014 4780
rect 10965 4777 10977 4780
rect 11011 4777 11023 4811
rect 10965 4771 11023 4777
rect 11333 4811 11391 4817
rect 11333 4777 11345 4811
rect 11379 4808 11391 4811
rect 12066 4808 12072 4820
rect 11379 4780 12072 4808
rect 11379 4777 11391 4780
rect 11333 4771 11391 4777
rect 12066 4768 12072 4780
rect 12124 4768 12130 4820
rect 13538 4808 13544 4820
rect 13499 4780 13544 4808
rect 13538 4768 13544 4780
rect 13596 4768 13602 4820
rect 15105 4811 15163 4817
rect 15105 4777 15117 4811
rect 15151 4777 15163 4811
rect 15105 4771 15163 4777
rect 9582 4740 9588 4752
rect 8404 4712 9588 4740
rect 9582 4700 9588 4712
rect 9640 4700 9646 4752
rect 9674 4700 9680 4752
rect 9732 4740 9738 4752
rect 11977 4743 12035 4749
rect 11977 4740 11989 4743
rect 9732 4712 11989 4740
rect 9732 4700 9738 4712
rect 11977 4709 11989 4712
rect 12023 4709 12035 4743
rect 13998 4740 14004 4752
rect 11977 4703 12035 4709
rect 12406 4712 14004 4740
rect 2593 4675 2651 4681
rect 2593 4641 2605 4675
rect 2639 4672 2651 4675
rect 2958 4672 2964 4684
rect 2639 4644 2964 4672
rect 2639 4641 2651 4644
rect 2593 4635 2651 4641
rect 2958 4632 2964 4644
rect 3016 4632 3022 4684
rect 3234 4632 3240 4684
rect 3292 4672 3298 4684
rect 3292 4644 3385 4672
rect 3292 4632 3298 4644
rect 3418 4632 3424 4684
rect 3476 4672 3482 4684
rect 4062 4672 4068 4684
rect 3476 4644 4068 4672
rect 3476 4632 3482 4644
rect 4062 4632 4068 4644
rect 4120 4632 4126 4684
rect 4172 4644 5396 4672
rect 1486 4564 1492 4616
rect 1544 4604 1550 4616
rect 2314 4604 2320 4616
rect 1544 4576 2320 4604
rect 1544 4564 1550 4576
rect 2314 4564 2320 4576
rect 2372 4564 2378 4616
rect 3252 4604 3280 4632
rect 4172 4604 4200 4644
rect 3252 4576 4200 4604
rect 4985 4607 5043 4613
rect 4985 4573 4997 4607
rect 5031 4573 5043 4607
rect 4985 4567 5043 4573
rect 5077 4607 5135 4613
rect 5077 4573 5089 4607
rect 5123 4604 5135 4607
rect 5258 4604 5264 4616
rect 5123 4576 5264 4604
rect 5123 4573 5135 4576
rect 5077 4567 5135 4573
rect 3510 4496 3516 4548
rect 3568 4536 3574 4548
rect 3970 4536 3976 4548
rect 3568 4508 3976 4536
rect 3568 4496 3574 4508
rect 3970 4496 3976 4508
rect 4028 4496 4034 4548
rect 5000 4536 5028 4567
rect 5258 4564 5264 4576
rect 5316 4564 5322 4616
rect 5368 4604 5396 4644
rect 6288 4644 9444 4672
rect 6288 4604 6316 4644
rect 5368 4576 6316 4604
rect 6365 4607 6423 4613
rect 6365 4573 6377 4607
rect 6411 4573 6423 4607
rect 6365 4567 6423 4573
rect 6270 4536 6276 4548
rect 5000 4508 6276 4536
rect 6270 4496 6276 4508
rect 6328 4536 6334 4548
rect 6380 4536 6408 4567
rect 6638 4564 6644 4616
rect 6696 4604 6702 4616
rect 7285 4607 7343 4613
rect 7285 4604 7297 4607
rect 6696 4576 7297 4604
rect 6696 4564 6702 4576
rect 7285 4573 7297 4576
rect 7331 4573 7343 4607
rect 7285 4567 7343 4573
rect 7377 4607 7435 4613
rect 7377 4573 7389 4607
rect 7423 4573 7435 4607
rect 7377 4567 7435 4573
rect 8113 4607 8171 4613
rect 8113 4573 8125 4607
rect 8159 4604 8171 4607
rect 8570 4604 8576 4616
rect 8159 4576 8576 4604
rect 8159 4573 8171 4576
rect 8113 4567 8171 4573
rect 7392 4536 7420 4567
rect 8570 4564 8576 4576
rect 8628 4564 8634 4616
rect 9306 4604 9312 4616
rect 9267 4576 9312 4604
rect 9306 4564 9312 4576
rect 9364 4564 9370 4616
rect 9416 4604 9444 4644
rect 9766 4632 9772 4684
rect 9824 4672 9830 4684
rect 9953 4675 10011 4681
rect 9953 4672 9965 4675
rect 9824 4644 9965 4672
rect 9824 4632 9830 4644
rect 9953 4641 9965 4644
rect 9999 4641 10011 4675
rect 12406 4672 12434 4712
rect 13998 4700 14004 4712
rect 14056 4700 14062 4752
rect 15120 4740 15148 4771
rect 15378 4768 15384 4820
rect 15436 4808 15442 4820
rect 18233 4811 18291 4817
rect 15436 4780 17816 4808
rect 15436 4768 15442 4780
rect 17788 4740 17816 4780
rect 18233 4777 18245 4811
rect 18279 4808 18291 4811
rect 18598 4808 18604 4820
rect 18279 4780 18604 4808
rect 18279 4777 18291 4780
rect 18233 4771 18291 4777
rect 18598 4768 18604 4780
rect 18656 4768 18662 4820
rect 19794 4768 19800 4820
rect 19852 4808 19858 4820
rect 20165 4811 20223 4817
rect 20165 4808 20177 4811
rect 19852 4780 20177 4808
rect 19852 4768 19858 4780
rect 20165 4777 20177 4780
rect 20211 4777 20223 4811
rect 20165 4771 20223 4777
rect 18325 4743 18383 4749
rect 18325 4740 18337 4743
rect 15120 4712 17724 4740
rect 17788 4712 18337 4740
rect 9953 4635 10011 4641
rect 10796 4644 12434 4672
rect 10229 4607 10287 4613
rect 10229 4604 10241 4607
rect 9416 4576 10241 4604
rect 10229 4573 10241 4576
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 6328 4508 7420 4536
rect 6328 4496 6334 4508
rect 7834 4496 7840 4548
rect 7892 4536 7898 4548
rect 8478 4536 8484 4548
rect 7892 4508 8484 4536
rect 7892 4496 7898 4508
rect 8478 4496 8484 4508
rect 8536 4496 8542 4548
rect 9490 4496 9496 4548
rect 9548 4536 9554 4548
rect 10796 4536 10824 4644
rect 12802 4632 12808 4684
rect 12860 4672 12866 4684
rect 12897 4675 12955 4681
rect 12897 4672 12909 4675
rect 12860 4644 12909 4672
rect 12860 4632 12866 4644
rect 12897 4641 12909 4644
rect 12943 4672 12955 4675
rect 13170 4672 13176 4684
rect 12943 4644 13176 4672
rect 12943 4641 12955 4644
rect 12897 4635 12955 4641
rect 13170 4632 13176 4644
rect 13228 4632 13234 4684
rect 13357 4675 13415 4681
rect 13357 4641 13369 4675
rect 13403 4672 13415 4675
rect 13630 4672 13636 4684
rect 13403 4644 13636 4672
rect 13403 4641 13415 4644
rect 13357 4635 13415 4641
rect 13630 4632 13636 4644
rect 13688 4632 13694 4684
rect 13814 4672 13820 4684
rect 13775 4644 13820 4672
rect 13814 4632 13820 4644
rect 13872 4632 13878 4684
rect 14645 4675 14703 4681
rect 14645 4641 14657 4675
rect 14691 4672 14703 4675
rect 14918 4672 14924 4684
rect 14691 4644 14924 4672
rect 14691 4641 14703 4644
rect 14645 4635 14703 4641
rect 14918 4632 14924 4644
rect 14976 4632 14982 4684
rect 15378 4672 15384 4684
rect 15339 4644 15384 4672
rect 15378 4632 15384 4644
rect 15436 4632 15442 4684
rect 15838 4672 15844 4684
rect 15799 4644 15844 4672
rect 15838 4632 15844 4644
rect 15896 4632 15902 4684
rect 16114 4681 16120 4684
rect 16108 4635 16120 4681
rect 16172 4672 16178 4684
rect 17696 4681 17724 4712
rect 18325 4709 18337 4712
rect 18371 4709 18383 4743
rect 18325 4703 18383 4709
rect 21269 4743 21327 4749
rect 21269 4709 21281 4743
rect 21315 4740 21327 4743
rect 21358 4740 21364 4752
rect 21315 4712 21364 4740
rect 21315 4709 21327 4712
rect 21269 4703 21327 4709
rect 21358 4700 21364 4712
rect 21416 4700 21422 4752
rect 17681 4675 17739 4681
rect 16172 4644 16208 4672
rect 16114 4632 16120 4635
rect 16172 4632 16178 4644
rect 17681 4641 17693 4675
rect 17727 4641 17739 4675
rect 17681 4635 17739 4641
rect 19061 4675 19119 4681
rect 19061 4641 19073 4675
rect 19107 4672 19119 4675
rect 19242 4672 19248 4684
rect 19107 4644 19248 4672
rect 19107 4641 19119 4644
rect 19061 4635 19119 4641
rect 19242 4632 19248 4644
rect 19300 4632 19306 4684
rect 11146 4564 11152 4616
rect 11204 4604 11210 4616
rect 11425 4607 11483 4613
rect 11425 4604 11437 4607
rect 11204 4576 11437 4604
rect 11204 4564 11210 4576
rect 11425 4573 11437 4576
rect 11471 4573 11483 4607
rect 11425 4567 11483 4573
rect 11609 4607 11667 4613
rect 11609 4573 11621 4607
rect 11655 4604 11667 4607
rect 11698 4604 11704 4616
rect 11655 4576 11704 4604
rect 11655 4573 11667 4576
rect 11609 4567 11667 4573
rect 11698 4564 11704 4576
rect 11756 4564 11762 4616
rect 15286 4604 15292 4616
rect 13096 4576 15292 4604
rect 9548 4508 10824 4536
rect 9548 4496 9554 4508
rect 10870 4496 10876 4548
rect 10928 4536 10934 4548
rect 13096 4545 13124 4576
rect 15286 4564 15292 4576
rect 15344 4564 15350 4616
rect 18138 4604 18144 4616
rect 18099 4576 18144 4604
rect 18138 4564 18144 4576
rect 18196 4564 18202 4616
rect 20257 4607 20315 4613
rect 20257 4604 20269 4607
rect 18708 4576 20269 4604
rect 12345 4539 12403 4545
rect 12345 4536 12357 4539
rect 10928 4508 12357 4536
rect 10928 4496 10934 4508
rect 12345 4505 12357 4508
rect 12391 4505 12403 4539
rect 12345 4499 12403 4505
rect 13081 4539 13139 4545
rect 13081 4505 13093 4539
rect 13127 4505 13139 4539
rect 13081 4499 13139 4505
rect 14001 4539 14059 4545
rect 14001 4505 14013 4539
rect 14047 4536 14059 4539
rect 15194 4536 15200 4548
rect 14047 4508 15200 4536
rect 14047 4505 14059 4508
rect 14001 4499 14059 4505
rect 15194 4496 15200 4508
rect 15252 4496 15258 4548
rect 17218 4536 17224 4548
rect 17179 4508 17224 4536
rect 17218 4496 17224 4508
rect 17276 4496 17282 4548
rect 18708 4545 18736 4576
rect 20257 4573 20269 4576
rect 20303 4573 20315 4607
rect 20257 4567 20315 4573
rect 20441 4607 20499 4613
rect 20441 4573 20453 4607
rect 20487 4604 20499 4607
rect 20530 4604 20536 4616
rect 20487 4576 20536 4604
rect 20487 4573 20499 4576
rect 20441 4567 20499 4573
rect 20530 4564 20536 4576
rect 20588 4564 20594 4616
rect 18693 4539 18751 4545
rect 18693 4505 18705 4539
rect 18739 4505 18751 4539
rect 21082 4536 21088 4548
rect 21043 4508 21088 4536
rect 18693 4499 18751 4505
rect 21082 4496 21088 4508
rect 21140 4496 21146 4548
rect 1765 4471 1823 4477
rect 1765 4437 1777 4471
rect 1811 4468 1823 4471
rect 4062 4468 4068 4480
rect 1811 4440 4068 4468
rect 1811 4437 1823 4440
rect 1765 4431 1823 4437
rect 4062 4428 4068 4440
rect 4120 4428 4126 4480
rect 4249 4471 4307 4477
rect 4249 4437 4261 4471
rect 4295 4468 4307 4471
rect 5350 4468 5356 4480
rect 4295 4440 5356 4468
rect 4295 4437 4307 4440
rect 4249 4431 4307 4437
rect 5350 4428 5356 4440
rect 5408 4428 5414 4480
rect 5534 4468 5540 4480
rect 5495 4440 5540 4468
rect 5534 4428 5540 4440
rect 5592 4428 5598 4480
rect 5810 4468 5816 4480
rect 5771 4440 5816 4468
rect 5810 4428 5816 4440
rect 5868 4428 5874 4480
rect 5994 4428 6000 4480
rect 6052 4468 6058 4480
rect 6825 4471 6883 4477
rect 6825 4468 6837 4471
rect 6052 4440 6837 4468
rect 6052 4428 6058 4440
rect 6825 4437 6837 4440
rect 6871 4437 6883 4471
rect 6825 4431 6883 4437
rect 7190 4428 7196 4480
rect 7248 4468 7254 4480
rect 7466 4468 7472 4480
rect 7248 4440 7472 4468
rect 7248 4428 7254 4440
rect 7466 4428 7472 4440
rect 7524 4428 7530 4480
rect 8294 4428 8300 4480
rect 8352 4468 8358 4480
rect 8665 4471 8723 4477
rect 8665 4468 8677 4471
rect 8352 4440 8677 4468
rect 8352 4428 8358 4440
rect 8665 4437 8677 4440
rect 8711 4437 8723 4471
rect 8665 4431 8723 4437
rect 9858 4428 9864 4480
rect 9916 4468 9922 4480
rect 10597 4471 10655 4477
rect 10597 4468 10609 4471
rect 9916 4440 10609 4468
rect 9916 4428 9922 4440
rect 10597 4437 10609 4440
rect 10643 4437 10655 4471
rect 10597 4431 10655 4437
rect 15565 4471 15623 4477
rect 15565 4437 15577 4471
rect 15611 4468 15623 4471
rect 17126 4468 17132 4480
rect 15611 4440 17132 4468
rect 15611 4437 15623 4440
rect 15565 4431 15623 4437
rect 17126 4428 17132 4440
rect 17184 4428 17190 4480
rect 17494 4468 17500 4480
rect 17455 4440 17500 4468
rect 17494 4428 17500 4440
rect 17552 4428 17558 4480
rect 19150 4428 19156 4480
rect 19208 4468 19214 4480
rect 19245 4471 19303 4477
rect 19245 4468 19257 4471
rect 19208 4440 19257 4468
rect 19208 4428 19214 4440
rect 19245 4437 19257 4440
rect 19291 4437 19303 4471
rect 19245 4431 19303 4437
rect 19797 4471 19855 4477
rect 19797 4437 19809 4471
rect 19843 4468 19855 4471
rect 20438 4468 20444 4480
rect 19843 4440 20444 4468
rect 19843 4437 19855 4440
rect 19797 4431 19855 4437
rect 20438 4428 20444 4440
rect 20496 4428 20502 4480
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 1486 4264 1492 4276
rect 1447 4236 1492 4264
rect 1486 4224 1492 4236
rect 1544 4224 1550 4276
rect 2958 4224 2964 4276
rect 3016 4264 3022 4276
rect 3145 4267 3203 4273
rect 3145 4264 3157 4267
rect 3016 4236 3157 4264
rect 3016 4224 3022 4236
rect 3145 4233 3157 4236
rect 3191 4233 3203 4267
rect 3145 4227 3203 4233
rect 4062 4224 4068 4276
rect 4120 4264 4126 4276
rect 8570 4264 8576 4276
rect 4120 4236 7328 4264
rect 4120 4224 4126 4236
rect 4246 4156 4252 4208
rect 4304 4196 4310 4208
rect 4341 4199 4399 4205
rect 4341 4196 4353 4199
rect 4304 4168 4353 4196
rect 4304 4156 4310 4168
rect 4341 4165 4353 4168
rect 4387 4165 4399 4199
rect 6730 4196 6736 4208
rect 4341 4159 4399 4165
rect 5276 4168 6736 4196
rect 3050 4128 3056 4140
rect 2792 4100 3056 4128
rect 2792 4060 2820 4100
rect 3050 4088 3056 4100
rect 3108 4128 3114 4140
rect 3697 4131 3755 4137
rect 3697 4128 3709 4131
rect 3108 4100 3709 4128
rect 3108 4088 3114 4100
rect 3697 4097 3709 4100
rect 3743 4097 3755 4131
rect 3697 4091 3755 4097
rect 2608 4032 2820 4060
rect 1670 3952 1676 4004
rect 1728 3992 1734 4004
rect 2608 4001 2636 4032
rect 2866 4020 2872 4072
rect 2924 4060 2930 4072
rect 3142 4060 3148 4072
rect 2924 4032 3148 4060
rect 2924 4020 2930 4032
rect 3142 4020 3148 4032
rect 3200 4020 3206 4072
rect 3786 4020 3792 4072
rect 3844 4060 3850 4072
rect 4157 4063 4215 4069
rect 4157 4060 4169 4063
rect 3844 4032 4169 4060
rect 3844 4020 3850 4032
rect 4157 4029 4169 4032
rect 4203 4060 4215 4063
rect 5276 4060 5304 4168
rect 6730 4156 6736 4168
rect 6788 4156 6794 4208
rect 5442 4128 5448 4140
rect 5403 4100 5448 4128
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 6914 4128 6920 4140
rect 6104 4100 6920 4128
rect 4203 4032 5304 4060
rect 5353 4063 5411 4069
rect 4203 4029 4215 4032
rect 4157 4023 4215 4029
rect 5353 4029 5365 4063
rect 5399 4060 5411 4063
rect 5534 4060 5540 4072
rect 5399 4032 5540 4060
rect 5399 4029 5411 4032
rect 5353 4023 5411 4029
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 6104 4069 6132 4100
rect 6914 4088 6920 4100
rect 6972 4088 6978 4140
rect 5721 4063 5779 4069
rect 5721 4029 5733 4063
rect 5767 4060 5779 4063
rect 6089 4063 6147 4069
rect 6089 4060 6101 4063
rect 5767 4032 6101 4060
rect 5767 4029 5779 4032
rect 5721 4023 5779 4029
rect 6089 4029 6101 4032
rect 6135 4029 6147 4063
rect 6089 4023 6147 4029
rect 6641 4063 6699 4069
rect 6641 4029 6653 4063
rect 6687 4060 6699 4063
rect 7006 4060 7012 4072
rect 6687 4032 7012 4060
rect 6687 4029 6699 4032
rect 6641 4023 6699 4029
rect 7006 4020 7012 4032
rect 7064 4020 7070 4072
rect 2602 3995 2660 4001
rect 2602 3992 2614 3995
rect 1728 3964 2614 3992
rect 1728 3952 1734 3964
rect 2602 3961 2614 3964
rect 2648 3961 2660 3995
rect 4706 3992 4712 4004
rect 2602 3955 2660 3961
rect 2746 3964 4712 3992
rect 1854 3884 1860 3936
rect 1912 3924 1918 3936
rect 2746 3924 2774 3964
rect 4706 3952 4712 3964
rect 4764 3952 4770 4004
rect 4798 3952 4804 4004
rect 4856 3992 4862 4004
rect 5261 3995 5319 4001
rect 4856 3964 5028 3992
rect 4856 3952 4862 3964
rect 3510 3924 3516 3936
rect 1912 3896 2774 3924
rect 3471 3896 3516 3924
rect 1912 3884 1918 3896
rect 3510 3884 3516 3896
rect 3568 3884 3574 3936
rect 3602 3884 3608 3936
rect 3660 3924 3666 3936
rect 4890 3924 4896 3936
rect 3660 3896 3705 3924
rect 4851 3896 4896 3924
rect 3660 3884 3666 3896
rect 4890 3884 4896 3896
rect 4948 3884 4954 3936
rect 5000 3924 5028 3964
rect 5261 3961 5273 3995
rect 5307 3992 5319 3995
rect 5994 3992 6000 4004
rect 5307 3964 6000 3992
rect 5307 3961 5319 3964
rect 5261 3955 5319 3961
rect 5994 3952 6000 3964
rect 6052 3952 6058 4004
rect 6454 3952 6460 4004
rect 6512 3992 6518 4004
rect 7098 3992 7104 4004
rect 6512 3964 7104 3992
rect 6512 3952 6518 3964
rect 7098 3952 7104 3964
rect 7156 3952 7162 4004
rect 7300 3992 7328 4236
rect 7484 4236 8576 4264
rect 7484 4196 7512 4236
rect 8570 4224 8576 4236
rect 8628 4224 8634 4276
rect 10042 4264 10048 4276
rect 10003 4236 10048 4264
rect 10042 4224 10048 4236
rect 10100 4224 10106 4276
rect 10410 4224 10416 4276
rect 10468 4224 10474 4276
rect 11974 4224 11980 4276
rect 12032 4264 12038 4276
rect 12069 4267 12127 4273
rect 12069 4264 12081 4267
rect 12032 4236 12081 4264
rect 12032 4224 12038 4236
rect 12069 4233 12081 4236
rect 12115 4233 12127 4267
rect 12342 4264 12348 4276
rect 12303 4236 12348 4264
rect 12069 4227 12127 4233
rect 12342 4224 12348 4236
rect 12400 4224 12406 4276
rect 14918 4224 14924 4276
rect 14976 4264 14982 4276
rect 19242 4264 19248 4276
rect 14976 4236 19248 4264
rect 14976 4224 14982 4236
rect 19242 4224 19248 4236
rect 19300 4224 19306 4276
rect 7392 4168 7512 4196
rect 7392 4137 7420 4168
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 7466 4088 7472 4140
rect 7524 4128 7530 4140
rect 8202 4128 8208 4140
rect 7524 4100 8208 4128
rect 7524 4088 7530 4100
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 10318 4088 10324 4140
rect 10376 4088 10382 4140
rect 8297 4063 8355 4069
rect 8297 4029 8309 4063
rect 8343 4060 8355 4063
rect 8386 4060 8392 4072
rect 8343 4032 8392 4060
rect 8343 4029 8355 4032
rect 8297 4023 8355 4029
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 9306 4060 9312 4072
rect 8496 4032 9312 4060
rect 7561 3995 7619 4001
rect 7561 3992 7573 3995
rect 7300 3964 7573 3992
rect 7561 3961 7573 3964
rect 7607 3961 7619 3995
rect 7561 3955 7619 3961
rect 7653 3995 7711 4001
rect 7653 3961 7665 3995
rect 7699 3992 7711 3995
rect 8496 3992 8524 4032
rect 9306 4020 9312 4032
rect 9364 4020 9370 4072
rect 10042 4020 10048 4072
rect 10100 4060 10106 4072
rect 10229 4063 10287 4069
rect 10229 4060 10241 4063
rect 10100 4032 10241 4060
rect 10100 4020 10106 4032
rect 10229 4029 10241 4032
rect 10275 4060 10287 4063
rect 10336 4060 10364 4088
rect 10275 4032 10364 4060
rect 10275 4029 10287 4032
rect 10229 4023 10287 4029
rect 8570 4001 8576 4004
rect 7699 3964 8524 3992
rect 7699 3961 7711 3964
rect 7653 3955 7711 3961
rect 8564 3955 8576 4001
rect 8628 3992 8634 4004
rect 8628 3964 8664 3992
rect 5721 3927 5779 3933
rect 5721 3924 5733 3927
rect 5000 3896 5733 3924
rect 5721 3893 5733 3896
rect 5767 3893 5779 3927
rect 5902 3924 5908 3936
rect 5863 3896 5908 3924
rect 5721 3887 5779 3893
rect 5902 3884 5908 3896
rect 5960 3884 5966 3936
rect 6825 3927 6883 3933
rect 6825 3893 6837 3927
rect 6871 3924 6883 3927
rect 7466 3924 7472 3936
rect 6871 3896 7472 3924
rect 6871 3893 6883 3896
rect 6825 3887 6883 3893
rect 7466 3884 7472 3896
rect 7524 3884 7530 3936
rect 7576 3924 7604 3955
rect 8570 3952 8576 3955
rect 8628 3952 8634 3964
rect 8754 3952 8760 4004
rect 8812 3992 8818 4004
rect 10428 3992 10456 4224
rect 18138 4196 18144 4208
rect 18099 4168 18144 4196
rect 18138 4156 18144 4168
rect 18196 4156 18202 4208
rect 10870 4088 10876 4140
rect 10928 4088 10934 4140
rect 12342 4088 12348 4140
rect 12400 4128 12406 4140
rect 15286 4128 15292 4140
rect 12400 4100 12756 4128
rect 15247 4100 15292 4128
rect 12400 4088 12406 4100
rect 10502 4020 10508 4072
rect 10560 4060 10566 4072
rect 10689 4063 10747 4069
rect 10689 4060 10701 4063
rect 10560 4032 10701 4060
rect 10560 4020 10566 4032
rect 10689 4029 10701 4032
rect 10735 4060 10747 4063
rect 10778 4060 10784 4072
rect 10735 4032 10784 4060
rect 10735 4029 10747 4032
rect 10689 4023 10747 4029
rect 10778 4020 10784 4032
rect 10836 4020 10842 4072
rect 10594 3992 10600 4004
rect 8812 3964 10600 3992
rect 8812 3952 8818 3964
rect 10594 3952 10600 3964
rect 10652 3952 10658 4004
rect 10888 3992 10916 4088
rect 12728 4072 12756 4100
rect 15286 4088 15292 4100
rect 15344 4088 15350 4140
rect 15381 4131 15439 4137
rect 15381 4097 15393 4131
rect 15427 4128 15439 4131
rect 15470 4128 15476 4140
rect 15427 4100 15476 4128
rect 15427 4097 15439 4100
rect 15381 4091 15439 4097
rect 15470 4088 15476 4100
rect 15528 4088 15534 4140
rect 18414 4088 18420 4140
rect 18472 4128 18478 4140
rect 19518 4128 19524 4140
rect 18472 4100 19524 4128
rect 18472 4088 18478 4100
rect 19518 4088 19524 4100
rect 19576 4088 19582 4140
rect 21085 4131 21143 4137
rect 21085 4097 21097 4131
rect 21131 4128 21143 4131
rect 21174 4128 21180 4140
rect 21131 4100 21180 4128
rect 21131 4097 21143 4100
rect 21085 4091 21143 4097
rect 21174 4088 21180 4100
rect 21232 4088 21238 4140
rect 11149 4063 11207 4069
rect 11149 4029 11161 4063
rect 11195 4060 11207 4063
rect 11238 4060 11244 4072
rect 11195 4032 11244 4060
rect 11195 4029 11207 4032
rect 11149 4023 11207 4029
rect 11238 4020 11244 4032
rect 11296 4020 11302 4072
rect 11790 4020 11796 4072
rect 11848 4060 11854 4072
rect 11885 4063 11943 4069
rect 11885 4060 11897 4063
rect 11848 4032 11897 4060
rect 11848 4020 11854 4032
rect 11885 4029 11897 4032
rect 11931 4029 11943 4063
rect 11885 4023 11943 4029
rect 11974 4020 11980 4072
rect 12032 4060 12038 4072
rect 12250 4060 12256 4072
rect 12032 4032 12256 4060
rect 12032 4020 12038 4032
rect 12250 4020 12256 4032
rect 12308 4060 12314 4072
rect 12529 4063 12587 4069
rect 12529 4060 12541 4063
rect 12308 4032 12541 4060
rect 12308 4020 12314 4032
rect 12529 4029 12541 4032
rect 12575 4029 12587 4063
rect 12529 4023 12587 4029
rect 12710 4020 12716 4072
rect 12768 4060 12774 4072
rect 12805 4063 12863 4069
rect 12805 4060 12817 4063
rect 12768 4032 12817 4060
rect 12768 4020 12774 4032
rect 12805 4029 12817 4032
rect 12851 4029 12863 4063
rect 13446 4060 13452 4072
rect 13407 4032 13452 4060
rect 12805 4023 12863 4029
rect 13446 4020 13452 4032
rect 13504 4020 13510 4072
rect 13716 4063 13774 4069
rect 13716 4029 13728 4063
rect 13762 4060 13774 4063
rect 14090 4060 14096 4072
rect 13762 4032 14096 4060
rect 13762 4029 13774 4032
rect 13716 4023 13774 4029
rect 14090 4020 14096 4032
rect 14148 4020 14154 4072
rect 14200 4032 15608 4060
rect 10796 3964 10916 3992
rect 10796 3936 10824 3964
rect 7742 3924 7748 3936
rect 7576 3896 7748 3924
rect 7742 3884 7748 3896
rect 7800 3884 7806 3936
rect 8021 3927 8079 3933
rect 8021 3893 8033 3927
rect 8067 3924 8079 3927
rect 8386 3924 8392 3936
rect 8067 3896 8392 3924
rect 8067 3893 8079 3896
rect 8021 3887 8079 3893
rect 8386 3884 8392 3896
rect 8444 3884 8450 3936
rect 8478 3884 8484 3936
rect 8536 3924 8542 3936
rect 9030 3924 9036 3936
rect 8536 3896 9036 3924
rect 8536 3884 8542 3896
rect 9030 3884 9036 3896
rect 9088 3924 9094 3936
rect 9306 3924 9312 3936
rect 9088 3896 9312 3924
rect 9088 3884 9094 3896
rect 9306 3884 9312 3896
rect 9364 3884 9370 3936
rect 9677 3927 9735 3933
rect 9677 3893 9689 3927
rect 9723 3924 9735 3927
rect 9858 3924 9864 3936
rect 9723 3896 9864 3924
rect 9723 3893 9735 3896
rect 9677 3887 9735 3893
rect 9858 3884 9864 3896
rect 9916 3884 9922 3936
rect 10134 3884 10140 3936
rect 10192 3924 10198 3936
rect 10505 3927 10563 3933
rect 10505 3924 10517 3927
rect 10192 3896 10517 3924
rect 10192 3884 10198 3896
rect 10505 3893 10517 3896
rect 10551 3893 10563 3927
rect 10505 3887 10563 3893
rect 10778 3884 10784 3936
rect 10836 3884 10842 3936
rect 10965 3927 11023 3933
rect 10965 3893 10977 3927
rect 11011 3924 11023 3927
rect 11146 3924 11152 3936
rect 11011 3896 11152 3924
rect 11011 3893 11023 3896
rect 10965 3887 11023 3893
rect 11146 3884 11152 3896
rect 11204 3884 11210 3936
rect 12986 3924 12992 3936
rect 12947 3896 12992 3924
rect 12986 3884 12992 3896
rect 13044 3884 13050 3936
rect 13538 3884 13544 3936
rect 13596 3924 13602 3936
rect 14200 3924 14228 4032
rect 14274 3952 14280 4004
rect 14332 3992 14338 4004
rect 15473 3995 15531 4001
rect 15473 3992 15485 3995
rect 14332 3964 15485 3992
rect 14332 3952 14338 3964
rect 15473 3961 15485 3964
rect 15519 3961 15531 3995
rect 15580 3992 15608 4032
rect 16574 4020 16580 4072
rect 16632 4060 16638 4072
rect 17865 4063 17923 4069
rect 17865 4060 17877 4063
rect 16632 4032 17877 4060
rect 16632 4020 16638 4032
rect 17865 4029 17877 4032
rect 17911 4029 17923 4063
rect 17865 4023 17923 4029
rect 18046 4020 18052 4072
rect 18104 4060 18110 4072
rect 18325 4063 18383 4069
rect 18325 4060 18337 4063
rect 18104 4032 18337 4060
rect 18104 4020 18110 4032
rect 18325 4029 18337 4032
rect 18371 4029 18383 4063
rect 18874 4060 18880 4072
rect 18835 4032 18880 4060
rect 18325 4023 18383 4029
rect 18874 4020 18880 4032
rect 18932 4020 18938 4072
rect 19334 4060 19340 4072
rect 19295 4032 19340 4060
rect 19334 4020 19340 4032
rect 19392 4020 19398 4072
rect 20530 4020 20536 4072
rect 20588 4060 20594 4072
rect 20818 4063 20876 4069
rect 20818 4060 20830 4063
rect 20588 4032 20830 4060
rect 20588 4020 20594 4032
rect 20818 4029 20830 4032
rect 20864 4029 20876 4063
rect 20818 4023 20876 4029
rect 15580 3964 16896 3992
rect 15473 3955 15531 3961
rect 13596 3896 14228 3924
rect 14829 3927 14887 3933
rect 13596 3884 13602 3896
rect 14829 3893 14841 3927
rect 14875 3924 14887 3927
rect 15286 3924 15292 3936
rect 14875 3896 15292 3924
rect 14875 3893 14887 3896
rect 14829 3887 14887 3893
rect 15286 3884 15292 3896
rect 15344 3884 15350 3936
rect 15838 3924 15844 3936
rect 15799 3896 15844 3924
rect 15838 3884 15844 3896
rect 15896 3884 15902 3936
rect 16390 3924 16396 3936
rect 16351 3896 16396 3924
rect 16390 3884 16396 3896
rect 16448 3884 16454 3936
rect 16868 3924 16896 3964
rect 16942 3952 16948 4004
rect 17000 3992 17006 4004
rect 17129 3995 17187 4001
rect 17129 3992 17141 3995
rect 17000 3964 17141 3992
rect 17000 3952 17006 3964
rect 17129 3961 17141 3964
rect 17175 3961 17187 3995
rect 17129 3955 17187 3961
rect 17313 3995 17371 4001
rect 17313 3961 17325 3995
rect 17359 3961 17371 3995
rect 17313 3955 17371 3961
rect 17034 3924 17040 3936
rect 16868 3896 17040 3924
rect 17034 3884 17040 3896
rect 17092 3884 17098 3936
rect 17328 3924 17356 3955
rect 17402 3952 17408 4004
rect 17460 3992 17466 4004
rect 17460 3964 19748 3992
rect 17460 3952 17466 3964
rect 17681 3927 17739 3933
rect 17681 3924 17693 3927
rect 17328 3896 17693 3924
rect 17681 3893 17693 3896
rect 17727 3893 17739 3927
rect 17681 3887 17739 3893
rect 17770 3884 17776 3936
rect 17828 3924 17834 3936
rect 18693 3927 18751 3933
rect 18693 3924 18705 3927
rect 17828 3896 18705 3924
rect 17828 3884 17834 3896
rect 18693 3893 18705 3896
rect 18739 3893 18751 3927
rect 18693 3887 18751 3893
rect 19153 3927 19211 3933
rect 19153 3893 19165 3927
rect 19199 3924 19211 3927
rect 19242 3924 19248 3936
rect 19199 3896 19248 3924
rect 19199 3893 19211 3896
rect 19153 3887 19211 3893
rect 19242 3884 19248 3896
rect 19300 3884 19306 3936
rect 19720 3933 19748 3964
rect 20070 3952 20076 4004
rect 20128 3992 20134 4004
rect 21818 3992 21824 4004
rect 20128 3964 21824 3992
rect 20128 3952 20134 3964
rect 21818 3952 21824 3964
rect 21876 3952 21882 4004
rect 19705 3927 19763 3933
rect 19705 3893 19717 3927
rect 19751 3893 19763 3927
rect 19705 3887 19763 3893
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 1670 3720 1676 3732
rect 1631 3692 1676 3720
rect 1670 3680 1676 3692
rect 1728 3680 1734 3732
rect 3510 3680 3516 3732
rect 3568 3720 3574 3732
rect 4249 3723 4307 3729
rect 4249 3720 4261 3723
rect 3568 3692 4261 3720
rect 3568 3680 3574 3692
rect 4249 3689 4261 3692
rect 4295 3720 4307 3723
rect 5721 3723 5779 3729
rect 4295 3692 5028 3720
rect 4295 3689 4307 3692
rect 4249 3683 4307 3689
rect 1946 3612 1952 3664
rect 2004 3652 2010 3664
rect 2004 3624 3740 3652
rect 2004 3612 2010 3624
rect 3712 3596 3740 3624
rect 3878 3612 3884 3664
rect 3936 3652 3942 3664
rect 3936 3624 4568 3652
rect 3936 3612 3942 3624
rect 2774 3544 2780 3596
rect 2832 3593 2838 3596
rect 2832 3584 2844 3593
rect 3326 3584 3332 3596
rect 2832 3556 2877 3584
rect 3287 3556 3332 3584
rect 2832 3547 2844 3556
rect 2832 3544 2838 3547
rect 3326 3544 3332 3556
rect 3384 3544 3390 3596
rect 3694 3544 3700 3596
rect 3752 3584 3758 3596
rect 4065 3587 4123 3593
rect 4065 3584 4077 3587
rect 3752 3556 4077 3584
rect 3752 3544 3758 3556
rect 4065 3553 4077 3556
rect 4111 3553 4123 3587
rect 4430 3584 4436 3596
rect 4391 3556 4436 3584
rect 4065 3547 4123 3553
rect 4430 3544 4436 3556
rect 4488 3544 4494 3596
rect 4540 3593 4568 3624
rect 4525 3587 4583 3593
rect 4525 3553 4537 3587
rect 4571 3553 4583 3587
rect 5000 3584 5028 3692
rect 5721 3689 5733 3723
rect 5767 3720 5779 3723
rect 5810 3720 5816 3732
rect 5767 3692 5816 3720
rect 5767 3689 5779 3692
rect 5721 3683 5779 3689
rect 5810 3680 5816 3692
rect 5868 3680 5874 3732
rect 6270 3680 6276 3732
rect 6328 3720 6334 3732
rect 6365 3723 6423 3729
rect 6365 3720 6377 3723
rect 6328 3692 6377 3720
rect 6328 3680 6334 3692
rect 6365 3689 6377 3692
rect 6411 3689 6423 3723
rect 8386 3720 8392 3732
rect 8347 3692 8392 3720
rect 6365 3683 6423 3689
rect 8386 3680 8392 3692
rect 8444 3680 8450 3732
rect 8570 3680 8576 3732
rect 8628 3720 8634 3732
rect 10965 3723 11023 3729
rect 10965 3720 10977 3723
rect 8628 3692 10977 3720
rect 8628 3680 8634 3692
rect 10965 3689 10977 3692
rect 11011 3689 11023 3723
rect 10965 3683 11023 3689
rect 11333 3723 11391 3729
rect 11333 3689 11345 3723
rect 11379 3720 11391 3723
rect 11606 3720 11612 3732
rect 11379 3692 11612 3720
rect 11379 3689 11391 3692
rect 11333 3683 11391 3689
rect 11606 3680 11612 3692
rect 11664 3680 11670 3732
rect 11716 3692 15424 3720
rect 5074 3612 5080 3664
rect 5132 3652 5138 3664
rect 7006 3652 7012 3664
rect 5132 3624 7012 3652
rect 5132 3612 5138 3624
rect 7006 3612 7012 3624
rect 7064 3612 7070 3664
rect 8294 3652 8300 3664
rect 7392 3624 8064 3652
rect 8255 3624 8300 3652
rect 5629 3587 5687 3593
rect 5000 3556 5580 3584
rect 4525 3547 4583 3553
rect 3053 3519 3111 3525
rect 3053 3485 3065 3519
rect 3099 3516 3111 3519
rect 3142 3516 3148 3528
rect 3099 3488 3148 3516
rect 3099 3485 3111 3488
rect 3053 3479 3111 3485
rect 3142 3476 3148 3488
rect 3200 3516 3206 3528
rect 4246 3516 4252 3528
rect 3200 3488 4252 3516
rect 3200 3476 3206 3488
rect 4246 3476 4252 3488
rect 4304 3476 4310 3528
rect 5552 3516 5580 3556
rect 5629 3553 5641 3587
rect 5675 3584 5687 3587
rect 6638 3584 6644 3596
rect 5675 3556 6644 3584
rect 5675 3553 5687 3556
rect 5629 3547 5687 3553
rect 6638 3544 6644 3556
rect 6696 3544 6702 3596
rect 7392 3584 7420 3624
rect 6748 3556 7420 3584
rect 7489 3587 7547 3593
rect 5810 3516 5816 3528
rect 5552 3488 5672 3516
rect 5771 3488 5816 3516
rect 3234 3448 3240 3460
rect 3068 3420 3240 3448
rect 1762 3340 1768 3392
rect 1820 3380 1826 3392
rect 3068 3380 3096 3420
rect 3234 3408 3240 3420
rect 3292 3408 3298 3460
rect 3510 3448 3516 3460
rect 3471 3420 3516 3448
rect 3510 3408 3516 3420
rect 3568 3408 3574 3460
rect 5644 3448 5672 3488
rect 5810 3476 5816 3488
rect 5868 3476 5874 3528
rect 6748 3448 6776 3556
rect 7489 3553 7501 3587
rect 7535 3584 7547 3587
rect 7926 3584 7932 3596
rect 7535 3556 7932 3584
rect 7535 3553 7547 3556
rect 7489 3547 7547 3553
rect 7926 3544 7932 3556
rect 7984 3544 7990 3596
rect 8036 3584 8064 3624
rect 8294 3612 8300 3624
rect 8352 3612 8358 3664
rect 10505 3655 10563 3661
rect 10505 3621 10517 3655
rect 10551 3652 10563 3655
rect 10870 3652 10876 3664
rect 10551 3624 10876 3652
rect 10551 3621 10563 3624
rect 10505 3615 10563 3621
rect 10870 3612 10876 3624
rect 10928 3612 10934 3664
rect 11054 3612 11060 3664
rect 11112 3652 11118 3664
rect 11112 3624 11652 3652
rect 11112 3612 11118 3624
rect 9398 3584 9404 3596
rect 8036 3556 9404 3584
rect 9398 3544 9404 3556
rect 9456 3544 9462 3596
rect 9582 3544 9588 3596
rect 9640 3584 9646 3596
rect 9769 3587 9827 3593
rect 9769 3584 9781 3587
rect 9640 3556 9781 3584
rect 9640 3544 9646 3556
rect 9769 3553 9781 3556
rect 9815 3584 9827 3587
rect 9815 3556 10272 3584
rect 9815 3553 9827 3556
rect 9769 3547 9827 3553
rect 7745 3519 7803 3525
rect 7745 3485 7757 3519
rect 7791 3516 7803 3519
rect 8110 3516 8116 3528
rect 7791 3488 8116 3516
rect 7791 3485 7803 3488
rect 7745 3479 7803 3485
rect 8110 3476 8116 3488
rect 8168 3476 8174 3528
rect 8205 3519 8263 3525
rect 8205 3485 8217 3519
rect 8251 3516 8263 3519
rect 9858 3516 9864 3528
rect 8251 3488 9864 3516
rect 8251 3485 8263 3488
rect 8205 3479 8263 3485
rect 9858 3476 9864 3488
rect 9916 3476 9922 3528
rect 9125 3451 9183 3457
rect 9125 3448 9137 3451
rect 3620 3420 5396 3448
rect 5644 3420 6776 3448
rect 7760 3420 9137 3448
rect 1820 3352 3096 3380
rect 1820 3340 1826 3352
rect 3142 3340 3148 3392
rect 3200 3380 3206 3392
rect 3620 3380 3648 3420
rect 3200 3352 3648 3380
rect 3200 3340 3206 3352
rect 3878 3340 3884 3392
rect 3936 3380 3942 3392
rect 4062 3380 4068 3392
rect 3936 3352 4068 3380
rect 3936 3340 3942 3352
rect 4062 3340 4068 3352
rect 4120 3340 4126 3392
rect 4433 3383 4491 3389
rect 4433 3349 4445 3383
rect 4479 3380 4491 3383
rect 4709 3383 4767 3389
rect 4709 3380 4721 3383
rect 4479 3352 4721 3380
rect 4479 3349 4491 3352
rect 4433 3343 4491 3349
rect 4709 3349 4721 3352
rect 4755 3349 4767 3383
rect 4709 3343 4767 3349
rect 4982 3340 4988 3392
rect 5040 3380 5046 3392
rect 5261 3383 5319 3389
rect 5261 3380 5273 3383
rect 5040 3352 5273 3380
rect 5040 3340 5046 3352
rect 5261 3349 5273 3352
rect 5307 3349 5319 3383
rect 5368 3380 5396 3420
rect 7760 3380 7788 3420
rect 9125 3417 9137 3420
rect 9171 3417 9183 3451
rect 9125 3411 9183 3417
rect 9490 3408 9496 3460
rect 9548 3448 9554 3460
rect 9585 3451 9643 3457
rect 9585 3448 9597 3451
rect 9548 3420 9597 3448
rect 9548 3408 9554 3420
rect 9585 3417 9597 3420
rect 9631 3417 9643 3451
rect 10244 3448 10272 3556
rect 10318 3544 10324 3596
rect 10376 3584 10382 3596
rect 10597 3587 10655 3593
rect 10597 3584 10609 3587
rect 10376 3556 10609 3584
rect 10376 3544 10382 3556
rect 10597 3553 10609 3556
rect 10643 3553 10655 3587
rect 10597 3547 10655 3553
rect 10686 3544 10692 3596
rect 10744 3584 10750 3596
rect 11624 3593 11652 3624
rect 11149 3587 11207 3593
rect 11149 3584 11161 3587
rect 10744 3556 11161 3584
rect 10744 3544 10750 3556
rect 11149 3553 11161 3556
rect 11195 3553 11207 3587
rect 11149 3547 11207 3553
rect 11609 3587 11667 3593
rect 11609 3553 11621 3587
rect 11655 3553 11667 3587
rect 11609 3547 11667 3553
rect 10781 3519 10839 3525
rect 10781 3485 10793 3519
rect 10827 3516 10839 3519
rect 10870 3516 10876 3528
rect 10827 3488 10876 3516
rect 10827 3485 10839 3488
rect 10781 3479 10839 3485
rect 10870 3476 10876 3488
rect 10928 3516 10934 3528
rect 10965 3519 11023 3525
rect 10965 3516 10977 3519
rect 10928 3488 10977 3516
rect 10928 3476 10934 3488
rect 10965 3485 10977 3488
rect 11011 3516 11023 3519
rect 11716 3516 11744 3692
rect 12529 3655 12587 3661
rect 12529 3621 12541 3655
rect 12575 3652 12587 3655
rect 12575 3624 13400 3652
rect 12575 3621 12587 3624
rect 12529 3615 12587 3621
rect 12158 3584 12164 3596
rect 12119 3556 12164 3584
rect 12158 3544 12164 3556
rect 12216 3544 12222 3596
rect 12618 3584 12624 3596
rect 12579 3556 12624 3584
rect 12618 3544 12624 3556
rect 12676 3544 12682 3596
rect 13372 3593 13400 3624
rect 13446 3612 13452 3664
rect 13504 3652 13510 3664
rect 13504 3624 14872 3652
rect 13504 3612 13510 3624
rect 14844 3593 14872 3624
rect 15286 3612 15292 3664
rect 15344 3612 15350 3664
rect 15396 3652 15424 3692
rect 16114 3680 16120 3732
rect 16172 3720 16178 3732
rect 16209 3723 16267 3729
rect 16209 3720 16221 3723
rect 16172 3692 16221 3720
rect 16172 3680 16178 3692
rect 16209 3689 16221 3692
rect 16255 3689 16267 3723
rect 16209 3683 16267 3689
rect 16390 3680 16396 3732
rect 16448 3720 16454 3732
rect 16853 3723 16911 3729
rect 16853 3720 16865 3723
rect 16448 3692 16865 3720
rect 16448 3680 16454 3692
rect 16853 3689 16865 3692
rect 16899 3689 16911 3723
rect 16853 3683 16911 3689
rect 18049 3723 18107 3729
rect 18049 3689 18061 3723
rect 18095 3689 18107 3723
rect 18049 3683 18107 3689
rect 17402 3652 17408 3664
rect 15396 3624 17408 3652
rect 17402 3612 17408 3624
rect 17460 3612 17466 3664
rect 17681 3655 17739 3661
rect 17681 3621 17693 3655
rect 17727 3652 17739 3655
rect 18064 3652 18092 3683
rect 18690 3680 18696 3732
rect 18748 3720 18754 3732
rect 19705 3723 19763 3729
rect 18748 3692 19012 3720
rect 18748 3680 18754 3692
rect 17727 3624 18092 3652
rect 17727 3621 17739 3624
rect 17681 3615 17739 3621
rect 13357 3587 13415 3593
rect 13357 3553 13369 3587
rect 13403 3553 13415 3587
rect 13357 3547 13415 3553
rect 13633 3587 13691 3593
rect 13633 3553 13645 3587
rect 13679 3553 13691 3587
rect 13633 3547 13691 3553
rect 14829 3587 14887 3593
rect 14829 3553 14841 3587
rect 14875 3553 14887 3587
rect 14829 3547 14887 3553
rect 15096 3587 15154 3593
rect 15096 3553 15108 3587
rect 15142 3584 15154 3587
rect 15304 3584 15332 3612
rect 15142 3556 17080 3584
rect 15142 3553 15154 3556
rect 15096 3547 15154 3553
rect 13648 3516 13676 3547
rect 11011 3488 11744 3516
rect 11808 3488 13676 3516
rect 11011 3485 11023 3488
rect 10965 3479 11023 3485
rect 11808 3457 11836 3488
rect 16666 3476 16672 3528
rect 16724 3516 16730 3528
rect 17052 3525 17080 3556
rect 17126 3544 17132 3596
rect 17184 3584 17190 3596
rect 18233 3587 18291 3593
rect 18233 3584 18245 3587
rect 17184 3556 18245 3584
rect 17184 3544 17190 3556
rect 18233 3553 18245 3556
rect 18279 3553 18291 3587
rect 18233 3547 18291 3553
rect 18693 3587 18751 3593
rect 18693 3553 18705 3587
rect 18739 3553 18751 3587
rect 18984 3584 19012 3692
rect 19705 3689 19717 3723
rect 19751 3720 19763 3723
rect 20622 3720 20628 3732
rect 19751 3692 20628 3720
rect 19751 3689 19763 3692
rect 19705 3683 19763 3689
rect 20622 3680 20628 3692
rect 20680 3680 20686 3732
rect 19058 3612 19064 3664
rect 19116 3652 19122 3664
rect 20165 3655 20223 3661
rect 20165 3652 20177 3655
rect 19116 3624 20177 3652
rect 19116 3612 19122 3624
rect 20165 3621 20177 3624
rect 20211 3621 20223 3655
rect 20165 3615 20223 3621
rect 19153 3587 19211 3593
rect 19153 3584 19165 3587
rect 18984 3556 19165 3584
rect 18693 3547 18751 3553
rect 19153 3553 19165 3556
rect 19199 3553 19211 3587
rect 19153 3547 19211 3553
rect 16945 3519 17003 3525
rect 16945 3516 16957 3519
rect 16724 3488 16957 3516
rect 16724 3476 16730 3488
rect 16945 3485 16957 3488
rect 16991 3485 17003 3519
rect 16945 3479 17003 3485
rect 17037 3519 17095 3525
rect 17037 3485 17049 3519
rect 17083 3485 17095 3519
rect 17037 3479 17095 3485
rect 17954 3476 17960 3528
rect 18012 3516 18018 3528
rect 18708 3516 18736 3547
rect 19518 3544 19524 3596
rect 19576 3584 19582 3596
rect 20809 3587 20867 3593
rect 20809 3584 20821 3587
rect 19576 3556 20821 3584
rect 19576 3544 19582 3556
rect 20809 3553 20821 3556
rect 20855 3553 20867 3587
rect 20809 3547 20867 3553
rect 20530 3516 20536 3528
rect 18012 3488 18736 3516
rect 19168 3488 20536 3516
rect 18012 3476 18018 3488
rect 11793 3451 11851 3457
rect 10244 3420 11652 3448
rect 9585 3411 9643 3417
rect 8754 3380 8760 3392
rect 5368 3352 7788 3380
rect 8715 3352 8760 3380
rect 5261 3343 5319 3349
rect 8754 3340 8760 3352
rect 8812 3340 8818 3392
rect 10042 3340 10048 3392
rect 10100 3380 10106 3392
rect 10137 3383 10195 3389
rect 10137 3380 10149 3383
rect 10100 3352 10149 3380
rect 10100 3340 10106 3352
rect 10137 3349 10149 3352
rect 10183 3349 10195 3383
rect 11624 3380 11652 3420
rect 11793 3417 11805 3451
rect 11839 3417 11851 3451
rect 14369 3451 14427 3457
rect 14369 3448 14381 3451
rect 11793 3411 11851 3417
rect 11900 3420 14381 3448
rect 11900 3380 11928 3420
rect 14369 3417 14381 3420
rect 14415 3417 14427 3451
rect 14369 3411 14427 3417
rect 16390 3408 16396 3460
rect 16448 3448 16454 3460
rect 17497 3451 17555 3457
rect 17497 3448 17509 3451
rect 16448 3420 17509 3448
rect 16448 3408 16454 3420
rect 17497 3417 17509 3420
rect 17543 3417 17555 3451
rect 19168 3448 19196 3488
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 19978 3448 19984 3460
rect 17497 3411 17555 3417
rect 17880 3420 19196 3448
rect 19939 3420 19984 3448
rect 11624 3352 11928 3380
rect 12345 3383 12403 3389
rect 10137 3343 10195 3349
rect 12345 3349 12357 3383
rect 12391 3380 12403 3383
rect 12529 3383 12587 3389
rect 12529 3380 12541 3383
rect 12391 3352 12541 3380
rect 12391 3349 12403 3352
rect 12345 3343 12403 3349
rect 12529 3349 12541 3352
rect 12575 3349 12587 3383
rect 12529 3343 12587 3349
rect 12805 3383 12863 3389
rect 12805 3349 12817 3383
rect 12851 3380 12863 3383
rect 12986 3380 12992 3392
rect 12851 3352 12992 3380
rect 12851 3349 12863 3352
rect 12805 3343 12863 3349
rect 12986 3340 12992 3352
rect 13044 3340 13050 3392
rect 13078 3340 13084 3392
rect 13136 3380 13142 3392
rect 13173 3383 13231 3389
rect 13173 3380 13185 3383
rect 13136 3352 13185 3380
rect 13136 3340 13142 3352
rect 13173 3349 13185 3352
rect 13219 3349 13231 3383
rect 13173 3343 13231 3349
rect 13817 3383 13875 3389
rect 13817 3349 13829 3383
rect 13863 3380 13875 3383
rect 16206 3380 16212 3392
rect 13863 3352 16212 3380
rect 13863 3349 13875 3352
rect 13817 3343 13875 3349
rect 16206 3340 16212 3352
rect 16264 3340 16270 3392
rect 16298 3340 16304 3392
rect 16356 3380 16362 3392
rect 16485 3383 16543 3389
rect 16485 3380 16497 3383
rect 16356 3352 16497 3380
rect 16356 3340 16362 3352
rect 16485 3349 16497 3352
rect 16531 3349 16543 3383
rect 16485 3343 16543 3349
rect 16574 3340 16580 3392
rect 16632 3380 16638 3392
rect 17880 3380 17908 3420
rect 19978 3408 19984 3420
rect 20036 3408 20042 3460
rect 16632 3352 17908 3380
rect 16632 3340 16638 3352
rect 17954 3340 17960 3392
rect 18012 3380 18018 3392
rect 18509 3383 18567 3389
rect 18509 3380 18521 3383
rect 18012 3352 18521 3380
rect 18012 3340 18018 3352
rect 18509 3349 18521 3352
rect 18555 3349 18567 3383
rect 18966 3380 18972 3392
rect 18927 3352 18972 3380
rect 18509 3343 18567 3349
rect 18966 3340 18972 3352
rect 19024 3340 19030 3392
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 1762 3176 1768 3188
rect 1723 3148 1768 3176
rect 1762 3136 1768 3148
rect 1820 3136 1826 3188
rect 6638 3176 6644 3188
rect 2746 3148 5856 3176
rect 6599 3148 6644 3176
rect 198 3000 204 3052
rect 256 3040 262 3052
rect 1670 3040 1676 3052
rect 256 3012 1676 3040
rect 256 3000 262 3012
rect 1670 3000 1676 3012
rect 1728 3040 1734 3052
rect 2746 3040 2774 3148
rect 5828 3108 5856 3148
rect 6638 3136 6644 3148
rect 6696 3136 6702 3188
rect 7926 3136 7932 3188
rect 7984 3176 7990 3188
rect 8021 3179 8079 3185
rect 8021 3176 8033 3179
rect 7984 3148 8033 3176
rect 7984 3136 7990 3148
rect 8021 3145 8033 3148
rect 8067 3176 8079 3179
rect 8202 3176 8208 3188
rect 8067 3148 8208 3176
rect 8067 3145 8079 3148
rect 8021 3139 8079 3145
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 8478 3136 8484 3188
rect 8536 3176 8542 3188
rect 12161 3179 12219 3185
rect 12161 3176 12173 3179
rect 8536 3148 12173 3176
rect 8536 3136 8542 3148
rect 12161 3145 12173 3148
rect 12207 3145 12219 3179
rect 14274 3176 14280 3188
rect 12161 3139 12219 3145
rect 12406 3148 14280 3176
rect 7653 3111 7711 3117
rect 7653 3108 7665 3111
rect 5828 3080 7665 3108
rect 7653 3077 7665 3080
rect 7699 3077 7711 3111
rect 7653 3071 7711 3077
rect 9398 3068 9404 3120
rect 9456 3108 9462 3120
rect 12406 3108 12434 3148
rect 14274 3136 14280 3148
rect 14332 3136 14338 3188
rect 15378 3176 15384 3188
rect 15339 3148 15384 3176
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 15930 3136 15936 3188
rect 15988 3176 15994 3188
rect 17773 3179 17831 3185
rect 17773 3176 17785 3179
rect 15988 3148 17785 3176
rect 15988 3136 15994 3148
rect 17773 3145 17785 3148
rect 17819 3145 17831 3179
rect 17773 3139 17831 3145
rect 17862 3136 17868 3188
rect 17920 3176 17926 3188
rect 17920 3148 20576 3176
rect 17920 3136 17926 3148
rect 12526 3108 12532 3120
rect 9456 3080 12434 3108
rect 12487 3080 12532 3108
rect 9456 3068 9462 3080
rect 4706 3040 4712 3052
rect 1728 3012 2774 3040
rect 4080 3012 4712 3040
rect 1728 3000 1734 3012
rect 2225 2975 2283 2981
rect 2225 2941 2237 2975
rect 2271 2972 2283 2975
rect 2958 2972 2964 2984
rect 2271 2944 2964 2972
rect 2271 2941 2283 2944
rect 2225 2935 2283 2941
rect 2958 2932 2964 2944
rect 3016 2932 3022 2984
rect 3602 2972 3608 2984
rect 3252 2944 3608 2972
rect 3252 2916 3280 2944
rect 3602 2932 3608 2944
rect 3660 2972 3666 2984
rect 4080 2972 4108 3012
rect 4706 3000 4712 3012
rect 4764 3000 4770 3052
rect 6270 3000 6276 3052
rect 6328 3040 6334 3052
rect 7193 3043 7251 3049
rect 7193 3040 7205 3043
rect 6328 3012 7205 3040
rect 6328 3000 6334 3012
rect 7193 3009 7205 3012
rect 7239 3009 7251 3043
rect 7193 3003 7251 3009
rect 9585 3043 9643 3049
rect 9585 3009 9597 3043
rect 9631 3040 9643 3043
rect 9858 3040 9864 3052
rect 9631 3012 9864 3040
rect 9631 3009 9643 3012
rect 9585 3003 9643 3009
rect 9858 3000 9864 3012
rect 9916 3000 9922 3052
rect 10594 3040 10600 3052
rect 10555 3012 10600 3040
rect 10594 3000 10600 3012
rect 10652 3000 10658 3052
rect 10781 3043 10839 3049
rect 10781 3009 10793 3043
rect 10827 3040 10839 3043
rect 10870 3040 10876 3052
rect 10827 3012 10876 3040
rect 10827 3009 10839 3012
rect 10781 3003 10839 3009
rect 10870 3000 10876 3012
rect 10928 3000 10934 3052
rect 3660 2944 4108 2972
rect 4157 2975 4215 2981
rect 3660 2932 3666 2944
rect 4157 2941 4169 2975
rect 4203 2972 4215 2975
rect 4246 2972 4252 2984
rect 4203 2944 4252 2972
rect 4203 2941 4215 2944
rect 4157 2935 4215 2941
rect 4246 2932 4252 2944
rect 4304 2932 4310 2984
rect 4614 2932 4620 2984
rect 4672 2972 4678 2984
rect 5166 2972 5172 2984
rect 4672 2944 5172 2972
rect 4672 2932 4678 2944
rect 5166 2932 5172 2944
rect 5224 2932 5230 2984
rect 5810 2972 5816 2984
rect 5771 2944 5816 2972
rect 5810 2932 5816 2944
rect 5868 2932 5874 2984
rect 6730 2932 6736 2984
rect 6788 2972 6794 2984
rect 7009 2975 7067 2981
rect 7009 2972 7021 2975
rect 6788 2944 7021 2972
rect 6788 2932 6794 2944
rect 7009 2941 7021 2944
rect 7055 2941 7067 2975
rect 7009 2935 7067 2941
rect 9145 2975 9203 2981
rect 9145 2941 9157 2975
rect 9191 2972 9203 2975
rect 9191 2944 9260 2972
rect 9191 2941 9203 2944
rect 9145 2935 9203 2941
rect 1673 2907 1731 2913
rect 1673 2873 1685 2907
rect 1719 2904 1731 2907
rect 1854 2904 1860 2916
rect 1719 2876 1860 2904
rect 1719 2873 1731 2876
rect 1673 2867 1731 2873
rect 1854 2864 1860 2876
rect 1912 2864 1918 2916
rect 2409 2907 2467 2913
rect 2409 2873 2421 2907
rect 2455 2904 2467 2907
rect 2866 2904 2872 2916
rect 2455 2876 2872 2904
rect 2455 2873 2467 2876
rect 2409 2867 2467 2873
rect 2866 2864 2872 2876
rect 2924 2864 2930 2916
rect 3234 2864 3240 2916
rect 3292 2864 3298 2916
rect 3912 2907 3970 2913
rect 3912 2873 3924 2907
rect 3958 2904 3970 2907
rect 5442 2904 5448 2916
rect 3958 2876 5448 2904
rect 3958 2873 3970 2876
rect 3912 2867 3970 2873
rect 2774 2796 2780 2848
rect 2832 2836 2838 2848
rect 4246 2836 4252 2848
rect 2832 2808 4252 2836
rect 2832 2796 2838 2808
rect 4246 2796 4252 2808
rect 4304 2796 4310 2848
rect 4448 2845 4476 2876
rect 5442 2864 5448 2876
rect 5500 2864 5506 2916
rect 5568 2907 5626 2913
rect 5568 2873 5580 2907
rect 5614 2904 5626 2907
rect 6270 2904 6276 2916
rect 5614 2876 6276 2904
rect 5614 2873 5626 2876
rect 5568 2867 5626 2873
rect 6270 2864 6276 2876
rect 6328 2864 6334 2916
rect 8662 2904 8668 2916
rect 6472 2876 8668 2904
rect 4433 2839 4491 2845
rect 4433 2805 4445 2839
rect 4479 2805 4491 2839
rect 4433 2799 4491 2805
rect 4706 2796 4712 2848
rect 4764 2836 4770 2848
rect 6472 2836 6500 2876
rect 8662 2864 8668 2876
rect 8720 2864 8726 2916
rect 4764 2808 6500 2836
rect 4764 2796 4770 2808
rect 6638 2796 6644 2848
rect 6696 2836 6702 2848
rect 6822 2836 6828 2848
rect 6696 2808 6828 2836
rect 6696 2796 6702 2808
rect 6822 2796 6828 2808
rect 6880 2836 6886 2848
rect 7101 2839 7159 2845
rect 7101 2836 7113 2839
rect 6880 2808 7113 2836
rect 6880 2796 6886 2808
rect 7101 2805 7113 2808
rect 7147 2805 7159 2839
rect 7101 2799 7159 2805
rect 7742 2796 7748 2848
rect 7800 2836 7806 2848
rect 9122 2836 9128 2848
rect 7800 2808 9128 2836
rect 7800 2796 7806 2808
rect 9122 2796 9128 2808
rect 9180 2796 9186 2848
rect 9232 2836 9260 2944
rect 9306 2932 9312 2984
rect 9364 2972 9370 2984
rect 9401 2975 9459 2981
rect 9401 2972 9413 2975
rect 9364 2944 9413 2972
rect 9364 2932 9370 2944
rect 9401 2941 9413 2944
rect 9447 2941 9459 2975
rect 9674 2972 9680 2984
rect 9635 2944 9680 2972
rect 9401 2935 9459 2941
rect 9674 2932 9680 2944
rect 9732 2932 9738 2984
rect 9766 2932 9772 2984
rect 9824 2972 9830 2984
rect 11149 2975 11207 2981
rect 11149 2972 11161 2975
rect 9824 2944 11161 2972
rect 9824 2932 9830 2944
rect 11149 2941 11161 2944
rect 11195 2941 11207 2975
rect 11149 2935 11207 2941
rect 9490 2864 9496 2916
rect 9548 2904 9554 2916
rect 9692 2904 9720 2932
rect 9548 2876 9720 2904
rect 10505 2907 10563 2913
rect 9548 2864 9554 2876
rect 10505 2873 10517 2907
rect 10551 2904 10563 2907
rect 11256 2904 11284 3080
rect 12526 3068 12532 3080
rect 12584 3068 12590 3120
rect 13081 3111 13139 3117
rect 13081 3077 13093 3111
rect 13127 3108 13139 3111
rect 14090 3108 14096 3120
rect 13127 3080 14096 3108
rect 13127 3077 13139 3080
rect 13081 3071 13139 3077
rect 14090 3068 14096 3080
rect 14148 3068 14154 3120
rect 15194 3068 15200 3120
rect 15252 3108 15258 3120
rect 16577 3111 16635 3117
rect 15252 3080 16436 3108
rect 15252 3068 15258 3080
rect 11698 3000 11704 3052
rect 11756 3040 11762 3052
rect 15838 3040 15844 3052
rect 11756 3012 13860 3040
rect 15799 3012 15844 3040
rect 11756 3000 11762 3012
rect 11885 2975 11943 2981
rect 11885 2972 11897 2975
rect 10551 2876 11284 2904
rect 11348 2944 11897 2972
rect 10551 2873 10563 2876
rect 10505 2867 10563 2873
rect 9585 2839 9643 2845
rect 9585 2836 9597 2839
rect 9232 2808 9597 2836
rect 9585 2805 9597 2808
rect 9631 2805 9643 2839
rect 9585 2799 9643 2805
rect 9861 2839 9919 2845
rect 9861 2805 9873 2839
rect 9907 2836 9919 2839
rect 9950 2836 9956 2848
rect 9907 2808 9956 2836
rect 9907 2805 9919 2808
rect 9861 2799 9919 2805
rect 9950 2796 9956 2808
rect 10008 2796 10014 2848
rect 10134 2836 10140 2848
rect 10095 2808 10140 2836
rect 10134 2796 10140 2808
rect 10192 2796 10198 2848
rect 11348 2845 11376 2944
rect 11885 2941 11897 2944
rect 11931 2941 11943 2975
rect 11885 2935 11943 2941
rect 12161 2975 12219 2981
rect 12161 2941 12173 2975
rect 12207 2972 12219 2975
rect 12345 2975 12403 2981
rect 12345 2972 12357 2975
rect 12207 2944 12357 2972
rect 12207 2941 12219 2944
rect 12161 2935 12219 2941
rect 12345 2941 12357 2944
rect 12391 2941 12403 2975
rect 12894 2972 12900 2984
rect 12855 2944 12900 2972
rect 12345 2935 12403 2941
rect 12894 2932 12900 2944
rect 12952 2932 12958 2984
rect 12986 2932 12992 2984
rect 13044 2972 13050 2984
rect 13832 2981 13860 3012
rect 15838 3000 15844 3012
rect 15896 3000 15902 3052
rect 16025 3043 16083 3049
rect 16025 3009 16037 3043
rect 16071 3040 16083 3043
rect 16114 3040 16120 3052
rect 16071 3012 16120 3040
rect 16071 3009 16083 3012
rect 16025 3003 16083 3009
rect 16114 3000 16120 3012
rect 16172 3000 16178 3052
rect 13541 2975 13599 2981
rect 13541 2972 13553 2975
rect 13044 2944 13553 2972
rect 13044 2932 13050 2944
rect 13541 2941 13553 2944
rect 13587 2941 13599 2975
rect 13541 2935 13599 2941
rect 13817 2975 13875 2981
rect 13817 2941 13829 2975
rect 13863 2941 13875 2975
rect 13817 2935 13875 2941
rect 15749 2975 15807 2981
rect 15749 2941 15761 2975
rect 15795 2972 15807 2975
rect 16298 2972 16304 2984
rect 15795 2944 16304 2972
rect 15795 2941 15807 2944
rect 15749 2935 15807 2941
rect 16298 2932 16304 2944
rect 16356 2932 16362 2984
rect 16408 2981 16436 3080
rect 16577 3077 16589 3111
rect 16623 3077 16635 3111
rect 16577 3071 16635 3077
rect 16393 2975 16451 2981
rect 16393 2941 16405 2975
rect 16439 2941 16451 2975
rect 16592 2972 16620 3071
rect 17218 3068 17224 3120
rect 17276 3108 17282 3120
rect 20438 3108 20444 3120
rect 17276 3080 20444 3108
rect 17276 3068 17282 3080
rect 20438 3068 20444 3080
rect 20496 3068 20502 3120
rect 17034 3000 17040 3052
rect 17092 3040 17098 3052
rect 17092 3012 19012 3040
rect 17092 3000 17098 3012
rect 17865 2975 17923 2981
rect 17865 2972 17877 2975
rect 16592 2944 17877 2972
rect 16393 2935 16451 2941
rect 17865 2941 17877 2944
rect 17911 2941 17923 2975
rect 17865 2935 17923 2941
rect 18601 2975 18659 2981
rect 18601 2941 18613 2975
rect 18647 2972 18659 2975
rect 18874 2972 18880 2984
rect 18647 2944 18880 2972
rect 18647 2941 18659 2944
rect 18601 2935 18659 2941
rect 18874 2932 18880 2944
rect 18932 2932 18938 2984
rect 18984 2972 19012 3012
rect 19150 3000 19156 3052
rect 19208 3040 19214 3052
rect 19208 3012 19840 3040
rect 19208 3000 19214 3012
rect 18984 2944 19196 2972
rect 12434 2864 12440 2916
rect 12492 2864 12498 2916
rect 14550 2904 14556 2916
rect 14511 2876 14556 2904
rect 14550 2864 14556 2876
rect 14608 2864 14614 2916
rect 14737 2907 14795 2913
rect 14737 2873 14749 2907
rect 14783 2873 14795 2907
rect 14737 2867 14795 2873
rect 11333 2839 11391 2845
rect 11333 2805 11345 2839
rect 11379 2805 11391 2839
rect 11333 2799 11391 2805
rect 12069 2839 12127 2845
rect 12069 2805 12081 2839
rect 12115 2836 12127 2839
rect 12452 2836 12480 2864
rect 13354 2836 13360 2848
rect 12115 2808 12480 2836
rect 13315 2808 13360 2836
rect 12115 2805 12127 2808
rect 12069 2799 12127 2805
rect 13354 2796 13360 2808
rect 13412 2796 13418 2848
rect 14001 2839 14059 2845
rect 14001 2805 14013 2839
rect 14047 2836 14059 2839
rect 14752 2836 14780 2867
rect 16206 2864 16212 2916
rect 16264 2904 16270 2916
rect 17313 2907 17371 2913
rect 17313 2904 17325 2907
rect 16264 2876 17325 2904
rect 16264 2864 16270 2876
rect 17313 2873 17325 2876
rect 17359 2873 17371 2907
rect 19058 2904 19064 2916
rect 19019 2876 19064 2904
rect 17313 2867 17371 2873
rect 19058 2864 19064 2876
rect 19116 2864 19122 2916
rect 19168 2904 19196 2944
rect 19242 2932 19248 2984
rect 19300 2981 19306 2984
rect 19812 2981 19840 3012
rect 19300 2975 19320 2981
rect 19308 2941 19320 2975
rect 19797 2975 19855 2981
rect 19300 2935 19320 2941
rect 19352 2944 19748 2972
rect 19300 2932 19306 2935
rect 19352 2904 19380 2944
rect 19168 2876 19380 2904
rect 19518 2864 19524 2916
rect 19576 2904 19582 2916
rect 19613 2907 19671 2913
rect 19613 2904 19625 2907
rect 19576 2876 19625 2904
rect 19576 2864 19582 2876
rect 19613 2873 19625 2876
rect 19659 2873 19671 2907
rect 19720 2904 19748 2944
rect 19797 2941 19809 2975
rect 19843 2941 19855 2975
rect 20548 2972 20576 3148
rect 21085 2975 21143 2981
rect 21085 2972 21097 2975
rect 20548 2944 21097 2972
rect 19797 2935 19855 2941
rect 21085 2941 21097 2944
rect 21131 2972 21143 2975
rect 22738 2972 22744 2984
rect 21131 2944 22744 2972
rect 21131 2941 21143 2944
rect 21085 2935 21143 2941
rect 22738 2932 22744 2944
rect 22796 2932 22802 2984
rect 20441 2907 20499 2913
rect 20441 2904 20453 2907
rect 19720 2876 20453 2904
rect 19613 2867 19671 2873
rect 20441 2873 20453 2876
rect 20487 2873 20499 2907
rect 20441 2867 20499 2873
rect 14047 2808 14780 2836
rect 14047 2805 14059 2808
rect 14001 2799 14059 2805
rect 15470 2796 15476 2848
rect 15528 2836 15534 2848
rect 17221 2839 17279 2845
rect 17221 2836 17233 2839
rect 15528 2808 17233 2836
rect 15528 2796 15534 2808
rect 17221 2805 17233 2808
rect 17267 2805 17279 2839
rect 17221 2799 17279 2805
rect 18693 2839 18751 2845
rect 18693 2805 18705 2839
rect 18739 2836 18751 2839
rect 20898 2836 20904 2848
rect 18739 2808 20904 2836
rect 18739 2805 18751 2808
rect 18693 2799 18751 2805
rect 20898 2796 20904 2808
rect 20956 2796 20962 2848
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 2869 2635 2927 2641
rect 2869 2601 2881 2635
rect 2915 2632 2927 2635
rect 3234 2632 3240 2644
rect 2915 2604 3240 2632
rect 2915 2601 2927 2604
rect 2869 2595 2927 2601
rect 3234 2592 3240 2604
rect 3292 2592 3298 2644
rect 3329 2635 3387 2641
rect 3329 2601 3341 2635
rect 3375 2632 3387 2635
rect 5445 2635 5503 2641
rect 3375 2604 5396 2632
rect 3375 2601 3387 2604
rect 3329 2595 3387 2601
rect 1670 2564 1676 2576
rect 1631 2536 1676 2564
rect 1670 2524 1676 2536
rect 1728 2524 1734 2576
rect 1857 2567 1915 2573
rect 1857 2533 1869 2567
rect 1903 2564 1915 2567
rect 2130 2564 2136 2576
rect 1903 2536 2136 2564
rect 1903 2533 1915 2536
rect 1857 2527 1915 2533
rect 2130 2524 2136 2536
rect 2188 2524 2194 2576
rect 2406 2564 2412 2576
rect 2367 2536 2412 2564
rect 2406 2524 2412 2536
rect 2464 2524 2470 2576
rect 3878 2524 3884 2576
rect 3936 2564 3942 2576
rect 4157 2567 4215 2573
rect 4157 2564 4169 2567
rect 3936 2536 4169 2564
rect 3936 2524 3942 2536
rect 4157 2533 4169 2536
rect 4203 2564 4215 2567
rect 4706 2564 4712 2576
rect 4203 2536 4712 2564
rect 4203 2533 4215 2536
rect 4157 2527 4215 2533
rect 4706 2524 4712 2536
rect 4764 2524 4770 2576
rect 4890 2524 4896 2576
rect 4948 2564 4954 2576
rect 5077 2567 5135 2573
rect 5077 2564 5089 2567
rect 4948 2536 5089 2564
rect 4948 2524 4954 2536
rect 5077 2533 5089 2536
rect 5123 2533 5135 2567
rect 5368 2564 5396 2604
rect 5445 2601 5457 2635
rect 5491 2632 5503 2635
rect 5629 2635 5687 2641
rect 5629 2632 5641 2635
rect 5491 2604 5641 2632
rect 5491 2601 5503 2604
rect 5445 2595 5503 2601
rect 5629 2601 5641 2604
rect 5675 2601 5687 2635
rect 5629 2595 5687 2601
rect 5905 2635 5963 2641
rect 5905 2601 5917 2635
rect 5951 2632 5963 2635
rect 6730 2632 6736 2644
rect 5951 2604 6736 2632
rect 5951 2601 5963 2604
rect 5905 2595 5963 2601
rect 6730 2592 6736 2604
rect 6788 2592 6794 2644
rect 7282 2592 7288 2644
rect 7340 2632 7346 2644
rect 7377 2635 7435 2641
rect 7377 2632 7389 2635
rect 7340 2604 7389 2632
rect 7340 2592 7346 2604
rect 7377 2601 7389 2604
rect 7423 2601 7435 2635
rect 7377 2595 7435 2601
rect 8481 2635 8539 2641
rect 8481 2601 8493 2635
rect 8527 2632 8539 2635
rect 8754 2632 8760 2644
rect 8527 2604 8760 2632
rect 8527 2601 8539 2604
rect 8481 2595 8539 2601
rect 8754 2592 8760 2604
rect 8812 2592 8818 2644
rect 8849 2635 8907 2641
rect 8849 2601 8861 2635
rect 8895 2632 8907 2635
rect 9766 2632 9772 2644
rect 8895 2604 9772 2632
rect 8895 2601 8907 2604
rect 8849 2595 8907 2601
rect 9766 2592 9772 2604
rect 9824 2592 9830 2644
rect 10042 2632 10048 2644
rect 10003 2604 10048 2632
rect 10042 2592 10048 2604
rect 10100 2592 10106 2644
rect 10318 2592 10324 2644
rect 10376 2632 10382 2644
rect 10597 2635 10655 2641
rect 10597 2632 10609 2635
rect 10376 2604 10609 2632
rect 10376 2592 10382 2604
rect 10597 2601 10609 2604
rect 10643 2601 10655 2635
rect 13354 2632 13360 2644
rect 10597 2595 10655 2601
rect 12360 2604 13360 2632
rect 6638 2564 6644 2576
rect 5368 2536 6644 2564
rect 5077 2527 5135 2533
rect 6638 2524 6644 2536
rect 6696 2524 6702 2576
rect 9953 2567 10011 2573
rect 6840 2536 8708 2564
rect 2222 2496 2228 2508
rect 2183 2468 2228 2496
rect 2222 2456 2228 2468
rect 2280 2456 2286 2508
rect 2682 2496 2688 2508
rect 2643 2468 2688 2496
rect 2682 2456 2688 2468
rect 2740 2456 2746 2508
rect 3142 2496 3148 2508
rect 3103 2468 3148 2496
rect 3142 2456 3148 2468
rect 3200 2456 3206 2508
rect 4341 2499 4399 2505
rect 4341 2465 4353 2499
rect 4387 2496 4399 2499
rect 5258 2496 5264 2508
rect 4387 2468 5264 2496
rect 4387 2465 4399 2468
rect 4341 2459 4399 2465
rect 5258 2456 5264 2468
rect 5316 2456 5322 2508
rect 5718 2496 5724 2508
rect 5679 2468 5724 2496
rect 5718 2456 5724 2468
rect 5776 2496 5782 2508
rect 6086 2496 6092 2508
rect 5776 2468 6092 2496
rect 5776 2456 5782 2468
rect 6086 2456 6092 2468
rect 6144 2456 6150 2508
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2465 6791 2499
rect 6733 2459 6791 2465
rect 1486 2388 1492 2440
rect 1544 2428 1550 2440
rect 3160 2428 3188 2456
rect 1544 2400 3188 2428
rect 1544 2388 1550 2400
rect 4246 2388 4252 2440
rect 4304 2428 4310 2440
rect 4801 2431 4859 2437
rect 4801 2428 4813 2431
rect 4304 2400 4813 2428
rect 4304 2388 4310 2400
rect 4801 2397 4813 2400
rect 4847 2397 4859 2431
rect 4982 2428 4988 2440
rect 4943 2400 4988 2428
rect 4801 2391 4859 2397
rect 4982 2388 4988 2400
rect 5040 2388 5046 2440
rect 5629 2431 5687 2437
rect 5629 2397 5641 2431
rect 5675 2428 5687 2431
rect 6748 2428 6776 2459
rect 5675 2400 6776 2428
rect 5675 2397 5687 2400
rect 5629 2391 5687 2397
rect 3694 2320 3700 2372
rect 3752 2360 3758 2372
rect 4614 2360 4620 2372
rect 3752 2332 4620 2360
rect 3752 2320 3758 2332
rect 4614 2320 4620 2332
rect 4672 2320 4678 2372
rect 4706 2320 4712 2372
rect 4764 2360 4770 2372
rect 6840 2360 6868 2536
rect 7193 2499 7251 2505
rect 7193 2465 7205 2499
rect 7239 2496 7251 2499
rect 7374 2496 7380 2508
rect 7239 2468 7380 2496
rect 7239 2465 7251 2468
rect 7193 2459 7251 2465
rect 7374 2456 7380 2468
rect 7432 2456 7438 2508
rect 7837 2499 7895 2505
rect 7837 2465 7849 2499
rect 7883 2496 7895 2499
rect 8570 2496 8576 2508
rect 7883 2468 8576 2496
rect 7883 2465 7895 2468
rect 7837 2459 7895 2465
rect 8570 2456 8576 2468
rect 8628 2456 8634 2508
rect 8680 2496 8708 2536
rect 9953 2533 9965 2567
rect 9999 2564 10011 2567
rect 10134 2564 10140 2576
rect 9999 2536 10140 2564
rect 9999 2533 10011 2536
rect 9953 2527 10011 2533
rect 10134 2524 10140 2536
rect 10192 2524 10198 2576
rect 12360 2573 12388 2604
rect 13354 2592 13360 2604
rect 13412 2592 13418 2644
rect 17770 2632 17776 2644
rect 16132 2604 17776 2632
rect 12345 2567 12403 2573
rect 12345 2533 12357 2567
rect 12391 2533 12403 2567
rect 12345 2527 12403 2533
rect 12434 2524 12440 2576
rect 12492 2564 12498 2576
rect 12989 2567 13047 2573
rect 12989 2564 13001 2567
rect 12492 2536 13001 2564
rect 12492 2524 12498 2536
rect 12989 2533 13001 2536
rect 13035 2533 13047 2567
rect 14090 2564 14096 2576
rect 14051 2536 14096 2564
rect 12989 2527 13047 2533
rect 14090 2524 14096 2536
rect 14148 2524 14154 2576
rect 16132 2573 16160 2604
rect 17770 2592 17776 2604
rect 17828 2592 17834 2644
rect 20073 2635 20131 2641
rect 20073 2632 20085 2635
rect 18800 2604 20085 2632
rect 16117 2567 16175 2573
rect 16117 2533 16129 2567
rect 16163 2533 16175 2567
rect 17494 2564 17500 2576
rect 16117 2527 16175 2533
rect 16592 2536 17500 2564
rect 8680 2468 10272 2496
rect 8202 2428 8208 2440
rect 8163 2400 8208 2428
rect 8202 2388 8208 2400
rect 8260 2388 8266 2440
rect 8389 2431 8447 2437
rect 8389 2397 8401 2431
rect 8435 2428 8447 2431
rect 8435 2400 9628 2428
rect 8435 2397 8447 2400
rect 8389 2391 8447 2397
rect 4764 2332 6868 2360
rect 7653 2363 7711 2369
rect 4764 2320 4770 2332
rect 7653 2329 7665 2363
rect 7699 2360 7711 2363
rect 9030 2360 9036 2372
rect 7699 2332 9036 2360
rect 7699 2329 7711 2332
rect 7653 2323 7711 2329
rect 9030 2320 9036 2332
rect 9088 2320 9094 2372
rect 9600 2369 9628 2400
rect 9858 2388 9864 2440
rect 9916 2428 9922 2440
rect 10137 2431 10195 2437
rect 10137 2428 10149 2431
rect 9916 2400 10149 2428
rect 9916 2388 9922 2400
rect 10137 2397 10149 2400
rect 10183 2397 10195 2431
rect 10244 2428 10272 2468
rect 10686 2456 10692 2508
rect 10744 2496 10750 2508
rect 10781 2499 10839 2505
rect 10781 2496 10793 2499
rect 10744 2468 10793 2496
rect 10744 2456 10750 2468
rect 10781 2465 10793 2468
rect 10827 2465 10839 2499
rect 10781 2459 10839 2465
rect 11333 2499 11391 2505
rect 11333 2465 11345 2499
rect 11379 2496 11391 2499
rect 11379 2468 12434 2496
rect 11379 2465 11391 2468
rect 11333 2459 11391 2465
rect 11885 2431 11943 2437
rect 11885 2428 11897 2431
rect 10244 2400 11897 2428
rect 10137 2391 10195 2397
rect 11885 2397 11897 2400
rect 11931 2397 11943 2431
rect 12406 2428 12434 2468
rect 12526 2456 12532 2508
rect 12584 2496 12590 2508
rect 13541 2499 13599 2505
rect 13541 2496 13553 2499
rect 12584 2468 13553 2496
rect 12584 2456 12590 2468
rect 13541 2465 13553 2468
rect 13587 2465 13599 2499
rect 15010 2496 15016 2508
rect 14971 2468 15016 2496
rect 13541 2459 13599 2465
rect 15010 2456 15016 2468
rect 15068 2456 15074 2508
rect 15565 2499 15623 2505
rect 15565 2465 15577 2499
rect 15611 2496 15623 2499
rect 16592 2496 16620 2536
rect 17494 2524 17500 2536
rect 17552 2524 17558 2576
rect 17589 2567 17647 2573
rect 17589 2533 17601 2567
rect 17635 2564 17647 2567
rect 17954 2564 17960 2576
rect 17635 2536 17960 2564
rect 17635 2533 17647 2536
rect 17589 2527 17647 2533
rect 17954 2524 17960 2536
rect 18012 2524 18018 2576
rect 18138 2564 18144 2576
rect 18099 2536 18144 2564
rect 18138 2524 18144 2536
rect 18196 2524 18202 2576
rect 18800 2573 18828 2604
rect 20073 2601 20085 2604
rect 20119 2601 20131 2635
rect 20073 2595 20131 2601
rect 18785 2567 18843 2573
rect 18785 2533 18797 2567
rect 18831 2533 18843 2567
rect 18785 2527 18843 2533
rect 19150 2524 19156 2576
rect 19208 2564 19214 2576
rect 19429 2567 19487 2573
rect 19429 2564 19441 2567
rect 19208 2536 19441 2564
rect 19208 2524 19214 2536
rect 19429 2533 19441 2536
rect 19475 2533 19487 2567
rect 19429 2527 19487 2533
rect 15611 2468 16620 2496
rect 16669 2499 16727 2505
rect 15611 2465 15623 2468
rect 15565 2459 15623 2465
rect 16669 2465 16681 2499
rect 16715 2496 16727 2499
rect 19242 2496 19248 2508
rect 16715 2468 18552 2496
rect 19203 2468 19248 2496
rect 16715 2465 16727 2468
rect 16669 2459 16727 2465
rect 13078 2428 13084 2440
rect 12406 2400 13084 2428
rect 11885 2391 11943 2397
rect 13078 2388 13084 2400
rect 13136 2388 13142 2440
rect 14090 2428 14096 2440
rect 13188 2400 14096 2428
rect 9585 2363 9643 2369
rect 9585 2329 9597 2363
rect 9631 2329 9643 2363
rect 9585 2323 9643 2329
rect 11517 2363 11575 2369
rect 11517 2329 11529 2363
rect 11563 2360 11575 2363
rect 12618 2360 12624 2372
rect 11563 2332 12624 2360
rect 11563 2329 11575 2332
rect 11517 2323 11575 2329
rect 12618 2320 12624 2332
rect 12676 2320 12682 2372
rect 12802 2360 12808 2372
rect 12763 2332 12808 2360
rect 12802 2320 12808 2332
rect 12860 2320 12866 2372
rect 6917 2295 6975 2301
rect 6917 2261 6929 2295
rect 6963 2292 6975 2295
rect 8478 2292 8484 2304
rect 6963 2264 8484 2292
rect 6963 2261 6975 2264
rect 6917 2255 6975 2261
rect 8478 2252 8484 2264
rect 8536 2252 8542 2304
rect 9214 2292 9220 2304
rect 9175 2264 9220 2292
rect 9214 2252 9220 2264
rect 9272 2252 9278 2304
rect 12437 2295 12495 2301
rect 12437 2261 12449 2295
rect 12483 2292 12495 2295
rect 13188 2292 13216 2400
rect 14090 2388 14096 2400
rect 14148 2388 14154 2440
rect 15749 2431 15807 2437
rect 15749 2397 15761 2431
rect 15795 2428 15807 2431
rect 17218 2428 17224 2440
rect 15795 2400 17224 2428
rect 15795 2397 15807 2400
rect 15749 2391 15807 2397
rect 17218 2388 17224 2400
rect 17276 2388 17282 2440
rect 18524 2428 18552 2468
rect 19242 2456 19248 2468
rect 19300 2456 19306 2508
rect 20254 2496 20260 2508
rect 20215 2468 20260 2496
rect 20254 2456 20260 2468
rect 20312 2456 20318 2508
rect 20806 2496 20812 2508
rect 20767 2468 20812 2496
rect 20806 2456 20812 2468
rect 20864 2456 20870 2508
rect 18874 2428 18880 2440
rect 18524 2400 18880 2428
rect 18874 2388 18880 2400
rect 18932 2388 18938 2440
rect 20530 2428 20536 2440
rect 20491 2400 20536 2428
rect 20530 2388 20536 2400
rect 20588 2388 20594 2440
rect 13262 2320 13268 2372
rect 13320 2360 13326 2372
rect 13357 2363 13415 2369
rect 13357 2360 13369 2363
rect 13320 2332 13369 2360
rect 13320 2320 13326 2332
rect 13357 2329 13369 2332
rect 13403 2329 13415 2363
rect 13357 2323 13415 2329
rect 13722 2320 13728 2372
rect 13780 2360 13786 2372
rect 13909 2363 13967 2369
rect 13909 2360 13921 2363
rect 13780 2332 13921 2360
rect 13780 2320 13786 2332
rect 13909 2329 13921 2332
rect 13955 2329 13967 2363
rect 15194 2360 15200 2372
rect 15155 2332 15200 2360
rect 13909 2323 13967 2329
rect 15194 2320 15200 2332
rect 15252 2320 15258 2372
rect 16301 2363 16359 2369
rect 16301 2329 16313 2363
rect 16347 2360 16359 2363
rect 17126 2360 17132 2372
rect 16347 2332 17132 2360
rect 16347 2329 16359 2332
rect 16301 2323 16359 2329
rect 17126 2320 17132 2332
rect 17184 2320 17190 2372
rect 17310 2320 17316 2372
rect 17368 2360 17374 2372
rect 17405 2363 17463 2369
rect 17405 2360 17417 2363
rect 17368 2332 17417 2360
rect 17368 2320 17374 2332
rect 17405 2329 17417 2332
rect 17451 2329 17463 2363
rect 17405 2323 17463 2329
rect 17770 2320 17776 2372
rect 17828 2360 17834 2372
rect 17957 2363 18015 2369
rect 17957 2360 17969 2363
rect 17828 2332 17969 2360
rect 17828 2320 17834 2332
rect 17957 2329 17969 2332
rect 18003 2329 18015 2363
rect 17957 2323 18015 2329
rect 18322 2320 18328 2372
rect 18380 2320 18386 2372
rect 18969 2363 19027 2369
rect 18969 2329 18981 2363
rect 19015 2360 19027 2363
rect 22278 2360 22284 2372
rect 19015 2332 22284 2360
rect 19015 2329 19027 2332
rect 18969 2323 19027 2329
rect 22278 2320 22284 2332
rect 22336 2320 22342 2372
rect 12483 2264 13216 2292
rect 12483 2261 12495 2264
rect 12437 2255 12495 2261
rect 13446 2252 13452 2304
rect 13504 2292 13510 2304
rect 14553 2295 14611 2301
rect 14553 2292 14565 2295
rect 13504 2264 14565 2292
rect 13504 2252 13510 2264
rect 14553 2261 14565 2264
rect 14599 2261 14611 2295
rect 14553 2255 14611 2261
rect 16761 2295 16819 2301
rect 16761 2261 16773 2295
rect 16807 2292 16819 2295
rect 18138 2292 18144 2304
rect 16807 2264 18144 2292
rect 16807 2261 16819 2264
rect 16761 2255 16819 2261
rect 18138 2252 18144 2264
rect 18196 2252 18202 2304
rect 18340 2292 18368 2320
rect 20530 2292 20536 2304
rect 18340 2264 20536 2292
rect 20530 2252 20536 2264
rect 20588 2252 20594 2304
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
rect 8294 2048 8300 2100
rect 8352 2088 8358 2100
rect 8570 2088 8576 2100
rect 8352 2060 8576 2088
rect 8352 2048 8358 2060
rect 8570 2048 8576 2060
rect 8628 2088 8634 2100
rect 13446 2088 13452 2100
rect 8628 2060 13452 2088
rect 8628 2048 8634 2060
rect 13446 2048 13452 2060
rect 13504 2048 13510 2100
rect 15010 2048 15016 2100
rect 15068 2088 15074 2100
rect 18782 2088 18788 2100
rect 15068 2060 18788 2088
rect 15068 2048 15074 2060
rect 18782 2048 18788 2060
rect 18840 2048 18846 2100
rect 566 1980 572 2032
rect 624 2020 630 2032
rect 2222 2020 2228 2032
rect 624 1992 2228 2020
rect 624 1980 630 1992
rect 2222 1980 2228 1992
rect 2280 2020 2286 2032
rect 9214 2020 9220 2032
rect 2280 1992 9220 2020
rect 2280 1980 2286 1992
rect 9214 1980 9220 1992
rect 9272 1980 9278 2032
rect 16666 1980 16672 2032
rect 16724 2020 16730 2032
rect 19150 2020 19156 2032
rect 16724 1992 19156 2020
rect 16724 1980 16730 1992
rect 19150 1980 19156 1992
rect 19208 1980 19214 2032
rect 1026 1912 1032 1964
rect 1084 1952 1090 1964
rect 2682 1952 2688 1964
rect 1084 1924 2688 1952
rect 1084 1912 1090 1924
rect 2682 1912 2688 1924
rect 2740 1912 2746 1964
rect 13538 1912 13544 1964
rect 13596 1952 13602 1964
rect 17954 1952 17960 1964
rect 13596 1924 17960 1952
rect 13596 1912 13602 1924
rect 17954 1912 17960 1924
rect 18012 1912 18018 1964
rect 2406 1844 2412 1896
rect 2464 1884 2470 1896
rect 5718 1884 5724 1896
rect 2464 1856 5724 1884
rect 2464 1844 2470 1856
rect 5718 1844 5724 1856
rect 5776 1844 5782 1896
rect 12986 1844 12992 1896
rect 13044 1884 13050 1896
rect 18046 1884 18052 1896
rect 13044 1856 18052 1884
rect 13044 1844 13050 1856
rect 18046 1844 18052 1856
rect 18104 1844 18110 1896
rect 4246 1776 4252 1828
rect 4304 1816 4310 1828
rect 7374 1816 7380 1828
rect 4304 1788 7380 1816
rect 4304 1776 4310 1788
rect 7374 1776 7380 1788
rect 7432 1776 7438 1828
rect 9214 1776 9220 1828
rect 9272 1816 9278 1828
rect 10686 1816 10692 1828
rect 9272 1788 10692 1816
rect 9272 1776 9278 1788
rect 10686 1776 10692 1788
rect 10744 1776 10750 1828
rect 3326 1572 3332 1624
rect 3384 1612 3390 1624
rect 4338 1612 4344 1624
rect 3384 1584 4344 1612
rect 3384 1572 3390 1584
rect 4338 1572 4344 1584
rect 4396 1572 4402 1624
rect 3326 1436 3332 1488
rect 3384 1476 3390 1488
rect 3878 1476 3884 1488
rect 3384 1448 3884 1476
rect 3384 1436 3390 1448
rect 3878 1436 3884 1448
rect 3936 1436 3942 1488
rect 8754 1436 8760 1488
rect 8812 1476 8818 1488
rect 9490 1476 9496 1488
rect 8812 1448 9496 1476
rect 8812 1436 8818 1448
rect 9490 1436 9496 1448
rect 9548 1436 9554 1488
rect 15194 1436 15200 1488
rect 15252 1476 15258 1488
rect 21358 1476 21364 1488
rect 15252 1448 21364 1476
rect 15252 1436 15258 1448
rect 21358 1436 21364 1448
rect 21416 1436 21422 1488
rect 12618 1368 12624 1420
rect 12676 1408 12682 1420
rect 15010 1408 15016 1420
rect 12676 1380 15016 1408
rect 12676 1368 12682 1380
rect 15010 1368 15016 1380
rect 15068 1368 15074 1420
rect 17126 1368 17132 1420
rect 17184 1408 17190 1420
rect 18598 1408 18604 1420
rect 17184 1380 18604 1408
rect 17184 1368 17190 1380
rect 18598 1368 18604 1380
rect 18656 1368 18662 1420
rect 15562 1300 15568 1352
rect 15620 1340 15626 1352
rect 18782 1340 18788 1352
rect 15620 1312 18788 1340
rect 15620 1300 15626 1312
rect 18782 1300 18788 1312
rect 18840 1300 18846 1352
rect 2866 1164 2872 1216
rect 2924 1204 2930 1216
rect 4062 1204 4068 1216
rect 2924 1176 4068 1204
rect 2924 1164 2930 1176
rect 4062 1164 4068 1176
rect 4120 1164 4126 1216
<< via1 >>
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 2228 20587 2280 20596
rect 2228 20553 2237 20587
rect 2237 20553 2271 20587
rect 2271 20553 2280 20587
rect 2228 20544 2280 20553
rect 2780 20476 2832 20528
rect 3240 20519 3292 20528
rect 3240 20485 3249 20519
rect 3249 20485 3283 20519
rect 3283 20485 3292 20519
rect 3240 20476 3292 20485
rect 4068 20519 4120 20528
rect 4068 20485 4077 20519
rect 4077 20485 4111 20519
rect 4111 20485 4120 20519
rect 4068 20476 4120 20485
rect 17224 20476 17276 20528
rect 18604 20476 18656 20528
rect 18972 20519 19024 20528
rect 18972 20485 18981 20519
rect 18981 20485 19015 20519
rect 19015 20485 19024 20519
rect 18972 20476 19024 20485
rect 19524 20519 19576 20528
rect 19524 20485 19533 20519
rect 19533 20485 19567 20519
rect 19567 20485 19576 20519
rect 19524 20476 19576 20485
rect 1584 20383 1636 20392
rect 1584 20349 1593 20383
rect 1593 20349 1627 20383
rect 1627 20349 1636 20383
rect 1584 20340 1636 20349
rect 2596 20340 2648 20392
rect 4160 20340 4212 20392
rect 5724 20383 5776 20392
rect 5724 20349 5733 20383
rect 5733 20349 5767 20383
rect 5767 20349 5776 20383
rect 5724 20340 5776 20349
rect 19708 20340 19760 20392
rect 20260 20383 20312 20392
rect 20260 20349 20269 20383
rect 20269 20349 20303 20383
rect 20303 20349 20312 20383
rect 20260 20340 20312 20349
rect 2320 20315 2372 20324
rect 2320 20281 2329 20315
rect 2329 20281 2363 20315
rect 2363 20281 2372 20315
rect 2320 20272 2372 20281
rect 2872 20315 2924 20324
rect 2872 20281 2881 20315
rect 2881 20281 2915 20315
rect 2915 20281 2924 20315
rect 2872 20272 2924 20281
rect 2964 20272 3016 20324
rect 4252 20315 4304 20324
rect 4252 20281 4261 20315
rect 4261 20281 4295 20315
rect 4295 20281 4304 20315
rect 4252 20272 4304 20281
rect 9680 20272 9732 20324
rect 18788 20315 18840 20324
rect 18788 20281 18797 20315
rect 18797 20281 18831 20315
rect 18831 20281 18840 20315
rect 18788 20272 18840 20281
rect 19340 20315 19392 20324
rect 19340 20281 19349 20315
rect 19349 20281 19383 20315
rect 19383 20281 19392 20315
rect 19340 20272 19392 20281
rect 20628 20315 20680 20324
rect 20628 20281 20637 20315
rect 20637 20281 20671 20315
rect 20671 20281 20680 20315
rect 20628 20272 20680 20281
rect 20812 20315 20864 20324
rect 20812 20281 20821 20315
rect 20821 20281 20855 20315
rect 20855 20281 20864 20315
rect 20812 20272 20864 20281
rect 4988 20204 5040 20256
rect 5908 20247 5960 20256
rect 5908 20213 5917 20247
rect 5917 20213 5951 20247
rect 5951 20213 5960 20247
rect 5908 20204 5960 20213
rect 8208 20204 8260 20256
rect 19524 20204 19576 20256
rect 20260 20204 20312 20256
rect 21456 20272 21508 20324
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 2320 20043 2372 20052
rect 2320 20009 2329 20043
rect 2329 20009 2363 20043
rect 2363 20009 2372 20043
rect 2320 20000 2372 20009
rect 2964 20043 3016 20052
rect 2964 20009 2973 20043
rect 2973 20009 3007 20043
rect 3007 20009 3016 20043
rect 2964 20000 3016 20009
rect 4252 20000 4304 20052
rect 8208 20000 8260 20052
rect 18788 20000 18840 20052
rect 20536 20000 20588 20052
rect 1768 19907 1820 19916
rect 1768 19873 1777 19907
rect 1777 19873 1811 19907
rect 1811 19873 1820 19907
rect 1768 19864 1820 19873
rect 5080 19932 5132 19984
rect 5908 19932 5960 19984
rect 20168 19932 20220 19984
rect 3056 19796 3108 19848
rect 1584 19771 1636 19780
rect 1584 19737 1593 19771
rect 1593 19737 1627 19771
rect 1627 19737 1636 19771
rect 1584 19728 1636 19737
rect 4160 19864 4212 19916
rect 4344 19907 4396 19916
rect 4344 19873 4378 19907
rect 4378 19873 4396 19907
rect 4344 19864 4396 19873
rect 17960 19864 18012 19916
rect 20352 19864 20404 19916
rect 21180 19907 21232 19916
rect 21180 19873 21189 19907
rect 21189 19873 21223 19907
rect 21223 19873 21232 19907
rect 21180 19864 21232 19873
rect 7656 19796 7708 19848
rect 10324 19839 10376 19848
rect 7840 19728 7892 19780
rect 10324 19805 10333 19839
rect 10333 19805 10367 19839
rect 10367 19805 10376 19839
rect 10324 19796 10376 19805
rect 21364 19771 21416 19780
rect 21364 19737 21373 19771
rect 21373 19737 21407 19771
rect 21407 19737 21416 19771
rect 21364 19728 21416 19737
rect 5264 19660 5316 19712
rect 7748 19703 7800 19712
rect 7748 19669 7757 19703
rect 7757 19669 7791 19703
rect 7791 19669 7800 19703
rect 7748 19660 7800 19669
rect 8208 19660 8260 19712
rect 11704 19703 11756 19712
rect 11704 19669 11713 19703
rect 11713 19669 11747 19703
rect 11747 19669 11756 19703
rect 11704 19660 11756 19669
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 1768 19456 1820 19508
rect 2596 19499 2648 19508
rect 2596 19465 2605 19499
rect 2605 19465 2639 19499
rect 2639 19465 2648 19499
rect 2596 19456 2648 19465
rect 4160 19456 4212 19508
rect 9680 19499 9732 19508
rect 1584 19295 1636 19304
rect 1584 19261 1593 19295
rect 1593 19261 1627 19295
rect 1627 19261 1636 19295
rect 1584 19252 1636 19261
rect 1768 19227 1820 19236
rect 1768 19193 1777 19227
rect 1777 19193 1811 19227
rect 1811 19193 1820 19227
rect 1768 19184 1820 19193
rect 3884 19252 3936 19304
rect 9680 19465 9689 19499
rect 9689 19465 9723 19499
rect 9723 19465 9732 19499
rect 9680 19456 9732 19465
rect 19340 19456 19392 19508
rect 20628 19499 20680 19508
rect 20628 19465 20637 19499
rect 20637 19465 20671 19499
rect 20671 19465 20680 19499
rect 20628 19456 20680 19465
rect 20352 19388 20404 19440
rect 4252 19184 4304 19236
rect 4528 19252 4580 19304
rect 5080 19295 5132 19304
rect 5080 19261 5089 19295
rect 5089 19261 5123 19295
rect 5123 19261 5132 19295
rect 5080 19252 5132 19261
rect 7748 19252 7800 19304
rect 9496 19252 9548 19304
rect 10324 19252 10376 19304
rect 13360 19252 13412 19304
rect 4344 19116 4396 19168
rect 5816 19116 5868 19168
rect 7288 19159 7340 19168
rect 7288 19125 7297 19159
rect 7297 19125 7331 19159
rect 7331 19125 7340 19159
rect 7288 19116 7340 19125
rect 7472 19116 7524 19168
rect 8208 19184 8260 19236
rect 13452 19184 13504 19236
rect 10140 19116 10192 19168
rect 14556 19116 14608 19168
rect 18052 19116 18104 19168
rect 18604 19227 18656 19236
rect 18604 19193 18613 19227
rect 18613 19193 18647 19227
rect 18647 19193 18656 19227
rect 19984 19252 20036 19304
rect 18604 19184 18656 19193
rect 19340 19116 19392 19168
rect 19708 19159 19760 19168
rect 19708 19125 19717 19159
rect 19717 19125 19751 19159
rect 19751 19125 19760 19159
rect 19708 19116 19760 19125
rect 20444 19184 20496 19236
rect 21364 19227 21416 19236
rect 21364 19193 21373 19227
rect 21373 19193 21407 19227
rect 21407 19193 21416 19227
rect 21364 19184 21416 19193
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 1768 18912 1820 18964
rect 2872 18912 2924 18964
rect 3056 18955 3108 18964
rect 3056 18921 3065 18955
rect 3065 18921 3099 18955
rect 3099 18921 3108 18955
rect 3056 18912 3108 18921
rect 1584 18819 1636 18828
rect 1584 18785 1593 18819
rect 1593 18785 1627 18819
rect 1627 18785 1636 18819
rect 1584 18776 1636 18785
rect 1768 18819 1820 18828
rect 1768 18785 1777 18819
rect 1777 18785 1811 18819
rect 1811 18785 1820 18819
rect 1768 18776 1820 18785
rect 6552 18912 6604 18964
rect 19984 18912 20036 18964
rect 20260 18912 20312 18964
rect 21180 18912 21232 18964
rect 7288 18844 7340 18896
rect 11704 18844 11756 18896
rect 14004 18844 14056 18896
rect 4160 18776 4212 18828
rect 5080 18776 5132 18828
rect 5264 18819 5316 18828
rect 5264 18785 5298 18819
rect 5298 18785 5316 18819
rect 5264 18776 5316 18785
rect 9036 18776 9088 18828
rect 12624 18776 12676 18828
rect 14556 18776 14608 18828
rect 21180 18819 21232 18828
rect 4528 18708 4580 18760
rect 3976 18615 4028 18624
rect 3976 18581 3985 18615
rect 3985 18581 4019 18615
rect 4019 18581 4028 18615
rect 3976 18572 4028 18581
rect 5356 18572 5408 18624
rect 13360 18708 13412 18760
rect 20536 18708 20588 18760
rect 21180 18785 21189 18819
rect 21189 18785 21223 18819
rect 21223 18785 21232 18819
rect 21180 18776 21232 18785
rect 21364 18683 21416 18692
rect 21364 18649 21373 18683
rect 21373 18649 21407 18683
rect 21407 18649 21416 18683
rect 21364 18640 21416 18649
rect 7564 18572 7616 18624
rect 8208 18572 8260 18624
rect 13360 18615 13412 18624
rect 13360 18581 13369 18615
rect 13369 18581 13403 18615
rect 13403 18581 13412 18615
rect 13360 18572 13412 18581
rect 15936 18572 15988 18624
rect 18696 18615 18748 18624
rect 18696 18581 18705 18615
rect 18705 18581 18739 18615
rect 18739 18581 18748 18615
rect 18696 18572 18748 18581
rect 19800 18615 19852 18624
rect 19800 18581 19809 18615
rect 19809 18581 19843 18615
rect 19843 18581 19852 18615
rect 19800 18572 19852 18581
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 2228 18411 2280 18420
rect 2228 18377 2237 18411
rect 2237 18377 2271 18411
rect 2271 18377 2280 18411
rect 2228 18368 2280 18377
rect 3976 18368 4028 18420
rect 7472 18411 7524 18420
rect 1768 18300 1820 18352
rect 4344 18300 4396 18352
rect 4896 18300 4948 18352
rect 7472 18377 7481 18411
rect 7481 18377 7515 18411
rect 7515 18377 7524 18411
rect 7472 18368 7524 18377
rect 10876 18368 10928 18420
rect 20444 18368 20496 18420
rect 21180 18368 21232 18420
rect 10692 18300 10744 18352
rect 18880 18300 18932 18352
rect 5264 18232 5316 18284
rect 8208 18232 8260 18284
rect 9036 18275 9088 18284
rect 9036 18241 9045 18275
rect 9045 18241 9079 18275
rect 9079 18241 9088 18275
rect 9036 18232 9088 18241
rect 9588 18232 9640 18284
rect 12348 18232 12400 18284
rect 14556 18275 14608 18284
rect 14556 18241 14565 18275
rect 14565 18241 14599 18275
rect 14599 18241 14608 18275
rect 14556 18232 14608 18241
rect 17684 18275 17736 18284
rect 17684 18241 17693 18275
rect 17693 18241 17727 18275
rect 17727 18241 17736 18275
rect 17684 18232 17736 18241
rect 6828 18164 6880 18216
rect 19432 18164 19484 18216
rect 1768 18139 1820 18148
rect 1768 18105 1777 18139
rect 1777 18105 1811 18139
rect 1811 18105 1820 18139
rect 1768 18096 1820 18105
rect 2320 18139 2372 18148
rect 2320 18105 2329 18139
rect 2329 18105 2363 18139
rect 2363 18105 2372 18139
rect 2320 18096 2372 18105
rect 3424 18139 3476 18148
rect 3424 18105 3433 18139
rect 3433 18105 3467 18139
rect 3467 18105 3476 18139
rect 3424 18096 3476 18105
rect 1676 18071 1728 18080
rect 1676 18037 1685 18071
rect 1685 18037 1719 18071
rect 1719 18037 1728 18071
rect 1676 18028 1728 18037
rect 3516 18071 3568 18080
rect 3516 18037 3525 18071
rect 3525 18037 3559 18071
rect 3559 18037 3568 18071
rect 3516 18028 3568 18037
rect 9128 18096 9180 18148
rect 11980 18096 12032 18148
rect 17500 18139 17552 18148
rect 17500 18105 17509 18139
rect 17509 18105 17543 18139
rect 17543 18105 17552 18139
rect 17500 18096 17552 18105
rect 4160 18071 4212 18080
rect 4160 18037 4169 18071
rect 4169 18037 4203 18071
rect 4203 18037 4212 18071
rect 4160 18028 4212 18037
rect 4620 18071 4672 18080
rect 4620 18037 4629 18071
rect 4629 18037 4663 18071
rect 4663 18037 4672 18071
rect 4620 18028 4672 18037
rect 5172 18071 5224 18080
rect 5172 18037 5181 18071
rect 5181 18037 5215 18071
rect 5215 18037 5224 18071
rect 5172 18028 5224 18037
rect 8852 18071 8904 18080
rect 8852 18037 8861 18071
rect 8861 18037 8895 18071
rect 8895 18037 8904 18071
rect 8852 18028 8904 18037
rect 8944 18071 8996 18080
rect 8944 18037 8953 18071
rect 8953 18037 8987 18071
rect 8987 18037 8996 18071
rect 8944 18028 8996 18037
rect 9404 18028 9456 18080
rect 11704 18028 11756 18080
rect 14648 18071 14700 18080
rect 14648 18037 14657 18071
rect 14657 18037 14691 18071
rect 14691 18037 14700 18071
rect 14648 18028 14700 18037
rect 14740 18071 14792 18080
rect 14740 18037 14749 18071
rect 14749 18037 14783 18071
rect 14783 18037 14792 18071
rect 14740 18028 14792 18037
rect 15200 18028 15252 18080
rect 15384 18071 15436 18080
rect 15384 18037 15393 18071
rect 15393 18037 15427 18071
rect 15427 18037 15436 18071
rect 15384 18028 15436 18037
rect 17592 18071 17644 18080
rect 17592 18037 17601 18071
rect 17601 18037 17635 18071
rect 17635 18037 17644 18071
rect 18972 18071 19024 18080
rect 17592 18028 17644 18037
rect 18972 18037 18981 18071
rect 18981 18037 19015 18071
rect 19015 18037 19024 18071
rect 18972 18028 19024 18037
rect 20444 18164 20496 18216
rect 20260 18096 20312 18148
rect 21364 18139 21416 18148
rect 21364 18105 21373 18139
rect 21373 18105 21407 18139
rect 21407 18105 21416 18139
rect 21364 18096 21416 18105
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 2320 17824 2372 17876
rect 3516 17867 3568 17876
rect 3516 17833 3525 17867
rect 3525 17833 3559 17867
rect 3559 17833 3568 17867
rect 3516 17824 3568 17833
rect 4620 17824 4672 17876
rect 6828 17824 6880 17876
rect 9404 17824 9456 17876
rect 10324 17824 10376 17876
rect 10600 17824 10652 17876
rect 14740 17824 14792 17876
rect 15384 17824 15436 17876
rect 5172 17756 5224 17808
rect 6000 17756 6052 17808
rect 6552 17756 6604 17808
rect 11060 17756 11112 17808
rect 2596 17620 2648 17672
rect 1676 17527 1728 17536
rect 1676 17493 1685 17527
rect 1685 17493 1719 17527
rect 1719 17493 1728 17527
rect 1676 17484 1728 17493
rect 4068 17688 4120 17740
rect 4344 17688 4396 17740
rect 6920 17688 6972 17740
rect 8300 17688 8352 17740
rect 9404 17688 9456 17740
rect 11244 17731 11296 17740
rect 11244 17697 11278 17731
rect 11278 17697 11296 17731
rect 11244 17688 11296 17697
rect 15476 17756 15528 17808
rect 15568 17756 15620 17808
rect 17684 17824 17736 17876
rect 19984 17824 20036 17876
rect 20260 17867 20312 17876
rect 20260 17833 20269 17867
rect 20269 17833 20303 17867
rect 20303 17833 20312 17867
rect 20260 17824 20312 17833
rect 13728 17688 13780 17740
rect 15108 17688 15160 17740
rect 15200 17688 15252 17740
rect 16488 17688 16540 17740
rect 17960 17688 18012 17740
rect 18144 17688 18196 17740
rect 2964 17663 3016 17672
rect 2964 17629 2973 17663
rect 2973 17629 3007 17663
rect 3007 17629 3016 17663
rect 2964 17620 3016 17629
rect 4804 17663 4856 17672
rect 4804 17629 4813 17663
rect 4813 17629 4847 17663
rect 4847 17629 4856 17663
rect 4804 17620 4856 17629
rect 4896 17663 4948 17672
rect 4896 17629 4905 17663
rect 4905 17629 4939 17663
rect 4939 17629 4948 17663
rect 4896 17620 4948 17629
rect 5356 17620 5408 17672
rect 8944 17552 8996 17604
rect 7012 17527 7064 17536
rect 7012 17493 7021 17527
rect 7021 17493 7055 17527
rect 7055 17493 7064 17527
rect 7012 17484 7064 17493
rect 8852 17484 8904 17536
rect 12072 17620 12124 17672
rect 13360 17663 13412 17672
rect 13360 17629 13369 17663
rect 13369 17629 13403 17663
rect 13403 17629 13412 17663
rect 13360 17620 13412 17629
rect 13544 17620 13596 17672
rect 15476 17663 15528 17672
rect 15476 17629 15485 17663
rect 15485 17629 15519 17663
rect 15519 17629 15528 17663
rect 15476 17620 15528 17629
rect 15936 17663 15988 17672
rect 15936 17629 15945 17663
rect 15945 17629 15979 17663
rect 15979 17629 15988 17663
rect 15936 17620 15988 17629
rect 16120 17663 16172 17672
rect 16120 17629 16129 17663
rect 16129 17629 16163 17663
rect 16163 17629 16172 17663
rect 16120 17620 16172 17629
rect 18788 17663 18840 17672
rect 18788 17629 18797 17663
rect 18797 17629 18831 17663
rect 18831 17629 18840 17663
rect 18788 17620 18840 17629
rect 18972 17620 19024 17672
rect 20352 17688 20404 17740
rect 21180 17731 21232 17740
rect 21180 17697 21189 17731
rect 21189 17697 21223 17731
rect 21223 17697 21232 17731
rect 21180 17688 21232 17697
rect 9496 17484 9548 17536
rect 10508 17484 10560 17536
rect 11244 17484 11296 17536
rect 12164 17484 12216 17536
rect 12348 17527 12400 17536
rect 12348 17493 12357 17527
rect 12357 17493 12391 17527
rect 12391 17493 12400 17527
rect 12348 17484 12400 17493
rect 13912 17527 13964 17536
rect 13912 17493 13921 17527
rect 13921 17493 13955 17527
rect 13955 17493 13964 17527
rect 13912 17484 13964 17493
rect 14096 17484 14148 17536
rect 19800 17552 19852 17604
rect 20812 17595 20864 17604
rect 20812 17561 20821 17595
rect 20821 17561 20855 17595
rect 20855 17561 20864 17595
rect 20812 17552 20864 17561
rect 21364 17595 21416 17604
rect 21364 17561 21373 17595
rect 21373 17561 21407 17595
rect 21407 17561 21416 17595
rect 21364 17552 21416 17561
rect 19708 17527 19760 17536
rect 19708 17493 19717 17527
rect 19717 17493 19751 17527
rect 19751 17493 19760 17527
rect 19708 17484 19760 17493
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 1768 17280 1820 17332
rect 3424 17280 3476 17332
rect 4804 17280 4856 17332
rect 6920 17323 6972 17332
rect 6920 17289 6929 17323
rect 6929 17289 6963 17323
rect 6963 17289 6972 17323
rect 6920 17280 6972 17289
rect 9128 17323 9180 17332
rect 9128 17289 9137 17323
rect 9137 17289 9171 17323
rect 9171 17289 9180 17323
rect 9128 17280 9180 17289
rect 2964 17212 3016 17264
rect 4252 17212 4304 17264
rect 4068 17187 4120 17196
rect 4068 17153 4077 17187
rect 4077 17153 4111 17187
rect 4111 17153 4120 17187
rect 4068 17144 4120 17153
rect 8852 17212 8904 17264
rect 11244 17280 11296 17332
rect 11704 17280 11756 17332
rect 13544 17280 13596 17332
rect 15660 17280 15712 17332
rect 17500 17280 17552 17332
rect 17592 17280 17644 17332
rect 18144 17323 18196 17332
rect 18144 17289 18153 17323
rect 18153 17289 18187 17323
rect 18187 17289 18196 17323
rect 18144 17280 18196 17289
rect 20352 17323 20404 17332
rect 20352 17289 20361 17323
rect 20361 17289 20395 17323
rect 20395 17289 20404 17323
rect 20352 17280 20404 17289
rect 21180 17280 21232 17332
rect 10508 17212 10560 17264
rect 7012 17144 7064 17196
rect 9588 17144 9640 17196
rect 12716 17212 12768 17264
rect 14004 17212 14056 17264
rect 10876 17187 10928 17196
rect 10876 17153 10885 17187
rect 10885 17153 10919 17187
rect 10919 17153 10928 17187
rect 10876 17144 10928 17153
rect 11428 17144 11480 17196
rect 12072 17187 12124 17196
rect 12072 17153 12081 17187
rect 12081 17153 12115 17187
rect 12115 17153 12124 17187
rect 12072 17144 12124 17153
rect 12256 17144 12308 17196
rect 13728 17144 13780 17196
rect 15476 17144 15528 17196
rect 1584 17119 1636 17128
rect 1584 17085 1593 17119
rect 1593 17085 1627 17119
rect 1627 17085 1636 17119
rect 1584 17076 1636 17085
rect 2320 17119 2372 17128
rect 2320 17085 2329 17119
rect 2329 17085 2363 17119
rect 2363 17085 2372 17119
rect 2320 17076 2372 17085
rect 2044 17008 2096 17060
rect 1860 16940 1912 16992
rect 4988 17076 5040 17128
rect 2872 17008 2924 17060
rect 10508 17076 10560 17128
rect 5908 17008 5960 17060
rect 9220 17008 9272 17060
rect 12992 17076 13044 17128
rect 18788 17076 18840 17128
rect 20076 17076 20128 17128
rect 20628 17119 20680 17128
rect 11244 17008 11296 17060
rect 5448 16983 5500 16992
rect 5448 16949 5457 16983
rect 5457 16949 5491 16983
rect 5491 16949 5500 16983
rect 5448 16940 5500 16949
rect 5632 16940 5684 16992
rect 7104 16940 7156 16992
rect 8392 16940 8444 16992
rect 10600 16940 10652 16992
rect 10968 16983 11020 16992
rect 10968 16949 10977 16983
rect 10977 16949 11011 16983
rect 11011 16949 11020 16983
rect 10968 16940 11020 16949
rect 17224 17008 17276 17060
rect 17316 17008 17368 17060
rect 19064 17008 19116 17060
rect 19708 17008 19760 17060
rect 20628 17085 20637 17119
rect 20637 17085 20671 17119
rect 20671 17085 20680 17119
rect 20628 17076 20680 17085
rect 20352 17008 20404 17060
rect 15384 16983 15436 16992
rect 15384 16949 15393 16983
rect 15393 16949 15427 16983
rect 15427 16949 15436 16983
rect 15384 16940 15436 16949
rect 16212 16940 16264 16992
rect 17408 16983 17460 16992
rect 17408 16949 17417 16983
rect 17417 16949 17451 16983
rect 17451 16949 17460 16983
rect 17408 16940 17460 16949
rect 19524 16940 19576 16992
rect 19800 16983 19852 16992
rect 19800 16949 19809 16983
rect 19809 16949 19843 16983
rect 19843 16949 19852 16983
rect 19800 16940 19852 16949
rect 21272 16983 21324 16992
rect 21272 16949 21281 16983
rect 21281 16949 21315 16983
rect 21315 16949 21324 16983
rect 21272 16940 21324 16949
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 2044 16736 2096 16788
rect 2320 16736 2372 16788
rect 5448 16779 5500 16788
rect 5448 16745 5457 16779
rect 5457 16745 5491 16779
rect 5491 16745 5500 16779
rect 5448 16736 5500 16745
rect 6552 16779 6604 16788
rect 6552 16745 6561 16779
rect 6561 16745 6595 16779
rect 6595 16745 6604 16779
rect 6552 16736 6604 16745
rect 2964 16668 3016 16720
rect 1584 16643 1636 16652
rect 1584 16609 1593 16643
rect 1593 16609 1627 16643
rect 1627 16609 1636 16643
rect 1584 16600 1636 16609
rect 5632 16668 5684 16720
rect 5908 16668 5960 16720
rect 10968 16736 11020 16788
rect 11980 16779 12032 16788
rect 11980 16745 11989 16779
rect 11989 16745 12023 16779
rect 12023 16745 12032 16779
rect 11980 16736 12032 16745
rect 14648 16736 14700 16788
rect 15384 16736 15436 16788
rect 16212 16779 16264 16788
rect 16212 16745 16221 16779
rect 16221 16745 16255 16779
rect 16255 16745 16264 16779
rect 16212 16736 16264 16745
rect 16764 16736 16816 16788
rect 17224 16779 17276 16788
rect 17224 16745 17233 16779
rect 17233 16745 17267 16779
rect 17267 16745 17276 16779
rect 17224 16736 17276 16745
rect 20260 16736 20312 16788
rect 20352 16779 20404 16788
rect 20352 16745 20361 16779
rect 20361 16745 20395 16779
rect 20395 16745 20404 16779
rect 20352 16736 20404 16745
rect 21180 16736 21232 16788
rect 9128 16668 9180 16720
rect 9220 16668 9272 16720
rect 10876 16668 10928 16720
rect 4160 16600 4212 16652
rect 3516 16532 3568 16584
rect 3608 16532 3660 16584
rect 8392 16600 8444 16652
rect 9312 16600 9364 16652
rect 10416 16600 10468 16652
rect 12716 16668 12768 16720
rect 12992 16600 13044 16652
rect 13912 16668 13964 16720
rect 6000 16575 6052 16584
rect 6000 16541 6009 16575
rect 6009 16541 6043 16575
rect 6043 16541 6052 16575
rect 6000 16532 6052 16541
rect 9404 16532 9456 16584
rect 11428 16532 11480 16584
rect 2596 16507 2648 16516
rect 2596 16473 2605 16507
rect 2605 16473 2639 16507
rect 2639 16473 2648 16507
rect 2596 16464 2648 16473
rect 13360 16575 13412 16584
rect 12164 16464 12216 16516
rect 13360 16541 13369 16575
rect 13369 16541 13403 16575
rect 13403 16541 13412 16575
rect 13360 16532 13412 16541
rect 13084 16464 13136 16516
rect 14556 16532 14608 16584
rect 16120 16600 16172 16652
rect 17408 16600 17460 16652
rect 17868 16600 17920 16652
rect 18880 16600 18932 16652
rect 19984 16668 20036 16720
rect 19800 16600 19852 16652
rect 2780 16396 2832 16448
rect 5264 16396 5316 16448
rect 14004 16396 14056 16448
rect 17316 16532 17368 16584
rect 19892 16532 19944 16584
rect 21364 16643 21416 16652
rect 21364 16609 21373 16643
rect 21373 16609 21407 16643
rect 21407 16609 21416 16643
rect 21364 16600 21416 16609
rect 15476 16396 15528 16448
rect 18604 16396 18656 16448
rect 19616 16396 19668 16448
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 2964 16192 3016 16244
rect 3516 16235 3568 16244
rect 3516 16201 3525 16235
rect 3525 16201 3559 16235
rect 3559 16201 3568 16235
rect 3516 16192 3568 16201
rect 1584 16099 1636 16108
rect 1584 16065 1593 16099
rect 1593 16065 1627 16099
rect 1627 16065 1636 16099
rect 1584 16056 1636 16065
rect 6000 16192 6052 16244
rect 7656 16192 7708 16244
rect 7288 16124 7340 16176
rect 2780 16031 2832 16040
rect 2780 15997 2789 16031
rect 2789 15997 2823 16031
rect 2823 15997 2832 16031
rect 2780 15988 2832 15997
rect 3608 15988 3660 16040
rect 4344 16031 4396 16040
rect 4344 15997 4353 16031
rect 4353 15997 4387 16031
rect 4387 15997 4396 16031
rect 4344 15988 4396 15997
rect 9588 16192 9640 16244
rect 13084 16192 13136 16244
rect 19616 16192 19668 16244
rect 19892 16235 19944 16244
rect 19892 16201 19901 16235
rect 19901 16201 19935 16235
rect 19935 16201 19944 16235
rect 19892 16192 19944 16201
rect 20628 16124 20680 16176
rect 11060 16056 11112 16108
rect 17040 16056 17092 16108
rect 18604 16056 18656 16108
rect 5724 15988 5776 16040
rect 6276 15988 6328 16040
rect 15292 15988 15344 16040
rect 2320 15852 2372 15904
rect 3792 15920 3844 15972
rect 4252 15920 4304 15972
rect 9496 15920 9548 15972
rect 9864 15920 9916 15972
rect 20260 15988 20312 16040
rect 11060 15852 11112 15904
rect 12256 15852 12308 15904
rect 13084 15895 13136 15904
rect 13084 15861 13093 15895
rect 13093 15861 13127 15895
rect 13127 15861 13136 15895
rect 13084 15852 13136 15861
rect 16764 15852 16816 15904
rect 17316 15852 17368 15904
rect 18604 15895 18656 15904
rect 18604 15861 18613 15895
rect 18613 15861 18647 15895
rect 18647 15861 18656 15895
rect 18604 15852 18656 15861
rect 18696 15852 18748 15904
rect 20352 15895 20404 15904
rect 20352 15861 20361 15895
rect 20361 15861 20395 15895
rect 20395 15861 20404 15895
rect 20352 15852 20404 15861
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 1860 15580 1912 15632
rect 2136 15623 2188 15632
rect 2136 15589 2145 15623
rect 2145 15589 2179 15623
rect 2179 15589 2188 15623
rect 2136 15580 2188 15589
rect 2320 15623 2372 15632
rect 2320 15589 2329 15623
rect 2329 15589 2363 15623
rect 2363 15589 2372 15623
rect 2320 15580 2372 15589
rect 4252 15648 4304 15700
rect 15292 15691 15344 15700
rect 15292 15657 15301 15691
rect 15301 15657 15335 15691
rect 15335 15657 15344 15691
rect 15292 15648 15344 15657
rect 4344 15580 4396 15632
rect 5356 15580 5408 15632
rect 12348 15623 12400 15632
rect 3056 15555 3108 15564
rect 3056 15521 3065 15555
rect 3065 15521 3099 15555
rect 3099 15521 3108 15555
rect 3056 15512 3108 15521
rect 5172 15555 5224 15564
rect 5172 15521 5190 15555
rect 5190 15521 5224 15555
rect 5172 15512 5224 15521
rect 12348 15589 12366 15623
rect 12366 15589 12400 15623
rect 12348 15580 12400 15589
rect 15936 15580 15988 15632
rect 20352 15580 20404 15632
rect 7288 15512 7340 15564
rect 8484 15512 8536 15564
rect 12624 15555 12676 15564
rect 12624 15521 12633 15555
rect 12633 15521 12667 15555
rect 12667 15521 12676 15555
rect 12624 15512 12676 15521
rect 14924 15555 14976 15564
rect 14924 15521 14933 15555
rect 14933 15521 14967 15555
rect 14967 15521 14976 15555
rect 14924 15512 14976 15521
rect 17960 15555 18012 15564
rect 17960 15521 17994 15555
rect 17994 15521 18012 15555
rect 17960 15512 18012 15521
rect 19616 15512 19668 15564
rect 20812 15555 20864 15564
rect 20812 15521 20821 15555
rect 20821 15521 20855 15555
rect 20855 15521 20864 15555
rect 20812 15512 20864 15521
rect 4068 15444 4120 15496
rect 5448 15487 5500 15496
rect 5448 15453 5457 15487
rect 5457 15453 5491 15487
rect 5491 15453 5500 15487
rect 5448 15444 5500 15453
rect 8392 15444 8444 15496
rect 14556 15444 14608 15496
rect 14740 15444 14792 15496
rect 15568 15487 15620 15496
rect 15568 15453 15577 15487
rect 15577 15453 15611 15487
rect 15611 15453 15620 15487
rect 15568 15444 15620 15453
rect 17132 15444 17184 15496
rect 1676 15351 1728 15360
rect 1676 15317 1685 15351
rect 1685 15317 1719 15351
rect 1719 15317 1728 15351
rect 1676 15308 1728 15317
rect 4252 15308 4304 15360
rect 6552 15351 6604 15360
rect 6552 15317 6561 15351
rect 6561 15317 6595 15351
rect 6595 15317 6604 15351
rect 6552 15308 6604 15317
rect 9496 15351 9548 15360
rect 9496 15317 9505 15351
rect 9505 15317 9539 15351
rect 9539 15317 9548 15351
rect 9496 15308 9548 15317
rect 11888 15308 11940 15360
rect 17592 15308 17644 15360
rect 19064 15351 19116 15360
rect 19064 15317 19073 15351
rect 19073 15317 19107 15351
rect 19107 15317 19116 15351
rect 19064 15308 19116 15317
rect 19340 15308 19392 15360
rect 19616 15351 19668 15360
rect 19616 15317 19625 15351
rect 19625 15317 19659 15351
rect 19659 15317 19668 15351
rect 19616 15308 19668 15317
rect 21272 15351 21324 15360
rect 21272 15317 21281 15351
rect 21281 15317 21315 15351
rect 21315 15317 21324 15351
rect 21272 15308 21324 15317
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 22008 15215 22060 15224
rect 22008 15181 22017 15215
rect 22017 15181 22051 15215
rect 22051 15181 22060 15215
rect 22008 15172 22060 15181
rect 4160 15147 4212 15156
rect 4160 15113 4169 15147
rect 4169 15113 4203 15147
rect 4203 15113 4212 15147
rect 4160 15104 4212 15113
rect 7104 15104 7156 15156
rect 8208 15104 8260 15156
rect 9864 15104 9916 15156
rect 12256 15104 12308 15156
rect 9680 15079 9732 15088
rect 9680 15045 9689 15079
rect 9689 15045 9723 15079
rect 9723 15045 9732 15079
rect 14924 15104 14976 15156
rect 19708 15104 19760 15156
rect 9680 15036 9732 15045
rect 4344 14968 4396 15020
rect 12624 14968 12676 15020
rect 6552 14900 6604 14952
rect 2596 14832 2648 14884
rect 3700 14832 3752 14884
rect 7564 14832 7616 14884
rect 8392 14900 8444 14952
rect 9496 14900 9548 14952
rect 11244 14900 11296 14952
rect 10692 14832 10744 14884
rect 13176 14900 13228 14952
rect 17960 15011 18012 15020
rect 17960 14977 17969 15011
rect 17969 14977 18003 15011
rect 18003 14977 18012 15011
rect 17960 14968 18012 14977
rect 19064 15036 19116 15088
rect 19248 14968 19300 15020
rect 13636 14832 13688 14884
rect 15292 14832 15344 14884
rect 1676 14807 1728 14816
rect 1676 14773 1685 14807
rect 1685 14773 1719 14807
rect 1719 14773 1728 14807
rect 1676 14764 1728 14773
rect 2504 14764 2556 14816
rect 6460 14764 6512 14816
rect 14556 14764 14608 14816
rect 14648 14764 14700 14816
rect 15384 14764 15436 14816
rect 16580 14764 16632 14816
rect 20352 14832 20404 14884
rect 21364 14875 21416 14884
rect 21364 14841 21373 14875
rect 21373 14841 21407 14875
rect 21407 14841 21416 14875
rect 21364 14832 21416 14841
rect 19156 14807 19208 14816
rect 19156 14773 19165 14807
rect 19165 14773 19199 14807
rect 19199 14773 19208 14807
rect 19156 14764 19208 14773
rect 19708 14764 19760 14816
rect 19800 14807 19852 14816
rect 19800 14773 19809 14807
rect 19809 14773 19843 14807
rect 19843 14773 19852 14807
rect 19800 14764 19852 14773
rect 19984 14764 20036 14816
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 3056 14560 3108 14612
rect 3240 14560 3292 14612
rect 3792 14560 3844 14612
rect 4068 14603 4120 14612
rect 4068 14569 4077 14603
rect 4077 14569 4111 14603
rect 4111 14569 4120 14603
rect 4068 14560 4120 14569
rect 5724 14603 5776 14612
rect 5724 14569 5733 14603
rect 5733 14569 5767 14603
rect 5767 14569 5776 14603
rect 5724 14560 5776 14569
rect 5448 14492 5500 14544
rect 8208 14560 8260 14612
rect 9680 14492 9732 14544
rect 9864 14560 9916 14612
rect 10692 14603 10744 14612
rect 10692 14569 10701 14603
rect 10701 14569 10735 14603
rect 10735 14569 10744 14603
rect 10692 14560 10744 14569
rect 12072 14560 12124 14612
rect 13176 14603 13228 14612
rect 13176 14569 13185 14603
rect 13185 14569 13219 14603
rect 13219 14569 13228 14603
rect 13176 14560 13228 14569
rect 13636 14603 13688 14612
rect 13636 14569 13645 14603
rect 13645 14569 13679 14603
rect 13679 14569 13688 14603
rect 13636 14560 13688 14569
rect 15292 14603 15344 14612
rect 15292 14569 15301 14603
rect 15301 14569 15335 14603
rect 15335 14569 15344 14603
rect 15292 14560 15344 14569
rect 17960 14560 18012 14612
rect 19156 14560 19208 14612
rect 19708 14560 19760 14612
rect 1768 14467 1820 14476
rect 1768 14433 1777 14467
rect 1777 14433 1811 14467
rect 1811 14433 1820 14467
rect 1768 14424 1820 14433
rect 2964 14424 3016 14476
rect 4344 14424 4396 14476
rect 6092 14467 6144 14476
rect 6092 14433 6101 14467
rect 6101 14433 6135 14467
rect 6135 14433 6144 14467
rect 6092 14424 6144 14433
rect 7104 14467 7156 14476
rect 7104 14433 7113 14467
rect 7113 14433 7147 14467
rect 7147 14433 7156 14467
rect 7104 14424 7156 14433
rect 8484 14424 8536 14476
rect 9956 14424 10008 14476
rect 12624 14492 12676 14544
rect 15384 14492 15436 14544
rect 15844 14535 15896 14544
rect 15844 14501 15878 14535
rect 15878 14501 15896 14535
rect 15844 14492 15896 14501
rect 19892 14492 19944 14544
rect 11888 14424 11940 14476
rect 13820 14467 13872 14476
rect 13820 14433 13829 14467
rect 13829 14433 13863 14467
rect 13863 14433 13872 14467
rect 13820 14424 13872 14433
rect 14832 14467 14884 14476
rect 14832 14433 14841 14467
rect 14841 14433 14875 14467
rect 14875 14433 14884 14467
rect 14832 14424 14884 14433
rect 15476 14424 15528 14476
rect 2504 14399 2556 14408
rect 2504 14365 2513 14399
rect 2513 14365 2547 14399
rect 2547 14365 2556 14399
rect 2504 14356 2556 14365
rect 3976 14356 4028 14408
rect 4160 14356 4212 14408
rect 5172 14356 5224 14408
rect 6552 14356 6604 14408
rect 7196 14399 7248 14408
rect 7196 14365 7205 14399
rect 7205 14365 7239 14399
rect 7239 14365 7248 14399
rect 7196 14356 7248 14365
rect 7288 14399 7340 14408
rect 7288 14365 7297 14399
rect 7297 14365 7331 14399
rect 7331 14365 7340 14399
rect 7288 14356 7340 14365
rect 6460 14288 6512 14340
rect 1676 14263 1728 14272
rect 1676 14229 1685 14263
rect 1685 14229 1719 14263
rect 1719 14229 1728 14263
rect 1676 14220 1728 14229
rect 9496 14220 9548 14272
rect 11152 14220 11204 14272
rect 11980 14220 12032 14272
rect 15568 14399 15620 14408
rect 15568 14365 15577 14399
rect 15577 14365 15611 14399
rect 15611 14365 15620 14399
rect 15568 14356 15620 14365
rect 15384 14288 15436 14340
rect 19616 14424 19668 14476
rect 17132 14356 17184 14408
rect 18604 14356 18656 14408
rect 20812 14424 20864 14476
rect 21456 14288 21508 14340
rect 16948 14263 17000 14272
rect 16948 14229 16957 14263
rect 16957 14229 16991 14263
rect 16991 14229 17000 14263
rect 16948 14220 17000 14229
rect 17408 14220 17460 14272
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 2964 14059 3016 14068
rect 2964 14025 2973 14059
rect 2973 14025 3007 14059
rect 3007 14025 3016 14059
rect 2964 14016 3016 14025
rect 4160 14059 4212 14068
rect 4160 14025 4169 14059
rect 4169 14025 4203 14059
rect 4203 14025 4212 14059
rect 4160 14016 4212 14025
rect 7196 14016 7248 14068
rect 8300 14059 8352 14068
rect 8300 14025 8309 14059
rect 8309 14025 8343 14059
rect 8343 14025 8352 14059
rect 8300 14016 8352 14025
rect 10508 14016 10560 14068
rect 10692 14059 10744 14068
rect 10692 14025 10701 14059
rect 10701 14025 10735 14059
rect 10735 14025 10744 14059
rect 10692 14016 10744 14025
rect 14740 14016 14792 14068
rect 19984 14016 20036 14068
rect 20352 14059 20404 14068
rect 20352 14025 20361 14059
rect 20361 14025 20395 14059
rect 20395 14025 20404 14059
rect 20352 14016 20404 14025
rect 20812 14059 20864 14068
rect 20812 14025 20821 14059
rect 20821 14025 20855 14059
rect 20855 14025 20864 14059
rect 20812 14016 20864 14025
rect 1768 13948 1820 14000
rect 5172 13880 5224 13932
rect 7564 13880 7616 13932
rect 14648 13948 14700 14000
rect 9772 13880 9824 13932
rect 9864 13923 9916 13932
rect 9864 13889 9873 13923
rect 9873 13889 9907 13923
rect 9907 13889 9916 13923
rect 9864 13880 9916 13889
rect 11888 13880 11940 13932
rect 13176 13880 13228 13932
rect 14832 13880 14884 13932
rect 17960 13923 18012 13932
rect 17960 13889 17969 13923
rect 17969 13889 18003 13923
rect 18003 13889 18012 13923
rect 17960 13880 18012 13889
rect 19248 13880 19300 13932
rect 1584 13855 1636 13864
rect 1584 13821 1593 13855
rect 1593 13821 1627 13855
rect 1627 13821 1636 13855
rect 1584 13812 1636 13821
rect 3700 13812 3752 13864
rect 3884 13855 3936 13864
rect 3884 13821 3893 13855
rect 3893 13821 3927 13855
rect 3927 13821 3936 13855
rect 3884 13812 3936 13821
rect 5080 13812 5132 13864
rect 1768 13787 1820 13796
rect 1768 13753 1777 13787
rect 1777 13753 1811 13787
rect 1811 13753 1820 13787
rect 1768 13744 1820 13753
rect 7748 13812 7800 13864
rect 2504 13719 2556 13728
rect 2504 13685 2513 13719
rect 2513 13685 2547 13719
rect 2547 13685 2556 13719
rect 2504 13676 2556 13685
rect 4620 13719 4672 13728
rect 4620 13685 4629 13719
rect 4629 13685 4663 13719
rect 4663 13685 4672 13719
rect 5356 13744 5408 13796
rect 8208 13812 8260 13864
rect 11796 13812 11848 13864
rect 12256 13855 12308 13864
rect 12256 13821 12265 13855
rect 12265 13821 12299 13855
rect 12299 13821 12308 13855
rect 12256 13812 12308 13821
rect 13820 13812 13872 13864
rect 16856 13812 16908 13864
rect 18604 13812 18656 13864
rect 18880 13812 18932 13864
rect 20168 13855 20220 13864
rect 20168 13821 20177 13855
rect 20177 13821 20211 13855
rect 20211 13821 20220 13855
rect 20168 13812 20220 13821
rect 20628 13855 20680 13864
rect 20628 13821 20637 13855
rect 20637 13821 20671 13855
rect 20671 13821 20680 13855
rect 20628 13812 20680 13821
rect 21180 13855 21232 13864
rect 21180 13821 21189 13855
rect 21189 13821 21223 13855
rect 21223 13821 21232 13855
rect 21180 13812 21232 13821
rect 21364 13855 21416 13864
rect 21364 13821 21373 13855
rect 21373 13821 21407 13855
rect 21407 13821 21416 13855
rect 21364 13812 21416 13821
rect 4620 13676 4672 13685
rect 5540 13719 5592 13728
rect 5540 13685 5549 13719
rect 5549 13685 5583 13719
rect 5583 13685 5592 13719
rect 5540 13676 5592 13685
rect 7656 13676 7708 13728
rect 9036 13676 9088 13728
rect 9680 13719 9732 13728
rect 9680 13685 9689 13719
rect 9689 13685 9723 13719
rect 9723 13685 9732 13719
rect 9680 13676 9732 13685
rect 9772 13719 9824 13728
rect 9772 13685 9781 13719
rect 9781 13685 9815 13719
rect 9815 13685 9824 13719
rect 10048 13744 10100 13796
rect 9772 13676 9824 13685
rect 10508 13676 10560 13728
rect 11704 13744 11756 13796
rect 15752 13744 15804 13796
rect 18788 13744 18840 13796
rect 19800 13744 19852 13796
rect 13912 13719 13964 13728
rect 13912 13685 13921 13719
rect 13921 13685 13955 13719
rect 13955 13685 13964 13719
rect 13912 13676 13964 13685
rect 14464 13676 14516 13728
rect 15568 13676 15620 13728
rect 17132 13676 17184 13728
rect 18236 13719 18288 13728
rect 18236 13685 18245 13719
rect 18245 13685 18279 13719
rect 18279 13685 18288 13719
rect 18236 13676 18288 13685
rect 19340 13719 19392 13728
rect 19340 13685 19349 13719
rect 19349 13685 19383 13719
rect 19383 13685 19392 13719
rect 19340 13676 19392 13685
rect 19524 13676 19576 13728
rect 20260 13676 20312 13728
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 2504 13472 2556 13524
rect 3240 13472 3292 13524
rect 3516 13472 3568 13524
rect 3884 13472 3936 13524
rect 4620 13472 4672 13524
rect 5264 13515 5316 13524
rect 5264 13481 5273 13515
rect 5273 13481 5307 13515
rect 5307 13481 5316 13515
rect 5264 13472 5316 13481
rect 6092 13472 6144 13524
rect 7656 13472 7708 13524
rect 8484 13472 8536 13524
rect 9772 13472 9824 13524
rect 11704 13515 11756 13524
rect 11704 13481 11713 13515
rect 11713 13481 11747 13515
rect 11747 13481 11756 13515
rect 11704 13472 11756 13481
rect 13912 13472 13964 13524
rect 16580 13515 16632 13524
rect 16580 13481 16589 13515
rect 16589 13481 16623 13515
rect 16623 13481 16632 13515
rect 16580 13472 16632 13481
rect 17500 13472 17552 13524
rect 4160 13404 4212 13456
rect 5080 13404 5132 13456
rect 5356 13404 5408 13456
rect 2136 13336 2188 13388
rect 4252 13379 4304 13388
rect 4252 13345 4261 13379
rect 4261 13345 4295 13379
rect 4295 13345 4304 13379
rect 4252 13336 4304 13345
rect 7012 13336 7064 13388
rect 7196 13379 7248 13388
rect 7196 13345 7205 13379
rect 7205 13345 7239 13379
rect 7239 13345 7248 13379
rect 7196 13336 7248 13345
rect 6460 13311 6512 13320
rect 1584 13243 1636 13252
rect 1584 13209 1593 13243
rect 1593 13209 1627 13243
rect 1627 13209 1636 13243
rect 1584 13200 1636 13209
rect 4160 13200 4212 13252
rect 5172 13200 5224 13252
rect 6460 13277 6469 13311
rect 6469 13277 6503 13311
rect 6503 13277 6512 13311
rect 6460 13268 6512 13277
rect 7288 13311 7340 13320
rect 7288 13277 7297 13311
rect 7297 13277 7331 13311
rect 7331 13277 7340 13311
rect 7288 13268 7340 13277
rect 7564 13268 7616 13320
rect 7748 13404 7800 13456
rect 10232 13404 10284 13456
rect 10968 13404 11020 13456
rect 8576 13379 8628 13388
rect 8576 13345 8585 13379
rect 8585 13345 8619 13379
rect 8619 13345 8628 13379
rect 8576 13336 8628 13345
rect 9772 13336 9824 13388
rect 10692 13336 10744 13388
rect 10232 13268 10284 13320
rect 9956 13200 10008 13252
rect 12808 13336 12860 13388
rect 15200 13379 15252 13388
rect 15200 13345 15209 13379
rect 15209 13345 15243 13379
rect 15243 13345 15252 13379
rect 15200 13336 15252 13345
rect 3424 13175 3476 13184
rect 3424 13141 3433 13175
rect 3433 13141 3467 13175
rect 3467 13141 3476 13175
rect 3424 13132 3476 13141
rect 5540 13132 5592 13184
rect 7472 13132 7524 13184
rect 11888 13200 11940 13252
rect 12624 13268 12676 13320
rect 12440 13200 12492 13252
rect 15384 13311 15436 13320
rect 15384 13277 15393 13311
rect 15393 13277 15427 13311
rect 15427 13277 15436 13311
rect 16948 13404 17000 13456
rect 18880 13404 18932 13456
rect 16212 13379 16264 13388
rect 16212 13345 16221 13379
rect 16221 13345 16255 13379
rect 16255 13345 16264 13379
rect 16212 13336 16264 13345
rect 16304 13336 16356 13388
rect 16764 13336 16816 13388
rect 19064 13379 19116 13388
rect 15384 13268 15436 13277
rect 16396 13268 16448 13320
rect 16948 13268 17000 13320
rect 17224 13311 17276 13320
rect 17224 13277 17233 13311
rect 17233 13277 17267 13311
rect 17267 13277 17276 13311
rect 17224 13268 17276 13277
rect 19064 13345 19073 13379
rect 19073 13345 19107 13379
rect 19107 13345 19116 13379
rect 19064 13336 19116 13345
rect 19340 13472 19392 13524
rect 20260 13515 20312 13524
rect 20260 13481 20269 13515
rect 20269 13481 20303 13515
rect 20303 13481 20312 13515
rect 20260 13472 20312 13481
rect 20628 13404 20680 13456
rect 19708 13268 19760 13320
rect 10508 13132 10560 13184
rect 14280 13132 14332 13184
rect 17500 13200 17552 13252
rect 16580 13132 16632 13184
rect 18604 13132 18656 13184
rect 20168 13200 20220 13252
rect 20352 13200 20404 13252
rect 21088 13243 21140 13252
rect 21088 13209 21097 13243
rect 21097 13209 21131 13243
rect 21131 13209 21140 13243
rect 21088 13200 21140 13209
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 1768 12928 1820 12980
rect 2596 12971 2648 12980
rect 2596 12937 2605 12971
rect 2605 12937 2639 12971
rect 2639 12937 2648 12971
rect 2596 12928 2648 12937
rect 4344 12971 4396 12980
rect 4344 12937 4353 12971
rect 4353 12937 4387 12971
rect 4387 12937 4396 12971
rect 4344 12928 4396 12937
rect 5264 12928 5316 12980
rect 7104 12928 7156 12980
rect 9036 12971 9088 12980
rect 9036 12937 9045 12971
rect 9045 12937 9079 12971
rect 9079 12937 9088 12971
rect 9036 12928 9088 12937
rect 9772 12928 9824 12980
rect 10140 12928 10192 12980
rect 10508 12860 10560 12912
rect 13820 12928 13872 12980
rect 15660 12928 15712 12980
rect 16396 12971 16448 12980
rect 16396 12937 16405 12971
rect 16405 12937 16439 12971
rect 16439 12937 16448 12971
rect 16396 12928 16448 12937
rect 18144 12928 18196 12980
rect 16028 12860 16080 12912
rect 20904 12860 20956 12912
rect 20996 12860 21048 12912
rect 3424 12792 3476 12844
rect 3700 12835 3752 12844
rect 3700 12801 3709 12835
rect 3709 12801 3743 12835
rect 3743 12801 3752 12835
rect 3700 12792 3752 12801
rect 5172 12835 5224 12844
rect 5172 12801 5181 12835
rect 5181 12801 5215 12835
rect 5215 12801 5224 12835
rect 5172 12792 5224 12801
rect 5448 12792 5500 12844
rect 7564 12792 7616 12844
rect 9036 12792 9088 12844
rect 9864 12792 9916 12844
rect 10692 12792 10744 12844
rect 12716 12792 12768 12844
rect 15844 12835 15896 12844
rect 15844 12801 15853 12835
rect 15853 12801 15887 12835
rect 15887 12801 15896 12835
rect 15844 12792 15896 12801
rect 1400 12767 1452 12776
rect 1400 12733 1409 12767
rect 1409 12733 1443 12767
rect 1443 12733 1452 12767
rect 1400 12724 1452 12733
rect 4436 12724 4488 12776
rect 5356 12724 5408 12776
rect 8208 12724 8260 12776
rect 2964 12656 3016 12708
rect 3056 12631 3108 12640
rect 3056 12597 3065 12631
rect 3065 12597 3099 12631
rect 3099 12597 3108 12631
rect 3056 12588 3108 12597
rect 4528 12588 4580 12640
rect 7104 12656 7156 12708
rect 8392 12656 8444 12708
rect 10048 12656 10100 12708
rect 4988 12631 5040 12640
rect 4988 12597 4997 12631
rect 4997 12597 5031 12631
rect 5031 12597 5040 12631
rect 4988 12588 5040 12597
rect 9404 12631 9456 12640
rect 9404 12597 9413 12631
rect 9413 12597 9447 12631
rect 9447 12597 9456 12631
rect 9404 12588 9456 12597
rect 9496 12631 9548 12640
rect 9496 12597 9505 12631
rect 9505 12597 9539 12631
rect 9539 12597 9548 12631
rect 12532 12724 12584 12776
rect 13360 12724 13412 12776
rect 15200 12724 15252 12776
rect 15292 12724 15344 12776
rect 12440 12656 12492 12708
rect 13268 12656 13320 12708
rect 17960 12724 18012 12776
rect 18880 12835 18932 12844
rect 18880 12801 18889 12835
rect 18889 12801 18923 12835
rect 18923 12801 18932 12835
rect 19892 12835 19944 12844
rect 18880 12792 18932 12801
rect 19892 12801 19901 12835
rect 19901 12801 19935 12835
rect 19935 12801 19944 12835
rect 19892 12792 19944 12801
rect 20352 12792 20404 12844
rect 20628 12767 20680 12776
rect 20628 12733 20637 12767
rect 20637 12733 20671 12767
rect 20671 12733 20680 12767
rect 20628 12724 20680 12733
rect 18420 12656 18472 12708
rect 19432 12656 19484 12708
rect 19524 12656 19576 12708
rect 21272 12699 21324 12708
rect 21272 12665 21281 12699
rect 21281 12665 21315 12699
rect 21315 12665 21324 12699
rect 21272 12656 21324 12665
rect 14188 12631 14240 12640
rect 9496 12588 9548 12597
rect 14188 12597 14197 12631
rect 14197 12597 14231 12631
rect 14231 12597 14240 12631
rect 14188 12588 14240 12597
rect 15660 12588 15712 12640
rect 16396 12588 16448 12640
rect 19708 12631 19760 12640
rect 19708 12597 19717 12631
rect 19717 12597 19751 12631
rect 19751 12597 19760 12631
rect 19708 12588 19760 12597
rect 20720 12631 20772 12640
rect 20720 12597 20729 12631
rect 20729 12597 20763 12631
rect 20763 12597 20772 12631
rect 20720 12588 20772 12597
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 22008 12495 22060 12504
rect 22008 12461 22017 12495
rect 22017 12461 22051 12495
rect 22051 12461 22060 12495
rect 22008 12452 22060 12461
rect 2688 12427 2740 12436
rect 2688 12393 2697 12427
rect 2697 12393 2731 12427
rect 2731 12393 2740 12427
rect 2688 12384 2740 12393
rect 2872 12384 2924 12436
rect 3516 12384 3568 12436
rect 4804 12384 4856 12436
rect 1676 12359 1728 12368
rect 1676 12325 1685 12359
rect 1685 12325 1719 12359
rect 1719 12325 1728 12359
rect 1676 12316 1728 12325
rect 3056 12316 3108 12368
rect 4160 12316 4212 12368
rect 6276 12384 6328 12436
rect 7012 12384 7064 12436
rect 9496 12384 9548 12436
rect 12164 12384 12216 12436
rect 12440 12427 12492 12436
rect 12440 12393 12449 12427
rect 12449 12393 12483 12427
rect 12483 12393 12492 12427
rect 12440 12384 12492 12393
rect 15476 12384 15528 12436
rect 15844 12384 15896 12436
rect 17132 12384 17184 12436
rect 18420 12427 18472 12436
rect 18420 12393 18429 12427
rect 18429 12393 18463 12427
rect 18463 12393 18472 12427
rect 18420 12384 18472 12393
rect 18512 12384 18564 12436
rect 18972 12384 19024 12436
rect 19800 12427 19852 12436
rect 19800 12393 19809 12427
rect 19809 12393 19843 12427
rect 19843 12393 19852 12427
rect 19800 12384 19852 12393
rect 20168 12427 20220 12436
rect 20168 12393 20177 12427
rect 20177 12393 20211 12427
rect 20211 12393 20220 12427
rect 20168 12384 20220 12393
rect 1860 12248 1912 12300
rect 2596 12223 2648 12232
rect 2596 12189 2605 12223
rect 2605 12189 2639 12223
rect 2639 12189 2648 12223
rect 2596 12180 2648 12189
rect 3516 12248 3568 12300
rect 4436 12248 4488 12300
rect 14188 12316 14240 12368
rect 14924 12316 14976 12368
rect 15752 12316 15804 12368
rect 17592 12359 17644 12368
rect 17592 12325 17610 12359
rect 17610 12325 17644 12359
rect 17592 12316 17644 12325
rect 18236 12316 18288 12368
rect 1768 12087 1820 12096
rect 1768 12053 1777 12087
rect 1777 12053 1811 12087
rect 1811 12053 1820 12087
rect 1768 12044 1820 12053
rect 4344 12112 4396 12164
rect 4620 12112 4672 12164
rect 4804 12112 4856 12164
rect 6000 12248 6052 12300
rect 8760 12248 8812 12300
rect 5264 12223 5316 12232
rect 5264 12189 5273 12223
rect 5273 12189 5307 12223
rect 5307 12189 5316 12223
rect 7748 12223 7800 12232
rect 5264 12180 5316 12189
rect 7748 12189 7757 12223
rect 7757 12189 7791 12223
rect 7791 12189 7800 12223
rect 7748 12180 7800 12189
rect 11152 12248 11204 12300
rect 11704 12248 11756 12300
rect 11796 12248 11848 12300
rect 9956 12223 10008 12232
rect 9956 12189 9965 12223
rect 9965 12189 9999 12223
rect 9999 12189 10008 12223
rect 9956 12180 10008 12189
rect 12900 12223 12952 12232
rect 12900 12189 12909 12223
rect 12909 12189 12943 12223
rect 12943 12189 12952 12223
rect 12900 12180 12952 12189
rect 13268 12223 13320 12232
rect 13268 12189 13277 12223
rect 13277 12189 13311 12223
rect 13311 12189 13320 12223
rect 13268 12180 13320 12189
rect 18144 12248 18196 12300
rect 18696 12248 18748 12300
rect 18788 12248 18840 12300
rect 20812 12248 20864 12300
rect 18236 12223 18288 12232
rect 8760 12112 8812 12164
rect 3424 12087 3476 12096
rect 3424 12053 3433 12087
rect 3433 12053 3467 12087
rect 3467 12053 3476 12087
rect 3424 12044 3476 12053
rect 4068 12044 4120 12096
rect 7012 12044 7064 12096
rect 7288 12044 7340 12096
rect 13176 12112 13228 12164
rect 11980 12044 12032 12096
rect 14188 12044 14240 12096
rect 14464 12112 14516 12164
rect 18236 12189 18245 12223
rect 18245 12189 18279 12223
rect 18279 12189 18288 12223
rect 18236 12180 18288 12189
rect 19156 12180 19208 12232
rect 20168 12180 20220 12232
rect 20352 12223 20404 12232
rect 20352 12189 20361 12223
rect 20361 12189 20395 12223
rect 20395 12189 20404 12223
rect 20352 12180 20404 12189
rect 20076 12112 20128 12164
rect 14924 12044 14976 12096
rect 15292 12044 15344 12096
rect 15844 12044 15896 12096
rect 17684 12044 17736 12096
rect 18788 12044 18840 12096
rect 18972 12044 19024 12096
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 1768 11840 1820 11892
rect 3700 11883 3752 11892
rect 1860 11815 1912 11824
rect 1860 11781 1869 11815
rect 1869 11781 1903 11815
rect 1903 11781 1912 11815
rect 1860 11772 1912 11781
rect 1676 11679 1728 11688
rect 1676 11645 1685 11679
rect 1685 11645 1719 11679
rect 1719 11645 1728 11679
rect 1676 11636 1728 11645
rect 2044 11636 2096 11688
rect 3424 11636 3476 11688
rect 2596 11611 2648 11620
rect 2596 11577 2630 11611
rect 2630 11577 2648 11611
rect 2596 11568 2648 11577
rect 3700 11849 3709 11883
rect 3709 11849 3743 11883
rect 3743 11849 3752 11883
rect 3700 11840 3752 11849
rect 3976 11883 4028 11892
rect 3976 11849 3985 11883
rect 3985 11849 4019 11883
rect 4019 11849 4028 11883
rect 3976 11840 4028 11849
rect 4252 11840 4304 11892
rect 7012 11840 7064 11892
rect 7288 11840 7340 11892
rect 7840 11840 7892 11892
rect 9404 11840 9456 11892
rect 9680 11840 9732 11892
rect 11796 11840 11848 11892
rect 12624 11883 12676 11892
rect 12624 11849 12633 11883
rect 12633 11849 12667 11883
rect 12667 11849 12676 11883
rect 12624 11840 12676 11849
rect 12808 11840 12860 11892
rect 4896 11772 4948 11824
rect 7748 11815 7800 11824
rect 7748 11781 7757 11815
rect 7757 11781 7791 11815
rect 7791 11781 7800 11815
rect 7748 11772 7800 11781
rect 7932 11772 7984 11824
rect 5172 11704 5224 11756
rect 5816 11704 5868 11756
rect 7656 11704 7708 11756
rect 9956 11704 10008 11756
rect 11704 11704 11756 11756
rect 14096 11772 14148 11824
rect 4160 11636 4212 11688
rect 9864 11636 9916 11688
rect 12900 11636 12952 11688
rect 13820 11568 13872 11620
rect 14188 11747 14240 11756
rect 14188 11713 14197 11747
rect 14197 11713 14231 11747
rect 14231 11713 14240 11747
rect 14188 11704 14240 11713
rect 14280 11679 14332 11688
rect 14280 11645 14289 11679
rect 14289 11645 14323 11679
rect 14323 11645 14332 11679
rect 14280 11636 14332 11645
rect 15292 11747 15344 11756
rect 15292 11713 15301 11747
rect 15301 11713 15335 11747
rect 15335 11713 15344 11747
rect 15292 11704 15344 11713
rect 16028 11840 16080 11892
rect 18144 11840 18196 11892
rect 18788 11840 18840 11892
rect 19432 11883 19484 11892
rect 19432 11849 19441 11883
rect 19441 11849 19475 11883
rect 19475 11849 19484 11883
rect 19432 11840 19484 11849
rect 16212 11772 16264 11824
rect 16856 11704 16908 11756
rect 19064 11772 19116 11824
rect 17040 11747 17092 11756
rect 17040 11713 17049 11747
rect 17049 11713 17083 11747
rect 17083 11713 17092 11747
rect 17592 11747 17644 11756
rect 17040 11704 17092 11713
rect 17592 11713 17601 11747
rect 17601 11713 17635 11747
rect 17635 11713 17644 11747
rect 17592 11704 17644 11713
rect 17684 11704 17736 11756
rect 20352 11704 20404 11756
rect 20720 11704 20772 11756
rect 17868 11636 17920 11688
rect 20904 11679 20956 11688
rect 20904 11645 20913 11679
rect 20913 11645 20947 11679
rect 20947 11645 20956 11679
rect 20904 11636 20956 11645
rect 20352 11568 20404 11620
rect 2688 11500 2740 11552
rect 3516 11500 3568 11552
rect 4344 11543 4396 11552
rect 4344 11509 4353 11543
rect 4353 11509 4387 11543
rect 4387 11509 4396 11543
rect 4344 11500 4396 11509
rect 4436 11543 4488 11552
rect 4436 11509 4445 11543
rect 4445 11509 4479 11543
rect 4479 11509 4488 11543
rect 4436 11500 4488 11509
rect 5080 11500 5132 11552
rect 5448 11543 5500 11552
rect 5448 11509 5457 11543
rect 5457 11509 5491 11543
rect 5491 11509 5500 11543
rect 5448 11500 5500 11509
rect 7196 11500 7248 11552
rect 8852 11543 8904 11552
rect 8852 11509 8861 11543
rect 8861 11509 8895 11543
rect 8895 11509 8904 11543
rect 8852 11500 8904 11509
rect 9864 11543 9916 11552
rect 9864 11509 9873 11543
rect 9873 11509 9907 11543
rect 9907 11509 9916 11543
rect 9864 11500 9916 11509
rect 10416 11500 10468 11552
rect 12164 11543 12216 11552
rect 12164 11509 12173 11543
rect 12173 11509 12207 11543
rect 12207 11509 12216 11543
rect 12164 11500 12216 11509
rect 12256 11543 12308 11552
rect 12256 11509 12265 11543
rect 12265 11509 12299 11543
rect 12299 11509 12308 11543
rect 12256 11500 12308 11509
rect 13176 11500 13228 11552
rect 15384 11543 15436 11552
rect 15384 11509 15393 11543
rect 15393 11509 15427 11543
rect 15427 11509 15436 11543
rect 15384 11500 15436 11509
rect 15476 11543 15528 11552
rect 15476 11509 15485 11543
rect 15485 11509 15519 11543
rect 15519 11509 15528 11543
rect 16580 11543 16632 11552
rect 15476 11500 15528 11509
rect 16580 11509 16589 11543
rect 16589 11509 16623 11543
rect 16623 11509 16632 11543
rect 16580 11500 16632 11509
rect 17592 11500 17644 11552
rect 17776 11500 17828 11552
rect 19064 11500 19116 11552
rect 20260 11500 20312 11552
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 4344 11296 4396 11348
rect 5264 11296 5316 11348
rect 6276 11339 6328 11348
rect 6276 11305 6285 11339
rect 6285 11305 6319 11339
rect 6319 11305 6328 11339
rect 6276 11296 6328 11305
rect 1676 11271 1728 11280
rect 1676 11237 1685 11271
rect 1685 11237 1719 11271
rect 1719 11237 1728 11271
rect 1676 11228 1728 11237
rect 3884 11228 3936 11280
rect 4160 11160 4212 11212
rect 5724 11160 5776 11212
rect 7012 11271 7064 11280
rect 7012 11237 7021 11271
rect 7021 11237 7055 11271
rect 7055 11237 7064 11271
rect 7012 11228 7064 11237
rect 7748 11228 7800 11280
rect 8208 11228 8260 11280
rect 8852 11296 8904 11348
rect 11244 11296 11296 11348
rect 12256 11296 12308 11348
rect 10876 11228 10928 11280
rect 15200 11296 15252 11348
rect 15844 11296 15896 11348
rect 15936 11296 15988 11348
rect 18052 11296 18104 11348
rect 20628 11296 20680 11348
rect 13452 11203 13504 11212
rect 13452 11169 13461 11203
rect 13461 11169 13495 11203
rect 13495 11169 13504 11203
rect 13452 11160 13504 11169
rect 18880 11228 18932 11280
rect 20352 11228 20404 11280
rect 17960 11203 18012 11212
rect 17960 11169 17969 11203
rect 17969 11169 18003 11203
rect 18003 11169 18012 11203
rect 17960 11160 18012 11169
rect 19064 11203 19116 11212
rect 19064 11169 19073 11203
rect 19073 11169 19107 11203
rect 19107 11169 19116 11203
rect 19064 11160 19116 11169
rect 20076 11160 20128 11212
rect 2596 11135 2648 11144
rect 2596 11101 2605 11135
rect 2605 11101 2639 11135
rect 2639 11101 2648 11135
rect 2596 11092 2648 11101
rect 4252 11092 4304 11144
rect 3792 10956 3844 11008
rect 8024 11024 8076 11076
rect 8852 11092 8904 11144
rect 9036 11092 9088 11144
rect 8576 11024 8628 11076
rect 11244 11092 11296 11144
rect 11980 11092 12032 11144
rect 15476 11092 15528 11144
rect 15384 11024 15436 11076
rect 16028 11092 16080 11144
rect 18052 11135 18104 11144
rect 7104 10956 7156 11008
rect 7656 10999 7708 11008
rect 7656 10965 7665 10999
rect 7665 10965 7699 10999
rect 7699 10965 7708 10999
rect 7656 10956 7708 10965
rect 10140 10956 10192 11008
rect 16212 11024 16264 11076
rect 16764 11024 16816 11076
rect 18052 11101 18061 11135
rect 18061 11101 18095 11135
rect 18095 11101 18104 11135
rect 18052 11092 18104 11101
rect 19156 11092 19208 11144
rect 18972 11024 19024 11076
rect 19892 11092 19944 11144
rect 19708 11067 19760 11076
rect 19708 11033 19717 11067
rect 19717 11033 19751 11067
rect 19751 11033 19760 11067
rect 19708 11024 19760 11033
rect 22008 11067 22060 11076
rect 22008 11033 22017 11067
rect 22017 11033 22051 11067
rect 22051 11033 22060 11067
rect 22008 11024 22060 11033
rect 16120 10956 16172 11008
rect 17224 10999 17276 11008
rect 17224 10965 17233 10999
rect 17233 10965 17267 10999
rect 17267 10965 17276 10999
rect 17224 10956 17276 10965
rect 21364 10999 21416 11008
rect 21364 10965 21373 10999
rect 21373 10965 21407 10999
rect 21407 10965 21416 10999
rect 21364 10956 21416 10965
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 2136 10795 2188 10804
rect 2136 10761 2145 10795
rect 2145 10761 2179 10795
rect 2179 10761 2188 10795
rect 2136 10752 2188 10761
rect 2964 10752 3016 10804
rect 4896 10752 4948 10804
rect 5172 10752 5224 10804
rect 5724 10752 5776 10804
rect 6092 10752 6144 10804
rect 10232 10752 10284 10804
rect 15568 10752 15620 10804
rect 16672 10752 16724 10804
rect 18052 10752 18104 10804
rect 20352 10752 20404 10804
rect 1676 10523 1728 10532
rect 1676 10489 1685 10523
rect 1685 10489 1719 10523
rect 1719 10489 1728 10523
rect 1676 10480 1728 10489
rect 3056 10548 3108 10600
rect 3608 10548 3660 10600
rect 3884 10591 3936 10600
rect 3884 10557 3893 10591
rect 3893 10557 3927 10591
rect 3927 10557 3936 10591
rect 3884 10548 3936 10557
rect 6276 10616 6328 10668
rect 6552 10480 6604 10532
rect 6184 10412 6236 10464
rect 6920 10412 6972 10464
rect 7564 10480 7616 10532
rect 8024 10480 8076 10532
rect 8300 10548 8352 10600
rect 8760 10616 8812 10668
rect 9680 10659 9732 10668
rect 9680 10625 9689 10659
rect 9689 10625 9723 10659
rect 9723 10625 9732 10659
rect 9680 10616 9732 10625
rect 9772 10616 9824 10668
rect 10692 10616 10744 10668
rect 10968 10616 11020 10668
rect 15476 10684 15528 10736
rect 16120 10684 16172 10736
rect 13176 10616 13228 10668
rect 13360 10616 13412 10668
rect 18052 10616 18104 10668
rect 14280 10548 14332 10600
rect 14556 10548 14608 10600
rect 16580 10548 16632 10600
rect 10876 10480 10928 10532
rect 17224 10480 17276 10532
rect 7196 10412 7248 10464
rect 7380 10412 7432 10464
rect 8668 10455 8720 10464
rect 8668 10421 8677 10455
rect 8677 10421 8711 10455
rect 8711 10421 8720 10455
rect 8668 10412 8720 10421
rect 9036 10455 9088 10464
rect 9036 10421 9045 10455
rect 9045 10421 9079 10455
rect 9079 10421 9088 10455
rect 9036 10412 9088 10421
rect 9220 10412 9272 10464
rect 10232 10455 10284 10464
rect 10232 10421 10241 10455
rect 10241 10421 10275 10455
rect 10275 10421 10284 10455
rect 10232 10412 10284 10421
rect 12716 10412 12768 10464
rect 13636 10455 13688 10464
rect 13636 10421 13645 10455
rect 13645 10421 13679 10455
rect 13679 10421 13688 10455
rect 13636 10412 13688 10421
rect 15384 10412 15436 10464
rect 16948 10412 17000 10464
rect 17132 10412 17184 10464
rect 19156 10480 19208 10532
rect 19708 10480 19760 10532
rect 21272 10523 21324 10532
rect 21272 10489 21281 10523
rect 21281 10489 21315 10523
rect 21315 10489 21324 10523
rect 21272 10480 21324 10489
rect 18420 10455 18472 10464
rect 18420 10421 18429 10455
rect 18429 10421 18463 10455
rect 18463 10421 18472 10455
rect 18420 10412 18472 10421
rect 18788 10412 18840 10464
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 3056 10251 3108 10260
rect 3056 10217 3065 10251
rect 3065 10217 3099 10251
rect 3099 10217 3108 10251
rect 3056 10208 3108 10217
rect 3608 10208 3660 10260
rect 7012 10208 7064 10260
rect 7104 10140 7156 10192
rect 1676 10115 1728 10124
rect 1676 10081 1685 10115
rect 1685 10081 1719 10115
rect 1719 10081 1728 10115
rect 1676 10072 1728 10081
rect 2504 10072 2556 10124
rect 3332 10115 3384 10124
rect 3332 10081 3341 10115
rect 3341 10081 3375 10115
rect 3375 10081 3384 10115
rect 3332 10072 3384 10081
rect 7012 10072 7064 10124
rect 7656 10140 7708 10192
rect 8208 10208 8260 10260
rect 8668 10208 8720 10260
rect 10876 10208 10928 10260
rect 10968 10208 11020 10260
rect 11704 10208 11756 10260
rect 12072 10208 12124 10260
rect 13820 10208 13872 10260
rect 15936 10208 15988 10260
rect 16672 10208 16724 10260
rect 18420 10208 18472 10260
rect 19156 10251 19208 10260
rect 19156 10217 19165 10251
rect 19165 10217 19199 10251
rect 19199 10217 19208 10251
rect 19156 10208 19208 10217
rect 20628 10251 20680 10260
rect 20628 10217 20637 10251
rect 20637 10217 20671 10251
rect 20671 10217 20680 10251
rect 20628 10208 20680 10217
rect 9680 10140 9732 10192
rect 10140 10140 10192 10192
rect 8208 10072 8260 10124
rect 8392 10072 8444 10124
rect 8576 10115 8628 10124
rect 8576 10081 8585 10115
rect 8585 10081 8619 10115
rect 8619 10081 8628 10115
rect 8576 10072 8628 10081
rect 9772 10072 9824 10124
rect 10784 10072 10836 10124
rect 21088 10140 21140 10192
rect 12348 10072 12400 10124
rect 12532 10115 12584 10124
rect 12532 10081 12566 10115
rect 12566 10081 12584 10115
rect 15200 10115 15252 10124
rect 12532 10072 12584 10081
rect 2780 10004 2832 10056
rect 5724 10004 5776 10056
rect 6368 10047 6420 10056
rect 6368 10013 6377 10047
rect 6377 10013 6411 10047
rect 6411 10013 6420 10047
rect 6368 10004 6420 10013
rect 6552 10047 6604 10056
rect 6552 10013 6561 10047
rect 6561 10013 6595 10047
rect 6595 10013 6604 10047
rect 6552 10004 6604 10013
rect 8760 10004 8812 10056
rect 15200 10081 15209 10115
rect 15209 10081 15243 10115
rect 15243 10081 15252 10115
rect 15200 10072 15252 10081
rect 15844 10115 15896 10124
rect 15844 10081 15853 10115
rect 15853 10081 15887 10115
rect 15887 10081 15896 10115
rect 15844 10072 15896 10081
rect 18052 10115 18104 10124
rect 15384 10047 15436 10056
rect 15384 10013 15393 10047
rect 15393 10013 15427 10047
rect 15427 10013 15436 10047
rect 18052 10081 18086 10115
rect 18086 10081 18104 10115
rect 18052 10072 18104 10081
rect 15384 10004 15436 10013
rect 3424 9936 3476 9988
rect 9220 9936 9272 9988
rect 11060 9979 11112 9988
rect 11060 9945 11069 9979
rect 11069 9945 11103 9979
rect 11103 9945 11112 9979
rect 11060 9936 11112 9945
rect 12072 9936 12124 9988
rect 17132 10004 17184 10056
rect 20812 10047 20864 10056
rect 20812 10013 20821 10047
rect 20821 10013 20855 10047
rect 20855 10013 20864 10047
rect 20812 10004 20864 10013
rect 21364 10004 21416 10056
rect 16488 9979 16540 9988
rect 16488 9945 16497 9979
rect 16497 9945 16531 9979
rect 16531 9945 16540 9979
rect 16488 9936 16540 9945
rect 17684 9936 17736 9988
rect 8300 9868 8352 9920
rect 8392 9911 8444 9920
rect 8392 9877 8401 9911
rect 8401 9877 8435 9911
rect 8435 9877 8444 9911
rect 8392 9868 8444 9877
rect 13728 9868 13780 9920
rect 13820 9868 13872 9920
rect 16120 9868 16172 9920
rect 16304 9868 16356 9920
rect 17960 9868 18012 9920
rect 19524 9868 19576 9920
rect 20168 9911 20220 9920
rect 20168 9877 20177 9911
rect 20177 9877 20211 9911
rect 20211 9877 20220 9911
rect 20168 9868 20220 9877
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 2044 9664 2096 9716
rect 3884 9664 3936 9716
rect 7012 9664 7064 9716
rect 3424 9639 3476 9648
rect 3424 9605 3433 9639
rect 3433 9605 3467 9639
rect 3467 9605 3476 9639
rect 3424 9596 3476 9605
rect 7840 9596 7892 9648
rect 10324 9596 10376 9648
rect 10968 9596 11020 9648
rect 11704 9664 11756 9716
rect 11796 9596 11848 9648
rect 14280 9664 14332 9716
rect 14648 9664 14700 9716
rect 17316 9664 17368 9716
rect 18052 9664 18104 9716
rect 19432 9596 19484 9648
rect 21088 9639 21140 9648
rect 21088 9605 21097 9639
rect 21097 9605 21131 9639
rect 21131 9605 21140 9639
rect 21088 9596 21140 9605
rect 1584 9503 1636 9512
rect 1584 9469 1593 9503
rect 1593 9469 1627 9503
rect 1627 9469 1636 9503
rect 1584 9460 1636 9469
rect 2044 9503 2096 9512
rect 2044 9469 2053 9503
rect 2053 9469 2087 9503
rect 2087 9469 2096 9503
rect 2044 9460 2096 9469
rect 7104 9528 7156 9580
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 7564 9528 7616 9580
rect 9588 9528 9640 9580
rect 11060 9528 11112 9580
rect 15200 9571 15252 9580
rect 15200 9537 15209 9571
rect 15209 9537 15243 9571
rect 15243 9537 15252 9571
rect 15200 9528 15252 9537
rect 16212 9571 16264 9580
rect 16212 9537 16221 9571
rect 16221 9537 16255 9571
rect 16255 9537 16264 9571
rect 16212 9528 16264 9537
rect 16304 9571 16356 9580
rect 16304 9537 16313 9571
rect 16313 9537 16347 9571
rect 16347 9537 16356 9571
rect 17132 9571 17184 9580
rect 16304 9528 16356 9537
rect 17132 9537 17141 9571
rect 17141 9537 17175 9571
rect 17175 9537 17184 9571
rect 17132 9528 17184 9537
rect 20260 9571 20312 9580
rect 3976 9460 4028 9512
rect 8392 9460 8444 9512
rect 10324 9503 10376 9512
rect 1860 9392 1912 9444
rect 2688 9392 2740 9444
rect 1676 9367 1728 9376
rect 1676 9333 1685 9367
rect 1685 9333 1719 9367
rect 1719 9333 1728 9367
rect 1676 9324 1728 9333
rect 3148 9324 3200 9376
rect 4344 9392 4396 9444
rect 7656 9392 7708 9444
rect 9956 9392 10008 9444
rect 4896 9324 4948 9376
rect 5080 9324 5132 9376
rect 5356 9324 5408 9376
rect 5816 9324 5868 9376
rect 7012 9324 7064 9376
rect 8300 9324 8352 9376
rect 8576 9324 8628 9376
rect 9772 9324 9824 9376
rect 10324 9469 10333 9503
rect 10333 9469 10367 9503
rect 10367 9469 10376 9503
rect 10324 9460 10376 9469
rect 16948 9460 17000 9512
rect 19524 9503 19576 9512
rect 19524 9469 19533 9503
rect 19533 9469 19567 9503
rect 19567 9469 19576 9503
rect 19524 9460 19576 9469
rect 20260 9537 20269 9571
rect 20269 9537 20303 9571
rect 20303 9537 20312 9571
rect 20260 9528 20312 9537
rect 20812 9528 20864 9580
rect 12072 9392 12124 9444
rect 12256 9392 12308 9444
rect 13728 9392 13780 9444
rect 17408 9435 17460 9444
rect 10692 9367 10744 9376
rect 10692 9333 10701 9367
rect 10701 9333 10735 9367
rect 10735 9333 10744 9367
rect 10692 9324 10744 9333
rect 11336 9324 11388 9376
rect 11888 9324 11940 9376
rect 13268 9367 13320 9376
rect 13268 9333 13277 9367
rect 13277 9333 13311 9367
rect 13311 9333 13320 9367
rect 13268 9324 13320 9333
rect 14740 9324 14792 9376
rect 15200 9324 15252 9376
rect 16120 9367 16172 9376
rect 16120 9333 16129 9367
rect 16129 9333 16163 9367
rect 16163 9333 16172 9367
rect 16120 9324 16172 9333
rect 17408 9401 17442 9435
rect 17442 9401 17460 9435
rect 17408 9392 17460 9401
rect 21272 9435 21324 9444
rect 21272 9401 21281 9435
rect 21281 9401 21315 9435
rect 21315 9401 21324 9435
rect 21272 9392 21324 9401
rect 19616 9324 19668 9376
rect 19800 9367 19852 9376
rect 19800 9333 19809 9367
rect 19809 9333 19843 9367
rect 19843 9333 19852 9367
rect 19800 9324 19852 9333
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 2504 9163 2556 9172
rect 2504 9129 2513 9163
rect 2513 9129 2547 9163
rect 2547 9129 2556 9163
rect 2504 9120 2556 9129
rect 2780 9163 2832 9172
rect 2780 9129 2789 9163
rect 2789 9129 2823 9163
rect 2823 9129 2832 9163
rect 2780 9120 2832 9129
rect 1952 9052 2004 9104
rect 3700 9120 3752 9172
rect 3424 9052 3476 9104
rect 2136 9027 2188 9036
rect 2136 8993 2145 9027
rect 2145 8993 2179 9027
rect 2179 8993 2188 9027
rect 2136 8984 2188 8993
rect 3608 8984 3660 9036
rect 1860 8959 1912 8968
rect 1860 8925 1869 8959
rect 1869 8925 1903 8959
rect 1903 8925 1912 8959
rect 1860 8916 1912 8925
rect 2044 8959 2096 8968
rect 2044 8925 2053 8959
rect 2053 8925 2087 8959
rect 2087 8925 2096 8959
rect 2044 8916 2096 8925
rect 2964 8916 3016 8968
rect 3424 8916 3476 8968
rect 3884 8916 3936 8968
rect 5816 8984 5868 9036
rect 6000 9120 6052 9172
rect 7564 9120 7616 9172
rect 7748 9163 7800 9172
rect 7748 9129 7757 9163
rect 7757 9129 7791 9163
rect 7791 9129 7800 9163
rect 7748 9120 7800 9129
rect 9588 9120 9640 9172
rect 10876 9120 10928 9172
rect 13820 9120 13872 9172
rect 15200 9120 15252 9172
rect 8300 9052 8352 9104
rect 16120 9052 16172 9104
rect 17776 9052 17828 9104
rect 7380 8984 7432 9036
rect 7196 8916 7248 8968
rect 8484 8984 8536 9036
rect 9680 9027 9732 9036
rect 9680 8993 9689 9027
rect 9689 8993 9723 9027
rect 9723 8993 9732 9027
rect 9680 8984 9732 8993
rect 9404 8959 9456 8968
rect 9404 8925 9413 8959
rect 9413 8925 9447 8959
rect 9447 8925 9456 8959
rect 9404 8916 9456 8925
rect 1400 8823 1452 8832
rect 1400 8789 1409 8823
rect 1409 8789 1443 8823
rect 1443 8789 1452 8823
rect 1400 8780 1452 8789
rect 2504 8780 2556 8832
rect 3792 8780 3844 8832
rect 7380 8823 7432 8832
rect 7380 8789 7389 8823
rect 7389 8789 7423 8823
rect 7423 8789 7432 8823
rect 7380 8780 7432 8789
rect 9680 8848 9732 8900
rect 11336 8984 11388 9036
rect 12440 9027 12492 9036
rect 12440 8993 12449 9027
rect 12449 8993 12483 9027
rect 12483 8993 12492 9027
rect 12440 8984 12492 8993
rect 10140 8848 10192 8900
rect 11244 8916 11296 8968
rect 12532 8916 12584 8968
rect 10968 8848 11020 8900
rect 11704 8780 11756 8832
rect 12808 8823 12860 8832
rect 12808 8789 12817 8823
rect 12817 8789 12851 8823
rect 12851 8789 12860 8823
rect 12808 8780 12860 8789
rect 16212 8984 16264 9036
rect 14740 8916 14792 8968
rect 18604 8984 18656 9036
rect 19800 9120 19852 9172
rect 20168 9052 20220 9104
rect 20812 9052 20864 9104
rect 19340 8984 19392 9036
rect 18880 8916 18932 8968
rect 21180 8959 21232 8968
rect 13728 8780 13780 8832
rect 17224 8780 17276 8832
rect 17960 8780 18012 8832
rect 18144 8823 18196 8832
rect 18144 8789 18153 8823
rect 18153 8789 18187 8823
rect 18187 8789 18196 8823
rect 18144 8780 18196 8789
rect 18604 8780 18656 8832
rect 19064 8848 19116 8900
rect 21180 8925 21189 8959
rect 21189 8925 21223 8959
rect 21223 8925 21232 8959
rect 21180 8916 21232 8925
rect 19248 8780 19300 8832
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 1676 8576 1728 8628
rect 1860 8551 1912 8560
rect 1860 8517 1869 8551
rect 1869 8517 1903 8551
rect 1903 8517 1912 8551
rect 1860 8508 1912 8517
rect 3056 8304 3108 8356
rect 1584 8279 1636 8288
rect 1584 8245 1593 8279
rect 1593 8245 1627 8279
rect 1627 8245 1636 8279
rect 1584 8236 1636 8245
rect 3608 8576 3660 8628
rect 6368 8576 6420 8628
rect 4068 8508 4120 8560
rect 4620 8440 4672 8492
rect 4988 8440 5040 8492
rect 3608 8415 3660 8424
rect 3608 8381 3617 8415
rect 3617 8381 3651 8415
rect 3651 8381 3660 8415
rect 3608 8372 3660 8381
rect 5448 8440 5500 8492
rect 6736 8440 6788 8492
rect 7380 8508 7432 8560
rect 11244 8576 11296 8628
rect 12440 8619 12492 8628
rect 12440 8585 12449 8619
rect 12449 8585 12483 8619
rect 12483 8585 12492 8619
rect 12440 8576 12492 8585
rect 12808 8576 12860 8628
rect 8484 8551 8536 8560
rect 7564 8440 7616 8492
rect 8484 8517 8493 8551
rect 8493 8517 8527 8551
rect 8527 8517 8536 8551
rect 8484 8508 8536 8517
rect 10140 8551 10192 8560
rect 10140 8517 10149 8551
rect 10149 8517 10183 8551
rect 10183 8517 10192 8551
rect 10140 8508 10192 8517
rect 8024 8483 8076 8492
rect 8024 8449 8033 8483
rect 8033 8449 8067 8483
rect 8067 8449 8076 8483
rect 8024 8440 8076 8449
rect 5724 8415 5776 8424
rect 5724 8381 5733 8415
rect 5733 8381 5767 8415
rect 5767 8381 5776 8415
rect 5724 8372 5776 8381
rect 7012 8415 7064 8424
rect 7012 8381 7021 8415
rect 7021 8381 7055 8415
rect 7055 8381 7064 8415
rect 7012 8372 7064 8381
rect 7656 8372 7708 8424
rect 8760 8415 8812 8424
rect 8760 8381 8769 8415
rect 8769 8381 8803 8415
rect 8803 8381 8812 8415
rect 8760 8372 8812 8381
rect 9404 8372 9456 8424
rect 9496 8372 9548 8424
rect 10324 8440 10376 8492
rect 11704 8508 11756 8560
rect 12900 8508 12952 8560
rect 14648 8508 14700 8560
rect 17408 8508 17460 8560
rect 14280 8440 14332 8492
rect 18052 8508 18104 8560
rect 18696 8508 18748 8560
rect 3424 8236 3476 8288
rect 3792 8236 3844 8288
rect 3884 8236 3936 8288
rect 4528 8236 4580 8288
rect 4896 8279 4948 8288
rect 4896 8245 4905 8279
rect 4905 8245 4939 8279
rect 4939 8245 4948 8279
rect 4896 8236 4948 8245
rect 4988 8236 5040 8288
rect 9220 8236 9272 8288
rect 10508 8304 10560 8356
rect 13268 8372 13320 8424
rect 11796 8236 11848 8288
rect 12072 8236 12124 8288
rect 14004 8304 14056 8356
rect 14464 8372 14516 8424
rect 18236 8440 18288 8492
rect 14556 8304 14608 8356
rect 14648 8236 14700 8288
rect 16580 8304 16632 8356
rect 16948 8372 17000 8424
rect 18696 8372 18748 8424
rect 19064 8415 19116 8424
rect 19064 8381 19098 8415
rect 19098 8381 19116 8415
rect 19064 8372 19116 8381
rect 21272 8415 21324 8424
rect 21272 8381 21281 8415
rect 21281 8381 21315 8415
rect 21315 8381 21324 8415
rect 21272 8372 21324 8381
rect 19248 8304 19300 8356
rect 20720 8347 20772 8356
rect 20720 8313 20729 8347
rect 20729 8313 20763 8347
rect 20763 8313 20772 8347
rect 20720 8304 20772 8313
rect 17132 8279 17184 8288
rect 17132 8245 17141 8279
rect 17141 8245 17175 8279
rect 17175 8245 17184 8279
rect 17132 8236 17184 8245
rect 17316 8236 17368 8288
rect 20168 8279 20220 8288
rect 20168 8245 20177 8279
rect 20177 8245 20211 8279
rect 20211 8245 20220 8279
rect 20168 8236 20220 8245
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 2044 8032 2096 8084
rect 1492 7964 1544 8016
rect 2872 7939 2924 7948
rect 2872 7905 2881 7939
rect 2881 7905 2915 7939
rect 2915 7905 2924 7939
rect 2872 7896 2924 7905
rect 3240 7896 3292 7948
rect 8484 8032 8536 8084
rect 9496 8032 9548 8084
rect 12072 8032 12124 8084
rect 14648 8032 14700 8084
rect 16948 8075 17000 8084
rect 16948 8041 16957 8075
rect 16957 8041 16991 8075
rect 16991 8041 17000 8075
rect 16948 8032 17000 8041
rect 17316 8075 17368 8084
rect 17316 8041 17325 8075
rect 17325 8041 17359 8075
rect 17359 8041 17368 8075
rect 17316 8032 17368 8041
rect 17684 8032 17736 8084
rect 18144 8032 18196 8084
rect 4068 7964 4120 8016
rect 6552 7964 6604 8016
rect 11704 7964 11756 8016
rect 13636 7964 13688 8016
rect 14280 7964 14332 8016
rect 14832 8007 14884 8016
rect 14832 7973 14866 8007
rect 14866 7973 14884 8007
rect 14832 7964 14884 7973
rect 17040 7964 17092 8016
rect 4988 7896 5040 7948
rect 5816 7896 5868 7948
rect 8392 7896 8444 7948
rect 9220 7896 9272 7948
rect 12348 7896 12400 7948
rect 13544 7896 13596 7948
rect 16212 7896 16264 7948
rect 16580 7896 16632 7948
rect 17868 7964 17920 8016
rect 17960 7964 18012 8016
rect 18880 7964 18932 8016
rect 20720 8007 20772 8016
rect 20720 7973 20729 8007
rect 20729 7973 20763 8007
rect 20763 7973 20772 8007
rect 20720 7964 20772 7973
rect 19156 7896 19208 7948
rect 20076 7939 20128 7948
rect 20076 7905 20085 7939
rect 20085 7905 20119 7939
rect 20119 7905 20128 7939
rect 20076 7896 20128 7905
rect 3056 7871 3108 7880
rect 3056 7837 3065 7871
rect 3065 7837 3099 7871
rect 3099 7837 3108 7871
rect 3056 7828 3108 7837
rect 4160 7828 4212 7880
rect 4804 7828 4856 7880
rect 1860 7803 1912 7812
rect 1860 7769 1869 7803
rect 1869 7769 1903 7803
rect 1903 7769 1912 7803
rect 1860 7760 1912 7769
rect 4528 7760 4580 7812
rect 5264 7828 5316 7880
rect 5632 7828 5684 7880
rect 7748 7828 7800 7880
rect 5724 7760 5776 7812
rect 8300 7760 8352 7812
rect 8392 7760 8444 7812
rect 9680 7760 9732 7812
rect 12256 7828 12308 7880
rect 3332 7692 3384 7744
rect 6920 7735 6972 7744
rect 6920 7701 6929 7735
rect 6929 7701 6963 7735
rect 6963 7701 6972 7735
rect 6920 7692 6972 7701
rect 7012 7692 7064 7744
rect 8760 7692 8812 7744
rect 10784 7692 10836 7744
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 14556 7871 14608 7880
rect 13360 7828 13412 7837
rect 14556 7837 14565 7871
rect 14565 7837 14599 7871
rect 14599 7837 14608 7871
rect 14556 7828 14608 7837
rect 17868 7871 17920 7880
rect 17868 7837 17877 7871
rect 17877 7837 17911 7871
rect 17911 7837 17920 7871
rect 17868 7828 17920 7837
rect 19616 7828 19668 7880
rect 16580 7760 16632 7812
rect 12808 7735 12860 7744
rect 12808 7701 12817 7735
rect 12817 7701 12851 7735
rect 12851 7701 12860 7735
rect 12808 7692 12860 7701
rect 13268 7692 13320 7744
rect 14464 7692 14516 7744
rect 15200 7692 15252 7744
rect 17040 7692 17092 7744
rect 17224 7692 17276 7744
rect 18144 7692 18196 7744
rect 19248 7735 19300 7744
rect 19248 7701 19257 7735
rect 19257 7701 19291 7735
rect 19291 7701 19300 7735
rect 19248 7692 19300 7701
rect 20260 7735 20312 7744
rect 20260 7701 20269 7735
rect 20269 7701 20303 7735
rect 20303 7701 20312 7735
rect 20260 7692 20312 7701
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 2136 7488 2188 7540
rect 3700 7488 3752 7540
rect 5264 7531 5316 7540
rect 1952 7420 2004 7472
rect 5264 7497 5273 7531
rect 5273 7497 5307 7531
rect 5307 7497 5316 7531
rect 5264 7488 5316 7497
rect 5448 7488 5500 7540
rect 3056 7352 3108 7404
rect 3700 7352 3752 7404
rect 3884 7352 3936 7404
rect 4436 7395 4488 7404
rect 4436 7361 4445 7395
rect 4445 7361 4479 7395
rect 4479 7361 4488 7395
rect 4436 7352 4488 7361
rect 4712 7352 4764 7404
rect 6736 7420 6788 7472
rect 6828 7420 6880 7472
rect 7748 7420 7800 7472
rect 9404 7488 9456 7540
rect 10876 7531 10928 7540
rect 10876 7497 10885 7531
rect 10885 7497 10919 7531
rect 10919 7497 10928 7531
rect 10876 7488 10928 7497
rect 14004 7531 14056 7540
rect 9680 7420 9732 7472
rect 5540 7352 5592 7404
rect 9036 7352 9088 7404
rect 1584 7284 1636 7336
rect 4804 7284 4856 7336
rect 6184 7284 6236 7336
rect 6368 7284 6420 7336
rect 3424 7259 3476 7268
rect 1584 7148 1636 7200
rect 3424 7225 3433 7259
rect 3433 7225 3467 7259
rect 3467 7225 3476 7259
rect 3424 7216 3476 7225
rect 9128 7284 9180 7336
rect 11152 7284 11204 7336
rect 12808 7395 12860 7404
rect 12808 7361 12817 7395
rect 12817 7361 12851 7395
rect 12851 7361 12860 7395
rect 12808 7352 12860 7361
rect 12900 7395 12952 7404
rect 12900 7361 12909 7395
rect 12909 7361 12943 7395
rect 12943 7361 12952 7395
rect 12900 7352 12952 7361
rect 14004 7497 14013 7531
rect 14013 7497 14047 7531
rect 14047 7497 14056 7531
rect 14004 7488 14056 7497
rect 16120 7488 16172 7540
rect 17500 7488 17552 7540
rect 17868 7488 17920 7540
rect 13176 7420 13228 7472
rect 16488 7420 16540 7472
rect 18328 7420 18380 7472
rect 20444 7488 20496 7540
rect 21272 7488 21324 7540
rect 18696 7420 18748 7472
rect 13544 7352 13596 7404
rect 16856 7284 16908 7336
rect 17040 7284 17092 7336
rect 19064 7327 19116 7336
rect 19064 7293 19073 7327
rect 19073 7293 19107 7327
rect 19107 7293 19116 7327
rect 19064 7284 19116 7293
rect 20168 7352 20220 7404
rect 21272 7327 21324 7336
rect 21272 7293 21281 7327
rect 21281 7293 21315 7327
rect 21315 7293 21324 7327
rect 21272 7284 21324 7293
rect 3884 7191 3936 7200
rect 3884 7157 3893 7191
rect 3893 7157 3927 7191
rect 3927 7157 3936 7191
rect 3884 7148 3936 7157
rect 4988 7191 5040 7200
rect 4988 7157 4997 7191
rect 4997 7157 5031 7191
rect 5031 7157 5040 7191
rect 4988 7148 5040 7157
rect 6092 7148 6144 7200
rect 6460 7191 6512 7200
rect 6460 7157 6469 7191
rect 6469 7157 6503 7191
rect 6503 7157 6512 7191
rect 6460 7148 6512 7157
rect 7380 7148 7432 7200
rect 7748 7148 7800 7200
rect 8760 7216 8812 7268
rect 9588 7216 9640 7268
rect 9680 7216 9732 7268
rect 16580 7216 16632 7268
rect 16672 7216 16724 7268
rect 9220 7148 9272 7200
rect 10876 7148 10928 7200
rect 11060 7148 11112 7200
rect 12348 7191 12400 7200
rect 12348 7157 12357 7191
rect 12357 7157 12391 7191
rect 12391 7157 12400 7191
rect 12348 7148 12400 7157
rect 12440 7148 12492 7200
rect 14648 7191 14700 7200
rect 14648 7157 14657 7191
rect 14657 7157 14691 7191
rect 14691 7157 14700 7191
rect 14648 7148 14700 7157
rect 16212 7148 16264 7200
rect 18880 7191 18932 7200
rect 18880 7157 18889 7191
rect 18889 7157 18923 7191
rect 18923 7157 18932 7191
rect 18880 7148 18932 7157
rect 18972 7148 19024 7200
rect 19708 7191 19760 7200
rect 19708 7157 19717 7191
rect 19717 7157 19751 7191
rect 19751 7157 19760 7191
rect 19708 7148 19760 7157
rect 19892 7216 19944 7268
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 2780 6987 2832 6996
rect 2780 6953 2789 6987
rect 2789 6953 2823 6987
rect 2823 6953 2832 6987
rect 2780 6944 2832 6953
rect 3332 6944 3384 6996
rect 3516 6876 3568 6928
rect 2320 6808 2372 6860
rect 3148 6808 3200 6860
rect 3700 6944 3752 6996
rect 4068 6944 4120 6996
rect 5724 6944 5776 6996
rect 7748 6987 7800 6996
rect 7748 6953 7757 6987
rect 7757 6953 7791 6987
rect 7791 6953 7800 6987
rect 7748 6944 7800 6953
rect 8300 6944 8352 6996
rect 8484 6944 8536 6996
rect 12348 6987 12400 6996
rect 4436 6876 4488 6928
rect 12348 6953 12357 6987
rect 12357 6953 12391 6987
rect 12391 6953 12400 6987
rect 12348 6944 12400 6953
rect 16672 6987 16724 6996
rect 16672 6953 16681 6987
rect 16681 6953 16715 6987
rect 16715 6953 16724 6987
rect 16672 6944 16724 6953
rect 17592 6987 17644 6996
rect 17592 6953 17601 6987
rect 17601 6953 17635 6987
rect 17635 6953 17644 6987
rect 17592 6944 17644 6953
rect 12440 6876 12492 6928
rect 6368 6851 6420 6860
rect 6368 6817 6377 6851
rect 6377 6817 6411 6851
rect 6411 6817 6420 6851
rect 6368 6808 6420 6817
rect 6644 6851 6696 6860
rect 6644 6817 6678 6851
rect 6678 6817 6696 6851
rect 6644 6808 6696 6817
rect 7564 6808 7616 6860
rect 9588 6808 9640 6860
rect 10784 6808 10836 6860
rect 3056 6740 3108 6792
rect 3792 6740 3844 6792
rect 7748 6740 7800 6792
rect 8300 6783 8352 6792
rect 8300 6749 8309 6783
rect 8309 6749 8343 6783
rect 8343 6749 8352 6783
rect 8300 6740 8352 6749
rect 8392 6740 8444 6792
rect 9036 6740 9088 6792
rect 9128 6740 9180 6792
rect 11796 6808 11848 6860
rect 15844 6808 15896 6860
rect 16212 6876 16264 6928
rect 18144 6944 18196 6996
rect 19064 6944 19116 6996
rect 16488 6808 16540 6860
rect 17592 6808 17644 6860
rect 18972 6876 19024 6928
rect 20168 6876 20220 6928
rect 22008 6919 22060 6928
rect 22008 6885 22017 6919
rect 22017 6885 22051 6919
rect 22051 6885 22060 6919
rect 22008 6876 22060 6885
rect 19156 6808 19208 6860
rect 21180 6808 21232 6860
rect 14556 6740 14608 6792
rect 15108 6740 15160 6792
rect 17500 6740 17552 6792
rect 1860 6604 1912 6656
rect 3700 6604 3752 6656
rect 4252 6604 4304 6656
rect 4804 6604 4856 6656
rect 5724 6604 5776 6656
rect 6644 6604 6696 6656
rect 7104 6604 7156 6656
rect 12624 6672 12676 6724
rect 19708 6740 19760 6792
rect 11704 6604 11756 6656
rect 12164 6604 12216 6656
rect 13176 6647 13228 6656
rect 13176 6613 13185 6647
rect 13185 6613 13219 6647
rect 13219 6613 13228 6647
rect 13176 6604 13228 6613
rect 13636 6647 13688 6656
rect 13636 6613 13645 6647
rect 13645 6613 13679 6647
rect 13679 6613 13688 6647
rect 13636 6604 13688 6613
rect 15568 6604 15620 6656
rect 19064 6604 19116 6656
rect 21088 6604 21140 6656
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 3240 6400 3292 6452
rect 4160 6400 4212 6452
rect 8300 6400 8352 6452
rect 4804 6332 4856 6384
rect 6368 6332 6420 6384
rect 2320 6264 2372 6316
rect 3056 6307 3108 6316
rect 3056 6273 3065 6307
rect 3065 6273 3099 6307
rect 3099 6273 3108 6307
rect 3056 6264 3108 6273
rect 3516 6307 3568 6316
rect 3516 6273 3525 6307
rect 3525 6273 3559 6307
rect 3559 6273 3568 6307
rect 3516 6264 3568 6273
rect 1860 6239 1912 6248
rect 1860 6205 1869 6239
rect 1869 6205 1903 6239
rect 1903 6205 1912 6239
rect 1860 6196 1912 6205
rect 1952 6196 2004 6248
rect 4252 6264 4304 6316
rect 5356 6264 5408 6316
rect 5724 6264 5776 6316
rect 2228 6103 2280 6112
rect 2228 6069 2237 6103
rect 2237 6069 2271 6103
rect 2271 6069 2280 6103
rect 2228 6060 2280 6069
rect 3516 6128 3568 6180
rect 6552 6196 6604 6248
rect 6736 6332 6788 6384
rect 12900 6400 12952 6452
rect 10324 6332 10376 6384
rect 7748 6264 7800 6316
rect 13360 6307 13412 6316
rect 13360 6273 13369 6307
rect 13369 6273 13403 6307
rect 13403 6273 13412 6307
rect 13360 6264 13412 6273
rect 6828 6196 6880 6248
rect 8392 6196 8444 6248
rect 9036 6196 9088 6248
rect 9588 6196 9640 6248
rect 9772 6196 9824 6248
rect 14004 6196 14056 6248
rect 15844 6332 15896 6384
rect 17224 6332 17276 6384
rect 16672 6264 16724 6316
rect 17408 6264 17460 6316
rect 18696 6332 18748 6384
rect 18788 6332 18840 6384
rect 19432 6332 19484 6384
rect 18052 6264 18104 6316
rect 18420 6264 18472 6316
rect 18512 6264 18564 6316
rect 17316 6196 17368 6248
rect 17500 6239 17552 6248
rect 17500 6205 17509 6239
rect 17509 6205 17543 6239
rect 17543 6205 17552 6239
rect 17500 6196 17552 6205
rect 18604 6196 18656 6248
rect 19156 6264 19208 6316
rect 4436 6060 4488 6112
rect 5172 6128 5224 6180
rect 5448 6128 5500 6180
rect 5724 6103 5776 6112
rect 5724 6069 5733 6103
rect 5733 6069 5767 6103
rect 5767 6069 5776 6103
rect 5724 6060 5776 6069
rect 6828 6060 6880 6112
rect 8668 6128 8720 6180
rect 9404 6171 9456 6180
rect 9404 6137 9422 6171
rect 9422 6137 9456 6171
rect 9404 6128 9456 6137
rect 8392 6060 8444 6112
rect 10324 6103 10376 6112
rect 10324 6069 10333 6103
rect 10333 6069 10367 6103
rect 10367 6069 10376 6103
rect 10324 6060 10376 6069
rect 10784 6103 10836 6112
rect 10784 6069 10793 6103
rect 10793 6069 10827 6103
rect 10827 6069 10836 6103
rect 10784 6060 10836 6069
rect 11244 6103 11296 6112
rect 11244 6069 11253 6103
rect 11253 6069 11287 6103
rect 11287 6069 11296 6103
rect 11244 6060 11296 6069
rect 11796 6103 11848 6112
rect 11796 6069 11805 6103
rect 11805 6069 11839 6103
rect 11839 6069 11848 6103
rect 11796 6060 11848 6069
rect 12256 6103 12308 6112
rect 12256 6069 12265 6103
rect 12265 6069 12299 6103
rect 12299 6069 12308 6103
rect 12256 6060 12308 6069
rect 12716 6103 12768 6112
rect 12716 6069 12725 6103
rect 12725 6069 12759 6103
rect 12759 6069 12768 6103
rect 12716 6060 12768 6069
rect 13912 6103 13964 6112
rect 13912 6069 13921 6103
rect 13921 6069 13955 6103
rect 13955 6069 13964 6103
rect 13912 6060 13964 6069
rect 14188 6103 14240 6112
rect 14188 6069 14197 6103
rect 14197 6069 14231 6103
rect 14231 6069 14240 6103
rect 14188 6060 14240 6069
rect 14556 6103 14608 6112
rect 14556 6069 14565 6103
rect 14565 6069 14599 6103
rect 14599 6069 14608 6103
rect 14556 6060 14608 6069
rect 15936 6060 15988 6112
rect 16304 6060 16356 6112
rect 16580 6103 16632 6112
rect 16580 6069 16589 6103
rect 16589 6069 16623 6103
rect 16623 6069 16632 6103
rect 16580 6060 16632 6069
rect 17684 6128 17736 6180
rect 21088 6239 21140 6248
rect 21088 6205 21106 6239
rect 21106 6205 21140 6239
rect 21088 6196 21140 6205
rect 21180 6128 21232 6180
rect 18788 6060 18840 6112
rect 18972 6060 19024 6112
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 1676 5831 1728 5840
rect 1676 5797 1685 5831
rect 1685 5797 1719 5831
rect 1719 5797 1728 5831
rect 1676 5788 1728 5797
rect 2780 5856 2832 5908
rect 5540 5856 5592 5908
rect 5724 5856 5776 5908
rect 3976 5788 4028 5840
rect 7472 5856 7524 5908
rect 8760 5899 8812 5908
rect 8760 5865 8769 5899
rect 8769 5865 8803 5899
rect 8803 5865 8812 5899
rect 8760 5856 8812 5865
rect 9772 5856 9824 5908
rect 2412 5763 2464 5772
rect 2412 5729 2446 5763
rect 2446 5729 2464 5763
rect 2412 5720 2464 5729
rect 2780 5720 2832 5772
rect 3792 5720 3844 5772
rect 5540 5652 5592 5704
rect 6184 5652 6236 5704
rect 6828 5788 6880 5840
rect 7564 5763 7616 5772
rect 7564 5729 7573 5763
rect 7573 5729 7607 5763
rect 7607 5729 7616 5763
rect 7564 5720 7616 5729
rect 9404 5788 9456 5840
rect 12900 5856 12952 5908
rect 14556 5899 14608 5908
rect 14556 5865 14565 5899
rect 14565 5865 14599 5899
rect 14599 5865 14608 5899
rect 14556 5856 14608 5865
rect 7748 5652 7800 5704
rect 9496 5720 9548 5772
rect 8300 5695 8352 5704
rect 8300 5661 8309 5695
rect 8309 5661 8343 5695
rect 8343 5661 8352 5695
rect 10508 5788 10560 5840
rect 11704 5788 11756 5840
rect 16028 5831 16080 5840
rect 8300 5652 8352 5661
rect 6092 5516 6144 5568
rect 6736 5584 6788 5636
rect 8576 5584 8628 5636
rect 13360 5720 13412 5772
rect 15568 5720 15620 5772
rect 16028 5797 16037 5831
rect 16037 5797 16071 5831
rect 16071 5797 16080 5831
rect 16028 5788 16080 5797
rect 16304 5856 16356 5908
rect 17316 5856 17368 5908
rect 17776 5788 17828 5840
rect 18328 5788 18380 5840
rect 20444 5788 20496 5840
rect 16764 5763 16816 5772
rect 16764 5729 16773 5763
rect 16773 5729 16807 5763
rect 16807 5729 16816 5763
rect 16764 5720 16816 5729
rect 17132 5720 17184 5772
rect 12072 5695 12124 5704
rect 12072 5661 12081 5695
rect 12081 5661 12115 5695
rect 12115 5661 12124 5695
rect 12072 5652 12124 5661
rect 15844 5695 15896 5704
rect 6644 5516 6696 5568
rect 10416 5559 10468 5568
rect 10416 5525 10425 5559
rect 10425 5525 10459 5559
rect 10459 5525 10468 5559
rect 10416 5516 10468 5525
rect 11888 5584 11940 5636
rect 15844 5661 15853 5695
rect 15853 5661 15887 5695
rect 15887 5661 15896 5695
rect 15844 5652 15896 5661
rect 18512 5720 18564 5772
rect 19064 5763 19116 5772
rect 19064 5729 19073 5763
rect 19073 5729 19107 5763
rect 19107 5729 19116 5763
rect 19064 5720 19116 5729
rect 20168 5763 20220 5772
rect 20168 5729 20177 5763
rect 20177 5729 20211 5763
rect 20211 5729 20220 5763
rect 20168 5720 20220 5729
rect 20628 5720 20680 5772
rect 11060 5516 11112 5568
rect 14648 5584 14700 5636
rect 17776 5652 17828 5704
rect 20352 5695 20404 5704
rect 20352 5661 20361 5695
rect 20361 5661 20395 5695
rect 20395 5661 20404 5695
rect 20352 5652 20404 5661
rect 18052 5584 18104 5636
rect 13268 5516 13320 5568
rect 14096 5516 14148 5568
rect 17960 5516 18012 5568
rect 18604 5559 18656 5568
rect 18604 5525 18613 5559
rect 18613 5525 18647 5559
rect 18647 5525 18656 5559
rect 18604 5516 18656 5525
rect 19064 5516 19116 5568
rect 19800 5559 19852 5568
rect 19800 5525 19809 5559
rect 19809 5525 19843 5559
rect 19843 5525 19852 5559
rect 19800 5516 19852 5525
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 2964 5312 3016 5364
rect 7656 5312 7708 5364
rect 4160 5244 4212 5296
rect 5724 5287 5776 5296
rect 5724 5253 5733 5287
rect 5733 5253 5767 5287
rect 5767 5253 5776 5287
rect 5724 5244 5776 5253
rect 6184 5244 6236 5296
rect 6368 5244 6420 5296
rect 8300 5244 8352 5296
rect 9312 5312 9364 5364
rect 10416 5312 10468 5364
rect 2872 5219 2924 5228
rect 2872 5185 2881 5219
rect 2881 5185 2915 5219
rect 2915 5185 2924 5219
rect 2872 5176 2924 5185
rect 3056 5219 3108 5228
rect 3056 5185 3065 5219
rect 3065 5185 3099 5219
rect 3099 5185 3108 5219
rect 3056 5176 3108 5185
rect 3976 5219 4028 5228
rect 3976 5185 3985 5219
rect 3985 5185 4019 5219
rect 4019 5185 4028 5219
rect 3976 5176 4028 5185
rect 8576 5219 8628 5228
rect 1400 5151 1452 5160
rect 1400 5117 1409 5151
rect 1409 5117 1443 5151
rect 1443 5117 1452 5151
rect 1400 5108 1452 5117
rect 1860 5151 1912 5160
rect 1860 5117 1869 5151
rect 1869 5117 1903 5151
rect 1903 5117 1912 5151
rect 1860 5108 1912 5117
rect 2504 5108 2556 5160
rect 2688 5108 2740 5160
rect 2136 5040 2188 5092
rect 2964 5040 3016 5092
rect 4160 5108 4212 5160
rect 4344 5108 4396 5160
rect 5448 5108 5500 5160
rect 8576 5185 8585 5219
rect 8585 5185 8619 5219
rect 8619 5185 8628 5219
rect 8576 5176 8628 5185
rect 5816 5108 5868 5160
rect 7104 5151 7156 5160
rect 7104 5117 7113 5151
rect 7113 5117 7147 5151
rect 7147 5117 7156 5151
rect 7104 5108 7156 5117
rect 7472 5108 7524 5160
rect 8392 5108 8444 5160
rect 8668 5040 8720 5092
rect 11060 5244 11112 5296
rect 9128 5108 9180 5160
rect 10416 5108 10468 5160
rect 1584 5015 1636 5024
rect 1584 4981 1593 5015
rect 1593 4981 1627 5015
rect 1627 4981 1636 5015
rect 1584 4972 1636 4981
rect 2044 5015 2096 5024
rect 2044 4981 2053 5015
rect 2053 4981 2087 5015
rect 2087 4981 2096 5015
rect 2044 4972 2096 4981
rect 2504 4972 2556 5024
rect 3332 4972 3384 5024
rect 3792 5015 3844 5024
rect 3792 4981 3801 5015
rect 3801 4981 3835 5015
rect 3835 4981 3844 5015
rect 3792 4972 3844 4981
rect 5264 5015 5316 5024
rect 5264 4981 5273 5015
rect 5273 4981 5307 5015
rect 5307 4981 5316 5015
rect 5264 4972 5316 4981
rect 7196 4972 7248 5024
rect 8760 4972 8812 5024
rect 9956 5015 10008 5024
rect 9956 4981 9965 5015
rect 9965 4981 9999 5015
rect 9999 4981 10008 5015
rect 9956 4972 10008 4981
rect 10416 4972 10468 5024
rect 10968 5108 11020 5160
rect 13360 5312 13412 5364
rect 17684 5312 17736 5364
rect 15844 5244 15896 5296
rect 11704 5176 11756 5228
rect 11888 5219 11940 5228
rect 11888 5185 11897 5219
rect 11897 5185 11931 5219
rect 11931 5185 11940 5219
rect 11888 5176 11940 5185
rect 13912 5176 13964 5228
rect 14096 5219 14148 5228
rect 14096 5185 14105 5219
rect 14105 5185 14139 5219
rect 14139 5185 14148 5219
rect 14096 5176 14148 5185
rect 15200 5176 15252 5228
rect 21180 5312 21232 5364
rect 14188 5040 14240 5092
rect 16580 5108 16632 5160
rect 17040 5108 17092 5160
rect 17776 5151 17828 5160
rect 17776 5117 17799 5151
rect 17799 5117 17828 5151
rect 17776 5108 17828 5117
rect 18144 5108 18196 5160
rect 18512 5108 18564 5160
rect 20168 5176 20220 5228
rect 13820 4972 13872 5024
rect 14004 4972 14056 5024
rect 15384 5015 15436 5024
rect 15384 4981 15393 5015
rect 15393 4981 15427 5015
rect 15427 4981 15436 5015
rect 15384 4972 15436 4981
rect 16580 5015 16632 5024
rect 16580 4981 16589 5015
rect 16589 4981 16623 5015
rect 16623 4981 16632 5015
rect 16580 4972 16632 4981
rect 17868 4972 17920 5024
rect 18144 4972 18196 5024
rect 20352 5108 20404 5160
rect 20536 5015 20588 5024
rect 20536 4981 20545 5015
rect 20545 4981 20579 5015
rect 20579 4981 20588 5015
rect 20536 4972 20588 4981
rect 21364 5015 21416 5024
rect 21364 4981 21373 5015
rect 21373 4981 21407 5015
rect 21407 4981 21416 5015
rect 21364 4972 21416 4981
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 2504 4811 2556 4820
rect 2504 4777 2513 4811
rect 2513 4777 2547 4811
rect 2547 4777 2556 4811
rect 2504 4768 2556 4777
rect 2964 4811 3016 4820
rect 2964 4777 2973 4811
rect 2973 4777 3007 4811
rect 3007 4777 3016 4811
rect 2964 4768 3016 4777
rect 5356 4768 5408 4820
rect 6000 4768 6052 4820
rect 6460 4768 6512 4820
rect 6552 4768 6604 4820
rect 1768 4700 1820 4752
rect 2412 4700 2464 4752
rect 6184 4743 6236 4752
rect 6184 4709 6193 4743
rect 6193 4709 6227 4743
rect 6227 4709 6236 4743
rect 6184 4700 6236 4709
rect 7196 4743 7248 4752
rect 7196 4709 7205 4743
rect 7205 4709 7239 4743
rect 7239 4709 7248 4743
rect 8300 4743 8352 4752
rect 7196 4700 7248 4709
rect 8300 4709 8309 4743
rect 8309 4709 8343 4743
rect 8343 4709 8352 4743
rect 8300 4700 8352 4709
rect 9404 4768 9456 4820
rect 9956 4768 10008 4820
rect 12072 4768 12124 4820
rect 13544 4811 13596 4820
rect 13544 4777 13553 4811
rect 13553 4777 13587 4811
rect 13587 4777 13596 4811
rect 13544 4768 13596 4777
rect 9588 4700 9640 4752
rect 9680 4700 9732 4752
rect 2964 4632 3016 4684
rect 3240 4675 3292 4684
rect 3240 4641 3249 4675
rect 3249 4641 3283 4675
rect 3283 4641 3292 4675
rect 3240 4632 3292 4641
rect 3424 4632 3476 4684
rect 4068 4675 4120 4684
rect 4068 4641 4077 4675
rect 4077 4641 4111 4675
rect 4111 4641 4120 4675
rect 4068 4632 4120 4641
rect 1492 4564 1544 4616
rect 2320 4607 2372 4616
rect 2320 4573 2329 4607
rect 2329 4573 2363 4607
rect 2363 4573 2372 4607
rect 2320 4564 2372 4573
rect 3516 4496 3568 4548
rect 3976 4496 4028 4548
rect 5264 4564 5316 4616
rect 6276 4496 6328 4548
rect 6644 4564 6696 4616
rect 8576 4564 8628 4616
rect 9312 4607 9364 4616
rect 9312 4573 9321 4607
rect 9321 4573 9355 4607
rect 9355 4573 9364 4607
rect 9312 4564 9364 4573
rect 9772 4632 9824 4684
rect 14004 4700 14056 4752
rect 15384 4768 15436 4820
rect 18604 4768 18656 4820
rect 19800 4768 19852 4820
rect 7840 4496 7892 4548
rect 8484 4496 8536 4548
rect 9496 4496 9548 4548
rect 12808 4632 12860 4684
rect 13176 4632 13228 4684
rect 13636 4632 13688 4684
rect 13820 4675 13872 4684
rect 13820 4641 13829 4675
rect 13829 4641 13863 4675
rect 13863 4641 13872 4675
rect 13820 4632 13872 4641
rect 14924 4675 14976 4684
rect 14924 4641 14933 4675
rect 14933 4641 14967 4675
rect 14967 4641 14976 4675
rect 14924 4632 14976 4641
rect 15384 4675 15436 4684
rect 15384 4641 15393 4675
rect 15393 4641 15427 4675
rect 15427 4641 15436 4675
rect 15384 4632 15436 4641
rect 15844 4675 15896 4684
rect 15844 4641 15853 4675
rect 15853 4641 15887 4675
rect 15887 4641 15896 4675
rect 15844 4632 15896 4641
rect 16120 4675 16172 4684
rect 16120 4641 16154 4675
rect 16154 4641 16172 4675
rect 21364 4700 21416 4752
rect 16120 4632 16172 4641
rect 19248 4632 19300 4684
rect 11152 4564 11204 4616
rect 11704 4564 11756 4616
rect 10876 4496 10928 4548
rect 15292 4564 15344 4616
rect 18144 4607 18196 4616
rect 18144 4573 18153 4607
rect 18153 4573 18187 4607
rect 18187 4573 18196 4607
rect 18144 4564 18196 4573
rect 15200 4496 15252 4548
rect 17224 4539 17276 4548
rect 17224 4505 17233 4539
rect 17233 4505 17267 4539
rect 17267 4505 17276 4539
rect 17224 4496 17276 4505
rect 20536 4564 20588 4616
rect 21088 4539 21140 4548
rect 21088 4505 21097 4539
rect 21097 4505 21131 4539
rect 21131 4505 21140 4539
rect 21088 4496 21140 4505
rect 4068 4428 4120 4480
rect 5356 4428 5408 4480
rect 5540 4471 5592 4480
rect 5540 4437 5549 4471
rect 5549 4437 5583 4471
rect 5583 4437 5592 4471
rect 5540 4428 5592 4437
rect 5816 4471 5868 4480
rect 5816 4437 5825 4471
rect 5825 4437 5859 4471
rect 5859 4437 5868 4471
rect 5816 4428 5868 4437
rect 6000 4428 6052 4480
rect 7196 4428 7248 4480
rect 7472 4428 7524 4480
rect 8300 4428 8352 4480
rect 9864 4428 9916 4480
rect 17132 4428 17184 4480
rect 17500 4471 17552 4480
rect 17500 4437 17509 4471
rect 17509 4437 17543 4471
rect 17543 4437 17552 4471
rect 17500 4428 17552 4437
rect 19156 4428 19208 4480
rect 20444 4428 20496 4480
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 1492 4267 1544 4276
rect 1492 4233 1501 4267
rect 1501 4233 1535 4267
rect 1535 4233 1544 4267
rect 1492 4224 1544 4233
rect 2964 4224 3016 4276
rect 4068 4224 4120 4276
rect 4252 4156 4304 4208
rect 3056 4088 3108 4140
rect 1676 3952 1728 4004
rect 2872 4063 2924 4072
rect 2872 4029 2881 4063
rect 2881 4029 2915 4063
rect 2915 4029 2924 4063
rect 2872 4020 2924 4029
rect 3148 4020 3200 4072
rect 3792 4020 3844 4072
rect 6736 4156 6788 4208
rect 5448 4131 5500 4140
rect 5448 4097 5457 4131
rect 5457 4097 5491 4131
rect 5491 4097 5500 4131
rect 5448 4088 5500 4097
rect 5540 4020 5592 4072
rect 6920 4088 6972 4140
rect 7012 4020 7064 4072
rect 1860 3884 1912 3936
rect 4712 3952 4764 4004
rect 4804 3952 4856 4004
rect 3516 3927 3568 3936
rect 3516 3893 3525 3927
rect 3525 3893 3559 3927
rect 3559 3893 3568 3927
rect 3516 3884 3568 3893
rect 3608 3927 3660 3936
rect 3608 3893 3617 3927
rect 3617 3893 3651 3927
rect 3651 3893 3660 3927
rect 4896 3927 4948 3936
rect 3608 3884 3660 3893
rect 4896 3893 4905 3927
rect 4905 3893 4939 3927
rect 4939 3893 4948 3927
rect 4896 3884 4948 3893
rect 6000 3952 6052 4004
rect 6460 3952 6512 4004
rect 7104 3952 7156 4004
rect 8576 4224 8628 4276
rect 10048 4267 10100 4276
rect 10048 4233 10057 4267
rect 10057 4233 10091 4267
rect 10091 4233 10100 4267
rect 10048 4224 10100 4233
rect 10416 4224 10468 4276
rect 11980 4224 12032 4276
rect 12348 4267 12400 4276
rect 12348 4233 12357 4267
rect 12357 4233 12391 4267
rect 12391 4233 12400 4267
rect 12348 4224 12400 4233
rect 14924 4224 14976 4276
rect 19248 4224 19300 4276
rect 7472 4088 7524 4140
rect 8208 4088 8260 4140
rect 10324 4088 10376 4140
rect 8392 4020 8444 4072
rect 9312 4020 9364 4072
rect 10048 4020 10100 4072
rect 8576 3995 8628 4004
rect 8576 3961 8610 3995
rect 8610 3961 8628 3995
rect 5908 3927 5960 3936
rect 5908 3893 5917 3927
rect 5917 3893 5951 3927
rect 5951 3893 5960 3927
rect 5908 3884 5960 3893
rect 7472 3884 7524 3936
rect 8576 3952 8628 3961
rect 8760 3952 8812 4004
rect 18144 4199 18196 4208
rect 18144 4165 18153 4199
rect 18153 4165 18187 4199
rect 18187 4165 18196 4199
rect 18144 4156 18196 4165
rect 10876 4088 10928 4140
rect 12348 4088 12400 4140
rect 15292 4131 15344 4140
rect 10508 4020 10560 4072
rect 10784 4020 10836 4072
rect 10600 3952 10652 4004
rect 15292 4097 15301 4131
rect 15301 4097 15335 4131
rect 15335 4097 15344 4131
rect 15292 4088 15344 4097
rect 15476 4088 15528 4140
rect 18420 4088 18472 4140
rect 19524 4088 19576 4140
rect 21180 4088 21232 4140
rect 11244 4020 11296 4072
rect 11796 4020 11848 4072
rect 11980 4020 12032 4072
rect 12256 4020 12308 4072
rect 12716 4020 12768 4072
rect 13452 4063 13504 4072
rect 13452 4029 13461 4063
rect 13461 4029 13495 4063
rect 13495 4029 13504 4063
rect 13452 4020 13504 4029
rect 14096 4020 14148 4072
rect 7748 3884 7800 3936
rect 8392 3884 8444 3936
rect 8484 3884 8536 3936
rect 9036 3884 9088 3936
rect 9312 3884 9364 3936
rect 9864 3884 9916 3936
rect 10140 3884 10192 3936
rect 10784 3884 10836 3936
rect 11152 3884 11204 3936
rect 12992 3927 13044 3936
rect 12992 3893 13001 3927
rect 13001 3893 13035 3927
rect 13035 3893 13044 3927
rect 12992 3884 13044 3893
rect 13544 3884 13596 3936
rect 14280 3952 14332 4004
rect 16580 4020 16632 4072
rect 18052 4020 18104 4072
rect 18880 4063 18932 4072
rect 18880 4029 18889 4063
rect 18889 4029 18923 4063
rect 18923 4029 18932 4063
rect 18880 4020 18932 4029
rect 19340 4063 19392 4072
rect 19340 4029 19349 4063
rect 19349 4029 19383 4063
rect 19383 4029 19392 4063
rect 19340 4020 19392 4029
rect 20536 4020 20588 4072
rect 15292 3884 15344 3936
rect 15844 3927 15896 3936
rect 15844 3893 15853 3927
rect 15853 3893 15887 3927
rect 15887 3893 15896 3927
rect 15844 3884 15896 3893
rect 16396 3927 16448 3936
rect 16396 3893 16405 3927
rect 16405 3893 16439 3927
rect 16439 3893 16448 3927
rect 16396 3884 16448 3893
rect 16948 3952 17000 4004
rect 17040 3884 17092 3936
rect 17408 3952 17460 4004
rect 17776 3884 17828 3936
rect 19248 3884 19300 3936
rect 20076 3952 20128 4004
rect 21824 3952 21876 4004
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 1676 3723 1728 3732
rect 1676 3689 1685 3723
rect 1685 3689 1719 3723
rect 1719 3689 1728 3723
rect 1676 3680 1728 3689
rect 3516 3680 3568 3732
rect 1952 3612 2004 3664
rect 3884 3612 3936 3664
rect 2780 3587 2832 3596
rect 2780 3553 2798 3587
rect 2798 3553 2832 3587
rect 3332 3587 3384 3596
rect 2780 3544 2832 3553
rect 3332 3553 3341 3587
rect 3341 3553 3375 3587
rect 3375 3553 3384 3587
rect 3332 3544 3384 3553
rect 3700 3544 3752 3596
rect 4436 3587 4488 3596
rect 4436 3553 4445 3587
rect 4445 3553 4479 3587
rect 4479 3553 4488 3587
rect 4436 3544 4488 3553
rect 5816 3680 5868 3732
rect 6276 3680 6328 3732
rect 8392 3723 8444 3732
rect 8392 3689 8401 3723
rect 8401 3689 8435 3723
rect 8435 3689 8444 3723
rect 8392 3680 8444 3689
rect 8576 3680 8628 3732
rect 11612 3680 11664 3732
rect 5080 3612 5132 3664
rect 7012 3612 7064 3664
rect 8300 3655 8352 3664
rect 3148 3476 3200 3528
rect 4252 3476 4304 3528
rect 6644 3544 6696 3596
rect 5816 3519 5868 3528
rect 1768 3340 1820 3392
rect 3240 3408 3292 3460
rect 3516 3451 3568 3460
rect 3516 3417 3525 3451
rect 3525 3417 3559 3451
rect 3559 3417 3568 3451
rect 3516 3408 3568 3417
rect 5816 3485 5825 3519
rect 5825 3485 5859 3519
rect 5859 3485 5868 3519
rect 5816 3476 5868 3485
rect 7932 3544 7984 3596
rect 8300 3621 8309 3655
rect 8309 3621 8343 3655
rect 8343 3621 8352 3655
rect 8300 3612 8352 3621
rect 10876 3612 10928 3664
rect 11060 3612 11112 3664
rect 9404 3544 9456 3596
rect 9588 3544 9640 3596
rect 8116 3476 8168 3528
rect 9864 3476 9916 3528
rect 3148 3340 3200 3392
rect 3884 3340 3936 3392
rect 4068 3340 4120 3392
rect 4988 3340 5040 3392
rect 9496 3408 9548 3460
rect 10324 3544 10376 3596
rect 10692 3544 10744 3596
rect 10876 3476 10928 3528
rect 12164 3587 12216 3596
rect 12164 3553 12173 3587
rect 12173 3553 12207 3587
rect 12207 3553 12216 3587
rect 12164 3544 12216 3553
rect 12624 3587 12676 3596
rect 12624 3553 12633 3587
rect 12633 3553 12667 3587
rect 12667 3553 12676 3587
rect 12624 3544 12676 3553
rect 13452 3612 13504 3664
rect 15292 3612 15344 3664
rect 16120 3680 16172 3732
rect 16396 3680 16448 3732
rect 17408 3612 17460 3664
rect 18696 3680 18748 3732
rect 16672 3476 16724 3528
rect 17132 3544 17184 3596
rect 20628 3680 20680 3732
rect 19064 3612 19116 3664
rect 17960 3476 18012 3528
rect 19524 3544 19576 3596
rect 20536 3519 20588 3528
rect 8760 3383 8812 3392
rect 8760 3349 8769 3383
rect 8769 3349 8803 3383
rect 8803 3349 8812 3383
rect 8760 3340 8812 3349
rect 10048 3340 10100 3392
rect 16396 3408 16448 3460
rect 20536 3485 20545 3519
rect 20545 3485 20579 3519
rect 20579 3485 20588 3519
rect 20536 3476 20588 3485
rect 19984 3451 20036 3460
rect 12992 3340 13044 3392
rect 13084 3340 13136 3392
rect 16212 3340 16264 3392
rect 16304 3340 16356 3392
rect 16580 3340 16632 3392
rect 19984 3417 19993 3451
rect 19993 3417 20027 3451
rect 20027 3417 20036 3451
rect 19984 3408 20036 3417
rect 17960 3340 18012 3392
rect 18972 3383 19024 3392
rect 18972 3349 18981 3383
rect 18981 3349 19015 3383
rect 19015 3349 19024 3383
rect 18972 3340 19024 3349
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 1768 3179 1820 3188
rect 1768 3145 1777 3179
rect 1777 3145 1811 3179
rect 1811 3145 1820 3179
rect 1768 3136 1820 3145
rect 6644 3179 6696 3188
rect 204 3000 256 3052
rect 1676 3000 1728 3052
rect 6644 3145 6653 3179
rect 6653 3145 6687 3179
rect 6687 3145 6696 3179
rect 6644 3136 6696 3145
rect 7932 3136 7984 3188
rect 8208 3136 8260 3188
rect 8484 3136 8536 3188
rect 9404 3068 9456 3120
rect 14280 3136 14332 3188
rect 15384 3179 15436 3188
rect 15384 3145 15393 3179
rect 15393 3145 15427 3179
rect 15427 3145 15436 3179
rect 15384 3136 15436 3145
rect 15936 3136 15988 3188
rect 17868 3136 17920 3188
rect 12532 3111 12584 3120
rect 2964 2932 3016 2984
rect 3608 2932 3660 2984
rect 4712 3000 4764 3052
rect 6276 3000 6328 3052
rect 9864 3000 9916 3052
rect 10600 3043 10652 3052
rect 10600 3009 10609 3043
rect 10609 3009 10643 3043
rect 10643 3009 10652 3043
rect 10600 3000 10652 3009
rect 10876 3000 10928 3052
rect 4252 2932 4304 2984
rect 4620 2932 4672 2984
rect 5172 2932 5224 2984
rect 5816 2975 5868 2984
rect 5816 2941 5825 2975
rect 5825 2941 5859 2975
rect 5859 2941 5868 2975
rect 5816 2932 5868 2941
rect 6736 2932 6788 2984
rect 1860 2864 1912 2916
rect 2872 2864 2924 2916
rect 3240 2864 3292 2916
rect 2780 2839 2832 2848
rect 2780 2805 2789 2839
rect 2789 2805 2823 2839
rect 2823 2805 2832 2839
rect 2780 2796 2832 2805
rect 4252 2796 4304 2848
rect 5448 2864 5500 2916
rect 6276 2864 6328 2916
rect 4712 2796 4764 2848
rect 8668 2864 8720 2916
rect 6644 2796 6696 2848
rect 6828 2796 6880 2848
rect 7748 2796 7800 2848
rect 9128 2796 9180 2848
rect 9312 2932 9364 2984
rect 9680 2975 9732 2984
rect 9680 2941 9689 2975
rect 9689 2941 9723 2975
rect 9723 2941 9732 2975
rect 9680 2932 9732 2941
rect 9772 2932 9824 2984
rect 9496 2864 9548 2916
rect 12532 3077 12541 3111
rect 12541 3077 12575 3111
rect 12575 3077 12584 3111
rect 12532 3068 12584 3077
rect 14096 3068 14148 3120
rect 15200 3068 15252 3120
rect 11704 3000 11756 3052
rect 15844 3043 15896 3052
rect 9956 2796 10008 2848
rect 10140 2839 10192 2848
rect 10140 2805 10149 2839
rect 10149 2805 10183 2839
rect 10183 2805 10192 2839
rect 10140 2796 10192 2805
rect 12900 2975 12952 2984
rect 12900 2941 12909 2975
rect 12909 2941 12943 2975
rect 12943 2941 12952 2975
rect 12900 2932 12952 2941
rect 12992 2932 13044 2984
rect 15844 3009 15853 3043
rect 15853 3009 15887 3043
rect 15887 3009 15896 3043
rect 15844 3000 15896 3009
rect 16120 3000 16172 3052
rect 16304 2932 16356 2984
rect 17224 3068 17276 3120
rect 20444 3068 20496 3120
rect 17040 3000 17092 3052
rect 18880 2932 18932 2984
rect 19156 3000 19208 3052
rect 12440 2864 12492 2916
rect 14556 2907 14608 2916
rect 14556 2873 14565 2907
rect 14565 2873 14599 2907
rect 14599 2873 14608 2907
rect 14556 2864 14608 2873
rect 13360 2839 13412 2848
rect 13360 2805 13369 2839
rect 13369 2805 13403 2839
rect 13403 2805 13412 2839
rect 13360 2796 13412 2805
rect 16212 2864 16264 2916
rect 19064 2907 19116 2916
rect 19064 2873 19073 2907
rect 19073 2873 19107 2907
rect 19107 2873 19116 2907
rect 19064 2864 19116 2873
rect 19248 2975 19300 2984
rect 19248 2941 19274 2975
rect 19274 2941 19300 2975
rect 19248 2932 19300 2941
rect 19524 2864 19576 2916
rect 22744 2932 22796 2984
rect 15476 2796 15528 2848
rect 20904 2796 20956 2848
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 3240 2592 3292 2644
rect 1676 2567 1728 2576
rect 1676 2533 1685 2567
rect 1685 2533 1719 2567
rect 1719 2533 1728 2567
rect 1676 2524 1728 2533
rect 2136 2524 2188 2576
rect 2412 2567 2464 2576
rect 2412 2533 2421 2567
rect 2421 2533 2455 2567
rect 2455 2533 2464 2567
rect 2412 2524 2464 2533
rect 3884 2524 3936 2576
rect 4712 2524 4764 2576
rect 4896 2524 4948 2576
rect 6736 2592 6788 2644
rect 7288 2592 7340 2644
rect 8760 2592 8812 2644
rect 9772 2592 9824 2644
rect 10048 2635 10100 2644
rect 10048 2601 10057 2635
rect 10057 2601 10091 2635
rect 10091 2601 10100 2635
rect 10048 2592 10100 2601
rect 10324 2592 10376 2644
rect 6644 2524 6696 2576
rect 2228 2499 2280 2508
rect 2228 2465 2237 2499
rect 2237 2465 2271 2499
rect 2271 2465 2280 2499
rect 2228 2456 2280 2465
rect 2688 2499 2740 2508
rect 2688 2465 2697 2499
rect 2697 2465 2731 2499
rect 2731 2465 2740 2499
rect 2688 2456 2740 2465
rect 3148 2499 3200 2508
rect 3148 2465 3157 2499
rect 3157 2465 3191 2499
rect 3191 2465 3200 2499
rect 3148 2456 3200 2465
rect 5264 2456 5316 2508
rect 5724 2499 5776 2508
rect 5724 2465 5733 2499
rect 5733 2465 5767 2499
rect 5767 2465 5776 2499
rect 5724 2456 5776 2465
rect 6092 2456 6144 2508
rect 1492 2388 1544 2440
rect 4252 2388 4304 2440
rect 4988 2431 5040 2440
rect 4988 2397 4997 2431
rect 4997 2397 5031 2431
rect 5031 2397 5040 2431
rect 4988 2388 5040 2397
rect 3700 2320 3752 2372
rect 4620 2320 4672 2372
rect 4712 2320 4764 2372
rect 7380 2456 7432 2508
rect 8576 2456 8628 2508
rect 10140 2524 10192 2576
rect 13360 2592 13412 2644
rect 12440 2524 12492 2576
rect 14096 2567 14148 2576
rect 14096 2533 14105 2567
rect 14105 2533 14139 2567
rect 14139 2533 14148 2567
rect 14096 2524 14148 2533
rect 17776 2592 17828 2644
rect 8208 2431 8260 2440
rect 8208 2397 8217 2431
rect 8217 2397 8251 2431
rect 8251 2397 8260 2431
rect 8208 2388 8260 2397
rect 9036 2320 9088 2372
rect 9864 2388 9916 2440
rect 10692 2456 10744 2508
rect 12532 2456 12584 2508
rect 15016 2499 15068 2508
rect 15016 2465 15025 2499
rect 15025 2465 15059 2499
rect 15059 2465 15068 2499
rect 15016 2456 15068 2465
rect 17500 2524 17552 2576
rect 17960 2524 18012 2576
rect 18144 2567 18196 2576
rect 18144 2533 18153 2567
rect 18153 2533 18187 2567
rect 18187 2533 18196 2567
rect 18144 2524 18196 2533
rect 19156 2524 19208 2576
rect 19248 2499 19300 2508
rect 13084 2388 13136 2440
rect 12624 2320 12676 2372
rect 12808 2363 12860 2372
rect 12808 2329 12817 2363
rect 12817 2329 12851 2363
rect 12851 2329 12860 2363
rect 12808 2320 12860 2329
rect 8484 2252 8536 2304
rect 9220 2295 9272 2304
rect 9220 2261 9229 2295
rect 9229 2261 9263 2295
rect 9263 2261 9272 2295
rect 9220 2252 9272 2261
rect 14096 2388 14148 2440
rect 17224 2388 17276 2440
rect 19248 2465 19257 2499
rect 19257 2465 19291 2499
rect 19291 2465 19300 2499
rect 19248 2456 19300 2465
rect 20260 2499 20312 2508
rect 20260 2465 20269 2499
rect 20269 2465 20303 2499
rect 20303 2465 20312 2499
rect 20260 2456 20312 2465
rect 20812 2499 20864 2508
rect 20812 2465 20821 2499
rect 20821 2465 20855 2499
rect 20855 2465 20864 2499
rect 20812 2456 20864 2465
rect 18880 2388 18932 2440
rect 20536 2431 20588 2440
rect 20536 2397 20545 2431
rect 20545 2397 20579 2431
rect 20579 2397 20588 2431
rect 20536 2388 20588 2397
rect 13268 2320 13320 2372
rect 13728 2320 13780 2372
rect 15200 2363 15252 2372
rect 15200 2329 15209 2363
rect 15209 2329 15243 2363
rect 15243 2329 15252 2363
rect 15200 2320 15252 2329
rect 17132 2320 17184 2372
rect 17316 2320 17368 2372
rect 17776 2320 17828 2372
rect 18328 2320 18380 2372
rect 22284 2320 22336 2372
rect 13452 2252 13504 2304
rect 18144 2252 18196 2304
rect 20536 2252 20588 2304
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
rect 8300 2048 8352 2100
rect 8576 2048 8628 2100
rect 13452 2048 13504 2100
rect 15016 2048 15068 2100
rect 18788 2048 18840 2100
rect 572 1980 624 2032
rect 2228 1980 2280 2032
rect 9220 1980 9272 2032
rect 16672 1980 16724 2032
rect 19156 1980 19208 2032
rect 1032 1912 1084 1964
rect 2688 1912 2740 1964
rect 13544 1912 13596 1964
rect 17960 1912 18012 1964
rect 2412 1844 2464 1896
rect 5724 1844 5776 1896
rect 12992 1844 13044 1896
rect 18052 1844 18104 1896
rect 4252 1776 4304 1828
rect 7380 1776 7432 1828
rect 9220 1776 9272 1828
rect 10692 1776 10744 1828
rect 3332 1572 3384 1624
rect 4344 1572 4396 1624
rect 3332 1436 3384 1488
rect 3884 1436 3936 1488
rect 8760 1436 8812 1488
rect 9496 1436 9548 1488
rect 15200 1436 15252 1488
rect 21364 1436 21416 1488
rect 12624 1368 12676 1420
rect 15016 1368 15068 1420
rect 17132 1368 17184 1420
rect 18604 1368 18656 1420
rect 15568 1300 15620 1352
rect 18788 1300 18840 1352
rect 2872 1164 2924 1216
rect 4068 1164 4120 1216
<< metal2 >>
rect 4158 22672 4214 22681
rect 4158 22607 4214 22616
rect 4066 22264 4122 22273
rect 4066 22199 4122 22208
rect 3238 21720 3294 21729
rect 3238 21655 3294 21664
rect 2778 21312 2834 21321
rect 2778 21247 2834 21256
rect 2226 20768 2282 20777
rect 2226 20703 2282 20712
rect 2240 20602 2268 20703
rect 2228 20596 2280 20602
rect 2228 20538 2280 20544
rect 2792 20534 2820 21247
rect 3252 20534 3280 21655
rect 4080 20534 4108 22199
rect 2780 20528 2832 20534
rect 2780 20470 2832 20476
rect 3240 20528 3292 20534
rect 3240 20470 3292 20476
rect 4068 20528 4120 20534
rect 4068 20470 4120 20476
rect 4172 20398 4200 22607
rect 5722 22200 5778 23000
rect 17222 22200 17278 23000
rect 20258 22672 20314 22681
rect 20258 22607 20314 22616
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 5736 20398 5764 22200
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 17236 20534 17264 22200
rect 18602 21720 18658 21729
rect 18602 21655 18658 21664
rect 18282 20700 18578 20720
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 18616 20534 18644 21655
rect 18970 21312 19026 21321
rect 18970 21247 19026 21256
rect 18984 20534 19012 21247
rect 19522 20768 19578 20777
rect 19522 20703 19578 20712
rect 19536 20534 19564 20703
rect 17224 20528 17276 20534
rect 17224 20470 17276 20476
rect 18604 20528 18656 20534
rect 18604 20470 18656 20476
rect 18972 20528 19024 20534
rect 18972 20470 19024 20476
rect 19524 20528 19576 20534
rect 19524 20470 19576 20476
rect 20272 20398 20300 22607
rect 20534 22264 20590 22273
rect 20534 22199 20590 22208
rect 1584 20392 1636 20398
rect 1582 20360 1584 20369
rect 2596 20392 2648 20398
rect 1636 20360 1638 20369
rect 2596 20334 2648 20340
rect 4160 20392 4212 20398
rect 4160 20334 4212 20340
rect 5724 20392 5776 20398
rect 5724 20334 5776 20340
rect 19708 20392 19760 20398
rect 20260 20392 20312 20398
rect 19708 20334 19760 20340
rect 20180 20340 20260 20346
rect 20180 20334 20312 20340
rect 1582 20295 1638 20304
rect 2320 20324 2372 20330
rect 2320 20266 2372 20272
rect 2332 20058 2360 20266
rect 2320 20052 2372 20058
rect 2320 19994 2372 20000
rect 1768 19916 1820 19922
rect 1768 19858 1820 19864
rect 1582 19816 1638 19825
rect 1582 19751 1584 19760
rect 1636 19751 1638 19760
rect 1584 19722 1636 19728
rect 1780 19514 1808 19858
rect 2608 19514 2636 20334
rect 2872 20324 2924 20330
rect 2872 20266 2924 20272
rect 2964 20324 3016 20330
rect 2964 20266 3016 20272
rect 4252 20324 4304 20330
rect 4252 20266 4304 20272
rect 9680 20324 9732 20330
rect 9680 20266 9732 20272
rect 18788 20324 18840 20330
rect 18788 20266 18840 20272
rect 19340 20324 19392 20330
rect 19340 20266 19392 20272
rect 1768 19508 1820 19514
rect 1768 19450 1820 19456
rect 2596 19508 2648 19514
rect 2596 19450 2648 19456
rect 1582 19408 1638 19417
rect 1582 19343 1638 19352
rect 1596 19310 1624 19343
rect 1584 19304 1636 19310
rect 1584 19246 1636 19252
rect 1768 19236 1820 19242
rect 1768 19178 1820 19184
rect 1780 18970 1808 19178
rect 2884 18970 2912 20266
rect 2976 20058 3004 20266
rect 4264 20058 4292 20266
rect 4988 20256 5040 20262
rect 4988 20198 5040 20204
rect 5908 20256 5960 20262
rect 5908 20198 5960 20204
rect 8208 20256 8260 20262
rect 8208 20198 8260 20204
rect 2964 20052 3016 20058
rect 2964 19994 3016 20000
rect 4252 20052 4304 20058
rect 4252 19994 4304 20000
rect 4160 19916 4212 19922
rect 4160 19858 4212 19864
rect 4344 19916 4396 19922
rect 4344 19858 4396 19864
rect 3056 19848 3108 19854
rect 3056 19790 3108 19796
rect 3068 18970 3096 19790
rect 4172 19514 4200 19858
rect 4160 19508 4212 19514
rect 4160 19450 4212 19456
rect 3884 19304 3936 19310
rect 3936 19252 4200 19258
rect 3884 19246 4200 19252
rect 3896 19230 4200 19246
rect 1768 18964 1820 18970
rect 1768 18906 1820 18912
rect 2872 18964 2924 18970
rect 2872 18906 2924 18912
rect 3056 18964 3108 18970
rect 3056 18906 3108 18912
rect 1582 18864 1638 18873
rect 4172 18834 4200 19230
rect 4252 19236 4304 19242
rect 4252 19178 4304 19184
rect 1582 18799 1584 18808
rect 1636 18799 1638 18808
rect 1768 18828 1820 18834
rect 1584 18770 1636 18776
rect 1768 18770 1820 18776
rect 4160 18828 4212 18834
rect 4160 18770 4212 18776
rect 1780 18358 1808 18770
rect 3976 18624 4028 18630
rect 3976 18566 4028 18572
rect 2226 18456 2282 18465
rect 3988 18426 4016 18566
rect 2226 18391 2228 18400
rect 2280 18391 2282 18400
rect 3976 18420 4028 18426
rect 2228 18362 2280 18368
rect 3976 18362 4028 18368
rect 1768 18352 1820 18358
rect 1768 18294 1820 18300
rect 1768 18148 1820 18154
rect 1768 18090 1820 18096
rect 2320 18148 2372 18154
rect 2320 18090 2372 18096
rect 3424 18148 3476 18154
rect 3424 18090 3476 18096
rect 1676 18080 1728 18086
rect 1674 18048 1676 18057
rect 1728 18048 1730 18057
rect 1674 17983 1730 17992
rect 1676 17536 1728 17542
rect 1674 17504 1676 17513
rect 1728 17504 1730 17513
rect 1674 17439 1730 17448
rect 1780 17338 1808 18090
rect 2332 17882 2360 18090
rect 2320 17876 2372 17882
rect 2320 17818 2372 17824
rect 2596 17672 2648 17678
rect 2596 17614 2648 17620
rect 2964 17672 3016 17678
rect 2964 17614 3016 17620
rect 1768 17332 1820 17338
rect 1768 17274 1820 17280
rect 1584 17128 1636 17134
rect 1582 17096 1584 17105
rect 2320 17128 2372 17134
rect 1636 17096 1638 17105
rect 2320 17070 2372 17076
rect 1582 17031 1638 17040
rect 2044 17060 2096 17066
rect 2044 17002 2096 17008
rect 1860 16992 1912 16998
rect 1860 16934 1912 16940
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1596 16561 1624 16594
rect 1582 16552 1638 16561
rect 1582 16487 1638 16496
rect 1582 16144 1638 16153
rect 1582 16079 1584 16088
rect 1636 16079 1638 16088
rect 1584 16050 1636 16056
rect 1872 15638 1900 16934
rect 2056 16794 2084 17002
rect 2332 16794 2360 17070
rect 2044 16788 2096 16794
rect 2044 16730 2096 16736
rect 2320 16788 2372 16794
rect 2320 16730 2372 16736
rect 2608 16522 2636 17614
rect 2976 17270 3004 17614
rect 3436 17338 3464 18090
rect 3516 18080 3568 18086
rect 3516 18022 3568 18028
rect 4160 18080 4212 18086
rect 4160 18022 4212 18028
rect 3528 17882 3556 18022
rect 3516 17876 3568 17882
rect 3516 17818 3568 17824
rect 4068 17740 4120 17746
rect 4068 17682 4120 17688
rect 3424 17332 3476 17338
rect 3424 17274 3476 17280
rect 2964 17264 3016 17270
rect 2964 17206 3016 17212
rect 4080 17202 4108 17682
rect 4068 17196 4120 17202
rect 4068 17138 4120 17144
rect 2872 17060 2924 17066
rect 2872 17002 2924 17008
rect 2596 16516 2648 16522
rect 2596 16458 2648 16464
rect 2780 16448 2832 16454
rect 2780 16390 2832 16396
rect 2792 16046 2820 16390
rect 2780 16040 2832 16046
rect 2780 15982 2832 15988
rect 2320 15904 2372 15910
rect 2320 15846 2372 15852
rect 2332 15638 2360 15846
rect 1860 15632 1912 15638
rect 2136 15632 2188 15638
rect 1860 15574 1912 15580
rect 2134 15600 2136 15609
rect 2320 15632 2372 15638
rect 2188 15600 2190 15609
rect 2320 15574 2372 15580
rect 2134 15535 2190 15544
rect 1676 15360 1728 15366
rect 1676 15302 1728 15308
rect 1688 15201 1716 15302
rect 1674 15192 1730 15201
rect 1674 15127 1730 15136
rect 2596 14884 2648 14890
rect 2596 14826 2648 14832
rect 1676 14816 1728 14822
rect 1676 14758 1728 14764
rect 2504 14816 2556 14822
rect 2504 14758 2556 14764
rect 1688 14657 1716 14758
rect 1674 14648 1730 14657
rect 1674 14583 1730 14592
rect 1768 14476 1820 14482
rect 1768 14418 1820 14424
rect 1676 14272 1728 14278
rect 1674 14240 1676 14249
rect 1728 14240 1730 14249
rect 1674 14175 1730 14184
rect 1780 14006 1808 14418
rect 2516 14414 2544 14758
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 1768 14000 1820 14006
rect 1768 13942 1820 13948
rect 1584 13864 1636 13870
rect 1582 13832 1584 13841
rect 1636 13832 1638 13841
rect 1582 13767 1638 13776
rect 1768 13796 1820 13802
rect 1768 13738 1820 13744
rect 1582 13288 1638 13297
rect 1582 13223 1584 13232
rect 1636 13223 1638 13232
rect 1584 13194 1636 13200
rect 1780 12986 1808 13738
rect 2504 13728 2556 13734
rect 2504 13670 2556 13676
rect 2516 13530 2544 13670
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2136 13388 2188 13394
rect 2136 13330 2188 13336
rect 1768 12980 1820 12986
rect 1768 12922 1820 12928
rect 1398 12880 1454 12889
rect 1398 12815 1454 12824
rect 1412 12782 1440 12815
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1676 12368 1728 12374
rect 1674 12336 1676 12345
rect 1728 12336 1730 12345
rect 1674 12271 1730 12280
rect 1860 12300 1912 12306
rect 1860 12242 1912 12248
rect 1768 12096 1820 12102
rect 1768 12038 1820 12044
rect 1674 11928 1730 11937
rect 1780 11898 1808 12038
rect 1674 11863 1730 11872
rect 1768 11892 1820 11898
rect 1688 11694 1716 11863
rect 1768 11834 1820 11840
rect 1872 11830 1900 12242
rect 1860 11824 1912 11830
rect 1860 11766 1912 11772
rect 1676 11688 1728 11694
rect 1676 11630 1728 11636
rect 2044 11688 2096 11694
rect 2044 11630 2096 11636
rect 1674 11384 1730 11393
rect 1674 11319 1730 11328
rect 1688 11286 1716 11319
rect 1676 11280 1728 11286
rect 1676 11222 1728 11228
rect 1676 10532 1728 10538
rect 1676 10474 1728 10480
rect 1688 10441 1716 10474
rect 1674 10432 1730 10441
rect 1674 10367 1730 10376
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 1688 10033 1716 10066
rect 1674 10024 1730 10033
rect 1674 9959 1730 9968
rect 2056 9722 2084 11630
rect 2148 10810 2176 13330
rect 2608 12986 2636 14826
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 2884 12442 2912 17002
rect 2964 16720 3016 16726
rect 2964 16662 3016 16668
rect 2976 16250 3004 16662
rect 4172 16658 4200 18022
rect 4264 17270 4292 19178
rect 4356 19174 4384 19858
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 4528 19304 4580 19310
rect 4528 19246 4580 19252
rect 4344 19168 4396 19174
rect 4344 19110 4396 19116
rect 4356 18358 4384 19110
rect 4540 18766 4568 19246
rect 4528 18760 4580 18766
rect 4528 18702 4580 18708
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4421 18448 4717 18468
rect 4344 18352 4396 18358
rect 4344 18294 4396 18300
rect 4896 18352 4948 18358
rect 4896 18294 4948 18300
rect 4620 18080 4672 18086
rect 4620 18022 4672 18028
rect 4632 17882 4660 18022
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 4344 17740 4396 17746
rect 4344 17682 4396 17688
rect 4252 17264 4304 17270
rect 4252 17206 4304 17212
rect 4160 16652 4212 16658
rect 4160 16594 4212 16600
rect 3516 16584 3568 16590
rect 3516 16526 3568 16532
rect 3608 16584 3660 16590
rect 3608 16526 3660 16532
rect 3528 16250 3556 16526
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 3516 16244 3568 16250
rect 3516 16186 3568 16192
rect 3620 16046 3648 16526
rect 4356 16130 4384 17682
rect 4908 17678 4936 18294
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 4896 17672 4948 17678
rect 4896 17614 4948 17620
rect 4421 17436 4717 17456
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 4816 17338 4844 17614
rect 4804 17332 4856 17338
rect 4804 17274 4856 17280
rect 5000 17134 5028 20198
rect 5920 19990 5948 20198
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 8220 20058 8248 20198
rect 8208 20052 8260 20058
rect 8208 19994 8260 20000
rect 5080 19984 5132 19990
rect 5080 19926 5132 19932
rect 5908 19984 5960 19990
rect 5908 19926 5960 19932
rect 5092 19310 5120 19926
rect 7656 19848 7708 19854
rect 7656 19790 7708 19796
rect 5264 19712 5316 19718
rect 5264 19654 5316 19660
rect 5080 19304 5132 19310
rect 5080 19246 5132 19252
rect 5276 18834 5304 19654
rect 5816 19168 5868 19174
rect 5816 19110 5868 19116
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 7472 19168 7524 19174
rect 7472 19110 7524 19116
rect 5080 18828 5132 18834
rect 5080 18770 5132 18776
rect 5264 18828 5316 18834
rect 5264 18770 5316 18776
rect 4988 17128 5040 17134
rect 4988 17070 5040 17076
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 4172 16102 4384 16130
rect 3608 16040 3660 16046
rect 3608 15982 3660 15988
rect 3792 15972 3844 15978
rect 3792 15914 3844 15920
rect 3056 15564 3108 15570
rect 3056 15506 3108 15512
rect 3068 14618 3096 15506
rect 3700 14884 3752 14890
rect 3700 14826 3752 14832
rect 3056 14612 3108 14618
rect 3056 14554 3108 14560
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 2964 14476 3016 14482
rect 2964 14418 3016 14424
rect 2976 14074 3004 14418
rect 2964 14068 3016 14074
rect 2964 14010 3016 14016
rect 3252 13530 3280 14554
rect 3712 13870 3740 14826
rect 3804 14618 3832 15914
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 4080 14618 4108 15438
rect 4172 15162 4200 16102
rect 4344 16040 4396 16046
rect 4344 15982 4396 15988
rect 4252 15972 4304 15978
rect 4252 15914 4304 15920
rect 4264 15706 4292 15914
rect 4252 15700 4304 15706
rect 4252 15642 4304 15648
rect 4356 15638 4384 15982
rect 4344 15632 4396 15638
rect 4344 15574 4396 15580
rect 4252 15360 4304 15366
rect 4252 15302 4304 15308
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 3792 14612 3844 14618
rect 3792 14554 3844 14560
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 4172 14498 4200 15098
rect 4080 14470 4200 14498
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 3700 13864 3752 13870
rect 3700 13806 3752 13812
rect 3884 13864 3936 13870
rect 3884 13806 3936 13812
rect 3240 13524 3292 13530
rect 3240 13466 3292 13472
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 3436 12850 3464 13126
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 2964 12708 3016 12714
rect 2964 12650 3016 12656
rect 2688 12436 2740 12442
rect 2688 12378 2740 12384
rect 2872 12436 2924 12442
rect 2872 12378 2924 12384
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2608 11626 2636 12174
rect 2596 11620 2648 11626
rect 2596 11562 2648 11568
rect 2608 11150 2636 11562
rect 2700 11558 2728 12378
rect 2688 11552 2740 11558
rect 2688 11494 2740 11500
rect 2596 11144 2648 11150
rect 2596 11086 2648 11092
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2044 9716 2096 9722
rect 2044 9658 2096 9664
rect 2056 9518 2084 9658
rect 1584 9512 1636 9518
rect 1582 9480 1584 9489
rect 2044 9512 2096 9518
rect 1636 9480 1638 9489
rect 2044 9454 2096 9460
rect 1582 9415 1638 9424
rect 1860 9444 1912 9450
rect 1860 9386 1912 9392
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1400 8832 1452 8838
rect 1400 8774 1452 8780
rect 1412 5166 1440 8774
rect 1490 8664 1546 8673
rect 1688 8634 1716 9318
rect 1872 8974 1900 9386
rect 2516 9178 2544 10066
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2688 9444 2740 9450
rect 2688 9386 2740 9392
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 1952 9104 2004 9110
rect 1952 9046 2004 9052
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 1490 8599 1546 8608
rect 1676 8628 1728 8634
rect 1504 8022 1532 8599
rect 1676 8570 1728 8576
rect 1872 8566 1900 8910
rect 1860 8560 1912 8566
rect 1860 8502 1912 8508
rect 1584 8288 1636 8294
rect 1584 8230 1636 8236
rect 1492 8016 1544 8022
rect 1492 7958 1544 7964
rect 1596 7342 1624 8230
rect 1860 7812 1912 7818
rect 1860 7754 1912 7760
rect 1584 7336 1636 7342
rect 1872 7313 1900 7754
rect 1964 7478 1992 9046
rect 2136 9036 2188 9042
rect 2136 8978 2188 8984
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 2056 8090 2084 8910
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 2148 7546 2176 8978
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 1952 7472 2004 7478
rect 1952 7414 2004 7420
rect 1584 7278 1636 7284
rect 1858 7304 1914 7313
rect 1858 7239 1914 7248
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 6225 1624 7142
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1674 6352 1730 6361
rect 1674 6287 1730 6296
rect 1582 6216 1638 6225
rect 1582 6151 1638 6160
rect 1688 5846 1716 6287
rect 1872 6254 1900 6598
rect 1964 6254 1992 7414
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 2332 6769 2360 6802
rect 2318 6760 2374 6769
rect 2318 6695 2374 6704
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 1860 6248 1912 6254
rect 1860 6190 1912 6196
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 2228 6112 2280 6118
rect 2228 6054 2280 6060
rect 1766 5944 1822 5953
rect 1766 5879 1822 5888
rect 1676 5840 1728 5846
rect 1674 5808 1676 5817
rect 1728 5808 1730 5817
rect 1674 5743 1730 5752
rect 1400 5160 1452 5166
rect 1400 5102 1452 5108
rect 1582 5128 1638 5137
rect 1412 3913 1440 5102
rect 1582 5063 1638 5072
rect 1596 5030 1624 5063
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 1780 4865 1808 5879
rect 2240 5409 2268 6054
rect 2332 5760 2360 6258
rect 2412 5772 2464 5778
rect 2332 5732 2412 5760
rect 2226 5400 2282 5409
rect 2226 5335 2282 5344
rect 1860 5160 1912 5166
rect 1860 5102 1912 5108
rect 1766 4856 1822 4865
rect 1766 4791 1822 4800
rect 1780 4758 1808 4791
rect 1768 4752 1820 4758
rect 1768 4694 1820 4700
rect 1492 4616 1544 4622
rect 1492 4558 1544 4564
rect 1504 4282 1532 4558
rect 1872 4457 1900 5102
rect 2136 5092 2188 5098
rect 2136 5034 2188 5040
rect 2044 5024 2096 5030
rect 2044 4966 2096 4972
rect 2056 4729 2084 4966
rect 2042 4720 2098 4729
rect 2042 4655 2098 4664
rect 1858 4448 1914 4457
rect 1858 4383 1914 4392
rect 1492 4276 1544 4282
rect 1492 4218 1544 4224
rect 1676 4004 1728 4010
rect 1676 3946 1728 3952
rect 1398 3904 1454 3913
rect 1398 3839 1454 3848
rect 1688 3738 1716 3946
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 1780 3194 1808 3334
rect 1768 3188 1820 3194
rect 1768 3130 1820 3136
rect 204 3052 256 3058
rect 204 2994 256 3000
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 216 800 244 2994
rect 1688 2582 1716 2994
rect 1872 2922 1900 3878
rect 1952 3664 2004 3670
rect 1952 3606 2004 3612
rect 1860 2916 1912 2922
rect 1860 2858 1912 2864
rect 1676 2576 1728 2582
rect 1676 2518 1728 2524
rect 1492 2440 1544 2446
rect 1492 2382 1544 2388
rect 572 2032 624 2038
rect 572 1974 624 1980
rect 584 800 612 1974
rect 1032 1964 1084 1970
rect 1032 1906 1084 1912
rect 1044 800 1072 1906
rect 1504 800 1532 2382
rect 1872 1057 1900 2858
rect 1858 1048 1914 1057
rect 1858 983 1914 992
rect 1964 800 1992 3606
rect 2148 2582 2176 5034
rect 2332 4622 2360 5732
rect 2412 5714 2464 5720
rect 2516 5166 2544 8774
rect 2700 6100 2728 9386
rect 2792 9178 2820 9998
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 2884 7954 2912 12378
rect 2976 10810 3004 12650
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 3068 12374 3096 12582
rect 3528 12442 3556 13466
rect 3712 12850 3740 13806
rect 3896 13530 3924 13806
rect 3884 13524 3936 13530
rect 3884 13466 3936 13472
rect 3700 12844 3752 12850
rect 3700 12786 3752 12792
rect 3516 12436 3568 12442
rect 3252 12406 3516 12434
rect 3056 12368 3108 12374
rect 3056 12310 3108 12316
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 3068 10266 3096 10542
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2872 7948 2924 7954
rect 2872 7890 2924 7896
rect 2778 7032 2834 7041
rect 2778 6967 2780 6976
rect 2832 6967 2834 6976
rect 2780 6938 2832 6944
rect 2700 6072 2912 6100
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 2792 5778 2820 5850
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 2504 5160 2556 5166
rect 2504 5102 2556 5108
rect 2688 5160 2740 5166
rect 2688 5102 2740 5108
rect 2504 5024 2556 5030
rect 2504 4966 2556 4972
rect 2516 4826 2544 4966
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2412 4752 2464 4758
rect 2412 4694 2464 4700
rect 2320 4616 2372 4622
rect 2320 4558 2372 4564
rect 2424 2582 2452 4694
rect 2136 2576 2188 2582
rect 2136 2518 2188 2524
rect 2412 2576 2464 2582
rect 2412 2518 2464 2524
rect 2700 2514 2728 5102
rect 2792 4060 2820 5714
rect 2884 5234 2912 6072
rect 2976 5370 3004 8910
rect 3056 8356 3108 8362
rect 3056 8298 3108 8304
rect 3068 7886 3096 8298
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 3068 7410 3096 7822
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 3160 6866 3188 9318
rect 3252 8265 3280 12406
rect 3516 12378 3568 12384
rect 3516 12300 3568 12306
rect 3516 12242 3568 12248
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3436 11694 3464 12038
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 3528 11558 3556 12242
rect 3712 11898 3740 12786
rect 3988 11898 4016 14350
rect 4080 13954 4108 14470
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 4172 14074 4200 14350
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4080 13926 4200 13954
rect 4172 13462 4200 13926
rect 4160 13456 4212 13462
rect 4160 13398 4212 13404
rect 4264 13394 4292 15302
rect 4356 15026 4384 15574
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 4344 15020 4396 15026
rect 4344 14962 4396 14968
rect 4344 14476 4396 14482
rect 4344 14418 4396 14424
rect 4252 13388 4304 13394
rect 4252 13330 4304 13336
rect 4160 13252 4212 13258
rect 4160 13194 4212 13200
rect 4172 12374 4200 13194
rect 4356 12986 4384 14418
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 4620 13728 4672 13734
rect 4620 13670 4672 13676
rect 4632 13530 4660 13670
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 4160 12368 4212 12374
rect 4160 12310 4212 12316
rect 4448 12306 4476 12718
rect 5000 12646 5028 17070
rect 5092 13870 5120 18770
rect 5276 18290 5304 18770
rect 5356 18624 5408 18630
rect 5356 18566 5408 18572
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 5172 18080 5224 18086
rect 5172 18022 5224 18028
rect 5184 17814 5212 18022
rect 5172 17808 5224 17814
rect 5172 17750 5224 17756
rect 5368 17678 5396 18566
rect 5356 17672 5408 17678
rect 5356 17614 5408 17620
rect 5264 16448 5316 16454
rect 5264 16390 5316 16396
rect 5172 15564 5224 15570
rect 5172 15506 5224 15512
rect 5184 14414 5212 15506
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 5172 13932 5224 13938
rect 5172 13874 5224 13880
rect 5080 13864 5132 13870
rect 5080 13806 5132 13812
rect 5080 13456 5132 13462
rect 5080 13398 5132 13404
rect 4528 12640 4580 12646
rect 4528 12582 4580 12588
rect 4988 12640 5040 12646
rect 4988 12582 5040 12588
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 4448 12209 4476 12242
rect 4434 12200 4490 12209
rect 4344 12164 4396 12170
rect 4540 12186 4568 12582
rect 4804 12436 4856 12442
rect 4856 12396 4936 12424
rect 4804 12378 4856 12384
rect 4540 12170 4660 12186
rect 4540 12164 4672 12170
rect 4540 12158 4620 12164
rect 4434 12135 4490 12144
rect 4344 12106 4396 12112
rect 4620 12106 4672 12112
rect 4804 12164 4856 12170
rect 4804 12106 4856 12112
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 3700 11892 3752 11898
rect 3700 11834 3752 11840
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 4080 11801 4108 12038
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 3698 11792 3754 11801
rect 3698 11727 3754 11736
rect 4066 11792 4122 11801
rect 4066 11727 4122 11736
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3330 10976 3386 10985
rect 3330 10911 3386 10920
rect 3344 10130 3372 10911
rect 3332 10124 3384 10130
rect 3332 10066 3384 10072
rect 3424 9988 3476 9994
rect 3424 9930 3476 9936
rect 3436 9654 3464 9930
rect 3424 9648 3476 9654
rect 3424 9590 3476 9596
rect 3436 9110 3464 9590
rect 3424 9104 3476 9110
rect 3424 9046 3476 9052
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3436 8294 3464 8910
rect 3424 8288 3476 8294
rect 3238 8256 3294 8265
rect 3424 8230 3476 8236
rect 3238 8191 3294 8200
rect 3422 7984 3478 7993
rect 3240 7948 3292 7954
rect 3422 7919 3478 7928
rect 3240 7890 3292 7896
rect 3148 6860 3200 6866
rect 3148 6802 3200 6808
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 3068 6322 3096 6734
rect 3252 6458 3280 7890
rect 3332 7744 3384 7750
rect 3436 7721 3464 7919
rect 3332 7686 3384 7692
rect 3422 7712 3478 7721
rect 3344 7177 3372 7686
rect 3422 7647 3478 7656
rect 3436 7274 3464 7647
rect 3424 7268 3476 7274
rect 3424 7210 3476 7216
rect 3330 7168 3386 7177
rect 3528 7154 3556 11494
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 3620 10266 3648 10542
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 3712 9178 3740 11727
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 3884 11280 3936 11286
rect 3884 11222 3936 11228
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 3700 9172 3752 9178
rect 3700 9114 3752 9120
rect 3608 9036 3660 9042
rect 3608 8978 3660 8984
rect 3620 8634 3648 8978
rect 3804 8838 3832 10950
rect 3896 10606 3924 11222
rect 4172 11218 4200 11630
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3896 9722 3924 10542
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3896 8974 3924 9658
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3884 8968 3936 8974
rect 3884 8910 3936 8916
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 3608 8424 3660 8430
rect 3608 8366 3660 8372
rect 3330 7103 3386 7112
rect 3436 7126 3556 7154
rect 3344 7002 3372 7103
rect 3332 6996 3384 7002
rect 3332 6938 3384 6944
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3436 6338 3464 7126
rect 3516 6928 3568 6934
rect 3516 6870 3568 6876
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 3160 6310 3464 6338
rect 3528 6322 3556 6870
rect 3516 6316 3568 6322
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 3068 5234 3096 6258
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 2964 5092 3016 5098
rect 2964 5034 3016 5040
rect 2976 4826 3004 5034
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 2976 4282 3004 4626
rect 2964 4276 3016 4282
rect 2964 4218 3016 4224
rect 3068 4146 3096 5170
rect 3160 4570 3188 6310
rect 3516 6258 3568 6264
rect 3516 6180 3568 6186
rect 3516 6122 3568 6128
rect 3238 5264 3294 5273
rect 3238 5199 3294 5208
rect 3252 4690 3280 5199
rect 3332 5024 3384 5030
rect 3332 4966 3384 4972
rect 3240 4684 3292 4690
rect 3240 4626 3292 4632
rect 3160 4542 3280 4570
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 2872 4072 2924 4078
rect 2792 4032 2872 4060
rect 2872 4014 2924 4020
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 2792 2854 2820 3538
rect 3160 3534 3188 4014
rect 3148 3528 3200 3534
rect 2870 3496 2926 3505
rect 3148 3470 3200 3476
rect 3252 3466 3280 4542
rect 3344 3602 3372 4966
rect 3424 4684 3476 4690
rect 3424 4626 3476 4632
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 2870 3431 2926 3440
rect 3240 3460 3292 3466
rect 2884 2922 2912 3431
rect 3240 3402 3292 3408
rect 3148 3392 3200 3398
rect 3148 3334 3200 3340
rect 2962 3088 3018 3097
rect 2962 3023 3018 3032
rect 2976 2990 3004 3023
rect 2964 2984 3016 2990
rect 2964 2926 3016 2932
rect 2872 2916 2924 2922
rect 2872 2858 2924 2864
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 3160 2514 3188 3334
rect 3240 2916 3292 2922
rect 3240 2858 3292 2864
rect 3252 2650 3280 2858
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 2228 2508 2280 2514
rect 2228 2450 2280 2456
rect 2688 2508 2740 2514
rect 2688 2450 2740 2456
rect 3148 2508 3200 2514
rect 3148 2450 3200 2456
rect 2240 2038 2268 2450
rect 2228 2032 2280 2038
rect 2228 1974 2280 1980
rect 2700 1970 2728 2450
rect 2688 1964 2740 1970
rect 2688 1906 2740 1912
rect 2412 1896 2464 1902
rect 2412 1838 2464 1844
rect 2424 800 2452 1838
rect 3332 1624 3384 1630
rect 3330 1592 3332 1601
rect 3384 1592 3386 1601
rect 3330 1527 3386 1536
rect 3332 1488 3384 1494
rect 3332 1430 3384 1436
rect 2872 1216 2924 1222
rect 2872 1158 2924 1164
rect 2884 800 2912 1158
rect 3344 800 3372 1430
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1490 0 1546 800
rect 1950 0 2006 800
rect 2410 0 2466 800
rect 2870 0 2926 800
rect 3330 0 3386 800
rect 3436 241 3464 4626
rect 3528 4554 3556 6122
rect 3516 4548 3568 4554
rect 3516 4490 3568 4496
rect 3620 4457 3648 8366
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3698 7848 3754 7857
rect 3698 7783 3754 7792
rect 3712 7546 3740 7783
rect 3700 7540 3752 7546
rect 3700 7482 3752 7488
rect 3700 7404 3752 7410
rect 3700 7346 3752 7352
rect 3712 7002 3740 7346
rect 3700 6996 3752 7002
rect 3700 6938 3752 6944
rect 3804 6798 3832 8230
rect 3896 7410 3924 8230
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3884 7200 3936 7206
rect 3884 7142 3936 7148
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3606 4448 3662 4457
rect 3606 4383 3662 4392
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 3608 3936 3660 3942
rect 3608 3878 3660 3884
rect 3528 3738 3556 3878
rect 3516 3732 3568 3738
rect 3516 3674 3568 3680
rect 3514 3496 3570 3505
rect 3514 3431 3516 3440
rect 3568 3431 3570 3440
rect 3516 3402 3568 3408
rect 3620 2990 3648 3878
rect 3712 3602 3740 6598
rect 3804 5778 3832 6734
rect 3792 5772 3844 5778
rect 3792 5714 3844 5720
rect 3790 5400 3846 5409
rect 3790 5335 3846 5344
rect 3804 5030 3832 5335
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 3700 3596 3752 3602
rect 3700 3538 3752 3544
rect 3608 2984 3660 2990
rect 3608 2926 3660 2932
rect 3700 2372 3752 2378
rect 3700 2314 3752 2320
rect 3712 2009 3740 2314
rect 3698 2000 3754 2009
rect 3698 1935 3754 1944
rect 3804 800 3832 4014
rect 3896 3670 3924 7142
rect 3988 5930 4016 9454
rect 4066 9072 4122 9081
rect 4066 9007 4122 9016
rect 4080 8566 4108 9007
rect 4068 8560 4120 8566
rect 4068 8502 4120 8508
rect 4066 8120 4122 8129
rect 4066 8055 4122 8064
rect 4080 8022 4108 8055
rect 4068 8016 4120 8022
rect 4068 7958 4120 7964
rect 4172 7886 4200 11154
rect 4264 11150 4292 11834
rect 4356 11642 4384 12106
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 4356 11614 4476 11642
rect 4448 11558 4476 11614
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4436 11552 4488 11558
rect 4436 11494 4488 11500
rect 4356 11354 4384 11494
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 4080 6338 4108 6938
rect 4172 6458 4200 7822
rect 4264 6662 4292 11086
rect 4421 10908 4717 10928
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 4344 9444 4396 9450
rect 4344 9386 4396 9392
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 4080 6310 4200 6338
rect 3988 5902 4108 5930
rect 3976 5840 4028 5846
rect 3976 5782 4028 5788
rect 3988 5234 4016 5782
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 4080 4690 4108 5902
rect 4172 5302 4200 6310
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4160 5296 4212 5302
rect 4160 5238 4212 5244
rect 4160 5160 4212 5166
rect 4160 5102 4212 5108
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 3976 4548 4028 4554
rect 3976 4490 4028 4496
rect 3884 3664 3936 3670
rect 3884 3606 3936 3612
rect 3896 3398 3924 3606
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3884 2576 3936 2582
rect 3988 2553 4016 4490
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 4080 4282 4108 4422
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 3884 2518 3936 2524
rect 3974 2544 4030 2553
rect 3896 1494 3924 2518
rect 3974 2479 4030 2488
rect 3884 1488 3936 1494
rect 3884 1430 3936 1436
rect 4080 1222 4108 3334
rect 4068 1216 4120 1222
rect 4068 1158 4120 1164
rect 3422 232 3478 241
rect 3422 167 3478 176
rect 3790 0 3846 800
rect 4066 640 4122 649
rect 4172 626 4200 5102
rect 4264 5012 4292 6258
rect 4356 5166 4384 9386
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4421 8656 4717 8676
rect 4816 8616 4844 12106
rect 4908 11830 4936 12396
rect 4896 11824 4948 11830
rect 4896 11766 4948 11772
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 4908 9382 4936 10746
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4540 8588 4844 8616
rect 4540 8294 4568 8588
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4632 8401 4660 8434
rect 4618 8392 4674 8401
rect 4908 8378 4936 9318
rect 5000 8498 5028 12582
rect 5092 11558 5120 13398
rect 5184 13258 5212 13874
rect 5276 13530 5304 16390
rect 5368 15638 5396 17614
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5632 16992 5684 16998
rect 5632 16934 5684 16940
rect 5460 16794 5488 16934
rect 5448 16788 5500 16794
rect 5448 16730 5500 16736
rect 5644 16726 5672 16934
rect 5632 16720 5684 16726
rect 5632 16662 5684 16668
rect 5724 16040 5776 16046
rect 5724 15982 5776 15988
rect 5356 15632 5408 15638
rect 5356 15574 5408 15580
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 5460 14550 5488 15438
rect 5736 14618 5764 15982
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 5448 14544 5500 14550
rect 5448 14486 5500 14492
rect 5356 13796 5408 13802
rect 5356 13738 5408 13744
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 5172 13252 5224 13258
rect 5172 13194 5224 13200
rect 5184 12850 5212 13194
rect 5276 12986 5304 13466
rect 5368 13462 5396 13738
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5356 13456 5408 13462
rect 5356 13398 5408 13404
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 5172 12844 5224 12850
rect 5172 12786 5224 12792
rect 5276 12322 5304 12922
rect 5368 12782 5396 13398
rect 5552 13190 5580 13670
rect 5540 13184 5592 13190
rect 5540 13126 5592 13132
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5184 12294 5304 12322
rect 5184 11762 5212 12294
rect 5264 12232 5316 12238
rect 5460 12220 5488 12786
rect 5316 12192 5488 12220
rect 5264 12174 5316 12180
rect 5172 11756 5224 11762
rect 5172 11698 5224 11704
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5184 10810 5212 11698
rect 5276 11354 5304 12174
rect 5828 11762 5856 19110
rect 6552 18964 6604 18970
rect 6552 18906 6604 18912
rect 6564 17814 6592 18906
rect 7300 18902 7328 19110
rect 7288 18896 7340 18902
rect 7288 18838 7340 18844
rect 7484 18426 7512 19110
rect 7564 18624 7616 18630
rect 7564 18566 7616 18572
rect 7472 18420 7524 18426
rect 7472 18362 7524 18368
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6840 17882 6868 18158
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 6000 17808 6052 17814
rect 6000 17750 6052 17756
rect 6552 17808 6604 17814
rect 6552 17750 6604 17756
rect 5908 17060 5960 17066
rect 5908 17002 5960 17008
rect 5920 16726 5948 17002
rect 5908 16720 5960 16726
rect 5908 16662 5960 16668
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 5356 9376 5408 9382
rect 5356 9318 5408 9324
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 4908 8350 5028 8378
rect 4618 8327 4674 8336
rect 4528 8288 4580 8294
rect 4528 8230 4580 8236
rect 4528 7812 4580 7818
rect 4632 7800 4660 8327
rect 5000 8294 5028 8350
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4580 7772 4660 7800
rect 4528 7754 4580 7760
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 4436 7404 4488 7410
rect 4436 7346 4488 7352
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 4448 6934 4476 7346
rect 4724 7154 4752 7346
rect 4816 7342 4844 7822
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4908 7154 4936 8230
rect 4988 7948 5040 7954
rect 4988 7890 5040 7896
rect 5000 7206 5028 7890
rect 4724 7126 4936 7154
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 4436 6928 4488 6934
rect 4436 6870 4488 6876
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 4816 6390 4844 6598
rect 4804 6384 4856 6390
rect 4804 6326 4856 6332
rect 4436 6112 4488 6118
rect 4488 6072 4844 6100
rect 4436 6054 4488 6060
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 4344 5160 4396 5166
rect 4344 5102 4396 5108
rect 4264 4984 4384 5012
rect 4250 4584 4306 4593
rect 4250 4519 4306 4528
rect 4264 4214 4292 4519
rect 4252 4208 4304 4214
rect 4252 4150 4304 4156
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4264 2990 4292 3470
rect 4252 2984 4304 2990
rect 4250 2952 4252 2961
rect 4304 2952 4306 2961
rect 4250 2887 4306 2896
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 4264 2446 4292 2790
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 4252 1828 4304 1834
rect 4252 1770 4304 1776
rect 4264 800 4292 1770
rect 4356 1630 4384 4984
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 4816 4321 4844 6072
rect 4802 4312 4858 4321
rect 4802 4247 4858 4256
rect 5092 4196 5120 9318
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5276 7546 5304 7822
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5368 6322 5396 9318
rect 5460 8498 5488 11494
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5736 10810 5764 11154
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5736 10062 5764 10746
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5828 9042 5856 9318
rect 5816 9036 5868 9042
rect 5816 8978 5868 8984
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5736 7993 5764 8366
rect 5722 7984 5778 7993
rect 5722 7919 5778 7928
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5460 6186 5488 7482
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5172 6180 5224 6186
rect 5172 6122 5224 6128
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 4434 4176 4490 4185
rect 4434 4111 4490 4120
rect 4724 4168 5120 4196
rect 4448 3602 4476 4111
rect 4724 4010 4752 4168
rect 4712 4004 4764 4010
rect 4712 3946 4764 3952
rect 4804 4004 4856 4010
rect 4804 3946 4856 3952
rect 4436 3596 4488 3602
rect 4436 3538 4488 3544
rect 4421 3292 4717 3312
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 4421 3216 4717 3236
rect 4712 3052 4764 3058
rect 4712 2994 4764 3000
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 4632 2378 4660 2926
rect 4724 2854 4752 2994
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 4724 2378 4752 2518
rect 4620 2372 4672 2378
rect 4620 2314 4672 2320
rect 4712 2372 4764 2378
rect 4712 2314 4764 2320
rect 4421 2204 4717 2224
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4421 2128 4717 2148
rect 4344 1624 4396 1630
rect 4344 1566 4396 1572
rect 4816 1442 4844 3946
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4908 2582 4936 3878
rect 5080 3664 5132 3670
rect 5080 3606 5132 3612
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 4896 2576 4948 2582
rect 4896 2518 4948 2524
rect 5000 2446 5028 3334
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 4724 1414 4844 1442
rect 4724 800 4752 1414
rect 5092 800 5120 3606
rect 5184 2990 5212 6122
rect 5552 5914 5580 7346
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5644 5794 5672 7822
rect 5724 7812 5776 7818
rect 5724 7754 5776 7760
rect 5736 7002 5764 7754
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 5736 6662 5764 6938
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5736 6322 5764 6598
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5736 5914 5764 6054
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 5460 5766 5672 5794
rect 5262 5400 5318 5409
rect 5262 5335 5318 5344
rect 5276 5030 5304 5335
rect 5460 5166 5488 5766
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 5552 4865 5580 5646
rect 5262 4856 5318 4865
rect 5538 4856 5594 4865
rect 5262 4791 5318 4800
rect 5356 4820 5408 4826
rect 5276 4622 5304 4791
rect 5538 4791 5594 4800
rect 5356 4762 5408 4768
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 5276 2514 5304 4558
rect 5368 4486 5396 4762
rect 5356 4480 5408 4486
rect 5356 4422 5408 4428
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5460 3369 5488 4082
rect 5552 4078 5580 4422
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5644 3584 5672 5766
rect 5722 5536 5778 5545
rect 5722 5471 5778 5480
rect 5736 5302 5764 5471
rect 5724 5296 5776 5302
rect 5724 5238 5776 5244
rect 5828 5166 5856 7890
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 5828 4570 5856 5102
rect 5736 4542 5856 4570
rect 5736 3618 5764 4542
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5828 3738 5856 4422
rect 5920 3942 5948 16662
rect 6012 16590 6040 17750
rect 6564 16794 6592 17750
rect 6920 17740 6972 17746
rect 6920 17682 6972 17688
rect 6932 17338 6960 17682
rect 7012 17536 7064 17542
rect 7012 17478 7064 17484
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 7024 17202 7052 17478
rect 7012 17196 7064 17202
rect 7012 17138 7064 17144
rect 7104 16992 7156 16998
rect 7104 16934 7156 16940
rect 6552 16788 6604 16794
rect 6552 16730 6604 16736
rect 6000 16584 6052 16590
rect 6000 16526 6052 16532
rect 6012 16250 6040 16526
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 6276 16040 6328 16046
rect 6276 15982 6328 15988
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 6104 13530 6132 14418
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6288 12442 6316 15982
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 6564 14958 6592 15302
rect 7116 15162 7144 16934
rect 7288 16176 7340 16182
rect 7340 16136 7420 16164
rect 7288 16118 7340 16124
rect 7288 15564 7340 15570
rect 7288 15506 7340 15512
rect 7104 15156 7156 15162
rect 7104 15098 7156 15104
rect 6552 14952 6604 14958
rect 6552 14894 6604 14900
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6472 14346 6500 14758
rect 6564 14414 6592 14894
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 6552 14408 6604 14414
rect 6552 14350 6604 14356
rect 6460 14340 6512 14346
rect 6460 14282 6512 14288
rect 6472 13326 6500 14282
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 7024 12442 7052 13330
rect 7116 12986 7144 14418
rect 7300 14414 7328 15506
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7208 14074 7236 14350
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7102 12744 7158 12753
rect 7102 12679 7104 12688
rect 7156 12679 7158 12688
rect 7104 12650 7156 12656
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 6012 9178 6040 12242
rect 6288 11354 6316 12378
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 7024 11898 7052 12038
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 7024 11286 7052 11834
rect 7208 11558 7236 13330
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7300 12102 7328 13262
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 6092 10804 6144 10810
rect 6092 10746 6144 10752
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 6012 4826 6040 9114
rect 6104 7206 6132 10746
rect 6276 10668 6328 10674
rect 6276 10610 6328 10616
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6196 7342 6224 10406
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 6104 7041 6132 7142
rect 6090 7032 6146 7041
rect 6090 6967 6146 6976
rect 6196 5710 6224 7278
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 6012 4010 6040 4422
rect 6000 4004 6052 4010
rect 6000 3946 6052 3952
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 5736 3590 6040 3618
rect 5552 3556 5672 3584
rect 5446 3360 5502 3369
rect 5446 3295 5502 3304
rect 5460 2922 5488 3295
rect 5448 2916 5500 2922
rect 5448 2858 5500 2864
rect 5264 2508 5316 2514
rect 5264 2450 5316 2456
rect 5552 800 5580 3556
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 5828 3369 5856 3470
rect 5814 3360 5870 3369
rect 5814 3295 5870 3304
rect 5816 2984 5868 2990
rect 5814 2952 5816 2961
rect 5868 2952 5870 2961
rect 5814 2887 5870 2896
rect 5724 2508 5776 2514
rect 5724 2450 5776 2456
rect 5736 1902 5764 2450
rect 5724 1896 5776 1902
rect 5724 1838 5776 1844
rect 6012 800 6040 3590
rect 6104 2514 6132 5510
rect 6184 5296 6236 5302
rect 6184 5238 6236 5244
rect 6196 4758 6224 5238
rect 6184 4752 6236 4758
rect 6184 4694 6236 4700
rect 6288 4706 6316 10610
rect 6552 10532 6604 10538
rect 6552 10474 6604 10480
rect 6564 10062 6592 10474
rect 6920 10464 6972 10470
rect 6972 10424 7052 10452
rect 6920 10406 6972 10412
rect 7024 10266 7052 10424
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 7116 10198 7144 10950
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 7104 10192 7156 10198
rect 7104 10134 7156 10140
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6380 8634 6408 9998
rect 7024 9722 7052 10066
rect 7012 9716 7064 9722
rect 7012 9658 7064 9664
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6552 8016 6604 8022
rect 6552 7958 6604 7964
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6380 6866 6408 7278
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6368 6860 6420 6866
rect 6368 6802 6420 6808
rect 6368 6384 6420 6390
rect 6472 6361 6500 7142
rect 6368 6326 6420 6332
rect 6458 6352 6514 6361
rect 6380 5302 6408 6326
rect 6458 6287 6514 6296
rect 6564 6254 6592 7958
rect 6748 7478 6776 8434
rect 7024 8430 7052 9318
rect 7116 8537 7144 9522
rect 7208 8974 7236 10406
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 7102 8528 7158 8537
rect 7102 8463 7158 8472
rect 7012 8424 7064 8430
rect 7012 8366 7064 8372
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6736 7472 6788 7478
rect 6736 7414 6788 7420
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6656 6662 6684 6802
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6748 6474 6776 7414
rect 6656 6446 6776 6474
rect 6552 6248 6604 6254
rect 6458 6216 6514 6225
rect 6552 6190 6604 6196
rect 6458 6151 6514 6160
rect 6368 5296 6420 5302
rect 6368 5238 6420 5244
rect 6472 4826 6500 6151
rect 6656 5681 6684 6446
rect 6736 6384 6788 6390
rect 6736 6326 6788 6332
rect 6748 5828 6776 6326
rect 6840 6254 6868 7414
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6840 5953 6868 6054
rect 6826 5944 6882 5953
rect 6826 5879 6882 5888
rect 6828 5840 6880 5846
rect 6748 5800 6828 5828
rect 6828 5782 6880 5788
rect 6642 5672 6698 5681
rect 6642 5607 6698 5616
rect 6736 5636 6788 5642
rect 6736 5578 6788 5584
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 6552 4820 6604 4826
rect 6552 4762 6604 4768
rect 6564 4706 6592 4762
rect 6288 4678 6592 4706
rect 6276 4548 6328 4554
rect 6276 4490 6328 4496
rect 6288 3738 6316 4490
rect 6564 4185 6592 4678
rect 6656 4622 6684 5510
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6748 4298 6776 5578
rect 6656 4270 6776 4298
rect 6550 4176 6606 4185
rect 6550 4111 6606 4120
rect 6460 4004 6512 4010
rect 6460 3946 6512 3952
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 6288 3058 6316 3674
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 6288 2922 6316 2994
rect 6276 2916 6328 2922
rect 6276 2858 6328 2864
rect 6092 2508 6144 2514
rect 6092 2450 6144 2456
rect 6472 800 6500 3946
rect 6656 3720 6684 4270
rect 6736 4208 6788 4214
rect 6734 4176 6736 4185
rect 6788 4176 6790 4185
rect 6734 4111 6790 4120
rect 6656 3692 6776 3720
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6656 3194 6684 3538
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6748 2990 6776 3692
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 6644 2848 6696 2854
rect 6644 2790 6696 2796
rect 6656 2582 6684 2790
rect 6748 2650 6776 2926
rect 6840 2854 6868 5782
rect 6932 4146 6960 7686
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 7024 4078 7052 7686
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7116 5166 7144 6598
rect 7208 6225 7236 8910
rect 7194 6216 7250 6225
rect 7194 6151 7250 6160
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 7024 3670 7052 4014
rect 7116 4010 7144 5102
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 7208 4758 7236 4966
rect 7196 4752 7248 4758
rect 7196 4694 7248 4700
rect 7196 4480 7248 4486
rect 7196 4422 7248 4428
rect 7104 4004 7156 4010
rect 7104 3946 7156 3952
rect 7012 3664 7064 3670
rect 7012 3606 7064 3612
rect 7208 3482 7236 4422
rect 6932 3454 7236 3482
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 6644 2576 6696 2582
rect 6644 2518 6696 2524
rect 6932 800 6960 3454
rect 7300 2650 7328 11834
rect 7392 10470 7420 16136
rect 7576 14890 7604 18566
rect 7668 16250 7696 19790
rect 7840 19780 7892 19786
rect 7840 19722 7892 19728
rect 7748 19712 7800 19718
rect 7748 19654 7800 19660
rect 7760 19310 7788 19654
rect 7748 19304 7800 19310
rect 7748 19246 7800 19252
rect 7852 19156 7880 19722
rect 8208 19712 8260 19718
rect 8208 19654 8260 19660
rect 8220 19242 8248 19654
rect 9692 19514 9720 20266
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 18800 20058 18828 20266
rect 18788 20052 18840 20058
rect 18788 19994 18840 20000
rect 17960 19916 18012 19922
rect 17960 19858 18012 19864
rect 10324 19848 10376 19854
rect 10324 19790 10376 19796
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 10336 19310 10364 19790
rect 11704 19712 11756 19718
rect 11704 19654 11756 19660
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 9496 19304 9548 19310
rect 9496 19246 9548 19252
rect 10324 19304 10376 19310
rect 10324 19246 10376 19252
rect 8208 19236 8260 19242
rect 8208 19178 8260 19184
rect 7760 19128 7880 19156
rect 7656 16244 7708 16250
rect 7656 16186 7708 16192
rect 7564 14884 7616 14890
rect 7564 14826 7616 14832
rect 7576 13938 7604 14826
rect 7760 13954 7788 19128
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 8220 18630 8248 19178
rect 9036 18828 9088 18834
rect 9036 18770 9088 18776
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 8220 18290 8248 18566
rect 9048 18290 9076 18770
rect 8208 18284 8260 18290
rect 8208 18226 8260 18232
rect 9036 18284 9088 18290
rect 9036 18226 9088 18232
rect 9128 18148 9180 18154
rect 9128 18090 9180 18096
rect 8852 18080 8904 18086
rect 8852 18022 8904 18028
rect 8944 18080 8996 18086
rect 8944 18022 8996 18028
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7886 15728 8182 15748
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 8220 14618 8248 15098
rect 8208 14612 8260 14618
rect 8208 14554 8260 14560
rect 7564 13932 7616 13938
rect 7564 13874 7616 13880
rect 7668 13926 7788 13954
rect 7576 13326 7604 13874
rect 7668 13734 7696 13926
rect 8220 13870 8248 14554
rect 8312 14074 8340 17682
rect 8864 17542 8892 18022
rect 8956 17610 8984 18022
rect 8944 17604 8996 17610
rect 8944 17546 8996 17552
rect 8852 17536 8904 17542
rect 8852 17478 8904 17484
rect 8864 17270 8892 17478
rect 9140 17338 9168 18090
rect 9404 18080 9456 18086
rect 9404 18022 9456 18028
rect 9416 17882 9444 18022
rect 9404 17876 9456 17882
rect 9404 17818 9456 17824
rect 9404 17740 9456 17746
rect 9404 17682 9456 17688
rect 9128 17332 9180 17338
rect 9128 17274 9180 17280
rect 8852 17264 8904 17270
rect 8852 17206 8904 17212
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 8404 16658 8432 16934
rect 8392 16652 8444 16658
rect 8392 16594 8444 16600
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 8392 15496 8444 15502
rect 8392 15438 8444 15444
rect 8404 14958 8432 15438
rect 8392 14952 8444 14958
rect 8392 14894 8444 14900
rect 8496 14482 8524 15506
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 7748 13864 7800 13870
rect 7748 13806 7800 13812
rect 8208 13864 8260 13870
rect 8208 13806 8260 13812
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7668 13530 7696 13670
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 7760 13462 7788 13806
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7886 13552 8182 13572
rect 8496 13530 8524 14418
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 7748 13456 7800 13462
rect 7748 13398 7800 13404
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7392 9042 7420 9522
rect 7380 9036 7432 9042
rect 7380 8978 7432 8984
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7392 8566 7420 8774
rect 7380 8560 7432 8566
rect 7380 8502 7432 8508
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 7392 2514 7420 7142
rect 7484 5914 7512 13126
rect 7576 12850 7604 13262
rect 7564 12844 7616 12850
rect 7616 12804 7696 12832
rect 7564 12786 7616 12792
rect 7668 12220 7696 12804
rect 7760 12434 7788 13398
rect 8576 13388 8628 13394
rect 8576 13330 8628 13336
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 8390 12744 8446 12753
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 7760 12406 7880 12434
rect 7748 12232 7800 12238
rect 7668 12192 7748 12220
rect 7748 12174 7800 12180
rect 7852 11898 7880 12406
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7748 11824 7800 11830
rect 7932 11824 7984 11830
rect 7748 11766 7800 11772
rect 7930 11792 7932 11801
rect 7984 11792 7986 11801
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 7668 11132 7696 11698
rect 7760 11286 7788 11766
rect 7930 11727 7986 11736
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 8220 11370 8248 12718
rect 8390 12679 8392 12688
rect 8444 12679 8446 12688
rect 8392 12650 8444 12656
rect 8220 11342 8432 11370
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 8208 11280 8260 11286
rect 8208 11222 8260 11228
rect 7668 11104 7788 11132
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 7564 10532 7616 10538
rect 7564 10474 7616 10480
rect 7576 9586 7604 10474
rect 7668 10198 7696 10950
rect 7656 10192 7708 10198
rect 7656 10134 7708 10140
rect 7760 9674 7788 11104
rect 8024 11076 8076 11082
rect 8024 11018 8076 11024
rect 8036 10538 8064 11018
rect 8024 10532 8076 10538
rect 8024 10474 8076 10480
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7886 10288 8182 10308
rect 8220 10266 8248 11222
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 7760 9654 7880 9674
rect 7760 9648 7892 9654
rect 7760 9646 7840 9648
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7576 9178 7604 9522
rect 7656 9444 7708 9450
rect 7656 9386 7708 9392
rect 7564 9172 7616 9178
rect 7564 9114 7616 9120
rect 7576 8498 7604 9114
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7668 8430 7696 9386
rect 7760 9178 7788 9646
rect 7840 9590 7892 9596
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 8022 8528 8078 8537
rect 8022 8463 8024 8472
rect 8076 8463 8078 8472
rect 8024 8434 8076 8440
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 7576 5778 7604 6802
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7484 4486 7512 5102
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7484 3942 7512 4082
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7576 2774 7604 5714
rect 7668 5370 7696 8366
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7886 8112 8182 8132
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 7760 7478 7788 7822
rect 7748 7472 7800 7478
rect 7748 7414 7800 7420
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7760 7002 7788 7142
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7760 6798 7788 6938
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7760 5710 7788 6258
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7656 5364 7708 5370
rect 7656 5306 7708 5312
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 7840 4548 7892 4554
rect 7840 4490 7892 4496
rect 7748 3936 7800 3942
rect 7852 3924 7880 4490
rect 8220 4146 8248 10066
rect 8312 9926 8340 10542
rect 8404 10130 8432 11342
rect 8588 11082 8616 13330
rect 8864 12434 8892 17206
rect 9220 17060 9272 17066
rect 9220 17002 9272 17008
rect 9232 16726 9260 17002
rect 9128 16720 9180 16726
rect 9128 16662 9180 16668
rect 9220 16720 9272 16726
rect 9220 16662 9272 16668
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 9048 12986 9076 13670
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 9036 12844 9088 12850
rect 9036 12786 9088 12792
rect 8864 12406 8984 12434
rect 8760 12300 8812 12306
rect 8760 12242 8812 12248
rect 8772 12170 8800 12242
rect 8760 12164 8812 12170
rect 8760 12106 8812 12112
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 8864 11354 8892 11494
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 8588 10130 8616 11018
rect 8760 10668 8812 10674
rect 8760 10610 8812 10616
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8680 10266 8708 10406
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8576 10124 8628 10130
rect 8576 10066 8628 10072
rect 8772 10062 8800 10610
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8404 9518 8432 9862
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8312 9110 8340 9318
rect 8300 9104 8352 9110
rect 8300 9046 8352 9052
rect 8404 7954 8432 9454
rect 8576 9376 8628 9382
rect 8576 9318 8628 9324
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8496 8566 8524 8978
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 8588 8265 8616 9318
rect 8772 8430 8800 9998
rect 8760 8424 8812 8430
rect 8666 8392 8722 8401
rect 8760 8366 8812 8372
rect 8666 8327 8722 8336
rect 8574 8256 8630 8265
rect 8574 8191 8630 8200
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8390 7848 8446 7857
rect 8300 7812 8352 7818
rect 8390 7783 8392 7792
rect 8300 7754 8352 7760
rect 8444 7783 8446 7792
rect 8392 7754 8444 7760
rect 8312 7002 8340 7754
rect 8496 7002 8524 8026
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 8588 6882 8616 8191
rect 8496 6854 8616 6882
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8312 6458 8340 6734
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8404 6254 8432 6734
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8312 5302 8340 5646
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 8404 5166 8432 6054
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8300 4752 8352 4758
rect 8298 4720 8300 4729
rect 8352 4720 8354 4729
rect 8298 4655 8354 4664
rect 8496 4554 8524 6854
rect 8680 6186 8708 8327
rect 8772 7750 8800 8366
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8772 7274 8800 7686
rect 8760 7268 8812 7274
rect 8760 7210 8812 7216
rect 8668 6180 8720 6186
rect 8668 6122 8720 6128
rect 8576 5636 8628 5642
rect 8576 5578 8628 5584
rect 8588 5234 8616 5578
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 8680 5098 8708 6122
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8668 5092 8720 5098
rect 8668 5034 8720 5040
rect 8772 5030 8800 5850
rect 8864 5250 8892 11086
rect 8956 5409 8984 12406
rect 9048 11150 9076 12786
rect 9036 11144 9088 11150
rect 9036 11086 9088 11092
rect 9036 10464 9088 10470
rect 9140 10452 9168 16662
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 9088 10424 9168 10452
rect 9220 10464 9272 10470
rect 9036 10406 9088 10412
rect 9220 10406 9272 10412
rect 9048 7410 9076 10406
rect 9232 9994 9260 10406
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 9232 7954 9260 8230
rect 9220 7948 9272 7954
rect 9220 7890 9272 7896
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 9048 6798 9076 7346
rect 9128 7336 9180 7342
rect 9126 7304 9128 7313
rect 9180 7304 9182 7313
rect 9126 7239 9182 7248
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 9036 6792 9088 6798
rect 9036 6734 9088 6740
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9036 6248 9088 6254
rect 9036 6190 9088 6196
rect 8942 5400 8998 5409
rect 8942 5335 8998 5344
rect 8864 5222 8984 5250
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8484 4548 8536 4554
rect 8484 4490 8536 4496
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 7800 3896 7880 3924
rect 7748 3878 7800 3884
rect 7886 3836 8182 3856
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7886 3760 8182 3780
rect 8312 3670 8340 4422
rect 8588 4282 8616 4558
rect 8576 4276 8628 4282
rect 8576 4218 8628 4224
rect 8392 4072 8444 4078
rect 8444 4032 8524 4060
rect 8392 4014 8444 4020
rect 8496 3942 8524 4032
rect 8588 4010 8616 4218
rect 8576 4004 8628 4010
rect 8576 3946 8628 3952
rect 8760 4004 8812 4010
rect 8760 3946 8812 3952
rect 8392 3936 8444 3942
rect 8392 3878 8444 3884
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8404 3738 8432 3878
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8300 3664 8352 3670
rect 8300 3606 8352 3612
rect 7932 3596 7984 3602
rect 7932 3538 7984 3544
rect 7944 3194 7972 3538
rect 8116 3528 8168 3534
rect 8496 3516 8524 3878
rect 8588 3738 8616 3946
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8772 3584 8800 3946
rect 8168 3488 8524 3516
rect 8680 3556 8800 3584
rect 8116 3470 8168 3476
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 7484 2746 7604 2774
rect 7380 2508 7432 2514
rect 7380 2450 7432 2456
rect 7392 1834 7420 2450
rect 7380 1828 7432 1834
rect 7380 1770 7432 1776
rect 7484 1442 7512 2746
rect 7392 1414 7512 1442
rect 7392 800 7420 1414
rect 7760 1170 7788 2790
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 8220 2446 8248 3130
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 8496 2310 8524 3130
rect 8680 2922 8708 3556
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8668 2916 8720 2922
rect 8668 2858 8720 2864
rect 8772 2650 8800 3334
rect 8956 2774 8984 5222
rect 9048 3942 9076 6190
rect 9140 5166 9168 6734
rect 9128 5160 9180 5166
rect 9128 5102 9180 5108
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 9140 2854 9168 5102
rect 9232 3097 9260 7142
rect 9324 5370 9352 16594
rect 9416 16590 9444 17682
rect 9508 17542 9536 19246
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 9496 17536 9548 17542
rect 9496 17478 9548 17484
rect 9404 16584 9456 16590
rect 9404 16526 9456 16532
rect 9508 15978 9536 17478
rect 9600 17202 9628 18226
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9600 16250 9628 17138
rect 9588 16244 9640 16250
rect 9588 16186 9640 16192
rect 9496 15972 9548 15978
rect 9496 15914 9548 15920
rect 9864 15972 9916 15978
rect 9864 15914 9916 15920
rect 9508 15366 9536 15914
rect 9496 15360 9548 15366
rect 9496 15302 9548 15308
rect 9508 14958 9536 15302
rect 9876 15162 9904 15914
rect 9864 15156 9916 15162
rect 9784 15116 9864 15144
rect 9680 15088 9732 15094
rect 9680 15030 9732 15036
rect 9496 14952 9548 14958
rect 9496 14894 9548 14900
rect 9508 14278 9536 14894
rect 9692 14550 9720 15030
rect 9680 14544 9732 14550
rect 9680 14486 9732 14492
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9784 13938 9812 15116
rect 9864 15098 9916 15104
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9876 13938 9904 14554
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9772 13932 9824 13938
rect 9772 13874 9824 13880
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 9680 13728 9732 13734
rect 9680 13670 9732 13676
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9416 11898 9444 12582
rect 9508 12442 9536 12582
rect 9496 12436 9548 12442
rect 9496 12378 9548 12384
rect 9586 12200 9642 12209
rect 9586 12135 9642 12144
rect 9404 11892 9456 11898
rect 9404 11834 9456 11840
rect 9600 11778 9628 12135
rect 9692 11898 9720 13670
rect 9784 13530 9812 13670
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9784 12986 9812 13330
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9876 12850 9904 13874
rect 9968 13258 9996 14418
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9968 12238 9996 13194
rect 10060 12714 10088 13738
rect 10152 12986 10180 19110
rect 11716 18902 11744 19654
rect 13360 19304 13412 19310
rect 13360 19246 13412 19252
rect 11704 18896 11756 18902
rect 11704 18838 11756 18844
rect 12624 18828 12676 18834
rect 12624 18770 12676 18776
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 10876 18420 10928 18426
rect 10876 18362 10928 18368
rect 10692 18352 10744 18358
rect 10692 18294 10744 18300
rect 10324 17876 10376 17882
rect 10324 17818 10376 17824
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10232 13456 10284 13462
rect 10230 13424 10232 13433
rect 10284 13424 10286 13433
rect 10230 13359 10286 13368
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 10048 12708 10100 12714
rect 10048 12650 10100 12656
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9600 11750 9812 11778
rect 9968 11762 9996 12174
rect 9784 10674 9812 11750
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 9864 11688 9916 11694
rect 9864 11630 9916 11636
rect 9876 11558 9904 11630
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9772 10668 9824 10674
rect 9772 10610 9824 10616
rect 9692 10198 9720 10610
rect 9680 10192 9732 10198
rect 9680 10134 9732 10140
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9678 9616 9734 9625
rect 9588 9580 9640 9586
rect 9678 9551 9734 9560
rect 9588 9522 9640 9528
rect 9600 9178 9628 9522
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9692 9042 9720 9551
rect 9784 9382 9812 10066
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9680 9036 9732 9042
rect 9600 8996 9680 9024
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9416 8430 9444 8910
rect 9404 8424 9456 8430
rect 9404 8366 9456 8372
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9416 7546 9444 8366
rect 9508 8265 9536 8366
rect 9494 8256 9550 8265
rect 9494 8191 9550 8200
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9404 6180 9456 6186
rect 9404 6122 9456 6128
rect 9416 5846 9444 6122
rect 9508 5930 9536 8026
rect 9600 7698 9628 8996
rect 9680 8978 9732 8984
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9692 7818 9720 8842
rect 9680 7812 9732 7818
rect 9680 7754 9732 7760
rect 9600 7670 9720 7698
rect 9692 7478 9720 7670
rect 9680 7472 9732 7478
rect 9680 7414 9732 7420
rect 9588 7268 9640 7274
rect 9588 7210 9640 7216
rect 9680 7268 9732 7274
rect 9680 7210 9732 7216
rect 9600 6866 9628 7210
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9600 6254 9628 6802
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 9508 5902 9628 5930
rect 9404 5840 9456 5846
rect 9404 5782 9456 5788
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9402 5672 9458 5681
rect 9402 5607 9458 5616
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 9416 4826 9444 5607
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9324 4078 9352 4558
rect 9508 4554 9536 5714
rect 9600 4758 9628 5902
rect 9692 5794 9720 7210
rect 9784 6254 9812 9318
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9784 5914 9812 6190
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9692 5766 9812 5794
rect 9588 4752 9640 4758
rect 9588 4694 9640 4700
rect 9680 4752 9732 4758
rect 9680 4694 9732 4700
rect 9496 4548 9548 4554
rect 9496 4490 9548 4496
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9218 3088 9274 3097
rect 9218 3023 9274 3032
rect 9324 2990 9352 3878
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9416 3126 9444 3538
rect 9508 3466 9536 4490
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 9496 3460 9548 3466
rect 9496 3402 9548 3408
rect 9404 3120 9456 3126
rect 9404 3062 9456 3068
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 9496 2916 9548 2922
rect 9496 2858 9548 2864
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 8956 2746 9076 2774
rect 8760 2644 8812 2650
rect 8760 2586 8812 2592
rect 8576 2508 8628 2514
rect 8576 2450 8628 2456
rect 8484 2304 8536 2310
rect 8484 2246 8536 2252
rect 8588 2106 8616 2450
rect 9048 2378 9076 2746
rect 9036 2372 9088 2378
rect 9036 2314 9088 2320
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 8300 2100 8352 2106
rect 8300 2042 8352 2048
rect 8576 2100 8628 2106
rect 8576 2042 8628 2048
rect 7760 1142 7880 1170
rect 7852 800 7880 1142
rect 8312 800 8340 2042
rect 9232 2038 9260 2246
rect 9220 2032 9272 2038
rect 9220 1974 9272 1980
rect 9220 1828 9272 1834
rect 9220 1770 9272 1776
rect 8760 1488 8812 1494
rect 8760 1430 8812 1436
rect 8772 800 8800 1430
rect 9232 800 9260 1770
rect 9508 1494 9536 2858
rect 9496 1488 9548 1494
rect 9496 1430 9548 1436
rect 9600 800 9628 3538
rect 9692 2990 9720 4694
rect 9784 4690 9812 5766
rect 9876 4706 9904 11494
rect 9956 9444 10008 9450
rect 9956 9386 10008 9392
rect 9968 8809 9996 9386
rect 9954 8800 10010 8809
rect 9954 8735 10010 8744
rect 9968 6236 9996 8735
rect 10060 6304 10088 12650
rect 10244 11744 10272 13262
rect 10152 11716 10272 11744
rect 10152 11014 10180 11716
rect 10230 11656 10286 11665
rect 10230 11591 10286 11600
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 10244 10810 10272 11591
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 10140 10192 10192 10198
rect 10140 10134 10192 10140
rect 10152 8906 10180 10134
rect 10244 9500 10272 10406
rect 10336 9654 10364 17818
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 10520 17270 10548 17478
rect 10508 17264 10560 17270
rect 10508 17206 10560 17212
rect 10508 17128 10560 17134
rect 10508 17070 10560 17076
rect 10416 16652 10468 16658
rect 10416 16594 10468 16600
rect 10428 11665 10456 16594
rect 10520 14074 10548 17070
rect 10612 16998 10640 17818
rect 10600 16992 10652 16998
rect 10600 16934 10652 16940
rect 10508 14068 10560 14074
rect 10508 14010 10560 14016
rect 10508 13728 10560 13734
rect 10508 13670 10560 13676
rect 10520 13190 10548 13670
rect 10508 13184 10560 13190
rect 10508 13126 10560 13132
rect 10508 12912 10560 12918
rect 10508 12854 10560 12860
rect 10414 11656 10470 11665
rect 10414 11591 10470 11600
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10324 9648 10376 9654
rect 10324 9590 10376 9596
rect 10324 9512 10376 9518
rect 10244 9472 10324 9500
rect 10324 9454 10376 9460
rect 10428 9058 10456 11494
rect 10244 9030 10456 9058
rect 10140 8900 10192 8906
rect 10140 8842 10192 8848
rect 10152 8566 10180 8842
rect 10140 8560 10192 8566
rect 10140 8502 10192 8508
rect 10060 6276 10180 6304
rect 9968 6208 10088 6236
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 9968 4826 9996 4966
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 9772 4684 9824 4690
rect 9876 4678 9996 4706
rect 9772 4626 9824 4632
rect 9784 3641 9812 4626
rect 9864 4480 9916 4486
rect 9864 4422 9916 4428
rect 9876 4185 9904 4422
rect 9862 4176 9918 4185
rect 9862 4111 9918 4120
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9770 3632 9826 3641
rect 9770 3567 9826 3576
rect 9876 3534 9904 3878
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 9876 3058 9904 3470
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 9680 2984 9732 2990
rect 9680 2926 9732 2932
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 9784 2650 9812 2926
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 9876 2446 9904 2994
rect 9968 2854 9996 4678
rect 10060 4282 10088 6208
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 10060 3754 10088 4014
rect 10152 3942 10180 6276
rect 10244 5545 10272 9030
rect 10414 8936 10470 8945
rect 10414 8871 10470 8880
rect 10322 8528 10378 8537
rect 10322 8463 10324 8472
rect 10376 8463 10378 8472
rect 10324 8434 10376 8440
rect 10324 6384 10376 6390
rect 10324 6326 10376 6332
rect 10336 6225 10364 6326
rect 10322 6216 10378 6225
rect 10322 6151 10378 6160
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10230 5536 10286 5545
rect 10230 5471 10286 5480
rect 10336 4146 10364 6054
rect 10428 5828 10456 8871
rect 10520 8362 10548 12854
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10508 5840 10560 5846
rect 10428 5800 10508 5828
rect 10508 5782 10560 5788
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10428 5370 10456 5510
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 10428 5166 10456 5306
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 10428 4282 10456 4966
rect 10520 4593 10548 5782
rect 10506 4584 10562 4593
rect 10506 4519 10562 4528
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10612 4162 10640 16934
rect 10704 16810 10732 18294
rect 10888 17202 10916 18362
rect 12348 18284 12400 18290
rect 12348 18226 12400 18232
rect 11980 18148 12032 18154
rect 11980 18090 12032 18096
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 11060 17808 11112 17814
rect 11060 17750 11112 17756
rect 10876 17196 10928 17202
rect 10876 17138 10928 17144
rect 10968 16992 11020 16998
rect 10968 16934 11020 16940
rect 10704 16782 10824 16810
rect 10980 16794 11008 16934
rect 10692 14884 10744 14890
rect 10692 14826 10744 14832
rect 10704 14618 10732 14826
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10704 13394 10732 14010
rect 10692 13388 10744 13394
rect 10692 13330 10744 13336
rect 10704 12850 10732 13330
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 10704 9489 10732 10610
rect 10796 10130 10824 16782
rect 10968 16788 11020 16794
rect 10968 16730 11020 16736
rect 10876 16720 10928 16726
rect 10874 16688 10876 16697
rect 10928 16688 10930 16697
rect 10874 16623 10930 16632
rect 11072 16114 11100 17750
rect 11244 17740 11296 17746
rect 11244 17682 11296 17688
rect 11256 17542 11284 17682
rect 11244 17536 11296 17542
rect 11244 17478 11296 17484
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 11716 17338 11744 18022
rect 11244 17332 11296 17338
rect 11244 17274 11296 17280
rect 11704 17332 11756 17338
rect 11704 17274 11756 17280
rect 11256 17066 11284 17274
rect 11428 17196 11480 17202
rect 11428 17138 11480 17144
rect 11244 17060 11296 17066
rect 11244 17002 11296 17008
rect 11440 16590 11468 17138
rect 11992 16794 12020 18090
rect 12072 17672 12124 17678
rect 12072 17614 12124 17620
rect 12084 17202 12112 17614
rect 12360 17542 12388 18226
rect 12164 17536 12216 17542
rect 12164 17478 12216 17484
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 12072 17196 12124 17202
rect 12072 17138 12124 17144
rect 11980 16788 12032 16794
rect 11980 16730 12032 16736
rect 11428 16584 11480 16590
rect 11428 16526 11480 16532
rect 12176 16522 12204 17478
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 12164 16516 12216 16522
rect 12164 16458 12216 16464
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 12268 15910 12296 17138
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 10968 13456 11020 13462
rect 10966 13424 10968 13433
rect 11020 13424 11022 13433
rect 10966 13359 11022 13368
rect 11072 12322 11100 15846
rect 12360 15638 12388 17478
rect 12348 15632 12400 15638
rect 12348 15574 12400 15580
rect 12636 15570 12664 18770
rect 13372 18766 13400 19246
rect 13452 19236 13504 19242
rect 13452 19178 13504 19184
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 13360 18624 13412 18630
rect 13464 18612 13492 19178
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 14004 18896 14056 18902
rect 14004 18838 14056 18844
rect 13412 18584 13492 18612
rect 13360 18566 13412 18572
rect 13372 17678 13400 18566
rect 13728 17740 13780 17746
rect 13728 17682 13780 17688
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 12716 17264 12768 17270
rect 12716 17206 12768 17212
rect 12728 16726 12756 17206
rect 12992 17128 13044 17134
rect 12992 17070 13044 17076
rect 12716 16720 12768 16726
rect 12716 16662 12768 16668
rect 13004 16658 13032 17070
rect 12992 16652 13044 16658
rect 12992 16594 13044 16600
rect 12624 15564 12676 15570
rect 12624 15506 12676 15512
rect 11888 15360 11940 15366
rect 11888 15302 11940 15308
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 11244 14952 11296 14958
rect 11164 14912 11244 14940
rect 11164 14278 11192 14912
rect 11244 14894 11296 14900
rect 11900 14482 11928 15302
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 12072 14612 12124 14618
rect 12072 14554 12124 14560
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 11900 14226 11928 14418
rect 11980 14272 12032 14278
rect 11900 14220 11980 14226
rect 11900 14214 12032 14220
rect 10888 12294 11100 12322
rect 11164 12306 11192 14214
rect 11900 14198 12020 14214
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 11900 13938 11928 14198
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11704 13796 11756 13802
rect 11704 13738 11756 13744
rect 11716 13530 11744 13738
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 11808 12434 11836 13806
rect 11900 13258 11928 13874
rect 11888 13252 11940 13258
rect 11888 13194 11940 13200
rect 11808 12406 11928 12434
rect 11152 12300 11204 12306
rect 10888 11286 10916 12294
rect 11152 12242 11204 12248
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11716 11762 11744 12242
rect 11808 11898 11836 12242
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11704 11756 11756 11762
rect 11704 11698 11756 11704
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 10876 11280 10928 11286
rect 10876 11222 10928 11228
rect 11256 11150 11284 11290
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 10876 10532 10928 10538
rect 10876 10474 10928 10480
rect 10888 10266 10916 10474
rect 10980 10266 11008 10610
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 10784 10124 10836 10130
rect 10784 10066 10836 10072
rect 10888 9602 10916 10202
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 10796 9574 10916 9602
rect 10968 9648 11020 9654
rect 10968 9590 11020 9596
rect 10690 9480 10746 9489
rect 10690 9415 10746 9424
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 10428 4134 10640 4162
rect 10322 4040 10378 4049
rect 10322 3975 10378 3984
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10060 3726 10272 3754
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 10060 2650 10088 3334
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 10152 2582 10180 2790
rect 10140 2576 10192 2582
rect 10140 2518 10192 2524
rect 9864 2440 9916 2446
rect 10244 2428 10272 3726
rect 10336 3602 10364 3975
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 10428 2774 10456 4134
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 10336 2746 10456 2774
rect 10336 2650 10364 2746
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 9864 2382 9916 2388
rect 10060 2400 10272 2428
rect 10060 800 10088 2400
rect 10520 800 10548 4014
rect 10600 4004 10652 4010
rect 10600 3946 10652 3952
rect 10612 3058 10640 3946
rect 10704 3602 10732 9318
rect 10796 7834 10824 9574
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 10888 8809 10916 9114
rect 10980 8906 11008 9590
rect 11072 9586 11100 9930
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11256 9160 11284 11086
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11716 9722 11744 10202
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11072 9132 11284 9160
rect 10968 8900 11020 8906
rect 10968 8842 11020 8848
rect 10874 8800 10930 8809
rect 10874 8735 10930 8744
rect 10796 7806 10916 7834
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 10796 6866 10824 7686
rect 10888 7546 10916 7806
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10784 6860 10836 6866
rect 10784 6802 10836 6808
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 10796 4078 10824 6054
rect 10888 5012 10916 7142
rect 10980 5166 11008 8842
rect 11072 7206 11100 9132
rect 11348 9042 11376 9318
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 11256 8634 11284 8910
rect 11716 8838 11744 9658
rect 11796 9648 11848 9654
rect 11794 9616 11796 9625
rect 11848 9616 11850 9625
rect 11794 9551 11850 9560
rect 11900 9382 11928 12406
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 11992 11150 12020 12038
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11704 8560 11756 8566
rect 11704 8502 11756 8508
rect 11716 8022 11744 8502
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11704 8016 11756 8022
rect 11704 7958 11756 7964
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11072 5574 11100 7142
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 11060 5296 11112 5302
rect 11060 5238 11112 5244
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 10888 4984 11008 5012
rect 10876 4548 10928 4554
rect 10876 4490 10928 4496
rect 10888 4146 10916 4490
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10796 2774 10824 3878
rect 10876 3664 10928 3670
rect 10980 3652 11008 4984
rect 11072 3670 11100 5238
rect 11164 4622 11192 7278
rect 11808 6866 11836 8230
rect 11796 6860 11848 6866
rect 11796 6802 11848 6808
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 11244 6112 11296 6118
rect 11244 6054 11296 6060
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 11256 4078 11284 6054
rect 11716 5846 11744 6598
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11704 5840 11756 5846
rect 11704 5782 11756 5788
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 11716 5234 11744 5782
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11716 4622 11744 5170
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 11808 4078 11836 6054
rect 11888 5636 11940 5642
rect 11888 5578 11940 5584
rect 11900 5234 11928 5578
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11992 4282 12020 11086
rect 12084 10266 12112 14554
rect 12268 13870 12296 15098
rect 12636 15026 12664 15506
rect 12624 15020 12676 15026
rect 12624 14962 12676 14968
rect 12636 14550 12664 14962
rect 12624 14544 12676 14550
rect 12624 14486 12676 14492
rect 12256 13864 12308 13870
rect 12256 13806 12308 13812
rect 12636 13410 12664 14486
rect 12544 13382 12664 13410
rect 12808 13388 12860 13394
rect 12440 13252 12492 13258
rect 12440 13194 12492 13200
rect 12452 12714 12480 13194
rect 12544 12782 12572 13382
rect 12808 13330 12860 13336
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12440 12708 12492 12714
rect 12440 12650 12492 12656
rect 12452 12442 12480 12650
rect 12164 12436 12216 12442
rect 12164 12378 12216 12384
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12176 11558 12204 12378
rect 12636 11898 12664 13262
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12624 11892 12676 11898
rect 12624 11834 12676 11840
rect 12164 11552 12216 11558
rect 12164 11494 12216 11500
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 12072 9988 12124 9994
rect 12072 9930 12124 9936
rect 12084 9450 12112 9930
rect 12072 9444 12124 9450
rect 12072 9386 12124 9392
rect 12072 8288 12124 8294
rect 12072 8230 12124 8236
rect 12084 8090 12112 8230
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12176 6780 12204 11494
rect 12268 11354 12296 11494
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 12728 10470 12756 12786
rect 12820 11898 12848 13330
rect 12900 12232 12952 12238
rect 12900 12174 12952 12180
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12912 11694 12940 12174
rect 12900 11688 12952 11694
rect 12900 11630 12952 11636
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12360 9674 12388 10066
rect 12268 9646 12388 9674
rect 12268 9450 12296 9646
rect 12256 9444 12308 9450
rect 12256 9386 12308 9392
rect 12268 7886 12296 9386
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12452 8634 12480 8978
rect 12544 8974 12572 10066
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12820 8634 12848 8774
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 12348 7948 12400 7954
rect 12348 7890 12400 7896
rect 12256 7880 12308 7886
rect 12360 7857 12388 7890
rect 12256 7822 12308 7828
rect 12346 7848 12402 7857
rect 12346 7783 12402 7792
rect 12452 7206 12480 8570
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12820 7410 12848 7686
rect 12912 7410 12940 8502
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 12348 7200 12400 7206
rect 12348 7142 12400 7148
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12360 7002 12388 7142
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12452 6934 12480 7142
rect 12440 6928 12492 6934
rect 12440 6870 12492 6876
rect 12176 6752 12388 6780
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 12084 4826 12112 5646
rect 12072 4820 12124 4826
rect 12072 4762 12124 4768
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11796 4072 11848 4078
rect 11796 4014 11848 4020
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 11152 3936 11204 3942
rect 11150 3904 11152 3913
rect 11204 3904 11206 3913
rect 11150 3839 11206 3848
rect 10928 3624 11008 3652
rect 11060 3664 11112 3670
rect 10876 3606 10928 3612
rect 11060 3606 11112 3612
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10888 3058 10916 3470
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 11256 2774 11284 4014
rect 11612 3732 11664 3738
rect 11664 3692 11744 3720
rect 11612 3674 11664 3680
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 11716 3058 11744 3692
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11808 2774 11836 4014
rect 11992 2774 12020 4014
rect 12176 3602 12204 6598
rect 12256 6112 12308 6118
rect 12256 6054 12308 6060
rect 12268 4078 12296 6054
rect 12360 4282 12388 6752
rect 12624 6724 12676 6730
rect 12624 6666 12676 6672
rect 12348 4276 12400 4282
rect 12348 4218 12400 4224
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12256 4072 12308 4078
rect 12256 4014 12308 4020
rect 12164 3596 12216 3602
rect 12164 3538 12216 3544
rect 10704 2746 10824 2774
rect 10980 2746 11284 2774
rect 11716 2746 11836 2774
rect 11900 2746 12020 2774
rect 10704 2514 10732 2746
rect 10692 2508 10744 2514
rect 10692 2450 10744 2456
rect 10704 1834 10732 2450
rect 10692 1828 10744 1834
rect 10692 1770 10744 1776
rect 10980 800 11008 2746
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 11716 1442 11744 2746
rect 11440 1414 11744 1442
rect 11440 800 11468 1414
rect 11900 800 11928 2746
rect 12360 800 12388 4082
rect 12636 3602 12664 6666
rect 12900 6452 12952 6458
rect 12900 6394 12952 6400
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12728 4078 12756 6054
rect 12912 5914 12940 6394
rect 12900 5908 12952 5914
rect 12900 5850 12952 5856
rect 12808 4684 12860 4690
rect 12808 4626 12860 4632
rect 12716 4072 12768 4078
rect 12716 4014 12768 4020
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 12532 3120 12584 3126
rect 12532 3062 12584 3068
rect 12440 2916 12492 2922
rect 12440 2858 12492 2864
rect 12452 2582 12480 2858
rect 12440 2576 12492 2582
rect 12440 2518 12492 2524
rect 12544 2514 12572 3062
rect 12820 2774 12848 4626
rect 13004 3942 13032 16594
rect 13372 16590 13400 17614
rect 13556 17338 13584 17614
rect 13544 17332 13596 17338
rect 13544 17274 13596 17280
rect 13740 17202 13768 17682
rect 13912 17536 13964 17542
rect 13912 17478 13964 17484
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 13924 16726 13952 17478
rect 14016 17270 14044 18838
rect 14568 18834 14596 19110
rect 14817 19068 15113 19088
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14817 18992 15113 19012
rect 14556 18828 14608 18834
rect 14556 18770 14608 18776
rect 14568 18290 14596 18770
rect 15936 18624 15988 18630
rect 15936 18566 15988 18572
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14096 17536 14148 17542
rect 14096 17478 14148 17484
rect 14004 17264 14056 17270
rect 14004 17206 14056 17212
rect 13912 16720 13964 16726
rect 13912 16662 13964 16668
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 13084 16516 13136 16522
rect 13084 16458 13136 16464
rect 13096 16250 13124 16458
rect 14016 16454 14044 17206
rect 14004 16448 14056 16454
rect 14004 16390 14056 16396
rect 14108 16266 14136 17478
rect 14568 16590 14596 18226
rect 14648 18080 14700 18086
rect 14648 18022 14700 18028
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 15200 18080 15252 18086
rect 15200 18022 15252 18028
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 14660 16794 14688 18022
rect 14752 17882 14780 18022
rect 14817 17980 15113 18000
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 14740 17876 14792 17882
rect 14740 17818 14792 17824
rect 15106 17776 15162 17785
rect 15212 17746 15240 18022
rect 15396 17882 15424 18022
rect 15384 17876 15436 17882
rect 15384 17818 15436 17824
rect 15476 17808 15528 17814
rect 15568 17808 15620 17814
rect 15476 17750 15528 17756
rect 15566 17776 15568 17785
rect 15620 17776 15622 17785
rect 15106 17711 15108 17720
rect 15160 17711 15162 17720
rect 15200 17740 15252 17746
rect 15108 17682 15160 17688
rect 15200 17682 15252 17688
rect 15488 17678 15516 17750
rect 15566 17711 15622 17720
rect 15948 17678 15976 18566
rect 17684 18284 17736 18290
rect 17684 18226 17736 18232
rect 17500 18148 17552 18154
rect 17500 18090 17552 18096
rect 16488 17740 16540 17746
rect 16488 17682 16540 17688
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 15936 17672 15988 17678
rect 15936 17614 15988 17620
rect 16120 17672 16172 17678
rect 16120 17614 16172 17620
rect 15488 17202 15516 17614
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 15396 16794 15424 16934
rect 14648 16788 14700 16794
rect 14648 16730 14700 16736
rect 15384 16788 15436 16794
rect 15384 16730 15436 16736
rect 14556 16584 14608 16590
rect 14556 16526 14608 16532
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 13084 16244 13136 16250
rect 13084 16186 13136 16192
rect 14016 16238 14136 16266
rect 13096 15910 13124 16186
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 13096 8537 13124 15846
rect 13176 14952 13228 14958
rect 13176 14894 13228 14900
rect 13188 14618 13216 14894
rect 13636 14884 13688 14890
rect 13636 14826 13688 14832
rect 13648 14618 13676 14826
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 13636 14612 13688 14618
rect 13636 14554 13688 14560
rect 13188 13938 13216 14554
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13176 13932 13228 13938
rect 13176 13874 13228 13880
rect 13832 13870 13860 14418
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13832 12986 13860 13806
rect 13912 13728 13964 13734
rect 13912 13670 13964 13676
rect 13924 13530 13952 13670
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 13268 12708 13320 12714
rect 13268 12650 13320 12656
rect 13280 12238 13308 12650
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 13176 12164 13228 12170
rect 13176 12106 13228 12112
rect 13188 11558 13216 12106
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 13188 10674 13216 11494
rect 13372 10674 13400 12718
rect 13820 11620 13872 11626
rect 13820 11562 13872 11568
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13082 8528 13138 8537
rect 13082 8463 13138 8472
rect 13188 7478 13216 10610
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 13280 8430 13308 9318
rect 13268 8424 13320 8430
rect 13320 8372 13400 8378
rect 13268 8366 13400 8372
rect 13280 8350 13400 8366
rect 13372 7886 13400 8350
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13268 7744 13320 7750
rect 13268 7686 13320 7692
rect 13176 7472 13228 7478
rect 13176 7414 13228 7420
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 13188 4690 13216 6598
rect 13280 5574 13308 7686
rect 13360 6316 13412 6322
rect 13360 6258 13412 6264
rect 13372 5778 13400 6258
rect 13360 5772 13412 5778
rect 13360 5714 13412 5720
rect 13268 5568 13320 5574
rect 13268 5510 13320 5516
rect 13176 4684 13228 4690
rect 13176 4626 13228 4632
rect 13280 4060 13308 5510
rect 13372 5370 13400 5714
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13464 4706 13492 11154
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13648 8022 13676 10406
rect 13832 10266 13860 11562
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 13740 9450 13768 9862
rect 13728 9444 13780 9450
rect 13728 9386 13780 9392
rect 13740 8838 13768 9386
rect 13832 9178 13860 9862
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 14016 8362 14044 16238
rect 15292 16040 15344 16046
rect 15292 15982 15344 15988
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 15304 15706 15332 15982
rect 15292 15700 15344 15706
rect 15292 15642 15344 15648
rect 14924 15564 14976 15570
rect 14924 15506 14976 15512
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14740 15496 14792 15502
rect 14740 15438 14792 15444
rect 14568 14822 14596 15438
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14648 14816 14700 14822
rect 14648 14758 14700 14764
rect 14464 13728 14516 13734
rect 14464 13670 14516 13676
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14188 12640 14240 12646
rect 14188 12582 14240 12588
rect 14200 12374 14228 12582
rect 14188 12368 14240 12374
rect 14108 12316 14188 12322
rect 14108 12310 14240 12316
rect 14108 12294 14228 12310
rect 14108 11830 14136 12294
rect 14200 12245 14228 12294
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14096 11824 14148 11830
rect 14096 11766 14148 11772
rect 14200 11762 14228 12038
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14292 11694 14320 13126
rect 14476 12170 14504 13670
rect 14464 12164 14516 12170
rect 14464 12106 14516 12112
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14568 10606 14596 14758
rect 14660 14006 14688 14758
rect 14752 14074 14780 15438
rect 14936 15162 14964 15506
rect 14924 15156 14976 15162
rect 14924 15098 14976 15104
rect 15292 14884 15344 14890
rect 15292 14826 15344 14832
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 15304 14618 15332 14826
rect 15384 14816 15436 14822
rect 15384 14758 15436 14764
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 15396 14550 15424 14758
rect 15384 14544 15436 14550
rect 15384 14486 15436 14492
rect 15488 14482 15516 16390
rect 15568 15496 15620 15502
rect 15568 15438 15620 15444
rect 14832 14476 14884 14482
rect 14832 14418 14884 14424
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 14648 14000 14700 14006
rect 14648 13942 14700 13948
rect 14844 13938 14872 14418
rect 15384 14340 15436 14346
rect 15384 14282 15436 14288
rect 14832 13932 14884 13938
rect 14832 13874 14884 13880
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 15212 12866 15240 13330
rect 15396 13326 15424 14282
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 15212 12838 15332 12866
rect 15304 12782 15332 12838
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15292 12776 15344 12782
rect 15292 12718 15344 12724
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14817 12464 15113 12484
rect 14924 12368 14976 12374
rect 14924 12310 14976 12316
rect 14936 12102 14964 12310
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 14817 11452 15113 11472
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 15212 11354 15240 12718
rect 15304 12186 15332 12718
rect 15488 12442 15516 14418
rect 15580 14414 15608 15438
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 15580 13734 15608 14350
rect 15568 13728 15620 13734
rect 15568 13670 15620 13676
rect 15672 12986 15700 17274
rect 15948 15638 15976 17614
rect 16132 16658 16160 17614
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 16224 16794 16252 16934
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16120 16652 16172 16658
rect 16120 16594 16172 16600
rect 15936 15632 15988 15638
rect 15936 15574 15988 15580
rect 15844 14544 15896 14550
rect 15844 14486 15896 14492
rect 15752 13796 15804 13802
rect 15752 13738 15804 13744
rect 15660 12980 15712 12986
rect 15660 12922 15712 12928
rect 15672 12646 15700 12922
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15304 12158 15424 12186
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15304 11762 15332 12038
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 15396 11642 15424 12158
rect 15304 11614 15424 11642
rect 15488 11642 15516 12378
rect 15764 12374 15792 13738
rect 15856 12850 15884 14486
rect 16212 13388 16264 13394
rect 16212 13330 16264 13336
rect 16304 13388 16356 13394
rect 16304 13330 16356 13336
rect 16028 12912 16080 12918
rect 16028 12854 16080 12860
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 15856 12442 15884 12786
rect 16040 12481 16068 12854
rect 16026 12472 16082 12481
rect 15844 12436 15896 12442
rect 16026 12407 16082 12416
rect 15844 12378 15896 12384
rect 15752 12368 15804 12374
rect 15752 12310 15804 12316
rect 15856 12102 15884 12378
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 16040 11898 16068 12407
rect 16028 11892 16080 11898
rect 16028 11834 16080 11840
rect 16224 11830 16252 13330
rect 16316 12345 16344 13330
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 16408 12986 16436 13262
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16396 12640 16448 12646
rect 16396 12582 16448 12588
rect 16302 12336 16358 12345
rect 16302 12271 16358 12280
rect 16212 11824 16264 11830
rect 16212 11766 16264 11772
rect 15488 11614 15608 11642
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14292 9722 14320 10542
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 14280 9716 14332 9722
rect 14280 9658 14332 9664
rect 14648 9716 14700 9722
rect 14648 9658 14700 9664
rect 14660 8566 14688 9658
rect 15212 9586 15240 10066
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 14752 8974 14780 9318
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 15212 9178 15240 9318
rect 15200 9172 15252 9178
rect 15200 9114 15252 9120
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 14648 8560 14700 8566
rect 14648 8502 14700 8508
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 14004 8356 14056 8362
rect 14004 8298 14056 8304
rect 13636 8016 13688 8022
rect 13636 7958 13688 7964
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 13556 7410 13584 7890
rect 14016 7546 14044 8298
rect 14292 8022 14320 8434
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 14280 8016 14332 8022
rect 14280 7958 14332 7964
rect 14476 7750 14504 8366
rect 14556 8356 14608 8362
rect 14556 8298 14608 8304
rect 14568 7886 14596 8298
rect 14648 8288 14700 8294
rect 14648 8230 14700 8236
rect 14660 8090 14688 8230
rect 14648 8084 14700 8090
rect 14648 8026 14700 8032
rect 14752 8004 14780 8910
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 14832 8016 14884 8022
rect 14752 7976 14832 8004
rect 14832 7958 14884 7964
rect 14556 7880 14608 7886
rect 14556 7822 14608 7828
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13542 5264 13598 5273
rect 13542 5199 13598 5208
rect 13556 4826 13584 5199
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 13464 4678 13584 4706
rect 13648 4690 13676 6598
rect 14016 6254 14044 7482
rect 14568 6798 14596 7822
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 14648 7200 14700 7206
rect 14648 7142 14700 7148
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 14004 6248 14056 6254
rect 14004 6190 14056 6196
rect 13912 6112 13964 6118
rect 13912 6054 13964 6060
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 13924 5234 13952 6054
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 14108 5234 14136 5510
rect 13912 5228 13964 5234
rect 13912 5170 13964 5176
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 13832 4690 13860 4966
rect 14016 4758 14044 4966
rect 14004 4752 14056 4758
rect 14004 4694 14056 4700
rect 13452 4072 13504 4078
rect 13280 4032 13452 4060
rect 13452 4014 13504 4020
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13464 3670 13492 4014
rect 13556 3942 13584 4678
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13452 3664 13504 3670
rect 13452 3606 13504 3612
rect 12898 3496 12954 3505
rect 12898 3431 12954 3440
rect 12912 2990 12940 3431
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 13084 3392 13136 3398
rect 13084 3334 13136 3340
rect 13004 2990 13032 3334
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 12992 2984 13044 2990
rect 12992 2926 13044 2932
rect 12820 2746 13032 2774
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 12624 2372 12676 2378
rect 12624 2314 12676 2320
rect 12808 2372 12860 2378
rect 12808 2314 12860 2320
rect 12636 1426 12664 2314
rect 12624 1420 12676 1426
rect 12624 1362 12676 1368
rect 12820 800 12848 2314
rect 13004 1902 13032 2746
rect 13096 2446 13124 3334
rect 13360 2848 13412 2854
rect 13360 2790 13412 2796
rect 13372 2650 13400 2790
rect 13648 2774 13676 4626
rect 14108 4078 14136 5170
rect 14200 5098 14228 6054
rect 14568 5914 14596 6054
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 14660 5642 14688 7142
rect 14817 7100 15113 7120
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 15108 6792 15160 6798
rect 15106 6760 15108 6769
rect 15160 6760 15162 6769
rect 15106 6695 15162 6704
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 14648 5636 14700 5642
rect 14648 5578 14700 5584
rect 14660 5137 14688 5578
rect 15212 5234 15240 7686
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 14646 5128 14702 5137
rect 14188 5092 14240 5098
rect 14646 5063 14702 5072
rect 14188 5034 14240 5040
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 14924 4684 14976 4690
rect 14924 4626 14976 4632
rect 14936 4282 14964 4626
rect 15304 4622 15332 11614
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15396 11082 15424 11494
rect 15488 11150 15516 11494
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15384 11076 15436 11082
rect 15384 11018 15436 11024
rect 15580 10810 15608 11614
rect 15844 11348 15896 11354
rect 15844 11290 15896 11296
rect 15936 11348 15988 11354
rect 15936 11290 15988 11296
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15476 10736 15528 10742
rect 15476 10678 15528 10684
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15396 10062 15424 10406
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15488 9625 15516 10678
rect 15856 10130 15884 11290
rect 15948 10266 15976 11290
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 15844 10124 15896 10130
rect 15844 10066 15896 10072
rect 15474 9616 15530 9625
rect 15474 9551 15530 9560
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15396 4826 15424 4966
rect 15384 4820 15436 4826
rect 15384 4762 15436 4768
rect 15384 4684 15436 4690
rect 15384 4626 15436 4632
rect 15292 4616 15344 4622
rect 15292 4558 15344 4564
rect 15200 4548 15252 4554
rect 15200 4490 15252 4496
rect 14924 4276 14976 4282
rect 14924 4218 14976 4224
rect 14096 4072 14148 4078
rect 14096 4014 14148 4020
rect 14280 4004 14332 4010
rect 14280 3946 14332 3952
rect 14292 3194 14320 3946
rect 14817 3836 15113 3856
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 15212 3126 15240 4490
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15304 3942 15332 4082
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 15304 3670 15332 3878
rect 15292 3664 15344 3670
rect 15292 3606 15344 3612
rect 15396 3194 15424 4626
rect 15488 4146 15516 9551
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15580 5778 15608 6598
rect 15856 6390 15884 6802
rect 15844 6384 15896 6390
rect 15844 6326 15896 6332
rect 15568 5772 15620 5778
rect 15568 5714 15620 5720
rect 15476 4140 15528 4146
rect 15476 4082 15528 4088
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 14096 3120 14148 3126
rect 14096 3062 14148 3068
rect 15200 3120 15252 3126
rect 15200 3062 15252 3068
rect 13556 2746 13676 2774
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 12992 1896 13044 1902
rect 12992 1838 13044 1844
rect 13280 800 13308 2314
rect 13452 2304 13504 2310
rect 13452 2246 13504 2252
rect 13464 2106 13492 2246
rect 13452 2100 13504 2106
rect 13452 2042 13504 2048
rect 13556 1970 13584 2746
rect 14108 2582 14136 3062
rect 14556 2916 14608 2922
rect 14556 2858 14608 2864
rect 14096 2576 14148 2582
rect 14096 2518 14148 2524
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 13728 2372 13780 2378
rect 13728 2314 13780 2320
rect 13544 1964 13596 1970
rect 13544 1906 13596 1912
rect 13740 800 13768 2314
rect 14108 800 14136 2382
rect 14568 800 14596 2858
rect 15476 2848 15528 2854
rect 15476 2790 15528 2796
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 15016 2508 15068 2514
rect 15016 2450 15068 2456
rect 15028 2106 15056 2450
rect 15200 2372 15252 2378
rect 15200 2314 15252 2320
rect 15016 2100 15068 2106
rect 15016 2042 15068 2048
rect 15212 1494 15240 2314
rect 15200 1488 15252 1494
rect 15200 1430 15252 1436
rect 15016 1420 15068 1426
rect 15016 1362 15068 1368
rect 15028 800 15056 1362
rect 15488 800 15516 2790
rect 15580 1358 15608 5714
rect 15856 5710 15884 6326
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15844 5704 15896 5710
rect 15844 5646 15896 5652
rect 15844 5296 15896 5302
rect 15844 5238 15896 5244
rect 15856 4690 15884 5238
rect 15844 4684 15896 4690
rect 15844 4626 15896 4632
rect 15844 3936 15896 3942
rect 15844 3878 15896 3884
rect 15856 3058 15884 3878
rect 15948 3641 15976 6054
rect 16040 5846 16068 11086
rect 16212 11076 16264 11082
rect 16316 11064 16344 12271
rect 16264 11036 16344 11064
rect 16212 11018 16264 11024
rect 16120 11008 16172 11014
rect 16120 10950 16172 10956
rect 16132 10742 16160 10950
rect 16120 10736 16172 10742
rect 16120 10678 16172 10684
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 16132 9466 16160 9862
rect 16224 9586 16252 11018
rect 16304 9920 16356 9926
rect 16304 9862 16356 9868
rect 16316 9586 16344 9862
rect 16212 9580 16264 9586
rect 16212 9522 16264 9528
rect 16304 9580 16356 9586
rect 16304 9522 16356 9528
rect 16132 9438 16252 9466
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16132 9110 16160 9318
rect 16120 9104 16172 9110
rect 16120 9046 16172 9052
rect 16224 9042 16252 9438
rect 16212 9036 16264 9042
rect 16212 8978 16264 8984
rect 16224 7954 16252 8978
rect 16212 7948 16264 7954
rect 16212 7890 16264 7896
rect 16120 7540 16172 7546
rect 16120 7482 16172 7488
rect 16132 7449 16160 7482
rect 16118 7440 16174 7449
rect 16118 7375 16174 7384
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 16224 6934 16252 7142
rect 16212 6928 16264 6934
rect 16212 6870 16264 6876
rect 16304 6112 16356 6118
rect 16304 6054 16356 6060
rect 16316 5914 16344 6054
rect 16304 5908 16356 5914
rect 16304 5850 16356 5856
rect 16028 5840 16080 5846
rect 16028 5782 16080 5788
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 16132 3738 16160 4626
rect 16408 4185 16436 12582
rect 16500 9994 16528 17682
rect 17512 17338 17540 18090
rect 17592 18080 17644 18086
rect 17592 18022 17644 18028
rect 17604 17338 17632 18022
rect 17696 17882 17724 18226
rect 17684 17876 17736 17882
rect 17684 17818 17736 17824
rect 17972 17746 18000 19858
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 19352 19514 19380 20266
rect 19524 20256 19576 20262
rect 19524 20198 19576 20204
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 18604 19236 18656 19242
rect 18604 19178 18656 19184
rect 18052 19168 18104 19174
rect 18052 19110 18104 19116
rect 17960 17740 18012 17746
rect 17960 17682 18012 17688
rect 17500 17332 17552 17338
rect 17500 17274 17552 17280
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17224 17060 17276 17066
rect 17224 17002 17276 17008
rect 17316 17060 17368 17066
rect 17316 17002 17368 17008
rect 17236 16794 17264 17002
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 17224 16788 17276 16794
rect 17224 16730 17276 16736
rect 16776 15910 16804 16730
rect 17328 16590 17356 17002
rect 17408 16992 17460 16998
rect 17408 16934 17460 16940
rect 17420 16658 17448 16934
rect 17408 16652 17460 16658
rect 17408 16594 17460 16600
rect 17868 16652 17920 16658
rect 17868 16594 17920 16600
rect 17316 16584 17368 16590
rect 17316 16526 17368 16532
rect 17040 16108 17092 16114
rect 17040 16050 17092 16056
rect 16764 15904 16816 15910
rect 16764 15846 16816 15852
rect 16580 14816 16632 14822
rect 16580 14758 16632 14764
rect 16592 13530 16620 14758
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16776 13394 16804 15846
rect 16948 14272 17000 14278
rect 16948 14214 17000 14220
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16764 13388 16816 13394
rect 16764 13330 16816 13336
rect 16580 13184 16632 13190
rect 16580 13126 16632 13132
rect 16592 12753 16620 13126
rect 16578 12744 16634 12753
rect 16578 12679 16634 12688
rect 16592 11558 16620 12679
rect 16868 11762 16896 13806
rect 16960 13462 16988 14214
rect 16948 13456 17000 13462
rect 17052 13433 17080 16050
rect 17328 15910 17356 16526
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17132 15496 17184 15502
rect 17132 15438 17184 15444
rect 17144 14414 17172 15438
rect 17132 14408 17184 14414
rect 17132 14350 17184 14356
rect 17144 13734 17172 14350
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 16948 13398 17000 13404
rect 17038 13424 17094 13433
rect 17038 13359 17094 13368
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 16580 11552 16632 11558
rect 16580 11494 16632 11500
rect 16592 10606 16620 11494
rect 16764 11076 16816 11082
rect 16764 11018 16816 11024
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16580 10600 16632 10606
rect 16580 10542 16632 10548
rect 16684 10266 16712 10746
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16488 9988 16540 9994
rect 16488 9930 16540 9936
rect 16580 8356 16632 8362
rect 16580 8298 16632 8304
rect 16592 7954 16620 8298
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16580 7812 16632 7818
rect 16580 7754 16632 7760
rect 16488 7472 16540 7478
rect 16488 7414 16540 7420
rect 16500 7154 16528 7414
rect 16592 7274 16620 7754
rect 16580 7268 16632 7274
rect 16580 7210 16632 7216
rect 16672 7268 16724 7274
rect 16672 7210 16724 7216
rect 16500 7126 16620 7154
rect 16488 6860 16540 6866
rect 16488 6802 16540 6808
rect 16394 4176 16450 4185
rect 16394 4111 16450 4120
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 16408 3738 16436 3878
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 16396 3732 16448 3738
rect 16396 3674 16448 3680
rect 15934 3632 15990 3641
rect 15934 3567 15990 3576
rect 15936 3188 15988 3194
rect 15936 3130 15988 3136
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 15568 1352 15620 1358
rect 15568 1294 15620 1300
rect 15948 800 15976 3130
rect 16132 3058 16160 3674
rect 16396 3460 16448 3466
rect 16396 3402 16448 3408
rect 16212 3392 16264 3398
rect 16212 3334 16264 3340
rect 16304 3392 16356 3398
rect 16304 3334 16356 3340
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 16224 2922 16252 3334
rect 16316 2990 16344 3334
rect 16304 2984 16356 2990
rect 16304 2926 16356 2932
rect 16212 2916 16264 2922
rect 16212 2858 16264 2864
rect 16408 800 16436 3402
rect 16500 3380 16528 6802
rect 16592 6202 16620 7126
rect 16684 7002 16712 7210
rect 16672 6996 16724 7002
rect 16672 6938 16724 6944
rect 16684 6322 16712 6938
rect 16672 6316 16724 6322
rect 16672 6258 16724 6264
rect 16592 6174 16712 6202
rect 16580 6112 16632 6118
rect 16580 6054 16632 6060
rect 16592 5166 16620 6054
rect 16580 5160 16632 5166
rect 16580 5102 16632 5108
rect 16580 5024 16632 5030
rect 16580 4966 16632 4972
rect 16592 4078 16620 4966
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 16684 3534 16712 6174
rect 16776 5778 16804 11018
rect 16960 10554 16988 13262
rect 17052 11762 17080 13359
rect 17144 12442 17172 13670
rect 17224 13320 17276 13326
rect 17222 13288 17224 13297
rect 17328 13308 17356 15846
rect 17592 15360 17644 15366
rect 17592 15302 17644 15308
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17276 13288 17356 13308
rect 17278 13280 17356 13288
rect 17222 13223 17278 13232
rect 17132 12436 17184 12442
rect 17132 12378 17184 12384
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 16868 10526 16988 10554
rect 16868 7426 16896 10526
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 16960 9518 16988 10406
rect 16948 9512 17000 9518
rect 16946 9480 16948 9489
rect 17000 9480 17002 9489
rect 16946 9415 17002 9424
rect 16948 8424 17000 8430
rect 16948 8366 17000 8372
rect 16960 8090 16988 8366
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 17052 8022 17080 11698
rect 17224 11008 17276 11014
rect 17224 10950 17276 10956
rect 17236 10538 17264 10950
rect 17224 10532 17276 10538
rect 17224 10474 17276 10480
rect 17132 10464 17184 10470
rect 17132 10406 17184 10412
rect 17144 10062 17172 10406
rect 17132 10056 17184 10062
rect 17132 9998 17184 10004
rect 17144 9586 17172 9998
rect 17316 9716 17368 9722
rect 17420 9704 17448 14214
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17512 13258 17540 13466
rect 17500 13252 17552 13258
rect 17500 13194 17552 13200
rect 17512 11540 17540 13194
rect 17604 12374 17632 15302
rect 17592 12368 17644 12374
rect 17592 12310 17644 12316
rect 17604 11762 17632 12310
rect 17880 12186 17908 16594
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 17972 15026 18000 15506
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 17972 14618 18000 14962
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 17972 13938 18000 14554
rect 17960 13932 18012 13938
rect 17960 13874 18012 13880
rect 17958 12880 18014 12889
rect 17958 12815 18014 12824
rect 17972 12782 18000 12815
rect 17960 12776 18012 12782
rect 17960 12718 18012 12724
rect 17788 12158 17908 12186
rect 17684 12096 17736 12102
rect 17684 12038 17736 12044
rect 17696 11762 17724 12038
rect 17592 11756 17644 11762
rect 17592 11698 17644 11704
rect 17684 11756 17736 11762
rect 17684 11698 17736 11704
rect 17788 11558 17816 12158
rect 17866 11792 17922 11801
rect 17866 11727 17922 11736
rect 17880 11694 17908 11727
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 17592 11552 17644 11558
rect 17512 11512 17592 11540
rect 17592 11494 17644 11500
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 17368 9676 17448 9704
rect 17316 9658 17368 9664
rect 17132 9580 17184 9586
rect 17132 9522 17184 9528
rect 17144 8820 17172 9522
rect 17224 8832 17276 8838
rect 17144 8792 17224 8820
rect 17224 8774 17276 8780
rect 17132 8288 17184 8294
rect 17132 8230 17184 8236
rect 17040 8016 17092 8022
rect 17040 7958 17092 7964
rect 17040 7744 17092 7750
rect 17040 7686 17092 7692
rect 16868 7398 16988 7426
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16764 5772 16816 5778
rect 16764 5714 16816 5720
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 16580 3392 16632 3398
rect 16500 3352 16580 3380
rect 16868 3380 16896 7278
rect 16960 5273 16988 7398
rect 17052 7342 17080 7686
rect 17040 7336 17092 7342
rect 17040 7278 17092 7284
rect 17052 6769 17080 7278
rect 17038 6760 17094 6769
rect 17038 6695 17094 6704
rect 16946 5264 17002 5273
rect 16946 5199 17002 5208
rect 17052 5166 17080 6695
rect 17144 5778 17172 8230
rect 17236 7750 17264 8774
rect 17328 8378 17356 9658
rect 17408 9444 17460 9450
rect 17408 9386 17460 9392
rect 17420 8566 17448 9386
rect 17408 8560 17460 8566
rect 17408 8502 17460 8508
rect 17328 8350 17448 8378
rect 17316 8288 17368 8294
rect 17316 8230 17368 8236
rect 17328 8090 17356 8230
rect 17316 8084 17368 8090
rect 17316 8026 17368 8032
rect 17224 7744 17276 7750
rect 17224 7686 17276 7692
rect 17224 6384 17276 6390
rect 17224 6326 17276 6332
rect 17132 5772 17184 5778
rect 17132 5714 17184 5720
rect 17040 5160 17092 5166
rect 17040 5102 17092 5108
rect 17236 4554 17264 6326
rect 17420 6322 17448 8350
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17512 6882 17540 7482
rect 17604 7002 17632 11494
rect 17684 9988 17736 9994
rect 17684 9930 17736 9936
rect 17696 8090 17724 9930
rect 17788 9110 17816 11494
rect 17776 9104 17828 9110
rect 17776 9046 17828 9052
rect 17788 8265 17816 9046
rect 17774 8256 17830 8265
rect 17774 8191 17830 8200
rect 17880 8106 17908 11630
rect 18064 11354 18092 19110
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 18144 17740 18196 17746
rect 18144 17682 18196 17688
rect 18156 17338 18184 17682
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 18144 17332 18196 17338
rect 18144 17274 18196 17280
rect 18616 16454 18644 19178
rect 19340 19168 19392 19174
rect 19340 19110 19392 19116
rect 18696 18624 18748 18630
rect 18696 18566 18748 18572
rect 18708 16640 18736 18566
rect 18880 18352 18932 18358
rect 18880 18294 18932 18300
rect 18788 17672 18840 17678
rect 18788 17614 18840 17620
rect 18800 17134 18828 17614
rect 18788 17128 18840 17134
rect 18788 17070 18840 17076
rect 18892 16658 18920 18294
rect 18972 18080 19024 18086
rect 18972 18022 19024 18028
rect 18984 17678 19012 18022
rect 18972 17672 19024 17678
rect 18972 17614 19024 17620
rect 18880 16652 18932 16658
rect 18708 16612 18828 16640
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18616 15910 18644 16050
rect 18604 15904 18656 15910
rect 18604 15846 18656 15852
rect 18696 15904 18748 15910
rect 18696 15846 18748 15852
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 18616 14414 18644 15846
rect 18604 14408 18656 14414
rect 18604 14350 18656 14356
rect 18282 14172 18578 14192
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18282 14096 18578 14116
rect 18616 13870 18644 14350
rect 18604 13864 18656 13870
rect 18604 13806 18656 13812
rect 18236 13728 18288 13734
rect 18156 13688 18236 13716
rect 18156 12986 18184 13688
rect 18236 13670 18288 13676
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 18420 12708 18472 12714
rect 18420 12650 18472 12656
rect 18432 12617 18460 12650
rect 18418 12608 18474 12617
rect 18418 12543 18474 12552
rect 18432 12442 18460 12543
rect 18420 12436 18472 12442
rect 18420 12378 18472 12384
rect 18512 12436 18564 12442
rect 18512 12378 18564 12384
rect 18236 12368 18288 12374
rect 18236 12310 18288 12316
rect 18144 12300 18196 12306
rect 18144 12242 18196 12248
rect 18156 11898 18184 12242
rect 18248 12238 18276 12310
rect 18236 12232 18288 12238
rect 18236 12174 18288 12180
rect 18524 12084 18552 12378
rect 18616 12209 18644 13126
rect 18708 12434 18736 15846
rect 18800 13802 18828 16612
rect 18880 16594 18932 16600
rect 18880 13864 18932 13870
rect 18880 13806 18932 13812
rect 18788 13796 18840 13802
rect 18788 13738 18840 13744
rect 18892 13462 18920 13806
rect 18880 13456 18932 13462
rect 18880 13398 18932 13404
rect 18892 12850 18920 13398
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 18984 12442 19012 17614
rect 19064 17060 19116 17066
rect 19064 17002 19116 17008
rect 19076 15366 19104 17002
rect 19352 15366 19380 19110
rect 19432 18216 19484 18222
rect 19432 18158 19484 18164
rect 19064 15360 19116 15366
rect 19064 15302 19116 15308
rect 19340 15360 19392 15366
rect 19340 15302 19392 15308
rect 19076 15094 19104 15302
rect 19064 15088 19116 15094
rect 19064 15030 19116 15036
rect 19248 15020 19300 15026
rect 19248 14962 19300 14968
rect 19156 14816 19208 14822
rect 19156 14758 19208 14764
rect 19168 14618 19196 14758
rect 19156 14612 19208 14618
rect 19156 14554 19208 14560
rect 19260 13938 19288 14962
rect 19248 13932 19300 13938
rect 19248 13874 19300 13880
rect 19340 13728 19392 13734
rect 19340 13670 19392 13676
rect 19352 13530 19380 13670
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19444 13410 19472 18158
rect 19536 16998 19564 20198
rect 19720 19174 19748 20334
rect 20180 20318 20300 20334
rect 20180 19990 20208 20318
rect 20260 20256 20312 20262
rect 20260 20198 20312 20204
rect 20168 19984 20220 19990
rect 20168 19926 20220 19932
rect 19984 19304 20036 19310
rect 19984 19246 20036 19252
rect 19708 19168 19760 19174
rect 19708 19110 19760 19116
rect 19996 18970 20024 19246
rect 20272 18970 20300 20198
rect 20548 20058 20576 22199
rect 20810 20360 20866 20369
rect 20628 20324 20680 20330
rect 20810 20295 20812 20304
rect 20628 20266 20680 20272
rect 20864 20295 20866 20304
rect 21456 20324 21508 20330
rect 20812 20266 20864 20272
rect 21456 20266 21508 20272
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 20352 19916 20404 19922
rect 20352 19858 20404 19864
rect 20364 19446 20392 19858
rect 20640 19514 20668 20266
rect 21180 19916 21232 19922
rect 21180 19858 21232 19864
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20352 19440 20404 19446
rect 20352 19382 20404 19388
rect 20444 19236 20496 19242
rect 20444 19178 20496 19184
rect 19984 18964 20036 18970
rect 19984 18906 20036 18912
rect 20260 18964 20312 18970
rect 20260 18906 20312 18912
rect 19800 18624 19852 18630
rect 19800 18566 19852 18572
rect 19812 17610 19840 18566
rect 20456 18426 20484 19178
rect 21192 18970 21220 19858
rect 21468 19825 21496 20266
rect 21454 19816 21510 19825
rect 21364 19780 21416 19786
rect 21454 19751 21510 19760
rect 21364 19722 21416 19728
rect 21376 19417 21404 19722
rect 21362 19408 21418 19417
rect 21362 19343 21418 19352
rect 21364 19236 21416 19242
rect 21364 19178 21416 19184
rect 21180 18964 21232 18970
rect 21180 18906 21232 18912
rect 21376 18873 21404 19178
rect 21362 18864 21418 18873
rect 21180 18828 21232 18834
rect 21362 18799 21418 18808
rect 21180 18770 21232 18776
rect 20536 18760 20588 18766
rect 20536 18702 20588 18708
rect 20444 18420 20496 18426
rect 20444 18362 20496 18368
rect 20444 18216 20496 18222
rect 20444 18158 20496 18164
rect 20260 18148 20312 18154
rect 20260 18090 20312 18096
rect 20272 17882 20300 18090
rect 19984 17876 20036 17882
rect 19984 17818 20036 17824
rect 20260 17876 20312 17882
rect 20260 17818 20312 17824
rect 19800 17604 19852 17610
rect 19800 17546 19852 17552
rect 19708 17536 19760 17542
rect 19708 17478 19760 17484
rect 19720 17066 19748 17478
rect 19708 17060 19760 17066
rect 19708 17002 19760 17008
rect 19524 16992 19576 16998
rect 19524 16934 19576 16940
rect 19536 13734 19564 16934
rect 19616 16448 19668 16454
rect 19616 16390 19668 16396
rect 19628 16250 19656 16390
rect 19616 16244 19668 16250
rect 19616 16186 19668 16192
rect 19628 15570 19656 16186
rect 19616 15564 19668 15570
rect 19616 15506 19668 15512
rect 19616 15360 19668 15366
rect 19616 15302 19668 15308
rect 19628 14482 19656 15302
rect 19720 15162 19748 17002
rect 19800 16992 19852 16998
rect 19800 16934 19852 16940
rect 19812 16658 19840 16934
rect 19996 16726 20024 17818
rect 20352 17740 20404 17746
rect 20352 17682 20404 17688
rect 20364 17338 20392 17682
rect 20352 17332 20404 17338
rect 20352 17274 20404 17280
rect 20076 17128 20128 17134
rect 20076 17070 20128 17076
rect 19984 16720 20036 16726
rect 19984 16662 20036 16668
rect 19800 16652 19852 16658
rect 19800 16594 19852 16600
rect 19892 16584 19944 16590
rect 19892 16526 19944 16532
rect 19904 16250 19932 16526
rect 19892 16244 19944 16250
rect 19892 16186 19944 16192
rect 19708 15156 19760 15162
rect 19708 15098 19760 15104
rect 19708 14816 19760 14822
rect 19708 14758 19760 14764
rect 19800 14816 19852 14822
rect 19800 14758 19852 14764
rect 19984 14816 20036 14822
rect 19984 14758 20036 14764
rect 19720 14618 19748 14758
rect 19708 14612 19760 14618
rect 19708 14554 19760 14560
rect 19616 14476 19668 14482
rect 19616 14418 19668 14424
rect 19812 13920 19840 14758
rect 19892 14544 19944 14550
rect 19892 14486 19944 14492
rect 19720 13892 19840 13920
rect 19524 13728 19576 13734
rect 19524 13670 19576 13676
rect 19064 13388 19116 13394
rect 19064 13330 19116 13336
rect 19352 13382 19472 13410
rect 18972 12436 19024 12442
rect 18708 12406 18920 12434
rect 18786 12336 18842 12345
rect 18696 12300 18748 12306
rect 18786 12271 18788 12280
rect 18696 12242 18748 12248
rect 18840 12271 18842 12280
rect 18788 12242 18840 12248
rect 18602 12200 18658 12209
rect 18602 12135 18658 12144
rect 18524 12056 18644 12084
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17972 9926 18000 11154
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 18064 10810 18092 11086
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 18064 10130 18092 10610
rect 18420 10464 18472 10470
rect 18420 10406 18472 10412
rect 18432 10266 18460 10406
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 18064 9722 18092 10066
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18282 9744 18578 9764
rect 18052 9716 18104 9722
rect 18052 9658 18104 9664
rect 18616 9042 18644 12056
rect 18708 11529 18736 12242
rect 18788 12096 18840 12102
rect 18788 12038 18840 12044
rect 18800 11898 18828 12038
rect 18788 11892 18840 11898
rect 18788 11834 18840 11840
rect 18694 11520 18750 11529
rect 18694 11455 18750 11464
rect 18604 9036 18656 9042
rect 18604 8978 18656 8984
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 18604 8832 18656 8838
rect 18604 8774 18656 8780
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17788 8078 17908 8106
rect 17592 6996 17644 7002
rect 17592 6938 17644 6944
rect 17512 6866 17632 6882
rect 17512 6860 17644 6866
rect 17512 6854 17592 6860
rect 17592 6802 17644 6808
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17408 6316 17460 6322
rect 17408 6258 17460 6264
rect 17512 6254 17540 6734
rect 17316 6248 17368 6254
rect 17316 6190 17368 6196
rect 17500 6248 17552 6254
rect 17500 6190 17552 6196
rect 17328 5914 17356 6190
rect 17316 5908 17368 5914
rect 17316 5850 17368 5856
rect 17224 4548 17276 4554
rect 17224 4490 17276 4496
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 17500 4480 17552 4486
rect 17500 4422 17552 4428
rect 16948 4004 17000 4010
rect 16948 3946 17000 3952
rect 16580 3334 16632 3340
rect 16684 3352 16896 3380
rect 16684 2038 16712 3352
rect 16960 2774 16988 3946
rect 17040 3936 17092 3942
rect 17040 3878 17092 3884
rect 17052 3058 17080 3878
rect 17144 3602 17172 4422
rect 17408 4004 17460 4010
rect 17408 3946 17460 3952
rect 17420 3670 17448 3946
rect 17408 3664 17460 3670
rect 17408 3606 17460 3612
rect 17132 3596 17184 3602
rect 17132 3538 17184 3544
rect 17224 3120 17276 3126
rect 17224 3062 17276 3068
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 16868 2746 16988 2774
rect 16672 2032 16724 2038
rect 16672 1974 16724 1980
rect 16868 800 16896 2746
rect 17236 2446 17264 3062
rect 17512 2582 17540 4422
rect 17604 2774 17632 6802
rect 17684 6180 17736 6186
rect 17684 6122 17736 6128
rect 17696 5370 17724 6122
rect 17788 5846 17816 8078
rect 17972 8022 18000 8774
rect 18052 8560 18104 8566
rect 18052 8502 18104 8508
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17960 8016 18012 8022
rect 17960 7958 18012 7964
rect 17880 7886 17908 7958
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17880 7546 17908 7822
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 18064 6322 18092 8502
rect 18156 8090 18184 8774
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18144 7744 18196 7750
rect 18248 7732 18276 8434
rect 18196 7704 18276 7732
rect 18144 7686 18196 7692
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18282 7568 18578 7588
rect 18328 7472 18380 7478
rect 18326 7440 18328 7449
rect 18380 7440 18382 7449
rect 18326 7375 18382 7384
rect 18144 6996 18196 7002
rect 18144 6938 18196 6944
rect 18052 6316 18104 6322
rect 18052 6258 18104 6264
rect 17776 5840 17828 5846
rect 17776 5782 17828 5788
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 17684 5364 17736 5370
rect 17684 5306 17736 5312
rect 17788 5166 17816 5646
rect 18052 5636 18104 5642
rect 18052 5578 18104 5584
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 17776 5160 17828 5166
rect 17776 5102 17828 5108
rect 17868 5024 17920 5030
rect 17868 4966 17920 4972
rect 17776 3936 17828 3942
rect 17880 3913 17908 4966
rect 17776 3878 17828 3884
rect 17866 3904 17922 3913
rect 17604 2746 17724 2774
rect 17500 2576 17552 2582
rect 17500 2518 17552 2524
rect 17224 2440 17276 2446
rect 17224 2382 17276 2388
rect 17132 2372 17184 2378
rect 17132 2314 17184 2320
rect 17316 2372 17368 2378
rect 17316 2314 17368 2320
rect 17144 1426 17172 2314
rect 17132 1420 17184 1426
rect 17132 1362 17184 1368
rect 17328 800 17356 2314
rect 4122 598 4200 626
rect 4066 575 4122 584
rect 4250 0 4306 800
rect 4710 0 4766 800
rect 5078 0 5134 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 6918 0 6974 800
rect 7378 0 7434 800
rect 7838 0 7894 800
rect 8298 0 8354 800
rect 8758 0 8814 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 10046 0 10102 800
rect 10506 0 10562 800
rect 10966 0 11022 800
rect 11426 0 11482 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12806 0 12862 800
rect 13266 0 13322 800
rect 13726 0 13782 800
rect 14094 0 14150 800
rect 14554 0 14610 800
rect 15014 0 15070 800
rect 15474 0 15530 800
rect 15934 0 15990 800
rect 16394 0 16450 800
rect 16854 0 16910 800
rect 17314 0 17370 800
rect 17696 241 17724 2746
rect 17788 2650 17816 3878
rect 17866 3839 17922 3848
rect 17866 3632 17922 3641
rect 17866 3567 17922 3576
rect 17880 3194 17908 3567
rect 17972 3534 18000 5510
rect 18064 4078 18092 5578
rect 18156 5166 18184 6938
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 18420 6316 18472 6322
rect 18420 6258 18472 6264
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18432 6202 18460 6258
rect 18340 6174 18460 6202
rect 18340 5846 18368 6174
rect 18328 5840 18380 5846
rect 18328 5782 18380 5788
rect 18524 5778 18552 6258
rect 18616 6254 18644 8774
rect 18708 8566 18736 11455
rect 18892 11286 18920 12406
rect 18972 12378 19024 12384
rect 18972 12096 19024 12102
rect 18972 12038 19024 12044
rect 18880 11280 18932 11286
rect 18880 11222 18932 11228
rect 18984 11082 19012 12038
rect 19076 11830 19104 13330
rect 19156 12232 19208 12238
rect 19156 12174 19208 12180
rect 19064 11824 19116 11830
rect 19168 11801 19196 12174
rect 19064 11766 19116 11772
rect 19154 11792 19210 11801
rect 19154 11727 19210 11736
rect 19064 11552 19116 11558
rect 19062 11520 19064 11529
rect 19116 11520 19118 11529
rect 19062 11455 19118 11464
rect 19064 11212 19116 11218
rect 19064 11154 19116 11160
rect 18972 11076 19024 11082
rect 18972 11018 19024 11024
rect 19076 10985 19104 11154
rect 19156 11144 19208 11150
rect 19156 11086 19208 11092
rect 19062 10976 19118 10985
rect 19062 10911 19118 10920
rect 19168 10538 19196 11086
rect 19156 10532 19208 10538
rect 19156 10474 19208 10480
rect 18788 10464 18840 10470
rect 18788 10406 18840 10412
rect 18696 8560 18748 8566
rect 18696 8502 18748 8508
rect 18696 8424 18748 8430
rect 18800 8378 18828 10406
rect 19168 10266 19196 10474
rect 19156 10260 19208 10266
rect 19156 10202 19208 10208
rect 19352 9042 19380 13382
rect 19720 13326 19748 13892
rect 19800 13796 19852 13802
rect 19800 13738 19852 13744
rect 19708 13320 19760 13326
rect 19522 13288 19578 13297
rect 19708 13262 19760 13268
rect 19522 13223 19578 13232
rect 19536 12714 19564 13223
rect 19432 12708 19484 12714
rect 19432 12650 19484 12656
rect 19524 12708 19576 12714
rect 19524 12650 19576 12656
rect 19444 11898 19472 12650
rect 19708 12640 19760 12646
rect 19706 12608 19708 12617
rect 19760 12608 19762 12617
rect 19706 12543 19762 12552
rect 19812 12442 19840 13738
rect 19904 12850 19932 14486
rect 19996 14074 20024 14758
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 19892 12844 19944 12850
rect 19892 12786 19944 12792
rect 19800 12436 19852 12442
rect 19800 12378 19852 12384
rect 20088 12170 20116 17070
rect 20352 17060 20404 17066
rect 20352 17002 20404 17008
rect 20364 16794 20392 17002
rect 20260 16788 20312 16794
rect 20260 16730 20312 16736
rect 20352 16788 20404 16794
rect 20352 16730 20404 16736
rect 20272 16046 20300 16730
rect 20260 16040 20312 16046
rect 20260 15982 20312 15988
rect 20352 15904 20404 15910
rect 20352 15846 20404 15852
rect 20364 15638 20392 15846
rect 20352 15632 20404 15638
rect 20352 15574 20404 15580
rect 20352 14884 20404 14890
rect 20352 14826 20404 14832
rect 20364 14074 20392 14826
rect 20352 14068 20404 14074
rect 20352 14010 20404 14016
rect 20168 13864 20220 13870
rect 20168 13806 20220 13812
rect 20180 13258 20208 13806
rect 20260 13728 20312 13734
rect 20260 13670 20312 13676
rect 20272 13530 20300 13670
rect 20260 13524 20312 13530
rect 20260 13466 20312 13472
rect 20168 13252 20220 13258
rect 20168 13194 20220 13200
rect 20352 13252 20404 13258
rect 20352 13194 20404 13200
rect 20364 12850 20392 13194
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20168 12436 20220 12442
rect 20168 12378 20220 12384
rect 20180 12238 20208 12378
rect 20364 12238 20392 12786
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 20352 12232 20404 12238
rect 20352 12174 20404 12180
rect 20076 12164 20128 12170
rect 20076 12106 20128 12112
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 20088 11218 20116 12106
rect 20364 11762 20392 12174
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 20352 11620 20404 11626
rect 20352 11562 20404 11568
rect 20260 11552 20312 11558
rect 20260 11494 20312 11500
rect 20076 11212 20128 11218
rect 20076 11154 20128 11160
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 19708 11076 19760 11082
rect 19708 11018 19760 11024
rect 19720 10538 19748 11018
rect 19708 10532 19760 10538
rect 19708 10474 19760 10480
rect 19524 9920 19576 9926
rect 19524 9862 19576 9868
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 18880 8968 18932 8974
rect 18880 8910 18932 8916
rect 18748 8372 18828 8378
rect 18696 8366 18828 8372
rect 18708 8350 18828 8366
rect 18694 7848 18750 7857
rect 18694 7783 18750 7792
rect 18708 7478 18736 7783
rect 18696 7472 18748 7478
rect 18696 7414 18748 7420
rect 18800 6390 18828 8350
rect 18892 8022 18920 8910
rect 19064 8900 19116 8906
rect 19064 8842 19116 8848
rect 19076 8430 19104 8842
rect 19248 8832 19300 8838
rect 19248 8774 19300 8780
rect 19064 8424 19116 8430
rect 19064 8366 19116 8372
rect 19260 8362 19288 8774
rect 19248 8356 19300 8362
rect 19248 8298 19300 8304
rect 18880 8016 18932 8022
rect 18880 7958 18932 7964
rect 19156 7948 19208 7954
rect 19156 7890 19208 7896
rect 19064 7336 19116 7342
rect 19064 7278 19116 7284
rect 18880 7200 18932 7206
rect 18880 7142 18932 7148
rect 18972 7200 19024 7206
rect 18972 7142 19024 7148
rect 18696 6384 18748 6390
rect 18696 6326 18748 6332
rect 18788 6384 18840 6390
rect 18788 6326 18840 6332
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 18512 5772 18564 5778
rect 18512 5714 18564 5720
rect 18604 5568 18656 5574
rect 18604 5510 18656 5516
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 18144 5160 18196 5166
rect 18144 5102 18196 5108
rect 18512 5160 18564 5166
rect 18512 5102 18564 5108
rect 18144 5024 18196 5030
rect 18144 4966 18196 4972
rect 18156 4622 18184 4966
rect 18144 4616 18196 4622
rect 18144 4558 18196 4564
rect 18524 4570 18552 5102
rect 18616 4826 18644 5510
rect 18604 4820 18656 4826
rect 18604 4762 18656 4768
rect 18524 4542 18644 4570
rect 18282 4380 18578 4400
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 18282 4304 18578 4324
rect 18144 4208 18196 4214
rect 18144 4150 18196 4156
rect 18418 4176 18474 4185
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 17960 3392 18012 3398
rect 17960 3334 18012 3340
rect 17868 3188 17920 3194
rect 17868 3130 17920 3136
rect 17776 2644 17828 2650
rect 17776 2586 17828 2592
rect 17972 2582 18000 3334
rect 18156 2582 18184 4150
rect 18418 4111 18420 4120
rect 18472 4111 18474 4120
rect 18420 4082 18472 4088
rect 18616 3618 18644 4542
rect 18708 3738 18736 6326
rect 18788 6112 18840 6118
rect 18788 6054 18840 6060
rect 18696 3732 18748 3738
rect 18696 3674 18748 3680
rect 18524 3590 18644 3618
rect 18524 3380 18552 3590
rect 18524 3352 18644 3380
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 18616 3074 18644 3352
rect 18340 3046 18644 3074
rect 17960 2576 18012 2582
rect 17960 2518 18012 2524
rect 18144 2576 18196 2582
rect 18144 2518 18196 2524
rect 18340 2378 18368 3046
rect 17776 2372 17828 2378
rect 17776 2314 17828 2320
rect 18328 2372 18380 2378
rect 18328 2314 18380 2320
rect 17788 800 17816 2314
rect 18144 2304 18196 2310
rect 18144 2246 18196 2252
rect 18050 2000 18106 2009
rect 17960 1964 18012 1970
rect 18050 1935 18106 1944
rect 17960 1906 18012 1912
rect 17972 1601 18000 1906
rect 18064 1902 18092 1935
rect 18052 1896 18104 1902
rect 18052 1838 18104 1844
rect 17958 1592 18014 1601
rect 17958 1527 18014 1536
rect 18156 1170 18184 2246
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 18800 2106 18828 6054
rect 18892 4078 18920 7142
rect 18984 6934 19012 7142
rect 19076 7002 19104 7278
rect 19168 7177 19196 7890
rect 19248 7744 19300 7750
rect 19248 7686 19300 7692
rect 19154 7168 19210 7177
rect 19154 7103 19210 7112
rect 19064 6996 19116 7002
rect 19064 6938 19116 6944
rect 18972 6928 19024 6934
rect 18972 6870 19024 6876
rect 18984 6225 19012 6870
rect 19156 6860 19208 6866
rect 19156 6802 19208 6808
rect 19064 6656 19116 6662
rect 19064 6598 19116 6604
rect 18970 6216 19026 6225
rect 18970 6151 19026 6160
rect 18972 6112 19024 6118
rect 18972 6054 19024 6060
rect 18880 4072 18932 4078
rect 18880 4014 18932 4020
rect 18984 3482 19012 6054
rect 19076 5778 19104 6598
rect 19168 6322 19196 6802
rect 19156 6316 19208 6322
rect 19156 6258 19208 6264
rect 19154 6216 19210 6225
rect 19154 6151 19210 6160
rect 19064 5772 19116 5778
rect 19064 5714 19116 5720
rect 19064 5568 19116 5574
rect 19064 5510 19116 5516
rect 19076 3670 19104 5510
rect 19168 5273 19196 6151
rect 19154 5264 19210 5273
rect 19154 5199 19210 5208
rect 19260 4690 19288 7686
rect 19444 6746 19472 9590
rect 19536 9518 19564 9862
rect 19524 9512 19576 9518
rect 19524 9454 19576 9460
rect 19536 9081 19564 9454
rect 19616 9376 19668 9382
rect 19616 9318 19668 9324
rect 19800 9376 19852 9382
rect 19800 9318 19852 9324
rect 19522 9072 19578 9081
rect 19522 9007 19578 9016
rect 19628 7886 19656 9318
rect 19812 9178 19840 9318
rect 19800 9172 19852 9178
rect 19800 9114 19852 9120
rect 19616 7880 19668 7886
rect 19616 7822 19668 7828
rect 19904 7274 19932 11086
rect 20168 9920 20220 9926
rect 20168 9862 20220 9868
rect 20180 9110 20208 9862
rect 20272 9586 20300 11494
rect 20364 11286 20392 11562
rect 20352 11280 20404 11286
rect 20352 11222 20404 11228
rect 20364 10810 20392 11222
rect 20352 10804 20404 10810
rect 20352 10746 20404 10752
rect 20260 9580 20312 9586
rect 20260 9522 20312 9528
rect 20168 9104 20220 9110
rect 20168 9046 20220 9052
rect 20168 8288 20220 8294
rect 20168 8230 20220 8236
rect 20076 7948 20128 7954
rect 20076 7890 20128 7896
rect 19892 7268 19944 7274
rect 19892 7210 19944 7216
rect 19708 7200 19760 7206
rect 19708 7142 19760 7148
rect 19720 6798 19748 7142
rect 19352 6718 19472 6746
rect 19708 6792 19760 6798
rect 19708 6734 19760 6740
rect 19248 4684 19300 4690
rect 19248 4626 19300 4632
rect 19156 4480 19208 4486
rect 19156 4422 19208 4428
rect 19246 4448 19302 4457
rect 19064 3664 19116 3670
rect 19064 3606 19116 3612
rect 18892 3454 19012 3482
rect 18892 2990 18920 3454
rect 18972 3392 19024 3398
rect 18972 3334 19024 3340
rect 18880 2984 18932 2990
rect 18880 2926 18932 2932
rect 18984 2666 19012 3334
rect 19168 3058 19196 4422
rect 19246 4383 19302 4392
rect 19260 4282 19288 4383
rect 19248 4276 19300 4282
rect 19248 4218 19300 4224
rect 19352 4078 19380 6718
rect 19432 6384 19484 6390
rect 19432 6326 19484 6332
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 19248 3936 19300 3942
rect 19248 3878 19300 3884
rect 19156 3052 19208 3058
rect 19156 2994 19208 3000
rect 19260 2990 19288 3878
rect 19248 2984 19300 2990
rect 19444 2961 19472 6326
rect 19800 5568 19852 5574
rect 19800 5510 19852 5516
rect 19812 4826 19840 5510
rect 19800 4820 19852 4826
rect 19800 4762 19852 4768
rect 19524 4140 19576 4146
rect 19524 4082 19576 4088
rect 19536 3602 19564 4082
rect 20088 4010 20116 7890
rect 20180 7410 20208 8230
rect 20260 7744 20312 7750
rect 20260 7686 20312 7692
rect 20168 7404 20220 7410
rect 20168 7346 20220 7352
rect 20180 6934 20208 7346
rect 20168 6928 20220 6934
rect 20168 6870 20220 6876
rect 20168 5772 20220 5778
rect 20168 5714 20220 5720
rect 20180 5234 20208 5714
rect 20168 5228 20220 5234
rect 20168 5170 20220 5176
rect 20076 4004 20128 4010
rect 20076 3946 20128 3952
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 19984 3460 20036 3466
rect 19984 3402 20036 3408
rect 19248 2926 19300 2932
rect 19430 2952 19486 2961
rect 19064 2916 19116 2922
rect 19430 2887 19486 2896
rect 19524 2916 19576 2922
rect 19064 2858 19116 2864
rect 19524 2858 19576 2864
rect 18892 2638 19012 2666
rect 18892 2446 18920 2638
rect 18880 2440 18932 2446
rect 18880 2382 18932 2388
rect 18788 2100 18840 2106
rect 18788 2042 18840 2048
rect 18604 1420 18656 1426
rect 18604 1362 18656 1368
rect 18156 1142 18276 1170
rect 18248 800 18276 1142
rect 18616 800 18644 1362
rect 18788 1352 18840 1358
rect 18788 1294 18840 1300
rect 18800 1057 18828 1294
rect 18786 1048 18842 1057
rect 18786 983 18842 992
rect 19076 800 19104 2858
rect 19246 2816 19302 2825
rect 19246 2751 19302 2760
rect 19156 2576 19208 2582
rect 19154 2544 19156 2553
rect 19208 2544 19210 2553
rect 19260 2514 19288 2751
rect 19154 2479 19210 2488
rect 19248 2508 19300 2514
rect 19168 2038 19196 2479
rect 19248 2450 19300 2456
rect 19156 2032 19208 2038
rect 19156 1974 19208 1980
rect 19536 800 19564 2858
rect 19996 800 20024 3402
rect 20272 2514 20300 7686
rect 20456 7546 20484 18158
rect 20444 7540 20496 7546
rect 20444 7482 20496 7488
rect 20456 5846 20484 7482
rect 20444 5840 20496 5846
rect 20444 5782 20496 5788
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 20364 5166 20392 5646
rect 20548 5250 20576 18702
rect 21192 18426 21220 18770
rect 21364 18692 21416 18698
rect 21364 18634 21416 18640
rect 21376 18465 21404 18634
rect 21362 18456 21418 18465
rect 21180 18420 21232 18426
rect 21362 18391 21418 18400
rect 21180 18362 21232 18368
rect 21364 18148 21416 18154
rect 21364 18090 21416 18096
rect 21376 18057 21404 18090
rect 21362 18048 21418 18057
rect 21362 17983 21418 17992
rect 21180 17740 21232 17746
rect 21180 17682 21232 17688
rect 20812 17604 20864 17610
rect 20812 17546 20864 17552
rect 20824 17513 20852 17546
rect 20810 17504 20866 17513
rect 20810 17439 20866 17448
rect 21192 17338 21220 17682
rect 21364 17604 21416 17610
rect 21364 17546 21416 17552
rect 21180 17332 21232 17338
rect 21180 17274 21232 17280
rect 20628 17128 20680 17134
rect 21376 17105 21404 17546
rect 20628 17070 20680 17076
rect 21362 17096 21418 17105
rect 20640 16182 20668 17070
rect 21362 17031 21418 17040
rect 21272 16992 21324 16998
rect 21272 16934 21324 16940
rect 21180 16788 21232 16794
rect 21180 16730 21232 16736
rect 20628 16176 20680 16182
rect 20628 16118 20680 16124
rect 20810 15600 20866 15609
rect 20810 15535 20812 15544
rect 20864 15535 20866 15544
rect 20812 15506 20864 15512
rect 20812 14476 20864 14482
rect 20812 14418 20864 14424
rect 20824 14074 20852 14418
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 21192 13870 21220 16730
rect 21284 16561 21312 16934
rect 21364 16652 21416 16658
rect 21364 16594 21416 16600
rect 21270 16552 21326 16561
rect 21270 16487 21326 16496
rect 21376 16153 21404 16594
rect 21362 16144 21418 16153
rect 21362 16079 21418 16088
rect 21272 15360 21324 15366
rect 21272 15302 21324 15308
rect 21284 14657 21312 15302
rect 22008 15224 22060 15230
rect 22006 15192 22008 15201
rect 22060 15192 22062 15201
rect 22006 15127 22062 15136
rect 21364 14884 21416 14890
rect 21364 14826 21416 14832
rect 21270 14648 21326 14657
rect 21270 14583 21326 14592
rect 21376 14249 21404 14826
rect 21456 14340 21508 14346
rect 21456 14282 21508 14288
rect 21362 14240 21418 14249
rect 21362 14175 21418 14184
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 21180 13864 21232 13870
rect 21180 13806 21232 13812
rect 21364 13864 21416 13870
rect 21468 13841 21496 14282
rect 21364 13806 21416 13812
rect 21454 13832 21510 13841
rect 20640 13462 20668 13806
rect 20628 13456 20680 13462
rect 20628 13398 20680 13404
rect 20994 13424 21050 13433
rect 20994 13359 21050 13368
rect 21008 12918 21036 13359
rect 21376 13297 21404 13806
rect 21454 13767 21510 13776
rect 21362 13288 21418 13297
rect 21088 13252 21140 13258
rect 21362 13223 21418 13232
rect 21088 13194 21140 13200
rect 20904 12912 20956 12918
rect 20904 12854 20956 12860
rect 20996 12912 21048 12918
rect 20996 12854 21048 12860
rect 20628 12776 20680 12782
rect 20628 12718 20680 12724
rect 20640 12345 20668 12718
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20732 12481 20760 12582
rect 20718 12472 20774 12481
rect 20718 12407 20774 12416
rect 20626 12336 20682 12345
rect 20626 12271 20682 12280
rect 20732 11762 20760 12407
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20824 11642 20852 12242
rect 20916 11694 20944 12854
rect 21100 12753 21128 13194
rect 21086 12744 21142 12753
rect 21086 12679 21142 12688
rect 21272 12708 21324 12714
rect 21272 12650 21324 12656
rect 21284 12209 21312 12650
rect 22008 12504 22060 12510
rect 22008 12446 22060 12452
rect 21270 12200 21326 12209
rect 21270 12135 21326 12144
rect 20732 11614 20852 11642
rect 20904 11688 20956 11694
rect 20904 11630 20956 11636
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20640 10266 20668 11290
rect 20628 10260 20680 10266
rect 20628 10202 20680 10208
rect 20732 8922 20760 11614
rect 21284 11393 21312 12135
rect 22020 11937 22048 12446
rect 22006 11928 22062 11937
rect 22006 11863 22062 11872
rect 21270 11384 21326 11393
rect 21270 11319 21326 11328
rect 22008 11076 22060 11082
rect 22008 11018 22060 11024
rect 21364 11008 21416 11014
rect 21364 10950 21416 10956
rect 21272 10532 21324 10538
rect 21272 10474 21324 10480
rect 21088 10192 21140 10198
rect 21088 10134 21140 10140
rect 20812 10056 20864 10062
rect 20812 9998 20864 10004
rect 20824 9586 20852 9998
rect 21100 9654 21128 10134
rect 21284 10033 21312 10474
rect 21376 10062 21404 10950
rect 22020 10441 22048 11018
rect 22006 10432 22062 10441
rect 22006 10367 22062 10376
rect 21364 10056 21416 10062
rect 21270 10024 21326 10033
rect 21364 9998 21416 10004
rect 21270 9959 21326 9968
rect 21088 9648 21140 9654
rect 21088 9590 21140 9596
rect 20812 9580 20864 9586
rect 20812 9522 20864 9528
rect 20824 9110 20852 9522
rect 21270 9480 21326 9489
rect 21270 9415 21272 9424
rect 21324 9415 21326 9424
rect 21272 9386 21324 9392
rect 20812 9104 20864 9110
rect 20812 9046 20864 9052
rect 21180 8968 21232 8974
rect 20732 8894 20852 8922
rect 21180 8910 21232 8916
rect 20720 8356 20772 8362
rect 20720 8298 20772 8304
rect 20732 8129 20760 8298
rect 20718 8120 20774 8129
rect 20718 8055 20774 8064
rect 20720 8016 20772 8022
rect 20720 7958 20772 7964
rect 20732 7721 20760 7958
rect 20718 7712 20774 7721
rect 20718 7647 20774 7656
rect 20626 5808 20682 5817
rect 20626 5743 20628 5752
rect 20680 5743 20682 5752
rect 20628 5714 20680 5720
rect 20456 5222 20576 5250
rect 20352 5160 20404 5166
rect 20352 5102 20404 5108
rect 20456 4486 20484 5222
rect 20536 5024 20588 5030
rect 20536 4966 20588 4972
rect 20548 4622 20576 4966
rect 20536 4616 20588 4622
rect 20536 4558 20588 4564
rect 20444 4480 20496 4486
rect 20444 4422 20496 4428
rect 20548 4078 20576 4558
rect 20536 4072 20588 4078
rect 20536 4014 20588 4020
rect 20640 3738 20668 5714
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 20536 3528 20588 3534
rect 20534 3496 20536 3505
rect 20588 3496 20590 3505
rect 20534 3431 20590 3440
rect 20444 3120 20496 3126
rect 20444 3062 20496 3068
rect 20260 2508 20312 2514
rect 20260 2450 20312 2456
rect 20456 800 20484 3062
rect 20824 2514 20852 8894
rect 21192 6866 21220 8910
rect 21270 8664 21326 8673
rect 21270 8599 21326 8608
rect 21284 8430 21312 8599
rect 21272 8424 21324 8430
rect 21272 8366 21324 8372
rect 21284 7546 21312 8366
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 21272 7336 21324 7342
rect 21272 7278 21324 7284
rect 21180 6860 21232 6866
rect 21180 6802 21232 6808
rect 21088 6656 21140 6662
rect 21088 6598 21140 6604
rect 21100 6254 21128 6598
rect 21088 6248 21140 6254
rect 21088 6190 21140 6196
rect 21192 6186 21220 6802
rect 21284 6225 21312 7278
rect 22008 6928 22060 6934
rect 22008 6870 22060 6876
rect 22020 6769 22048 6870
rect 22006 6760 22062 6769
rect 22006 6695 22062 6704
rect 21270 6216 21326 6225
rect 21180 6180 21232 6186
rect 21270 6151 21326 6160
rect 21180 6122 21232 6128
rect 21192 5370 21220 6122
rect 21180 5364 21232 5370
rect 21180 5306 21232 5312
rect 21086 4584 21142 4593
rect 21086 4519 21088 4528
rect 21140 4519 21142 4528
rect 21088 4490 21140 4496
rect 21192 4146 21220 5306
rect 21364 5024 21416 5030
rect 21364 4966 21416 4972
rect 21376 4865 21404 4966
rect 21362 4856 21418 4865
rect 21362 4791 21418 4800
rect 21376 4758 21404 4791
rect 21364 4752 21416 4758
rect 21364 4694 21416 4700
rect 21180 4140 21232 4146
rect 21180 4082 21232 4088
rect 21824 4004 21876 4010
rect 21824 3946 21876 3952
rect 20904 2848 20956 2854
rect 20904 2790 20956 2796
rect 20812 2508 20864 2514
rect 20812 2450 20864 2456
rect 20536 2440 20588 2446
rect 20536 2382 20588 2388
rect 20548 2310 20576 2382
rect 20536 2304 20588 2310
rect 20536 2246 20588 2252
rect 17682 232 17738 241
rect 17682 167 17738 176
rect 17774 0 17830 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 19062 0 19118 800
rect 19522 0 19578 800
rect 19982 0 20038 800
rect 20442 0 20498 800
rect 20548 649 20576 2246
rect 20916 800 20944 2790
rect 21364 1488 21416 1494
rect 21364 1430 21416 1436
rect 21376 800 21404 1430
rect 21836 800 21864 3946
rect 22744 2984 22796 2990
rect 22744 2926 22796 2932
rect 22284 2372 22336 2378
rect 22284 2314 22336 2320
rect 22296 800 22324 2314
rect 22756 800 22784 2926
rect 20534 640 20590 649
rect 20534 575 20590 584
rect 20902 0 20958 800
rect 21362 0 21418 800
rect 21822 0 21878 800
rect 22282 0 22338 800
rect 22742 0 22798 800
<< via2 >>
rect 4158 22616 4214 22672
rect 4066 22208 4122 22264
rect 3238 21664 3294 21720
rect 2778 21256 2834 21312
rect 2226 20712 2282 20768
rect 20258 22616 20314 22672
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 18602 21664 18658 21720
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 18970 21256 19026 21312
rect 19522 20712 19578 20768
rect 20534 22208 20590 22264
rect 1582 20340 1584 20360
rect 1584 20340 1636 20360
rect 1636 20340 1638 20360
rect 1582 20304 1638 20340
rect 1582 19780 1638 19816
rect 1582 19760 1584 19780
rect 1584 19760 1636 19780
rect 1636 19760 1638 19780
rect 1582 19352 1638 19408
rect 1582 18828 1638 18864
rect 1582 18808 1584 18828
rect 1584 18808 1636 18828
rect 1636 18808 1638 18828
rect 2226 18420 2282 18456
rect 2226 18400 2228 18420
rect 2228 18400 2280 18420
rect 2280 18400 2282 18420
rect 1674 18028 1676 18048
rect 1676 18028 1728 18048
rect 1728 18028 1730 18048
rect 1674 17992 1730 18028
rect 1674 17484 1676 17504
rect 1676 17484 1728 17504
rect 1728 17484 1730 17504
rect 1674 17448 1730 17484
rect 1582 17076 1584 17096
rect 1584 17076 1636 17096
rect 1636 17076 1638 17096
rect 1582 17040 1638 17076
rect 1582 16496 1638 16552
rect 1582 16108 1638 16144
rect 1582 16088 1584 16108
rect 1584 16088 1636 16108
rect 1636 16088 1638 16108
rect 2134 15580 2136 15600
rect 2136 15580 2188 15600
rect 2188 15580 2190 15600
rect 2134 15544 2190 15580
rect 1674 15136 1730 15192
rect 1674 14592 1730 14648
rect 1674 14220 1676 14240
rect 1676 14220 1728 14240
rect 1728 14220 1730 14240
rect 1674 14184 1730 14220
rect 1582 13812 1584 13832
rect 1584 13812 1636 13832
rect 1636 13812 1638 13832
rect 1582 13776 1638 13812
rect 1582 13252 1638 13288
rect 1582 13232 1584 13252
rect 1584 13232 1636 13252
rect 1636 13232 1638 13252
rect 1398 12824 1454 12880
rect 1674 12316 1676 12336
rect 1676 12316 1728 12336
rect 1728 12316 1730 12336
rect 1674 12280 1730 12316
rect 1674 11872 1730 11928
rect 1674 11328 1730 11384
rect 1674 10376 1730 10432
rect 1674 9968 1730 10024
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 1582 9460 1584 9480
rect 1584 9460 1636 9480
rect 1636 9460 1638 9480
rect 1582 9424 1638 9460
rect 1490 8608 1546 8664
rect 1858 7248 1914 7304
rect 1674 6296 1730 6352
rect 1582 6160 1638 6216
rect 2318 6704 2374 6760
rect 1766 5888 1822 5944
rect 1674 5788 1676 5808
rect 1676 5788 1728 5808
rect 1728 5788 1730 5808
rect 1674 5752 1730 5788
rect 1582 5072 1638 5128
rect 2226 5344 2282 5400
rect 1766 4800 1822 4856
rect 2042 4664 2098 4720
rect 1858 4392 1914 4448
rect 1398 3848 1454 3904
rect 1858 992 1914 1048
rect 2778 6996 2834 7032
rect 2778 6976 2780 6996
rect 2780 6976 2832 6996
rect 2832 6976 2834 6996
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 4434 12144 4490 12200
rect 3698 11736 3754 11792
rect 4066 11736 4122 11792
rect 3330 10920 3386 10976
rect 3238 8200 3294 8256
rect 3422 7928 3478 7984
rect 3422 7656 3478 7712
rect 3330 7112 3386 7168
rect 3238 5208 3294 5264
rect 2870 3440 2926 3496
rect 2962 3032 3018 3088
rect 3330 1572 3332 1592
rect 3332 1572 3384 1592
rect 3384 1572 3386 1592
rect 3330 1536 3386 1572
rect 3698 7792 3754 7848
rect 3606 4392 3662 4448
rect 3514 3460 3570 3496
rect 3514 3440 3516 3460
rect 3516 3440 3568 3460
rect 3568 3440 3570 3460
rect 3790 5344 3846 5400
rect 3698 1944 3754 2000
rect 4066 9016 4122 9072
rect 4066 8064 4122 8120
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 3974 2488 4030 2544
rect 3422 176 3478 232
rect 4066 584 4122 640
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 4618 8336 4674 8392
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 4250 4528 4306 4584
rect 4250 2932 4252 2952
rect 4252 2932 4304 2952
rect 4304 2932 4306 2952
rect 4250 2896 4306 2932
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 4802 4256 4858 4312
rect 5722 7928 5778 7984
rect 4434 4120 4490 4176
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 5262 5344 5318 5400
rect 5262 4800 5318 4856
rect 5538 4800 5594 4856
rect 5722 5480 5778 5536
rect 7102 12708 7158 12744
rect 7102 12688 7104 12708
rect 7104 12688 7156 12708
rect 7156 12688 7158 12708
rect 6090 6976 6146 7032
rect 5446 3304 5502 3360
rect 5814 3304 5870 3360
rect 5814 2932 5816 2952
rect 5816 2932 5868 2952
rect 5868 2932 5870 2952
rect 5814 2896 5870 2932
rect 6458 6296 6514 6352
rect 7102 8472 7158 8528
rect 6458 6160 6514 6216
rect 6826 5888 6882 5944
rect 6642 5616 6698 5672
rect 6550 4120 6606 4176
rect 6734 4156 6736 4176
rect 6736 4156 6788 4176
rect 6788 4156 6790 4176
rect 6734 4120 6790 4156
rect 7194 6160 7250 6216
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 7930 11772 7932 11792
rect 7932 11772 7984 11792
rect 7984 11772 7986 11792
rect 7930 11736 7986 11772
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 8390 12708 8446 12744
rect 8390 12688 8392 12708
rect 8392 12688 8444 12708
rect 8444 12688 8446 12708
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 8022 8492 8078 8528
rect 8022 8472 8024 8492
rect 8024 8472 8076 8492
rect 8076 8472 8078 8492
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 8666 8336 8722 8392
rect 8574 8200 8630 8256
rect 8390 7812 8446 7848
rect 8390 7792 8392 7812
rect 8392 7792 8444 7812
rect 8444 7792 8446 7812
rect 8298 4700 8300 4720
rect 8300 4700 8352 4720
rect 8352 4700 8354 4720
rect 8298 4664 8354 4700
rect 9126 7284 9128 7304
rect 9128 7284 9180 7304
rect 9180 7284 9182 7304
rect 9126 7248 9182 7284
rect 8942 5344 8998 5400
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 9586 12144 9642 12200
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 10230 13404 10232 13424
rect 10232 13404 10284 13424
rect 10284 13404 10286 13424
rect 10230 13368 10286 13404
rect 9678 9560 9734 9616
rect 9494 8200 9550 8256
rect 9402 5616 9458 5672
rect 9218 3032 9274 3088
rect 9954 8744 10010 8800
rect 10230 11600 10286 11656
rect 10414 11600 10470 11656
rect 9862 4120 9918 4176
rect 9770 3576 9826 3632
rect 10414 8880 10470 8936
rect 10322 8492 10378 8528
rect 10322 8472 10324 8492
rect 10324 8472 10376 8492
rect 10376 8472 10378 8492
rect 10322 6160 10378 6216
rect 10230 5480 10286 5536
rect 10506 4528 10562 4584
rect 10874 16668 10876 16688
rect 10876 16668 10928 16688
rect 10928 16668 10930 16688
rect 10874 16632 10930 16668
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 10966 13404 10968 13424
rect 10968 13404 11020 13424
rect 11020 13404 11022 13424
rect 10966 13368 11022 13404
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 10690 9424 10746 9480
rect 10322 3984 10378 4040
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 10874 8744 10930 8800
rect 11794 9596 11796 9616
rect 11796 9596 11848 9616
rect 11848 9596 11850 9616
rect 11794 9560 11850 9596
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 12346 7792 12402 7848
rect 11150 3884 11152 3904
rect 11152 3884 11204 3904
rect 11204 3884 11206 3904
rect 11150 3848 11206 3884
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 15106 17740 15162 17776
rect 15566 17756 15568 17776
rect 15568 17756 15620 17776
rect 15620 17756 15622 17776
rect 15106 17720 15108 17740
rect 15108 17720 15160 17740
rect 15160 17720 15162 17740
rect 15566 17720 15622 17756
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 13082 8472 13138 8528
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 16026 12416 16082 12472
rect 16302 12280 16358 12336
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 13542 5208 13598 5264
rect 12898 3440 12954 3496
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 15106 6740 15108 6760
rect 15108 6740 15160 6760
rect 15160 6740 15162 6760
rect 15106 6704 15162 6740
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 14646 5072 14702 5128
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 15474 9560 15530 9616
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 16118 7384 16174 7440
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 16578 12688 16634 12744
rect 17038 13368 17094 13424
rect 16394 4120 16450 4176
rect 15934 3576 15990 3632
rect 17222 13268 17224 13288
rect 17224 13268 17276 13288
rect 17276 13268 17278 13288
rect 17222 13232 17278 13268
rect 16946 9460 16948 9480
rect 16948 9460 17000 9480
rect 17000 9460 17002 9480
rect 16946 9424 17002 9460
rect 17958 12824 18014 12880
rect 17866 11736 17922 11792
rect 17038 6704 17094 6760
rect 16946 5208 17002 5264
rect 17774 8200 17830 8256
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 18418 12552 18474 12608
rect 20810 20324 20866 20360
rect 20810 20304 20812 20324
rect 20812 20304 20864 20324
rect 20864 20304 20866 20324
rect 21454 19760 21510 19816
rect 21362 19352 21418 19408
rect 21362 18808 21418 18864
rect 18786 12300 18842 12336
rect 18786 12280 18788 12300
rect 18788 12280 18840 12300
rect 18840 12280 18842 12300
rect 18602 12144 18658 12200
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 18694 11464 18750 11520
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 18326 7420 18328 7440
rect 18328 7420 18380 7440
rect 18380 7420 18382 7440
rect 18326 7384 18382 7420
rect 17866 3848 17922 3904
rect 17866 3576 17922 3632
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 19154 11736 19210 11792
rect 19062 11500 19064 11520
rect 19064 11500 19116 11520
rect 19116 11500 19118 11520
rect 19062 11464 19118 11500
rect 19062 10920 19118 10976
rect 19522 13232 19578 13288
rect 19706 12588 19708 12608
rect 19708 12588 19760 12608
rect 19760 12588 19762 12608
rect 19706 12552 19762 12588
rect 18694 7792 18750 7848
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 18418 4140 18474 4176
rect 18418 4120 18420 4140
rect 18420 4120 18472 4140
rect 18472 4120 18474 4140
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 18050 1944 18106 2000
rect 17958 1536 18014 1592
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 19154 7112 19210 7168
rect 18970 6160 19026 6216
rect 19154 6160 19210 6216
rect 19154 5208 19210 5264
rect 19522 9016 19578 9072
rect 19246 4392 19302 4448
rect 19430 2896 19486 2952
rect 18786 992 18842 1048
rect 19246 2760 19302 2816
rect 19154 2524 19156 2544
rect 19156 2524 19208 2544
rect 19208 2524 19210 2544
rect 19154 2488 19210 2524
rect 21362 18400 21418 18456
rect 21362 17992 21418 18048
rect 20810 17448 20866 17504
rect 21362 17040 21418 17096
rect 20810 15564 20866 15600
rect 20810 15544 20812 15564
rect 20812 15544 20864 15564
rect 20864 15544 20866 15564
rect 21270 16496 21326 16552
rect 21362 16088 21418 16144
rect 22006 15172 22008 15192
rect 22008 15172 22060 15192
rect 22060 15172 22062 15192
rect 22006 15136 22062 15172
rect 21270 14592 21326 14648
rect 21362 14184 21418 14240
rect 20994 13368 21050 13424
rect 21454 13776 21510 13832
rect 21362 13232 21418 13288
rect 20718 12416 20774 12472
rect 20626 12280 20682 12336
rect 21086 12688 21142 12744
rect 21270 12144 21326 12200
rect 22006 11872 22062 11928
rect 21270 11328 21326 11384
rect 22006 10376 22062 10432
rect 21270 9968 21326 10024
rect 21270 9444 21326 9480
rect 21270 9424 21272 9444
rect 21272 9424 21324 9444
rect 21324 9424 21326 9444
rect 20718 8064 20774 8120
rect 20718 7656 20774 7712
rect 20626 5772 20682 5808
rect 20626 5752 20628 5772
rect 20628 5752 20680 5772
rect 20680 5752 20682 5772
rect 20534 3476 20536 3496
rect 20536 3476 20588 3496
rect 20588 3476 20590 3496
rect 20534 3440 20590 3476
rect 21270 8608 21326 8664
rect 22006 6704 22062 6760
rect 21270 6160 21326 6216
rect 21086 4548 21142 4584
rect 21086 4528 21088 4548
rect 21088 4528 21140 4548
rect 21140 4528 21142 4548
rect 21362 4800 21418 4856
rect 17682 176 17738 232
rect 20534 584 20590 640
<< metal3 >>
rect 0 22674 800 22704
rect 4153 22674 4219 22677
rect 0 22672 4219 22674
rect 0 22616 4158 22672
rect 4214 22616 4219 22672
rect 0 22614 4219 22616
rect 0 22584 800 22614
rect 4153 22611 4219 22614
rect 20253 22674 20319 22677
rect 22200 22674 23000 22704
rect 20253 22672 23000 22674
rect 20253 22616 20258 22672
rect 20314 22616 23000 22672
rect 20253 22614 23000 22616
rect 20253 22611 20319 22614
rect 22200 22584 23000 22614
rect 0 22266 800 22296
rect 4061 22266 4127 22269
rect 0 22264 4127 22266
rect 0 22208 4066 22264
rect 4122 22208 4127 22264
rect 0 22206 4127 22208
rect 0 22176 800 22206
rect 4061 22203 4127 22206
rect 20529 22266 20595 22269
rect 22200 22266 23000 22296
rect 20529 22264 23000 22266
rect 20529 22208 20534 22264
rect 20590 22208 23000 22264
rect 20529 22206 23000 22208
rect 20529 22203 20595 22206
rect 22200 22176 23000 22206
rect 0 21722 800 21752
rect 3233 21722 3299 21725
rect 0 21720 3299 21722
rect 0 21664 3238 21720
rect 3294 21664 3299 21720
rect 0 21662 3299 21664
rect 0 21632 800 21662
rect 3233 21659 3299 21662
rect 18597 21722 18663 21725
rect 22200 21722 23000 21752
rect 18597 21720 23000 21722
rect 18597 21664 18602 21720
rect 18658 21664 23000 21720
rect 18597 21662 23000 21664
rect 18597 21659 18663 21662
rect 22200 21632 23000 21662
rect 0 21314 800 21344
rect 2773 21314 2839 21317
rect 0 21312 2839 21314
rect 0 21256 2778 21312
rect 2834 21256 2839 21312
rect 0 21254 2839 21256
rect 0 21224 800 21254
rect 2773 21251 2839 21254
rect 18965 21314 19031 21317
rect 22200 21314 23000 21344
rect 18965 21312 23000 21314
rect 18965 21256 18970 21312
rect 19026 21256 23000 21312
rect 18965 21254 23000 21256
rect 18965 21251 19031 21254
rect 22200 21224 23000 21254
rect 0 20770 800 20800
rect 2221 20770 2287 20773
rect 0 20768 2287 20770
rect 0 20712 2226 20768
rect 2282 20712 2287 20768
rect 0 20710 2287 20712
rect 0 20680 800 20710
rect 2221 20707 2287 20710
rect 19517 20770 19583 20773
rect 22200 20770 23000 20800
rect 19517 20768 23000 20770
rect 19517 20712 19522 20768
rect 19578 20712 23000 20768
rect 19517 20710 23000 20712
rect 19517 20707 19583 20710
rect 4409 20704 4729 20705
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 22200 20680 23000 20710
rect 18270 20639 18590 20640
rect 0 20362 800 20392
rect 1577 20362 1643 20365
rect 0 20360 1643 20362
rect 0 20304 1582 20360
rect 1638 20304 1643 20360
rect 0 20302 1643 20304
rect 0 20272 800 20302
rect 1577 20299 1643 20302
rect 20805 20362 20871 20365
rect 22200 20362 23000 20392
rect 20805 20360 23000 20362
rect 20805 20304 20810 20360
rect 20866 20304 23000 20360
rect 20805 20302 23000 20304
rect 20805 20299 20871 20302
rect 22200 20272 23000 20302
rect 7874 20160 8194 20161
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 20095 15125 20096
rect 0 19818 800 19848
rect 1577 19818 1643 19821
rect 0 19816 1643 19818
rect 0 19760 1582 19816
rect 1638 19760 1643 19816
rect 0 19758 1643 19760
rect 0 19728 800 19758
rect 1577 19755 1643 19758
rect 21449 19818 21515 19821
rect 22200 19818 23000 19848
rect 21449 19816 23000 19818
rect 21449 19760 21454 19816
rect 21510 19760 23000 19816
rect 21449 19758 23000 19760
rect 21449 19755 21515 19758
rect 22200 19728 23000 19758
rect 4409 19616 4729 19617
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 19551 18590 19552
rect 0 19410 800 19440
rect 1577 19410 1643 19413
rect 0 19408 1643 19410
rect 0 19352 1582 19408
rect 1638 19352 1643 19408
rect 0 19350 1643 19352
rect 0 19320 800 19350
rect 1577 19347 1643 19350
rect 21357 19410 21423 19413
rect 22200 19410 23000 19440
rect 21357 19408 23000 19410
rect 21357 19352 21362 19408
rect 21418 19352 23000 19408
rect 21357 19350 23000 19352
rect 21357 19347 21423 19350
rect 22200 19320 23000 19350
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 19007 15125 19008
rect 0 18866 800 18896
rect 1577 18866 1643 18869
rect 0 18864 1643 18866
rect 0 18808 1582 18864
rect 1638 18808 1643 18864
rect 0 18806 1643 18808
rect 0 18776 800 18806
rect 1577 18803 1643 18806
rect 21357 18866 21423 18869
rect 22200 18866 23000 18896
rect 21357 18864 23000 18866
rect 21357 18808 21362 18864
rect 21418 18808 23000 18864
rect 21357 18806 23000 18808
rect 21357 18803 21423 18806
rect 22200 18776 23000 18806
rect 4409 18528 4729 18529
rect 0 18458 800 18488
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 18463 18590 18464
rect 2221 18458 2287 18461
rect 0 18456 2287 18458
rect 0 18400 2226 18456
rect 2282 18400 2287 18456
rect 0 18398 2287 18400
rect 0 18368 800 18398
rect 2221 18395 2287 18398
rect 21357 18458 21423 18461
rect 22200 18458 23000 18488
rect 21357 18456 23000 18458
rect 21357 18400 21362 18456
rect 21418 18400 23000 18456
rect 21357 18398 23000 18400
rect 21357 18395 21423 18398
rect 22200 18368 23000 18398
rect 0 18050 800 18080
rect 1669 18050 1735 18053
rect 0 18048 1735 18050
rect 0 17992 1674 18048
rect 1730 17992 1735 18048
rect 0 17990 1735 17992
rect 0 17960 800 17990
rect 1669 17987 1735 17990
rect 21357 18050 21423 18053
rect 22200 18050 23000 18080
rect 21357 18048 23000 18050
rect 21357 17992 21362 18048
rect 21418 17992 23000 18048
rect 21357 17990 23000 17992
rect 21357 17987 21423 17990
rect 7874 17984 8194 17985
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 22200 17960 23000 17990
rect 14805 17919 15125 17920
rect 15101 17778 15167 17781
rect 15561 17778 15627 17781
rect 15101 17776 15627 17778
rect 15101 17720 15106 17776
rect 15162 17720 15566 17776
rect 15622 17720 15627 17776
rect 15101 17718 15627 17720
rect 15101 17715 15167 17718
rect 15561 17715 15627 17718
rect 0 17506 800 17536
rect 1669 17506 1735 17509
rect 0 17504 1735 17506
rect 0 17448 1674 17504
rect 1730 17448 1735 17504
rect 0 17446 1735 17448
rect 0 17416 800 17446
rect 1669 17443 1735 17446
rect 20805 17506 20871 17509
rect 22200 17506 23000 17536
rect 20805 17504 23000 17506
rect 20805 17448 20810 17504
rect 20866 17448 23000 17504
rect 20805 17446 23000 17448
rect 20805 17443 20871 17446
rect 4409 17440 4729 17441
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 22200 17416 23000 17446
rect 18270 17375 18590 17376
rect 0 17098 800 17128
rect 1577 17098 1643 17101
rect 0 17096 1643 17098
rect 0 17040 1582 17096
rect 1638 17040 1643 17096
rect 0 17038 1643 17040
rect 0 17008 800 17038
rect 1577 17035 1643 17038
rect 21357 17098 21423 17101
rect 22200 17098 23000 17128
rect 21357 17096 23000 17098
rect 21357 17040 21362 17096
rect 21418 17040 23000 17096
rect 21357 17038 23000 17040
rect 21357 17035 21423 17038
rect 22200 17008 23000 17038
rect 7874 16896 8194 16897
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 16831 15125 16832
rect 10726 16628 10732 16692
rect 10796 16690 10802 16692
rect 10869 16690 10935 16693
rect 10796 16688 10935 16690
rect 10796 16632 10874 16688
rect 10930 16632 10935 16688
rect 10796 16630 10935 16632
rect 10796 16628 10802 16630
rect 10869 16627 10935 16630
rect 0 16554 800 16584
rect 1577 16554 1643 16557
rect 0 16552 1643 16554
rect 0 16496 1582 16552
rect 1638 16496 1643 16552
rect 0 16494 1643 16496
rect 0 16464 800 16494
rect 1577 16491 1643 16494
rect 21265 16554 21331 16557
rect 22200 16554 23000 16584
rect 21265 16552 23000 16554
rect 21265 16496 21270 16552
rect 21326 16496 23000 16552
rect 21265 16494 23000 16496
rect 21265 16491 21331 16494
rect 22200 16464 23000 16494
rect 4409 16352 4729 16353
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 16287 18590 16288
rect 0 16146 800 16176
rect 1577 16146 1643 16149
rect 0 16144 1643 16146
rect 0 16088 1582 16144
rect 1638 16088 1643 16144
rect 0 16086 1643 16088
rect 0 16056 800 16086
rect 1577 16083 1643 16086
rect 21357 16146 21423 16149
rect 22200 16146 23000 16176
rect 21357 16144 23000 16146
rect 21357 16088 21362 16144
rect 21418 16088 23000 16144
rect 21357 16086 23000 16088
rect 21357 16083 21423 16086
rect 22200 16056 23000 16086
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 15743 15125 15744
rect 0 15602 800 15632
rect 2129 15602 2195 15605
rect 0 15600 2195 15602
rect 0 15544 2134 15600
rect 2190 15544 2195 15600
rect 0 15542 2195 15544
rect 0 15512 800 15542
rect 2129 15539 2195 15542
rect 20805 15602 20871 15605
rect 22200 15602 23000 15632
rect 20805 15600 23000 15602
rect 20805 15544 20810 15600
rect 20866 15544 23000 15600
rect 20805 15542 23000 15544
rect 20805 15539 20871 15542
rect 22200 15512 23000 15542
rect 4409 15264 4729 15265
rect 0 15194 800 15224
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 15199 18590 15200
rect 1669 15194 1735 15197
rect 0 15192 1735 15194
rect 0 15136 1674 15192
rect 1730 15136 1735 15192
rect 0 15134 1735 15136
rect 0 15104 800 15134
rect 1669 15131 1735 15134
rect 22001 15194 22067 15197
rect 22200 15194 23000 15224
rect 22001 15192 23000 15194
rect 22001 15136 22006 15192
rect 22062 15136 23000 15192
rect 22001 15134 23000 15136
rect 22001 15131 22067 15134
rect 22200 15104 23000 15134
rect 7874 14720 8194 14721
rect 0 14650 800 14680
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 1669 14650 1735 14653
rect 0 14648 1735 14650
rect 0 14592 1674 14648
rect 1730 14592 1735 14648
rect 0 14590 1735 14592
rect 0 14560 800 14590
rect 1669 14587 1735 14590
rect 21265 14650 21331 14653
rect 22200 14650 23000 14680
rect 21265 14648 23000 14650
rect 21265 14592 21270 14648
rect 21326 14592 23000 14648
rect 21265 14590 23000 14592
rect 21265 14587 21331 14590
rect 22200 14560 23000 14590
rect 0 14242 800 14272
rect 1669 14242 1735 14245
rect 0 14240 1735 14242
rect 0 14184 1674 14240
rect 1730 14184 1735 14240
rect 0 14182 1735 14184
rect 0 14152 800 14182
rect 1669 14179 1735 14182
rect 21357 14242 21423 14245
rect 22200 14242 23000 14272
rect 21357 14240 23000 14242
rect 21357 14184 21362 14240
rect 21418 14184 23000 14240
rect 21357 14182 23000 14184
rect 21357 14179 21423 14182
rect 4409 14176 4729 14177
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 22200 14152 23000 14182
rect 18270 14111 18590 14112
rect 0 13834 800 13864
rect 1577 13834 1643 13837
rect 0 13832 1643 13834
rect 0 13776 1582 13832
rect 1638 13776 1643 13832
rect 0 13774 1643 13776
rect 0 13744 800 13774
rect 1577 13771 1643 13774
rect 21449 13834 21515 13837
rect 22200 13834 23000 13864
rect 21449 13832 23000 13834
rect 21449 13776 21454 13832
rect 21510 13776 23000 13832
rect 21449 13774 23000 13776
rect 21449 13771 21515 13774
rect 22200 13744 23000 13774
rect 7874 13632 8194 13633
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 13567 15125 13568
rect 10225 13426 10291 13429
rect 10961 13426 11027 13429
rect 10225 13424 11027 13426
rect 10225 13368 10230 13424
rect 10286 13368 10966 13424
rect 11022 13368 11027 13424
rect 10225 13366 11027 13368
rect 10225 13363 10291 13366
rect 10961 13363 11027 13366
rect 17033 13426 17099 13429
rect 20989 13426 21055 13429
rect 17033 13424 21055 13426
rect 17033 13368 17038 13424
rect 17094 13368 20994 13424
rect 21050 13368 21055 13424
rect 17033 13366 21055 13368
rect 17033 13363 17099 13366
rect 20989 13363 21055 13366
rect 0 13290 800 13320
rect 1577 13290 1643 13293
rect 0 13288 1643 13290
rect 0 13232 1582 13288
rect 1638 13232 1643 13288
rect 0 13230 1643 13232
rect 0 13200 800 13230
rect 1577 13227 1643 13230
rect 17217 13290 17283 13293
rect 19517 13290 19583 13293
rect 17217 13288 19583 13290
rect 17217 13232 17222 13288
rect 17278 13232 19522 13288
rect 19578 13232 19583 13288
rect 17217 13230 19583 13232
rect 17217 13227 17283 13230
rect 19517 13227 19583 13230
rect 21357 13290 21423 13293
rect 22200 13290 23000 13320
rect 21357 13288 23000 13290
rect 21357 13232 21362 13288
rect 21418 13232 23000 13288
rect 21357 13230 23000 13232
rect 21357 13227 21423 13230
rect 22200 13200 23000 13230
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 13023 18590 13024
rect 0 12882 800 12912
rect 1393 12882 1459 12885
rect 0 12880 1459 12882
rect 0 12824 1398 12880
rect 1454 12824 1459 12880
rect 0 12822 1459 12824
rect 0 12792 800 12822
rect 1393 12819 1459 12822
rect 17953 12882 18019 12885
rect 22200 12882 23000 12912
rect 17953 12880 23000 12882
rect 17953 12824 17958 12880
rect 18014 12824 23000 12880
rect 17953 12822 23000 12824
rect 17953 12819 18019 12822
rect 22200 12792 23000 12822
rect 7097 12746 7163 12749
rect 8385 12746 8451 12749
rect 7097 12744 8451 12746
rect 7097 12688 7102 12744
rect 7158 12688 8390 12744
rect 8446 12688 8451 12744
rect 7097 12686 8451 12688
rect 7097 12683 7163 12686
rect 8385 12683 8451 12686
rect 16573 12746 16639 12749
rect 21081 12746 21147 12749
rect 16573 12744 21147 12746
rect 16573 12688 16578 12744
rect 16634 12688 21086 12744
rect 21142 12688 21147 12744
rect 16573 12686 21147 12688
rect 16573 12683 16639 12686
rect 21081 12683 21147 12686
rect 18413 12610 18479 12613
rect 19701 12610 19767 12613
rect 18413 12608 19767 12610
rect 18413 12552 18418 12608
rect 18474 12552 19706 12608
rect 19762 12552 19767 12608
rect 18413 12550 19767 12552
rect 18413 12547 18479 12550
rect 19701 12547 19767 12550
rect 7874 12544 8194 12545
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 12479 15125 12480
rect 16021 12474 16087 12477
rect 20713 12474 20779 12477
rect 16021 12472 20779 12474
rect 16021 12416 16026 12472
rect 16082 12416 20718 12472
rect 20774 12416 20779 12472
rect 16021 12414 20779 12416
rect 16021 12411 16087 12414
rect 20713 12411 20779 12414
rect 0 12338 800 12368
rect 1669 12338 1735 12341
rect 0 12336 1735 12338
rect 0 12280 1674 12336
rect 1730 12280 1735 12336
rect 0 12278 1735 12280
rect 0 12248 800 12278
rect 1669 12275 1735 12278
rect 16297 12338 16363 12341
rect 18781 12338 18847 12341
rect 16297 12336 18847 12338
rect 16297 12280 16302 12336
rect 16358 12280 18786 12336
rect 18842 12280 18847 12336
rect 16297 12278 18847 12280
rect 16297 12275 16363 12278
rect 18781 12275 18847 12278
rect 20621 12338 20687 12341
rect 22200 12338 23000 12368
rect 20621 12336 23000 12338
rect 20621 12280 20626 12336
rect 20682 12280 23000 12336
rect 20621 12278 23000 12280
rect 20621 12275 20687 12278
rect 22200 12248 23000 12278
rect 4429 12202 4495 12205
rect 9581 12202 9647 12205
rect 4429 12200 9647 12202
rect 4429 12144 4434 12200
rect 4490 12144 9586 12200
rect 9642 12144 9647 12200
rect 4429 12142 9647 12144
rect 4429 12139 4495 12142
rect 9581 12139 9647 12142
rect 18597 12202 18663 12205
rect 21265 12202 21331 12205
rect 18597 12200 21331 12202
rect 18597 12144 18602 12200
rect 18658 12144 21270 12200
rect 21326 12144 21331 12200
rect 18597 12142 21331 12144
rect 18597 12139 18663 12142
rect 21265 12139 21331 12142
rect 4409 12000 4729 12001
rect 0 11930 800 11960
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 11935 18590 11936
rect 1669 11930 1735 11933
rect 0 11928 1735 11930
rect 0 11872 1674 11928
rect 1730 11872 1735 11928
rect 0 11870 1735 11872
rect 0 11840 800 11870
rect 1669 11867 1735 11870
rect 22001 11930 22067 11933
rect 22200 11930 23000 11960
rect 22001 11928 23000 11930
rect 22001 11872 22006 11928
rect 22062 11872 23000 11928
rect 22001 11870 23000 11872
rect 22001 11867 22067 11870
rect 22200 11840 23000 11870
rect 3693 11794 3759 11797
rect 4061 11794 4127 11797
rect 7925 11794 7991 11797
rect 3693 11792 7991 11794
rect 3693 11736 3698 11792
rect 3754 11736 4066 11792
rect 4122 11736 7930 11792
rect 7986 11736 7991 11792
rect 3693 11734 7991 11736
rect 3693 11731 3759 11734
rect 4061 11731 4127 11734
rect 7925 11731 7991 11734
rect 17861 11794 17927 11797
rect 19149 11794 19215 11797
rect 17861 11792 19215 11794
rect 17861 11736 17866 11792
rect 17922 11736 19154 11792
rect 19210 11736 19215 11792
rect 17861 11734 19215 11736
rect 17861 11731 17927 11734
rect 19149 11731 19215 11734
rect 10225 11658 10291 11661
rect 10409 11658 10475 11661
rect 10225 11656 10475 11658
rect 10225 11600 10230 11656
rect 10286 11600 10414 11656
rect 10470 11600 10475 11656
rect 10225 11598 10475 11600
rect 10225 11595 10291 11598
rect 10409 11595 10475 11598
rect 18689 11522 18755 11525
rect 19057 11522 19123 11525
rect 18689 11520 19123 11522
rect 18689 11464 18694 11520
rect 18750 11464 19062 11520
rect 19118 11464 19123 11520
rect 18689 11462 19123 11464
rect 18689 11459 18755 11462
rect 19057 11459 19123 11462
rect 7874 11456 8194 11457
rect 0 11386 800 11416
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 11391 15125 11392
rect 1669 11386 1735 11389
rect 0 11384 1735 11386
rect 0 11328 1674 11384
rect 1730 11328 1735 11384
rect 0 11326 1735 11328
rect 0 11296 800 11326
rect 1669 11323 1735 11326
rect 21265 11386 21331 11389
rect 22200 11386 23000 11416
rect 21265 11384 23000 11386
rect 21265 11328 21270 11384
rect 21326 11328 23000 11384
rect 21265 11326 23000 11328
rect 21265 11323 21331 11326
rect 22200 11296 23000 11326
rect 0 10978 800 11008
rect 3325 10978 3391 10981
rect 0 10976 3391 10978
rect 0 10920 3330 10976
rect 3386 10920 3391 10976
rect 0 10918 3391 10920
rect 0 10888 800 10918
rect 3325 10915 3391 10918
rect 19057 10978 19123 10981
rect 22200 10978 23000 11008
rect 19057 10976 23000 10978
rect 19057 10920 19062 10976
rect 19118 10920 23000 10976
rect 19057 10918 23000 10920
rect 19057 10915 19123 10918
rect 4409 10912 4729 10913
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 22200 10888 23000 10918
rect 18270 10847 18590 10848
rect 0 10434 800 10464
rect 1669 10434 1735 10437
rect 0 10432 1735 10434
rect 0 10376 1674 10432
rect 1730 10376 1735 10432
rect 0 10374 1735 10376
rect 0 10344 800 10374
rect 1669 10371 1735 10374
rect 22001 10434 22067 10437
rect 22200 10434 23000 10464
rect 22001 10432 23000 10434
rect 22001 10376 22006 10432
rect 22062 10376 23000 10432
rect 22001 10374 23000 10376
rect 22001 10371 22067 10374
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 22200 10344 23000 10374
rect 14805 10303 15125 10304
rect 0 10026 800 10056
rect 1669 10026 1735 10029
rect 0 10024 1735 10026
rect 0 9968 1674 10024
rect 1730 9968 1735 10024
rect 0 9966 1735 9968
rect 0 9936 800 9966
rect 1669 9963 1735 9966
rect 21265 10026 21331 10029
rect 22200 10026 23000 10056
rect 21265 10024 23000 10026
rect 21265 9968 21270 10024
rect 21326 9968 23000 10024
rect 21265 9966 23000 9968
rect 21265 9963 21331 9966
rect 22200 9936 23000 9966
rect 4409 9824 4729 9825
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 9759 18590 9760
rect 9673 9618 9739 9621
rect 11789 9618 11855 9621
rect 15469 9618 15535 9621
rect 9673 9616 10978 9618
rect 9673 9560 9678 9616
rect 9734 9560 10978 9616
rect 9673 9558 10978 9560
rect 9673 9555 9739 9558
rect 0 9482 800 9512
rect 1577 9482 1643 9485
rect 10685 9482 10751 9485
rect 0 9480 1643 9482
rect 0 9424 1582 9480
rect 1638 9424 1643 9480
rect 0 9422 1643 9424
rect 0 9392 800 9422
rect 1577 9419 1643 9422
rect 10412 9480 10751 9482
rect 10412 9424 10690 9480
rect 10746 9424 10751 9480
rect 10412 9422 10751 9424
rect 10918 9482 10978 9558
rect 11789 9616 15535 9618
rect 11789 9560 11794 9616
rect 11850 9560 15474 9616
rect 15530 9560 15535 9616
rect 11789 9558 15535 9560
rect 11789 9555 11855 9558
rect 15469 9555 15535 9558
rect 16941 9482 17007 9485
rect 10918 9480 17007 9482
rect 10918 9424 16946 9480
rect 17002 9424 17007 9480
rect 10918 9422 17007 9424
rect 7874 9280 8194 9281
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 0 9074 800 9104
rect 4061 9074 4127 9077
rect 0 9072 4127 9074
rect 0 9016 4066 9072
rect 4122 9016 4127 9072
rect 0 9014 4127 9016
rect 0 8984 800 9014
rect 4061 9011 4127 9014
rect 10412 8941 10472 9422
rect 10685 9419 10751 9422
rect 16941 9419 17007 9422
rect 21265 9482 21331 9485
rect 22200 9482 23000 9512
rect 21265 9480 23000 9482
rect 21265 9424 21270 9480
rect 21326 9424 23000 9480
rect 21265 9422 23000 9424
rect 21265 9419 21331 9422
rect 22200 9392 23000 9422
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 9215 15125 9216
rect 19517 9074 19583 9077
rect 22200 9074 23000 9104
rect 19517 9072 23000 9074
rect 19517 9016 19522 9072
rect 19578 9016 23000 9072
rect 19517 9014 23000 9016
rect 19517 9011 19583 9014
rect 22200 8984 23000 9014
rect 10409 8936 10475 8941
rect 10409 8880 10414 8936
rect 10470 8880 10475 8936
rect 10409 8875 10475 8880
rect 9949 8802 10015 8805
rect 10869 8802 10935 8805
rect 9949 8800 10935 8802
rect 9949 8744 9954 8800
rect 10010 8744 10874 8800
rect 10930 8744 10935 8800
rect 9949 8742 10935 8744
rect 9949 8739 10015 8742
rect 10869 8739 10935 8742
rect 4409 8736 4729 8737
rect 0 8666 800 8696
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 8671 18590 8672
rect 1485 8666 1551 8669
rect 0 8664 1551 8666
rect 0 8608 1490 8664
rect 1546 8608 1551 8664
rect 0 8606 1551 8608
rect 0 8576 800 8606
rect 1485 8603 1551 8606
rect 21265 8666 21331 8669
rect 22200 8666 23000 8696
rect 21265 8664 23000 8666
rect 21265 8608 21270 8664
rect 21326 8608 23000 8664
rect 21265 8606 23000 8608
rect 21265 8603 21331 8606
rect 22200 8576 23000 8606
rect 7097 8530 7163 8533
rect 7598 8530 7604 8532
rect 7097 8528 7604 8530
rect 7097 8472 7102 8528
rect 7158 8472 7604 8528
rect 7097 8470 7604 8472
rect 7097 8467 7163 8470
rect 7598 8468 7604 8470
rect 7668 8530 7674 8532
rect 8017 8530 8083 8533
rect 7668 8528 8083 8530
rect 7668 8472 8022 8528
rect 8078 8472 8083 8528
rect 7668 8470 8083 8472
rect 7668 8468 7674 8470
rect 8017 8467 8083 8470
rect 10317 8530 10383 8533
rect 13077 8530 13143 8533
rect 10317 8528 13143 8530
rect 10317 8472 10322 8528
rect 10378 8472 13082 8528
rect 13138 8472 13143 8528
rect 10317 8470 13143 8472
rect 10317 8467 10383 8470
rect 13077 8467 13143 8470
rect 4613 8394 4679 8397
rect 8661 8394 8727 8397
rect 4613 8392 8727 8394
rect 4613 8336 4618 8392
rect 4674 8336 8666 8392
rect 8722 8336 8727 8392
rect 4613 8334 8727 8336
rect 4613 8331 4679 8334
rect 8661 8331 8727 8334
rect 3233 8260 3299 8261
rect 3182 8196 3188 8260
rect 3252 8258 3299 8260
rect 8569 8258 8635 8261
rect 9489 8258 9555 8261
rect 3252 8256 3344 8258
rect 3294 8200 3344 8256
rect 3252 8198 3344 8200
rect 8569 8256 9555 8258
rect 8569 8200 8574 8256
rect 8630 8200 9494 8256
rect 9550 8200 9555 8256
rect 8569 8198 9555 8200
rect 3252 8196 3299 8198
rect 3233 8195 3299 8196
rect 8569 8195 8635 8198
rect 9489 8195 9555 8198
rect 17769 8258 17835 8261
rect 17902 8258 17908 8260
rect 17769 8256 17908 8258
rect 17769 8200 17774 8256
rect 17830 8200 17908 8256
rect 17769 8198 17908 8200
rect 17769 8195 17835 8198
rect 17902 8196 17908 8198
rect 17972 8196 17978 8260
rect 7874 8192 8194 8193
rect 0 8122 800 8152
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 8127 15125 8128
rect 4061 8122 4127 8125
rect 0 8120 4127 8122
rect 0 8064 4066 8120
rect 4122 8064 4127 8120
rect 0 8062 4127 8064
rect 0 8032 800 8062
rect 4061 8059 4127 8062
rect 20713 8122 20779 8125
rect 22200 8122 23000 8152
rect 20713 8120 23000 8122
rect 20713 8064 20718 8120
rect 20774 8064 23000 8120
rect 20713 8062 23000 8064
rect 20713 8059 20779 8062
rect 22200 8032 23000 8062
rect 3417 7986 3483 7989
rect 5717 7986 5783 7989
rect 3417 7984 5783 7986
rect 3417 7928 3422 7984
rect 3478 7928 5722 7984
rect 5778 7928 5783 7984
rect 3417 7926 5783 7928
rect 3417 7923 3483 7926
rect 5717 7923 5783 7926
rect 3693 7850 3759 7853
rect 8385 7850 8451 7853
rect 3693 7848 8451 7850
rect 3693 7792 3698 7848
rect 3754 7792 8390 7848
rect 8446 7792 8451 7848
rect 3693 7790 8451 7792
rect 3693 7787 3759 7790
rect 8385 7787 8451 7790
rect 12341 7850 12407 7853
rect 18689 7850 18755 7853
rect 12341 7848 18755 7850
rect 12341 7792 12346 7848
rect 12402 7792 18694 7848
rect 18750 7792 18755 7848
rect 12341 7790 18755 7792
rect 12341 7787 12407 7790
rect 18689 7787 18755 7790
rect 0 7714 800 7744
rect 3417 7714 3483 7717
rect 0 7712 3483 7714
rect 0 7656 3422 7712
rect 3478 7656 3483 7712
rect 0 7654 3483 7656
rect 0 7624 800 7654
rect 3417 7651 3483 7654
rect 20713 7714 20779 7717
rect 22200 7714 23000 7744
rect 20713 7712 23000 7714
rect 20713 7656 20718 7712
rect 20774 7656 23000 7712
rect 20713 7654 23000 7656
rect 20713 7651 20779 7654
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 22200 7624 23000 7654
rect 18270 7583 18590 7584
rect 16113 7442 16179 7445
rect 18321 7442 18387 7445
rect 16113 7440 18387 7442
rect 16113 7384 16118 7440
rect 16174 7384 18326 7440
rect 18382 7384 18387 7440
rect 16113 7382 18387 7384
rect 16113 7379 16179 7382
rect 18321 7379 18387 7382
rect 1853 7306 1919 7309
rect 9121 7306 9187 7309
rect 1853 7304 9187 7306
rect 1853 7248 1858 7304
rect 1914 7248 9126 7304
rect 9182 7248 9187 7304
rect 1853 7246 9187 7248
rect 1853 7243 1919 7246
rect 9121 7243 9187 7246
rect 0 7170 800 7200
rect 3325 7170 3391 7173
rect 0 7168 3391 7170
rect 0 7112 3330 7168
rect 3386 7112 3391 7168
rect 0 7110 3391 7112
rect 0 7080 800 7110
rect 3325 7107 3391 7110
rect 19149 7170 19215 7173
rect 22200 7170 23000 7200
rect 19149 7168 23000 7170
rect 19149 7112 19154 7168
rect 19210 7112 23000 7168
rect 19149 7110 23000 7112
rect 19149 7107 19215 7110
rect 7874 7104 8194 7105
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 22200 7080 23000 7110
rect 14805 7039 15125 7040
rect 2773 7034 2839 7037
rect 6085 7034 6151 7037
rect 2773 7032 6151 7034
rect 2773 6976 2778 7032
rect 2834 6976 6090 7032
rect 6146 6976 6151 7032
rect 2773 6974 6151 6976
rect 2773 6971 2839 6974
rect 6085 6971 6151 6974
rect 0 6762 800 6792
rect 2313 6762 2379 6765
rect 0 6760 2379 6762
rect 0 6704 2318 6760
rect 2374 6704 2379 6760
rect 0 6702 2379 6704
rect 0 6672 800 6702
rect 2313 6699 2379 6702
rect 15101 6762 15167 6765
rect 17033 6762 17099 6765
rect 15101 6760 17099 6762
rect 15101 6704 15106 6760
rect 15162 6704 17038 6760
rect 17094 6704 17099 6760
rect 15101 6702 17099 6704
rect 15101 6699 15167 6702
rect 17033 6699 17099 6702
rect 22001 6762 22067 6765
rect 22200 6762 23000 6792
rect 22001 6760 23000 6762
rect 22001 6704 22006 6760
rect 22062 6704 23000 6760
rect 22001 6702 23000 6704
rect 22001 6699 22067 6702
rect 22200 6672 23000 6702
rect 4409 6560 4729 6561
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 6495 18590 6496
rect 1669 6354 1735 6357
rect 6453 6354 6519 6357
rect 1669 6352 6519 6354
rect 1669 6296 1674 6352
rect 1730 6296 6458 6352
rect 6514 6296 6519 6352
rect 1669 6294 6519 6296
rect 1669 6291 1735 6294
rect 6453 6291 6519 6294
rect 0 6218 800 6248
rect 1577 6218 1643 6221
rect 0 6216 1643 6218
rect 0 6160 1582 6216
rect 1638 6160 1643 6216
rect 0 6158 1643 6160
rect 0 6128 800 6158
rect 1577 6155 1643 6158
rect 6453 6218 6519 6221
rect 7189 6218 7255 6221
rect 10317 6218 10383 6221
rect 6453 6216 10383 6218
rect 6453 6160 6458 6216
rect 6514 6160 7194 6216
rect 7250 6160 10322 6216
rect 10378 6160 10383 6216
rect 6453 6158 10383 6160
rect 6453 6155 6519 6158
rect 7189 6155 7255 6158
rect 10317 6155 10383 6158
rect 18965 6218 19031 6221
rect 19149 6218 19215 6221
rect 18965 6216 19215 6218
rect 18965 6160 18970 6216
rect 19026 6160 19154 6216
rect 19210 6160 19215 6216
rect 18965 6158 19215 6160
rect 18965 6155 19031 6158
rect 19149 6155 19215 6158
rect 21265 6218 21331 6221
rect 22200 6218 23000 6248
rect 21265 6216 23000 6218
rect 21265 6160 21270 6216
rect 21326 6160 23000 6216
rect 21265 6158 23000 6160
rect 21265 6155 21331 6158
rect 22200 6128 23000 6158
rect 7874 6016 8194 6017
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 5951 15125 5952
rect 1761 5946 1827 5949
rect 6821 5946 6887 5949
rect 1761 5944 6887 5946
rect 1761 5888 1766 5944
rect 1822 5888 6826 5944
rect 6882 5888 6887 5944
rect 1761 5886 6887 5888
rect 1761 5883 1827 5886
rect 6821 5883 6887 5886
rect 0 5810 800 5840
rect 1669 5810 1735 5813
rect 0 5808 1735 5810
rect 0 5752 1674 5808
rect 1730 5752 1735 5808
rect 0 5750 1735 5752
rect 0 5720 800 5750
rect 1669 5747 1735 5750
rect 20621 5810 20687 5813
rect 22200 5810 23000 5840
rect 20621 5808 23000 5810
rect 20621 5752 20626 5808
rect 20682 5752 23000 5808
rect 20621 5750 23000 5752
rect 20621 5747 20687 5750
rect 22200 5720 23000 5750
rect 6637 5674 6703 5677
rect 9397 5674 9463 5677
rect 6637 5672 9463 5674
rect 6637 5616 6642 5672
rect 6698 5616 9402 5672
rect 9458 5616 9463 5672
rect 6637 5614 9463 5616
rect 6637 5611 6703 5614
rect 9397 5611 9463 5614
rect 5717 5538 5783 5541
rect 10225 5538 10291 5541
rect 5717 5536 10291 5538
rect 5717 5480 5722 5536
rect 5778 5480 10230 5536
rect 10286 5480 10291 5536
rect 5717 5478 10291 5480
rect 5717 5475 5783 5478
rect 10225 5475 10291 5478
rect 4409 5472 4729 5473
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 2221 5402 2287 5405
rect 3785 5402 3851 5405
rect 2221 5400 3851 5402
rect 2221 5344 2226 5400
rect 2282 5344 3790 5400
rect 3846 5344 3851 5400
rect 2221 5342 3851 5344
rect 2221 5339 2287 5342
rect 3785 5339 3851 5342
rect 5257 5402 5323 5405
rect 8937 5402 9003 5405
rect 5257 5400 9003 5402
rect 5257 5344 5262 5400
rect 5318 5344 8942 5400
rect 8998 5344 9003 5400
rect 5257 5342 9003 5344
rect 5257 5339 5323 5342
rect 8937 5339 9003 5342
rect 0 5266 800 5296
rect 3233 5266 3299 5269
rect 0 5264 3299 5266
rect 0 5208 3238 5264
rect 3294 5208 3299 5264
rect 0 5206 3299 5208
rect 0 5176 800 5206
rect 3233 5203 3299 5206
rect 13537 5266 13603 5269
rect 16941 5266 17007 5269
rect 13537 5264 17007 5266
rect 13537 5208 13542 5264
rect 13598 5208 16946 5264
rect 17002 5208 17007 5264
rect 13537 5206 17007 5208
rect 13537 5203 13603 5206
rect 16941 5203 17007 5206
rect 19149 5266 19215 5269
rect 22200 5266 23000 5296
rect 19149 5264 23000 5266
rect 19149 5208 19154 5264
rect 19210 5208 23000 5264
rect 19149 5206 23000 5208
rect 19149 5203 19215 5206
rect 22200 5176 23000 5206
rect 1577 5130 1643 5133
rect 14641 5130 14707 5133
rect 1577 5128 14707 5130
rect 1577 5072 1582 5128
rect 1638 5072 14646 5128
rect 14702 5072 14707 5128
rect 1577 5070 14707 5072
rect 1577 5067 1643 5070
rect 14641 5067 14707 5070
rect 7874 4928 8194 4929
rect 0 4858 800 4888
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 4863 15125 4864
rect 1761 4858 1827 4861
rect 0 4856 1827 4858
rect 0 4800 1766 4856
rect 1822 4800 1827 4856
rect 0 4798 1827 4800
rect 0 4768 800 4798
rect 1761 4795 1827 4798
rect 5257 4858 5323 4861
rect 5533 4858 5599 4861
rect 5257 4856 5599 4858
rect 5257 4800 5262 4856
rect 5318 4800 5538 4856
rect 5594 4800 5599 4856
rect 5257 4798 5599 4800
rect 5257 4795 5323 4798
rect 5533 4795 5599 4798
rect 21357 4858 21423 4861
rect 22200 4858 23000 4888
rect 21357 4856 23000 4858
rect 21357 4800 21362 4856
rect 21418 4800 23000 4856
rect 21357 4798 23000 4800
rect 21357 4795 21423 4798
rect 22200 4768 23000 4798
rect 2037 4722 2103 4725
rect 8293 4722 8359 4725
rect 2037 4720 8359 4722
rect 2037 4664 2042 4720
rect 2098 4664 8298 4720
rect 8354 4664 8359 4720
rect 2037 4662 8359 4664
rect 2037 4659 2103 4662
rect 8293 4659 8359 4662
rect 4245 4586 4311 4589
rect 7598 4586 7604 4588
rect 4245 4584 7604 4586
rect 4245 4528 4250 4584
rect 4306 4528 7604 4584
rect 4245 4526 7604 4528
rect 4245 4523 4311 4526
rect 7598 4524 7604 4526
rect 7668 4524 7674 4588
rect 10501 4586 10567 4589
rect 21081 4586 21147 4589
rect 10320 4584 21147 4586
rect 10320 4528 10506 4584
rect 10562 4528 21086 4584
rect 21142 4528 21147 4584
rect 10320 4526 21147 4528
rect 0 4450 800 4480
rect 1853 4450 1919 4453
rect 3601 4450 3667 4453
rect 0 4448 3667 4450
rect 0 4392 1858 4448
rect 1914 4392 3606 4448
rect 3662 4392 3667 4448
rect 0 4390 3667 4392
rect 0 4360 800 4390
rect 1853 4387 1919 4390
rect 3601 4387 3667 4390
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 4797 4314 4863 4317
rect 4797 4312 4906 4314
rect 4797 4256 4802 4312
rect 4858 4256 4906 4312
rect 4797 4251 4906 4256
rect 4429 4178 4495 4181
rect 4846 4178 4906 4251
rect 6545 4178 6611 4181
rect 4429 4176 6611 4178
rect 4429 4120 4434 4176
rect 4490 4120 6550 4176
rect 6606 4120 6611 4176
rect 4429 4118 6611 4120
rect 4429 4115 4495 4118
rect 6545 4115 6611 4118
rect 6729 4178 6795 4181
rect 9857 4178 9923 4181
rect 6729 4176 9923 4178
rect 6729 4120 6734 4176
rect 6790 4120 9862 4176
rect 9918 4120 9923 4176
rect 6729 4118 9923 4120
rect 6729 4115 6795 4118
rect 9857 4115 9923 4118
rect 10320 4045 10380 4526
rect 10501 4523 10567 4526
rect 21081 4523 21147 4526
rect 19241 4450 19307 4453
rect 22200 4450 23000 4480
rect 19241 4448 23000 4450
rect 19241 4392 19246 4448
rect 19302 4392 23000 4448
rect 19241 4390 23000 4392
rect 19241 4387 19307 4390
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 22200 4360 23000 4390
rect 18270 4319 18590 4320
rect 16389 4178 16455 4181
rect 18413 4178 18479 4181
rect 16389 4176 18479 4178
rect 16389 4120 16394 4176
rect 16450 4120 18418 4176
rect 18474 4120 18479 4176
rect 16389 4118 18479 4120
rect 16389 4115 16455 4118
rect 18413 4115 18479 4118
rect 10317 4040 10383 4045
rect 10317 3984 10322 4040
rect 10378 3984 10383 4040
rect 10317 3979 10383 3984
rect 0 3906 800 3936
rect 1393 3906 1459 3909
rect 0 3904 1459 3906
rect 0 3848 1398 3904
rect 1454 3848 1459 3904
rect 0 3846 1459 3848
rect 0 3816 800 3846
rect 1393 3843 1459 3846
rect 10726 3844 10732 3908
rect 10796 3906 10802 3908
rect 11145 3906 11211 3909
rect 10796 3904 11211 3906
rect 10796 3848 11150 3904
rect 11206 3848 11211 3904
rect 10796 3846 11211 3848
rect 10796 3844 10802 3846
rect 11145 3843 11211 3846
rect 17861 3906 17927 3909
rect 22200 3906 23000 3936
rect 17861 3904 23000 3906
rect 17861 3848 17866 3904
rect 17922 3848 23000 3904
rect 17861 3846 23000 3848
rect 17861 3843 17927 3846
rect 7874 3840 8194 3841
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 22200 3816 23000 3846
rect 14805 3775 15125 3776
rect 9765 3634 9831 3637
rect 2730 3632 9831 3634
rect 2730 3576 9770 3632
rect 9826 3576 9831 3632
rect 2730 3574 9831 3576
rect 0 3498 800 3528
rect 2730 3498 2790 3574
rect 9765 3571 9831 3574
rect 15929 3634 15995 3637
rect 17861 3634 17927 3637
rect 15929 3632 17927 3634
rect 15929 3576 15934 3632
rect 15990 3576 17866 3632
rect 17922 3576 17927 3632
rect 15929 3574 17927 3576
rect 15929 3571 15995 3574
rect 17861 3571 17927 3574
rect 0 3438 2790 3498
rect 2865 3498 2931 3501
rect 3182 3498 3188 3500
rect 2865 3496 3188 3498
rect 2865 3440 2870 3496
rect 2926 3440 3188 3496
rect 2865 3438 3188 3440
rect 0 3408 800 3438
rect 2865 3435 2931 3438
rect 3182 3436 3188 3438
rect 3252 3436 3258 3500
rect 3509 3498 3575 3501
rect 12893 3498 12959 3501
rect 3509 3496 12959 3498
rect 3509 3440 3514 3496
rect 3570 3440 12898 3496
rect 12954 3440 12959 3496
rect 3509 3438 12959 3440
rect 3509 3435 3575 3438
rect 12893 3435 12959 3438
rect 20529 3498 20595 3501
rect 22200 3498 23000 3528
rect 20529 3496 23000 3498
rect 20529 3440 20534 3496
rect 20590 3440 23000 3496
rect 20529 3438 23000 3440
rect 20529 3435 20595 3438
rect 22200 3408 23000 3438
rect 5441 3362 5507 3365
rect 5809 3362 5875 3365
rect 5441 3360 5875 3362
rect 5441 3304 5446 3360
rect 5502 3304 5814 3360
rect 5870 3304 5875 3360
rect 5441 3302 5875 3304
rect 5441 3299 5507 3302
rect 5809 3299 5875 3302
rect 4409 3296 4729 3297
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 3231 18590 3232
rect 2957 3090 3023 3093
rect 9213 3090 9279 3093
rect 2730 3088 9279 3090
rect 2730 3032 2962 3088
rect 3018 3032 9218 3088
rect 9274 3032 9279 3088
rect 2730 3030 9279 3032
rect 0 2954 800 2984
rect 2730 2954 2790 3030
rect 2957 3027 3023 3030
rect 9213 3027 9279 3030
rect 0 2894 2790 2954
rect 4245 2954 4311 2957
rect 5809 2954 5875 2957
rect 4245 2952 5875 2954
rect 4245 2896 4250 2952
rect 4306 2896 5814 2952
rect 5870 2896 5875 2952
rect 4245 2894 5875 2896
rect 0 2864 800 2894
rect 4245 2891 4311 2894
rect 5809 2891 5875 2894
rect 19425 2954 19491 2957
rect 22200 2954 23000 2984
rect 19425 2952 23000 2954
rect 19425 2896 19430 2952
rect 19486 2896 23000 2952
rect 19425 2894 23000 2896
rect 19425 2891 19491 2894
rect 22200 2864 23000 2894
rect 17902 2756 17908 2820
rect 17972 2818 17978 2820
rect 19241 2818 19307 2821
rect 17972 2816 19307 2818
rect 17972 2760 19246 2816
rect 19302 2760 19307 2816
rect 17972 2758 19307 2760
rect 17972 2756 17978 2758
rect 19241 2755 19307 2758
rect 7874 2752 8194 2753
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 0 2546 800 2576
rect 3969 2546 4035 2549
rect 0 2544 4035 2546
rect 0 2488 3974 2544
rect 4030 2488 4035 2544
rect 0 2486 4035 2488
rect 0 2456 800 2486
rect 3969 2483 4035 2486
rect 19149 2546 19215 2549
rect 22200 2546 23000 2576
rect 19149 2544 23000 2546
rect 19149 2488 19154 2544
rect 19210 2488 23000 2544
rect 19149 2486 23000 2488
rect 19149 2483 19215 2486
rect 22200 2456 23000 2486
rect 4409 2208 4729 2209
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2143 18590 2144
rect 0 2002 800 2032
rect 3693 2002 3759 2005
rect 0 2000 3759 2002
rect 0 1944 3698 2000
rect 3754 1944 3759 2000
rect 0 1942 3759 1944
rect 0 1912 800 1942
rect 3693 1939 3759 1942
rect 18045 2002 18111 2005
rect 22200 2002 23000 2032
rect 18045 2000 23000 2002
rect 18045 1944 18050 2000
rect 18106 1944 23000 2000
rect 18045 1942 23000 1944
rect 18045 1939 18111 1942
rect 22200 1912 23000 1942
rect 0 1594 800 1624
rect 3325 1594 3391 1597
rect 0 1592 3391 1594
rect 0 1536 3330 1592
rect 3386 1536 3391 1592
rect 0 1534 3391 1536
rect 0 1504 800 1534
rect 3325 1531 3391 1534
rect 17953 1594 18019 1597
rect 22200 1594 23000 1624
rect 17953 1592 23000 1594
rect 17953 1536 17958 1592
rect 18014 1536 23000 1592
rect 17953 1534 23000 1536
rect 17953 1531 18019 1534
rect 22200 1504 23000 1534
rect 0 1050 800 1080
rect 1853 1050 1919 1053
rect 0 1048 1919 1050
rect 0 992 1858 1048
rect 1914 992 1919 1048
rect 0 990 1919 992
rect 0 960 800 990
rect 1853 987 1919 990
rect 18781 1050 18847 1053
rect 22200 1050 23000 1080
rect 18781 1048 23000 1050
rect 18781 992 18786 1048
rect 18842 992 23000 1048
rect 18781 990 23000 992
rect 18781 987 18847 990
rect 22200 960 23000 990
rect 0 642 800 672
rect 4061 642 4127 645
rect 0 640 4127 642
rect 0 584 4066 640
rect 4122 584 4127 640
rect 0 582 4127 584
rect 0 552 800 582
rect 4061 579 4127 582
rect 20529 642 20595 645
rect 22200 642 23000 672
rect 20529 640 23000 642
rect 20529 584 20534 640
rect 20590 584 23000 640
rect 20529 582 23000 584
rect 20529 579 20595 582
rect 22200 552 23000 582
rect 0 234 800 264
rect 3417 234 3483 237
rect 0 232 3483 234
rect 0 176 3422 232
rect 3478 176 3483 232
rect 0 174 3483 176
rect 0 144 800 174
rect 3417 171 3483 174
rect 17677 234 17743 237
rect 22200 234 23000 264
rect 17677 232 23000 234
rect 17677 176 17682 232
rect 17738 176 23000 232
rect 17677 174 23000 176
rect 17677 171 17743 174
rect 22200 144 23000 174
<< via3 >>
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 10732 16628 10796 16692
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 7604 8468 7668 8532
rect 3188 8256 3252 8260
rect 3188 8200 3238 8256
rect 3238 8200 3252 8256
rect 3188 8196 3252 8200
rect 17908 8196 17972 8260
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 7604 4524 7668 4588
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 10732 3844 10796 3908
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 3188 3436 3252 3500
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 17908 2756 17972 2820
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
<< metal4 >>
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 17440 4729 18464
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 14176 4729 15200
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 13088 4729 14112
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 12000 4729 13024
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 10912 4729 11936
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 9824 4729 10848
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 8736 4729 9760
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 3187 8260 3253 8261
rect 3187 8196 3188 8260
rect 3252 8196 3253 8260
rect 3187 8195 3253 8196
rect 3190 3501 3250 8195
rect 4409 7648 4729 8672
rect 7874 20160 8195 20720
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 7874 19072 8195 20096
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 7874 17984 8195 19008
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7874 16896 8195 17920
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7874 15808 8195 16832
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 10731 16692 10797 16693
rect 10731 16628 10732 16692
rect 10796 16628 10797 16692
rect 10731 16627 10797 16628
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7874 14720 8195 15744
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7874 12544 8195 13568
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 7874 11456 8195 12480
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7874 10368 8195 11392
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 7874 9280 8195 10304
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 7603 8532 7669 8533
rect 7603 8468 7604 8532
rect 7668 8468 7669 8532
rect 7603 8467 7669 8468
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 6560 4729 7584
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 4384 4729 5408
rect 7606 4589 7666 8467
rect 7874 8192 8195 9216
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 7874 7104 8195 8128
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 7874 4928 8195 5952
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7603 4588 7669 4589
rect 7603 4524 7604 4588
rect 7668 4524 7669 4588
rect 7603 4523 7669 4524
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 3187 3500 3253 3501
rect 3187 3436 3188 3500
rect 3252 3436 3253 3500
rect 3187 3435 3253 3436
rect 4409 3296 4729 4320
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 2208 4729 3232
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 7874 3840 8195 4864
rect 10734 3909 10794 16627
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 10731 3908 10797 3909
rect 10731 3844 10732 3908
rect 10796 3844 10797 3908
rect 10731 3843 10797 3844
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 7874 2752 8195 3776
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 7874 2128 8195 2688
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 17984 15125 19008
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 16896 15125 17920
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 15808 15125 16832
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 14720 15125 15744
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 13632 15125 14656
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 12544 15125 13568
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 11456 15125 12480
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 10368 15125 11392
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 9280 15125 10304
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 8192 15125 9216
rect 18270 20704 18591 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18591 20704
rect 18270 19616 18591 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18591 19616
rect 18270 18528 18591 19552
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18591 18528
rect 18270 17440 18591 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18591 17440
rect 18270 16352 18591 17376
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18591 16352
rect 18270 15264 18591 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18591 15264
rect 18270 14176 18591 15200
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18591 14176
rect 18270 13088 18591 14112
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18591 13088
rect 18270 12000 18591 13024
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18591 12000
rect 18270 10912 18591 11936
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18591 10912
rect 18270 9824 18591 10848
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18591 9824
rect 18270 8736 18591 9760
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18591 8736
rect 17907 8260 17973 8261
rect 17907 8196 17908 8260
rect 17972 8196 17973 8260
rect 17907 8195 17973 8196
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 7104 15125 8128
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 6016 15125 7040
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 4928 15125 5952
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 3840 15125 4864
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 2752 15125 3776
rect 17910 2821 17970 8195
rect 18270 7648 18591 8672
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18591 7648
rect 18270 6560 18591 7584
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18591 6560
rect 18270 5472 18591 6496
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18591 5472
rect 18270 4384 18591 5408
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18591 4384
rect 18270 3296 18591 4320
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18591 3296
rect 17907 2820 17973 2821
rect 17907 2756 17908 2820
rect 17972 2756 17973 2820
rect 17907 2755 17973 2756
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2128 15125 2688
rect 18270 2208 18591 3232
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18591 2208
rect 18270 2128 18591 2144
use sky130_fd_sc_hd__fill_2  FILLER_1_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1624635492
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9
timestamp 1624635492
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3
timestamp 1624635492
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input73 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1564 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1624635492
transform 1 0 1564 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1624635492
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_15
timestamp 1624635492
transform 1 0 2484 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20
timestamp 1624635492
transform 1 0 2944 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15
timestamp 1624635492
transform 1 0 2484 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input77
timestamp 1624635492
transform 1 0 2116 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2668 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1624635492
transform 1 0 2116 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 4232 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 5888 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 5520 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1624635492
transform 1 0 3128 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1624635492
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3404 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30
timestamp 1624635492
transform 1 0 3864 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36
timestamp 1624635492
transform 1 0 4416 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_34
timestamp 1624635492
transform 1 0 4232 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48
timestamp 1624635492
transform 1 0 5520 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1624635492
transform 1 0 5704 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53
timestamp 1624635492
transform 1 0 5980 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1624635492
transform 1 0 5888 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 6256 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 6992 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1624635492
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1624635492
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1624635492
transform 1 0 6348 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59
timestamp 1624635492
transform 1 0 6532 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_58
timestamp 1624635492
transform 1 0 6440 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1624635492
transform 1 0 6624 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_69
timestamp 1624635492
transform 1 0 7452 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69
timestamp 1624635492
transform 1 0 7452 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64
timestamp 1624635492
transform 1 0 6992 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 7820 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input62
timestamp 1624635492
transform 1 0 7176 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input52
timestamp 1624635492
transform -1 0 7912 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_73
timestamp 1624635492
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74
timestamp 1624635492
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1624635492
transform -1 0 8924 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 9476 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_1_91
timestamp 1624635492
transform 1 0 9476 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_90
timestamp 1624635492
transform 1 0 9384 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1624635492
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1624635492
transform -1 0 9384 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 1624635492
transform 1 0 9660 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1624635492
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9568 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_96
timestamp 1624635492
transform 1 0 9936 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_101
timestamp 1624635492
transform 1 0 10396 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input54
timestamp 1624635492
transform -1 0 10856 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1624635492
transform 1 0 10120 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_107
timestamp 1624635492
transform 1 0 10948 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_106
timestamp 1624635492
transform 1 0 10856 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 11408 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_112
timestamp 1624635492
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output146
timestamp 1624635492
transform 1 0 11224 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_115
timestamp 1624635492
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114
timestamp 1624635492
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1624635492
transform -1 0 12052 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1624635492
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1624635492
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1624635492
transform -1 0 12144 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1624635492
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_119
timestamp 1624635492
transform 1 0 12052 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output144
timestamp 1624635492
transform 1 0 12236 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1624635492
transform -1 0 12604 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_125
timestamp 1624635492
transform 1 0 12604 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_125
timestamp 1624635492
transform 1 0 12604 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output131
timestamp 1624635492
transform -1 0 13156 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1624635492
transform -1 0 13156 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_131
timestamp 1624635492
transform 1 0 13156 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_131
timestamp 1624635492
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output142
timestamp 1624635492
transform -1 0 13708 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1624635492
transform 1 0 13340 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_136
timestamp 1624635492
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_137
timestamp 1624635492
transform 1 0 13708 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output143
timestamp 1624635492
transform -1 0 14260 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1624635492
transform -1 0 14076 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_141
timestamp 1624635492
transform 1 0 14076 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_143
timestamp 1624635492
transform 1 0 14260 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_145
timestamp 1624635492
transform 1 0 14444 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1624635492
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_154
timestamp 1624635492
transform 1 0 15272 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_150
timestamp 1624635492
transform 1 0 14904 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_154
timestamp 1624635492
transform 1 0 15272 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_148
timestamp 1624635492
transform 1 0 14720 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1624635492
transform -1 0 14720 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output145
timestamp 1624635492
transform -1 0 14904 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output141
timestamp 1624635492
transform 1 0 14904 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1624635492
transform 1 0 15364 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_164
timestamp 1624635492
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_160
timestamp 1624635492
transform 1 0 15824 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output139
timestamp 1624635492
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output135
timestamp 1624635492
transform 1 0 16008 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1624635492
transform 1 0 16376 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1624635492
transform -1 0 16652 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1624635492
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output134
timestamp 1624635492
transform 1 0 16560 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1624635492
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_172
timestamp 1624635492
transform 1 0 16928 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_175
timestamp 1624635492
transform 1 0 17204 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_172
timestamp 1624635492
transform 1 0 16928 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output147
timestamp 1624635492
transform -1 0 17480 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1624635492
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_178
timestamp 1624635492
transform 1 0 17480 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_181
timestamp 1624635492
transform 1 0 17756 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output148
timestamp 1624635492
transform -1 0 18032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output132
timestamp 1624635492
transform -1 0 17756 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_184
timestamp 1624635492
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output133
timestamp 1624635492
transform -1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1624635492
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_193
timestamp 1624635492
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_188
timestamp 1624635492
transform 1 0 18400 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_195
timestamp 1624635492
transform 1 0 19044 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output140
timestamp 1624635492
transform 1 0 18492 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output136
timestamp 1624635492
transform -1 0 19412 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output89
timestamp 1624635492
transform 1 0 18676 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1624635492
transform -1 0 19596 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_205
timestamp 1624635492
transform 1 0 19964 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_199
timestamp 1624635492
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_204
timestamp 1624635492
transform 1 0 19872 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_201
timestamp 1624635492
transform 1 0 19596 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output137
timestamp 1624635492
transform -1 0 19964 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1624635492
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _056_
timestamp 1624635492
transform 1 0 20056 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 21344 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624635492
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624635492
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 20516 0 -1 2720
box -38 -48 958 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1624635492
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1624635492
transform 1 0 21436 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_220
timestamp 1624635492
transform 1 0 21344 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 3128 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624635492
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1624635492
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 3588 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1624635492
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1624635492
transform 1 0 4048 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1624635492
transform 1 0 4508 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_22
timestamp 1624635492
transform 1 0 3128 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1624635492
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_30
timestamp 1624635492
transform 1 0 3864 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_35
timestamp 1624635492
transform 1 0 4324 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_40
timestamp 1624635492
transform 1 0 4784 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 7820 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1624635492
transform 1 0 5244 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_44
timestamp 1624635492
transform 1 0 5152 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_54
timestamp 1624635492
transform 1 0 6072 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1624635492
transform -1 0 8832 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_73
timestamp 1624635492
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1624635492
transform 1 0 10120 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1624635492
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input55
timestamp 1624635492
transform -1 0 9844 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1624635492
transform -1 0 9292 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_84
timestamp 1624635492
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_89
timestamp 1624635492
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_95
timestamp 1624635492
transform 1 0 9844 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 12420 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 11868 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 12880 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 11408 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_107
timestamp 1624635492
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_112
timestamp 1624635492
transform 1 0 11408 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_117
timestamp 1624635492
transform 1 0 11868 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_123
timestamp 1624635492
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1624635492
transform 1 0 13156 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1624635492
transform -1 0 13892 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1624635492
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1624635492
transform -1 0 14536 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_128
timestamp 1624635492
transform 1 0 12880 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_134
timestamp 1624635492
transform 1 0 13432 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_139
timestamp 1624635492
transform 1 0 13892 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 14812 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_2_146
timestamp 1624635492
transform 1 0 14536 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_165
timestamp 1624635492
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1624635492
transform 1 0 18032 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1624635492
transform 1 0 16468 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output149
timestamp 1624635492
transform -1 0 17848 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_176
timestamp 1624635492
transform 1 0 17296 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_182
timestamp 1624635492
transform 1 0 17848 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_187
timestamp 1624635492
transform 1 0 18308 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1624635492
transform 1 0 18492 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1624635492
transform 1 0 18952 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1624635492
transform 1 0 19504 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output138
timestamp 1624635492
transform -1 0 20332 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1624635492
transform -1 0 19780 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_192
timestamp 1624635492
transform 1 0 18768 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp 1624635492
transform 1 0 19228 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_203
timestamp 1624635492
transform 1 0 19780 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624635492
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input87
timestamp 1624635492
transform 1 0 20516 0 -1 3808
box -38 -48 958 592
use sky130_fd_sc_hd__fill_2  FILLER_2_209
timestamp 1624635492
transform 1 0 20332 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1624635492
transform 1 0 21436 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 2944 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624635492
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1624635492
transform 1 0 1380 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_20
timestamp 1624635492
transform 1 0 2944 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1624635492
transform 1 0 4876 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1624635492
transform 1 0 3128 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1624635492
transform 1 0 4140 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_31
timestamp 1624635492
transform 1 0 3956 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_36
timestamp 1624635492
transform 1 0 4416 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_40
timestamp 1624635492
transform 1 0 4784 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1624635492
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input63
timestamp 1624635492
transform -1 0 6164 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input64
timestamp 1624635492
transform 1 0 6624 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_50
timestamp 1624635492
transform 1 0 5704 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_55
timestamp 1624635492
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_58
timestamp 1624635492
transform 1 0 6440 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 8280 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1624635492
transform -1 0 8096 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_63
timestamp 1624635492
transform 1 0 6900 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_76
timestamp 1624635492
transform 1 0 8096 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input56
timestamp 1624635492
transform -1 0 10304 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 1624635492
transform -1 0 10764 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_94
timestamp 1624635492
transform 1 0 9752 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_100
timestamp 1624635492
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1624635492
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input58
timestamp 1624635492
transform -1 0 11224 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input59
timestamp 1624635492
transform 1 0 11868 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input60
timestamp 1624635492
transform -1 0 12604 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_105
timestamp 1624635492
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_110
timestamp 1624635492
transform 1 0 11224 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_115
timestamp 1624635492
transform 1 0 11684 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1624635492
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_125
timestamp 1624635492
transform 1 0 12604 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 13432 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1624635492
transform 1 0 12788 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_130
timestamp 1624635492
transform 1 0 13064 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _048_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 16468 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1624635492
transform -1 0 15916 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_150
timestamp 1624635492
transform 1 0 14904 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_161
timestamp 1624635492
transform 1 0 15916 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1624635492
transform 1 0 17664 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1624635492
transform 1 0 18124 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1624635492
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output150
timestamp 1624635492
transform -1 0 17480 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_167
timestamp 1624635492
transform 1 0 16468 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_172
timestamp 1624635492
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_178
timestamp 1624635492
transform 1 0 17480 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_183
timestamp 1624635492
transform 1 0 17940 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1624635492
transform 1 0 18676 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1624635492
transform 1 0 19136 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 21160 0 1 3808
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_3_188
timestamp 1624635492
transform 1 0 18400 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_194
timestamp 1624635492
transform 1 0 18952 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_199
timestamp 1624635492
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624635492
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_218
timestamp 1624635492
transform 1 0 21160 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_222
timestamp 1624635492
transform 1 0 21528 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1624635492
transform -1 0 3036 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624635492
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1624635492
transform 1 0 1564 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1624635492
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_9
timestamp 1624635492
transform 1 0 1932 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1624635492
transform -1 0 5612 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1624635492
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1624635492
transform -1 0 3496 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input71
timestamp 1624635492
transform 1 0 4048 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_21
timestamp 1624635492
transform 1 0 3036 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_26
timestamp 1624635492
transform 1 0 3496 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_30
timestamp 1624635492
transform 1 0 3864 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_35
timestamp 1624635492
transform 1 0 4324 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_39
timestamp 1624635492
transform 1 0 4692 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1624635492
transform 1 0 5796 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1624635492
transform 1 0 6808 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_49
timestamp 1624635492
transform 1 0 5612 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_60
timestamp 1624635492
transform 1 0 6624 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1624635492
transform -1 0 8740 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_4_71
timestamp 1624635492
transform 1 0 7636 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_83
timestamp 1624635492
transform 1 0 8740 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1624635492
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1624635492
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input78
timestamp 1624635492
transform -1 0 10028 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1624635492
transform -1 0 10396 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1624635492
transform -1 0 10764 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_87
timestamp 1624635492
transform 1 0 9108 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_92
timestamp 1624635492
transform 1 0 9568 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_97
timestamp 1624635492
transform 1 0 10028 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_101
timestamp 1624635492
transform 1 0 10396 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_1_
timestamp 1624635492
transform 1 0 10948 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1624635492
transform -1 0 12144 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1624635492
transform -1 0 12512 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_105
timestamp 1624635492
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_116
timestamp 1624635492
transform 1 0 11776 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_120
timestamp 1624635492
transform 1 0 12144 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_124
timestamp 1624635492
transform 1 0 12512 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 14076 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1624635492
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input83
timestamp 1624635492
transform 1 0 13340 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input84
timestamp 1624635492
transform 1 0 12880 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_131
timestamp 1624635492
transform 1 0 13156 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_136
timestamp 1624635492
transform 1 0 13616 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1624635492
transform 1 0 14076 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_144
timestamp 1624635492
transform 1 0 14352 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 15824 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 15640 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1624635492
transform -1 0 15180 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1624635492
transform -1 0 14720 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_148
timestamp 1624635492
transform 1 0 14720 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_153
timestamp 1624635492
transform 1 0 15180 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_158
timestamp 1624635492
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1624635492
transform 1 0 17480 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1624635492
transform -1 0 18768 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_176
timestamp 1624635492
transform 1 0 17296 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_181
timestamp 1624635492
transform 1 0 17756 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1624635492
transform -1 0 19320 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1624635492
transform 1 0 19780 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1624635492
transform 1 0 19504 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_192
timestamp 1624635492
transform 1 0 18768 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_198
timestamp 1624635492
transform 1 0 19320 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_201
timestamp 1624635492
transform 1 0 19596 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624635492
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1624635492
transform -1 0 21436 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_212
timestamp 1624635492
transform 1 0 20608 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_216
timestamp 1624635492
transform 1 0 20976 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1624635492
transform 1 0 21436 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1624635492
transform 1 0 2392 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1624635492
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1624635492
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1624635492
transform -1 0 2116 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_6
timestamp 1624635492
transform 1 0 1656 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_11
timestamp 1624635492
transform 1 0 2116 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1624635492
transform 1 0 3404 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input72
timestamp 1624635492
transform -1 0 4692 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_23
timestamp 1624635492
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_34
timestamp 1624635492
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_39
timestamp 1624635492
transform 1 0 4692 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1624635492
transform -1 0 6900 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1624635492
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input65
timestamp 1624635492
transform 1 0 5520 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input66
timestamp 1624635492
transform 1 0 5060 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1624635492
transform -1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_46
timestamp 1624635492
transform 1 0 5336 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_51
timestamp 1624635492
transform 1 0 5796 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_55
timestamp 1624635492
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_58
timestamp 1624635492
transform 1 0 6440 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1624635492
transform 1 0 8096 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 1624635492
transform 1 0 7084 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1624635492
transform -1 0 7820 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_63
timestamp 1624635492
transform 1 0 6900 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_68
timestamp 1624635492
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_73
timestamp 1624635492
transform 1 0 7820 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1624635492
transform 1 0 10580 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1624635492
transform -1 0 10396 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input70
timestamp 1624635492
transform -1 0 9384 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_85
timestamp 1624635492
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_90
timestamp 1624635492
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_101
timestamp 1624635492
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 11868 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1624635492
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_112
timestamp 1624635492
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_115
timestamp 1624635492
transform 1 0 11684 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1624635492
transform 1 0 13524 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_133
timestamp 1624635492
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_144
timestamp 1624635492
transform 1 0 14352 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 16652 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1624635492
transform -1 0 15456 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1624635492
transform -1 0 16192 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_156
timestamp 1624635492
transform 1 0 15456 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_160
timestamp 1624635492
transform 1 0 15824 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_164
timestamp 1624635492
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 17480 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1624635492
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1624635492
transform -1 0 17112 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1624635492
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_174
timestamp 1624635492
transform 1 0 17112 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 19136 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_194
timestamp 1624635492
transform 1 0 18952 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1624635492
transform 1 0 20792 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1624635492
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1624635492
transform -1 0 21436 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_212
timestamp 1624635492
transform 1 0 20608 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_217
timestamp 1624635492
transform 1 0 21068 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_221
timestamp 1624635492
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1624635492
transform 1 0 1380 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_9
timestamp 1624635492
transform 1 0 1932 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1624635492
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1624635492
transform 1 0 1564 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1624635492
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1624635492
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1624635492
transform -1 0 2300 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_13
timestamp 1624635492
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1624635492
transform 1 0 2484 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 2116 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_29
timestamp 1624635492
transform 1 0 3772 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_24
timestamp 1624635492
transform 1 0 3312 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_30
timestamp 1624635492
transform 1 0 3864 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1624635492
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input74
timestamp 1624635492
transform -1 0 4232 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1624635492
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1624635492
transform 1 0 3496 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_39
timestamp 1624635492
transform 1 0 4692 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_34
timestamp 1624635492
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input76
timestamp 1624635492
transform -1 0 5152 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input75
timestamp 1624635492
transform -1 0 4692 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4048 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_44
timestamp 1624635492
transform 1 0 5152 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_48
timestamp 1624635492
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1624635492
transform -1 0 5888 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1624635492
transform -1 0 6164 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_58
timestamp 1624635492
transform 1 0 6440 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_55
timestamp 1624635492
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_52
timestamp 1624635492
transform 1 0 5888 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1624635492
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1624635492
transform 1 0 6072 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1624635492
transform 1 0 6624 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 9752 0 1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1624635492
transform -1 0 8832 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input69
timestamp 1624635492
transform -1 0 7636 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1624635492
transform -1 0 7820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_63
timestamp 1624635492
transform 1 0 6900 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_67
timestamp 1624635492
transform 1 0 7268 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_71
timestamp 1624635492
transform 1 0 7636 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_69
timestamp 1624635492
transform 1 0 7452 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_73
timestamp 1624635492
transform 1 0 7820 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_87
timestamp 1624635492
transform 1 0 9108 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_84
timestamp 1624635492
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1624635492
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9292 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_7_102
timestamp 1624635492
transform 1 0 10488 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_98
timestamp 1624635492
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_94
timestamp 1624635492
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_98
timestamp 1624635492
transform 1 0 10120 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1624635492
transform -1 0 10120 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1624635492
transform -1 0 10488 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 11868 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_112
timestamp 1624635492
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_107
timestamp 1624635492
transform 1 0 10948 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1624635492
transform -1 0 11408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1624635492
transform -1 0 10948 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1624635492
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_122
timestamp 1624635492
transform 1 0 12328 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_117
timestamp 1624635492
transform 1 0 11868 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_122
timestamp 1624635492
transform 1 0 12328 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_117
timestamp 1624635492
transform 1 0 11868 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1624635492
transform -1 0 12788 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1624635492
transform -1 0 12328 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1624635492
transform -1 0 11868 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1624635492
transform 1 0 12052 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 12604 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1624635492
transform -1 0 13984 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_1_
timestamp 1624635492
transform 1 0 14168 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1624635492
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1624635492
transform 1 0 14076 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_144
timestamp 1624635492
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_127
timestamp 1624635492
transform 1 0 12788 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_140
timestamp 1624635492
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_155
timestamp 1624635492
transform 1 0 15364 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_151
timestamp 1624635492
transform 1 0 14996 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_153
timestamp 1624635492
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_149
timestamp 1624635492
transform 1 0 14812 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input82
timestamp 1624635492
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1624635492
transform 1 0 14536 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_158
timestamp 1624635492
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_157
timestamp 1624635492
transform 1 0 15548 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1624635492
transform -1 0 15640 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1624635492
transform -1 0 16652 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1624635492
transform -1 0 16560 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_172
timestamp 1624635492
transform 1 0 16928 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1624635492
transform 1 0 16652 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_173
timestamp 1624635492
transform 1 0 17020 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_168
timestamp 1624635492
transform 1 0 16560 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1624635492
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 17020 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 17480 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_1_
timestamp 1624635492
transform 1 0 17112 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_183
timestamp 1624635492
transform 1 0 17940 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_178
timestamp 1624635492
transform 1 0 17480 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1624635492
transform -1 0 18676 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 18400 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_193
timestamp 1624635492
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_188
timestamp 1624635492
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_191
timestamp 1624635492
transform 1 0 18676 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1624635492
transform 1 0 18584 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1624635492
transform 1 0 19044 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1624635492
transform -1 0 19320 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_203
timestamp 1624635492
transform 1 0 19780 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_198
timestamp 1624635492
transform 1 0 19320 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_201
timestamp 1624635492
transform 1 0 19596 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_198
timestamp 1624635492
transform 1 0 19320 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1624635492
transform 1 0 19504 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1624635492
transform 1 0 19780 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1624635492
transform 1 0 19504 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 21436 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1624635492
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1624635492
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1624635492
transform -1 0 21436 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_212
timestamp 1624635492
transform 1 0 20608 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_216
timestamp 1624635492
transform 1 0 20976 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_221
timestamp 1624635492
transform 1 0 21436 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1624635492
transform 1 0 21436 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1624635492
transform 1 0 1564 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1624635492
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1624635492
transform 1 0 2576 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1624635492
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_14
timestamp 1624635492
transform 1 0 2392 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_20
timestamp 1624635492
transform 1 0 2944 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 4416 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1624635492
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1624635492
transform 1 0 3128 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1624635492
transform -1 0 4048 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_25
timestamp 1624635492
transform 1 0 3404 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_32
timestamp 1624635492
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 6348 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_52
timestamp 1624635492
transform 1 0 5888 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_56
timestamp 1624635492
transform 1 0 6256 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1624635492
transform -1 0 8832 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_73
timestamp 1624635492
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 10212 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1624635492
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1624635492
transform -1 0 9292 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1624635492
transform -1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1624635492
transform -1 0 10028 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_84
timestamp 1624635492
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_89
timestamp 1624635492
transform 1 0 9292 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1624635492
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_97
timestamp 1624635492
transform 1 0 10028 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l3_in_0_
timestamp 1624635492
transform 1 0 11868 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_115
timestamp 1624635492
transform 1 0 11684 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1624635492
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1624635492
transform -1 0 13800 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1624635492
transform -1 0 13340 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_126
timestamp 1624635492
transform 1 0 12696 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_130
timestamp 1624635492
transform 1 0 13064 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_133
timestamp 1624635492
transform 1 0 13340 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_138
timestamp 1624635492
transform 1 0 13800 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_142
timestamp 1624635492
transform 1 0 14168 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_144
timestamp 1624635492
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 15272 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1624635492
transform -1 0 15088 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1624635492
transform -1 0 14720 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_148
timestamp 1624635492
transform 1 0 14720 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_152
timestamp 1624635492
transform 1 0 15088 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1624635492
transform -1 0 17296 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1624635492
transform -1 0 18308 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input80
timestamp 1624635492
transform -1 0 17848 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_170
timestamp 1624635492
transform 1 0 16744 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_176
timestamp 1624635492
transform 1 0 17296 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_182
timestamp 1624635492
transform 1 0 17848 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_187
timestamp 1624635492
transform 1 0 18308 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 19780 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1624635492
transform -1 0 19320 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1624635492
transform 1 0 19504 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_198
timestamp 1624635492
transform 1 0 19320 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_201
timestamp 1624635492
transform 1 0 19596 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1624635492
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_219
timestamp 1624635492
transform 1 0 21252 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1624635492
transform 1 0 2300 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1624635492
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1624635492
transform 1 0 1564 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1624635492
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_9
timestamp 1624635492
transform 1 0 1932 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_3_
timestamp 1624635492
transform -1 0 5060 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1624635492
transform 1 0 3312 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1624635492
transform -1 0 4048 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_22
timestamp 1624635492
transform 1 0 3128 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_28
timestamp 1624635492
transform 1 0 3680 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_32
timestamp 1624635492
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_2_
timestamp 1624635492
transform 1 0 5244 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1624635492
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1624635492
transform -1 0 6624 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1624635492
transform -1 0 6992 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_43
timestamp 1624635492
transform 1 0 5060 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_54
timestamp 1624635492
transform 1 0 6072 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_60
timestamp 1624635492
transform 1 0 6624 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 7728 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1624635492
transform -1 0 7360 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_64
timestamp 1624635492
transform 1 0 6992 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_68
timestamp 1624635492
transform 1 0 7360 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1624635492
transform -1 0 9568 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1624635492
transform -1 0 9936 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1624635492
transform -1 0 10304 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_88
timestamp 1624635492
transform 1 0 9200 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_92
timestamp 1624635492
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_96
timestamp 1624635492
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_100
timestamp 1624635492
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_104
timestamp 1624635492
transform 1 0 10672 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1624635492
transform 1 0 12328 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1624635492
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 10856 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 11224 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A1
timestamp 1624635492
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_108
timestamp 1624635492
transform 1 0 11040 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_112
timestamp 1624635492
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_117
timestamp 1624635492
transform 1 0 11868 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1624635492
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 14260 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 13892 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 13524 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_131
timestamp 1624635492
transform 1 0 13156 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_137
timestamp 1624635492
transform 1 0 13708 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_141
timestamp 1624635492
transform 1 0 14076 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_145
timestamp 1624635492
transform 1 0 14444 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1624635492
transform -1 0 14812 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_149
timestamp 1624635492
transform 1 0 14812 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 14996 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_153
timestamp 1624635492
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_157
timestamp 1624635492
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1624635492
transform -1 0 15548 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1624635492
transform -1 0 15916 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_161
timestamp 1624635492
transform 1 0 15916 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_165
timestamp 1624635492
transform 1 0 16284 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1624635492
transform -1 0 16284 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 17112 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1624635492
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1624635492
transform -1 0 16652 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1624635492
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_172
timestamp 1624635492
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1624635492
transform 1 0 19688 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 18860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1624635492
transform -1 0 19504 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_190
timestamp 1624635492
transform 1 0 18584 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_196
timestamp 1624635492
transform 1 0 19136 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_200
timestamp 1624635492
transform 1 0 19504 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1624635492
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1624635492
transform -1 0 21436 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1624635492
transform -1 0 20884 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_211
timestamp 1624635492
transform 1 0 20516 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_215
timestamp 1624635492
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_221
timestamp 1624635492
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1624635492
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1624635492
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1624635492
transform 1 0 1564 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1624635492
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_9
timestamp 1624635492
transform 1 0 1932 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_13
timestamp 1624635492
transform 1 0 2300 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1624635492
transform 1 0 4600 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1624635492
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1624635492
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1624635492
transform -1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_23
timestamp 1624635492
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1624635492
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_30
timestamp 1624635492
transform 1 0 3864 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_36
timestamp 1624635492
transform 1 0 4416 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_41
timestamp 1624635492
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1624635492
transform -1 0 5888 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1624635492
transform -1 0 6256 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1624635492
transform -1 0 6624 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1624635492
transform -1 0 6992 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_52
timestamp 1624635492
transform 1 0 5888 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_56
timestamp 1624635492
transform 1 0 6256 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_60
timestamp 1624635492
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 8740 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1624635492
transform -1 0 7360 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1624635492
transform -1 0 7728 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1624635492
transform -1 0 8096 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_64
timestamp 1624635492
transform 1 0 6992 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_68
timestamp 1624635492
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_72
timestamp 1624635492
transform 1 0 7728 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_76
timestamp 1624635492
transform 1 0 8096 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_83
timestamp 1624635492
transform 1 0 8740 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1624635492
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_89
timestamp 1624635492
transform 1 0 9292 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 9476 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1624635492
transform -1 0 9292 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1624635492
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_101
timestamp 1624635492
transform 1 0 10396 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_97
timestamp 1624635492
transform 1 0 10028 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 10212 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 9844 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 12144 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_120
timestamp 1624635492
transform 1 0 12144 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_125
timestamp 1624635492
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1624635492
transform 1 0 12788 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1624635492
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 13800 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_136
timestamp 1624635492
transform 1 0 13616 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1624635492
transform 1 0 14076 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_144
timestamp 1624635492
transform 1 0 14352 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 14536 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1624635492
transform -1 0 17020 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_162
timestamp 1624635492
transform 1 0 16008 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1624635492
transform 1 0 18308 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_1_
timestamp 1624635492
transform 1 0 17296 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_10_173
timestamp 1624635492
transform 1 0 17020 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_185
timestamp 1624635492
transform 1 0 18124 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1624635492
transform 1 0 19504 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1624635492
transform -1 0 20332 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1624635492
transform -1 0 19320 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1624635492
transform -1 0 19872 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_190
timestamp 1624635492
transform 1 0 18584 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_194
timestamp 1624635492
transform 1 0 18952 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_198
timestamp 1624635492
transform 1 0 19320 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_201
timestamp 1624635492
transform 1 0 19596 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_204
timestamp 1624635492
transform 1 0 19872 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1624635492
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1624635492
transform -1 0 21436 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1624635492
transform -1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_209
timestamp 1624635492
transform 1 0 20332 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_215
timestamp 1624635492
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_221
timestamp 1624635492
transform 1 0 21436 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1624635492
transform -1 0 1656 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 3312 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1624635492
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_6
timestamp 1624635492
transform 1 0 1656 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1624635492
transform 1 0 3864 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1624635492
transform 1 0 4876 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1624635492
transform -1 0 3680 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_24
timestamp 1624635492
transform 1 0 3312 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_28
timestamp 1624635492
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_39
timestamp 1624635492
transform 1 0 4692 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1624635492
transform 1 0 6624 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1624635492
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1624635492
transform -1 0 5520 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1624635492
transform -1 0 5888 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_44
timestamp 1624635492
transform 1 0 5152 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_48
timestamp 1624635492
transform 1 0 5520 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1624635492
transform 1 0 5888 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_56
timestamp 1624635492
transform 1 0 6256 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_58
timestamp 1624635492
transform 1 0 6440 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 8740 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1624635492
transform -1 0 8556 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_11_69
timestamp 1624635492
transform 1 0 7452 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_81
timestamp 1624635492
transform 1 0 8556 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_1_
timestamp 1624635492
transform -1 0 11408 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_99
timestamp 1624635492
transform 1 0 10212 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1624635492
transform 1 0 11868 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1624635492
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 12328 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_112
timestamp 1624635492
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_115
timestamp 1624635492
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1624635492
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_124
timestamp 1624635492
transform 1 0 12512 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 14168 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 14444 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_142
timestamp 1624635492
transform 1 0 14168 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 15180 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 14812 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_147
timestamp 1624635492
transform 1 0 14628 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_151
timestamp 1624635492
transform 1 0 14996 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1624635492
transform 1 0 17112 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1624635492
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input86
timestamp 1624635492
transform -1 0 18584 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1624635492
transform 1 0 16652 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_172
timestamp 1624635492
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_183
timestamp 1624635492
transform 1 0 17940 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 18768 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_190
timestamp 1624635492
transform 1 0 18584 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_208
timestamp 1624635492
transform 1 0 20240 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1624635492
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1624635492
transform -1 0 21436 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1624635492
transform -1 0 20884 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_215
timestamp 1624635492
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_221
timestamp 1624635492
transform 1 0 21436 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1624635492
transform 1 0 2760 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1624635492
transform -1 0 2576 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1624635492
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1624635492
transform -1 0 1564 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_5
timestamp 1624635492
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_16
timestamp 1624635492
transform 1 0 2576 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4048 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1624635492
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1624635492
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_30
timestamp 1624635492
transform 1 0 3864 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 5704 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_48
timestamp 1624635492
transform 1 0 5520 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1624635492
transform 1 0 7360 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 8648 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_66
timestamp 1624635492
transform 1 0 7176 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_77
timestamp 1624635492
transform 1 0 8188 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_81
timestamp 1624635492
transform 1 0 8556 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1624635492
transform -1 0 10120 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1624635492
transform 1 0 10304 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1624635492
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_84
timestamp 1624635492
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_87
timestamp 1624635492
transform 1 0 9108 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_98
timestamp 1624635492
transform 1 0 10120 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1624635492
transform -1 0 12144 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 12328 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_109
timestamp 1624635492
transform 1 0 11132 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_120
timestamp 1624635492
transform 1 0 12144 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_124
timestamp 1624635492
transform 1 0 12512 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1624635492
transform -1 0 14076 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1624635492
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 12696 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_128
timestamp 1624635492
transform 1 0 12880 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1624635492
transform 1 0 14076 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_144
timestamp 1624635492
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1624635492
transform -1 0 15364 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1624635492
transform -1 0 16376 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_155
timestamp 1624635492
transform 1 0 15364 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_166
timestamp 1624635492
transform 1 0 16376 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 16836 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_171
timestamp 1624635492
transform 1 0 16836 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1624635492
transform -1 0 17204 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_175
timestamp 1624635492
transform 1 0 17204 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1624635492
transform -1 0 17572 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_179
timestamp 1624635492
transform 1 0 17572 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1624635492
transform -1 0 17940 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_183
timestamp 1624635492
transform 1 0 17940 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1624635492
transform -1 0 18308 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_187
timestamp 1624635492
transform 1 0 18308 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 21252 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1624635492
transform 1 0 18492 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1624635492
transform 1 0 19504 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_198
timestamp 1624635492
transform 1 0 19320 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_201
timestamp 1624635492
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1624635492
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_219
timestamp 1624635492
transform 1 0 21252 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_9
timestamp 1624635492
transform 1 0 1932 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1624635492
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_8
timestamp 1624635492
transform 1 0 1840 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1624635492
transform 1 0 1380 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1624635492
transform 1 0 1564 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1624635492
transform 1 0 1472 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1624635492
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1624635492
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1624635492
transform -1 0 3128 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 2024 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1624635492
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_22
timestamp 1624635492
transform 1 0 3128 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_30
timestamp 1624635492
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_26
timestamp 1624635492
transform 1 0 3496 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1624635492
transform -1 0 4048 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1624635492
transform -1 0 3864 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1624635492
transform -1 0 3588 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1624635492
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_40
timestamp 1624635492
transform 1 0 4784 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_36
timestamp 1624635492
transform 1 0 4416 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_32
timestamp 1624635492
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_38
timestamp 1624635492
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_34
timestamp 1624635492
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1624635492
transform -1 0 4968 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1624635492
transform -1 0 4600 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1624635492
transform -1 0 4232 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1624635492
transform -1 0 4416 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1624635492
transform 1 0 4876 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_50
timestamp 1624635492
transform 1 0 5704 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_50
timestamp 1624635492
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_46
timestamp 1624635492
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_42
timestamp 1624635492
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1624635492
transform -1 0 5704 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1624635492
transform -1 0 5336 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_61
timestamp 1624635492
transform 1 0 6716 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_58
timestamp 1624635492
transform 1 0 6440 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_55
timestamp 1624635492
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 5888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1624635492
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1624635492
transform 1 0 5888 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1624635492
transform 1 0 6716 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_72
timestamp 1624635492
transform 1 0 7728 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_70
timestamp 1624635492
transform 1 0 7544 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1624635492
transform 1 0 6900 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1624635492
transform 1 0 7728 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_82
timestamp 1624635492
transform 1 0 8648 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_77
timestamp 1624635492
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_81
timestamp 1624635492
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 8372 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1624635492
transform -1 0 8188 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A1
timestamp 1624635492
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_89
timestamp 1624635492
transform 1 0 9292 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_89
timestamp 1624635492
transform 1 0 9292 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_85
timestamp 1624635492
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 9108 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1624635492
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_94
timestamp 1624635492
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1624635492
transform -1 0 10764 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 9660 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_113
timestamp 1624635492
transform 1 0 11500 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_109
timestamp 1624635492
transform 1 0 11132 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_113
timestamp 1624635492
transform 1 0 11500 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_109
timestamp 1624635492
transform 1 0 11132 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_105
timestamp 1624635492
transform 1 0 10764 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 11316 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 10948 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1624635492
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_117
timestamp 1624635492
transform 1 0 11868 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_115
timestamp 1624635492
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 11684 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 12236 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 11868 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 13524 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1624635492
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__A1
timestamp 1624635492
transform -1 0 14628 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 13892 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_133
timestamp 1624635492
transform 1 0 13340 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_137
timestamp 1624635492
transform 1 0 13708 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1624635492
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_144
timestamp 1624635492
transform 1 0 14352 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_147
timestamp 1624635492
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_151
timestamp 1624635492
transform 1 0 14996 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_3_
timestamp 1624635492
transform 1 0 14812 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1624635492
transform 1 0 15180 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_163
timestamp 1624635492
transform 1 0 16100 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_158
timestamp 1624635492
transform 1 0 15640 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_156
timestamp 1624635492
transform 1 0 15456 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 16100 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1624635492
transform 1 0 15732 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 16376 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 17112 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 17756 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_1_
timestamp 1624635492
transform -1 0 17572 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1624635492
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_168
timestamp 1624635492
transform 1 0 16560 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_172
timestamp 1624635492
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_168
timestamp 1624635492
transform 1 0 16560 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_179
timestamp 1624635492
transform 1 0 17572 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_197
timestamp 1624635492
transform 1 0 19228 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_196
timestamp 1624635492
transform 1 0 19136 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_190
timestamp 1624635492
transform 1 0 18584 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1624635492
transform -1 0 19136 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_203
timestamp 1624635492
transform 1 0 19780 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_201
timestamp 1624635492
transform 1 0 19596 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1624635492
transform -1 0 19780 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1624635492
transform 1 0 19320 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1624635492
transform 1 0 19504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1624635492
transform 1 0 20148 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1624635492
transform 1 0 19780 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1624635492
transform 1 0 21160 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1624635492
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1624635492
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1624635492
transform -1 0 21436 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_212
timestamp 1624635492
transform 1 0 20608 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_216
timestamp 1624635492
transform 1 0 20976 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1624635492
transform 1 0 21436 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_216
timestamp 1624635492
transform 1 0 20976 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_221
timestamp 1624635492
transform 1 0 21436 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _057_
timestamp 1624635492
transform 1 0 2116 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2576 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1624635492
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1624635492
transform 1 0 1564 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1624635492
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_9
timestamp 1624635492
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_14
timestamp 1624635492
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_19
timestamp 1624635492
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 3864 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3036 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1624635492
transform -1 0 3680 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_24
timestamp 1624635492
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_28
timestamp 1624635492
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1624635492
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1624635492
transform -1 0 5704 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 5888 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 6440 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_46
timestamp 1624635492
transform 1 0 5336 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_50
timestamp 1624635492
transform 1 0 5704 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_54
timestamp 1624635492
transform 1 0 6072 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_60
timestamp 1624635492
transform 1 0 6624 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 8464 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_80
timestamp 1624635492
transform 1 0 8464 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1624635492
transform 1 0 10488 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1624635492
transform -1 0 10304 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_84
timestamp 1624635492
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_88
timestamp 1624635492
transform 1 0 9200 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_100
timestamp 1624635492
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1624635492
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_105
timestamp 1624635492
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_109
timestamp 1624635492
transform 1 0 11132 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1624635492
transform 1 0 11500 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_115 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 11684 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_123
timestamp 1624635492
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 14444 0 1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 12696 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_128
timestamp 1624635492
transform 1 0 12880 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_138 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 13800 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_144
timestamp 1624635492
transform 1 0 14352 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_162
timestamp 1624635492
transform 1 0 16008 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_166
timestamp 1624635492
transform 1 0 16376 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1624635492
transform -1 0 18216 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1624635492
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 16468 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1624635492
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_172
timestamp 1624635492
transform 1 0 16928 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_175
timestamp 1624635492
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_186
timestamp 1624635492
transform 1 0 18216 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1624635492
transform 1 0 18400 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 19228 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1624635492
transform -1 0 19044 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_191
timestamp 1624635492
transform 1 0 18676 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_195
timestamp 1624635492
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1624635492
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1624635492
transform -1 0 21436 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_213
timestamp 1624635492
transform 1 0 20700 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_221
timestamp 1624635492
transform 1 0 21436 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_5_
timestamp 1624635492
transform -1 0 3220 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1624635492
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1624635492
transform 1 0 1564 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1624635492
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_9
timestamp 1624635492
transform 1 0 1932 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_13
timestamp 1624635492
transform 1 0 2300 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 5888 0 -1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1624635492
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1624635492
transform -1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 4048 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_23
timestamp 1624635492
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1624635492
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_32
timestamp 1624635492
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1624635492
transform -1 0 7452 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 6256 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_52
timestamp 1624635492
transform 1 0 5888 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_58
timestamp 1624635492
transform 1 0 6440 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1624635492
transform 1 0 7636 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_69
timestamp 1624635492
transform 1 0 7452 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_80
timestamp 1624635492
transform 1 0 8464 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1624635492
transform 1 0 9384 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1624635492
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 9844 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_87
timestamp 1624635492
transform 1 0 9108 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_93
timestamp 1624635492
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_98 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 10120 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 13524 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 11316 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_110
timestamp 1624635492
transform 1 0 11224 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_113
timestamp 1624635492
transform 1 0 11500 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1624635492
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 13984 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_135
timestamp 1624635492
transform 1 0 13524 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_140
timestamp 1624635492
transform 1 0 13984 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_144
timestamp 1624635492
transform 1 0 14352 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 15916 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__A1
timestamp 1624635492
transform 1 0 14904 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 15732 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_152
timestamp 1624635492
transform 1 0 15088 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_156
timestamp 1624635492
transform 1 0 15456 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_159
timestamp 1624635492
transform 1 0 15732 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_163
timestamp 1624635492
transform 1 0 16100 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1624635492
transform 1 0 17572 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 17388 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 16836 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 16468 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_169
timestamp 1624635492
transform 1 0 16652 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_173
timestamp 1624635492
transform 1 0 17020 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_177
timestamp 1624635492
transform 1 0 17388 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 19964 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1624635492
transform 1 0 19504 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1624635492
transform -1 0 19320 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1624635492
transform -1 0 19780 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1624635492
transform -1 0 18860 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_188
timestamp 1624635492
transform 1 0 18400 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_193
timestamp 1624635492
transform 1 0 18860 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_198
timestamp 1624635492
transform 1 0 19320 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_203
timestamp 1624635492
transform 1 0 19780 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1624635492
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1624635492
transform 1 0 21436 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 2300 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1624635492
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1624635492
transform 1 0 1564 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1624635492
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_9
timestamp 1624635492
transform 1 0 1932 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1624635492
transform 1 0 3956 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_29
timestamp 1624635492
transform 1 0 3772 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_40
timestamp 1624635492
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1624635492
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 5336 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_44
timestamp 1624635492
transform 1 0 5152 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_48
timestamp 1624635492
transform 1 0 5520 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_56
timestamp 1624635492
transform 1 0 6256 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_58
timestamp 1624635492
transform 1 0 6440 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1624635492
transform 1 0 7268 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_3_
timestamp 1624635492
transform -1 0 9292 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 7728 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_66
timestamp 1624635492
transform 1 0 7176 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_70
timestamp 1624635492
transform 1 0 7544 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_74
timestamp 1624635492
transform 1 0 7912 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1624635492
transform 1 0 9476 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1624635492
transform -1 0 11316 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_89
timestamp 1624635492
transform 1 0 9292 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_100
timestamp 1624635492
transform 1 0 10304 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1624635492
transform -1 0 12696 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1624635492
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_111
timestamp 1624635492
transform 1 0 11316 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_115
timestamp 1624635492
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1624635492
transform 1 0 12880 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1624635492
transform -1 0 14720 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_126
timestamp 1624635492
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_137
timestamp 1624635492
transform 1 0 13708 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_5_
timestamp 1624635492
transform -1 0 15916 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 16100 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_148
timestamp 1624635492
transform 1 0 14720 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_161
timestamp 1624635492
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_165
timestamp 1624635492
transform 1 0 16284 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1624635492
transform -1 0 18216 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1624635492
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 16468 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1624635492
transform 1 0 16652 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_172
timestamp 1624635492
transform 1 0 16928 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1624635492
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_186
timestamp 1624635492
transform 1 0 18216 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1624635492
transform 1 0 18400 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1624635492
transform 1 0 19412 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_197
timestamp 1624635492
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_208
timestamp 1624635492
transform 1 0 20240 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1624635492
transform 1 0 20516 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1624635492
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_220
timestamp 1624635492
transform 1 0 21344 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_4_
timestamp 1624635492
transform -1 0 3220 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1624635492
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1624635492
transform 1 0 1564 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1624635492
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_9
timestamp 1624635492
transform 1 0 1932 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_13
timestamp 1624635492
transform 1 0 2300 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1624635492
transform 1 0 4692 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1624635492
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1624635492
transform -1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 3864 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A
timestamp 1624635492
transform 1 0 4232 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1624635492
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1624635492
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_32
timestamp 1624635492
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_36
timestamp 1624635492
transform 1 0 4416 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__A1
timestamp 1624635492
transform 1 0 5704 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_48
timestamp 1624635492
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_52
timestamp 1624635492
transform 1 0 5888 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1624635492
transform 1 0 7176 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_64
timestamp 1624635492
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_75
timestamp 1624635492
transform 1 0 8004 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_83
timestamp 1624635492
transform 1 0 8740 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1624635492
transform 1 0 9384 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1624635492
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_87
timestamp 1624635492
transform 1 0 9108 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_99
timestamp 1624635492
transform 1 0 10212 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 11040 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_18_107
timestamp 1624635492
transform 1 0 10948 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_124
timestamp 1624635492
transform 1 0 12512 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1624635492
transform -1 0 12972 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1624635492
transform -1 0 13984 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1624635492
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_129
timestamp 1624635492
transform 1 0 12972 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_140
timestamp 1624635492
transform 1 0 13984 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_144
timestamp 1624635492
transform 1 0 14352 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 14536 0 -1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_18_163
timestamp 1624635492
transform 1 0 16100 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 17940 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1624635492
transform -1 0 18952 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_183
timestamp 1624635492
transform 1 0 17940 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1624635492
transform 1 0 19780 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1624635492
transform 1 0 19504 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1624635492
transform -1 0 19320 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1624635492
transform 1 0 18952 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_198
timestamp 1624635492
transform 1 0 19320 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_201
timestamp 1624635492
transform 1 0 19596 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1624635492
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1624635492
transform -1 0 21436 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_212
timestamp 1624635492
transform 1 0 20608 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_216
timestamp 1624635492
transform 1 0 20976 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 1624635492
transform 1 0 21436 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_9
timestamp 1624635492
transform 1 0 1932 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1624635492
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_6
timestamp 1624635492
transform 1 0 1656 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output91
timestamp 1624635492
transform -1 0 1932 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1624635492
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1624635492
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1624635492
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_13
timestamp 1624635492
transform 1 0 2300 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_19
timestamp 1624635492
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_14
timestamp 1624635492
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_10
timestamp 1624635492
transform 1 0 2024 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_6_
timestamp 1624635492
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp 1624635492
transform 1 0 2576 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _058_
timestamp 1624635492
transform 1 0 2116 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_30
timestamp 1624635492
transform 1 0 3864 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1624635492
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_23
timestamp 1624635492
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_23
timestamp 1624635492
transform 1 0 3220 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1624635492
transform -1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1624635492
transform -1 0 3220 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1624635492
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1624635492
transform -1 0 4416 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_39
timestamp 1624635492
transform 1 0 4692 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_35
timestamp 1624635492
transform 1 0 4324 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_36
timestamp 1624635492
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1624635492
transform 1 0 4600 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1624635492
transform 1 0 4784 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_49
timestamp 1624635492
transform 1 0 5612 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_51
timestamp 1624635492
transform 1 0 5796 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_47
timestamp 1624635492
transform 1 0 5428 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 5612 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1624635492
transform 1 0 5796 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_60
timestamp 1624635492
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_58
timestamp 1624635492
transform 1 0 6440 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_55
timestamp 1624635492
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1624635492
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1624635492
transform 1 0 6808 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_71
timestamp 1624635492
transform 1 0 7636 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_66
timestamp 1624635492
transform 1 0 7176 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1624635492
transform 1 0 7360 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_80
timestamp 1624635492
transform 1 0 8464 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_76
timestamp 1624635492
transform 1 0 8096 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_81
timestamp 1624635492
transform 1 0 8556 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_77
timestamp 1624635492
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1624635492
transform -1 0 8556 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 7912 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 8832 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_87
timestamp 1624635492
transform 1 0 9108 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1624635492
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_85
timestamp 1624635492
transform 1 0 8924 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1624635492
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1624635492
transform 1 0 9016 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_102
timestamp 1624635492
transform 1 0 10488 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_101
timestamp 1624635492
transform 1 0 10396 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_95
timestamp 1624635492
transform 1 0 9844 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 10488 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_104
timestamp 1624635492
transform 1 0 10672 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1624635492
transform -1 0 11776 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1624635492
transform -1 0 12880 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1624635492
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_112
timestamp 1624635492
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_115
timestamp 1624635492
transform 1 0 11684 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_106
timestamp 1624635492
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_116
timestamp 1624635492
transform 1 0 11776 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 12788 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1624635492
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_143
timestamp 1624635492
transform 1 0 14260 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_128
timestamp 1624635492
transform 1 0 12880 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_140
timestamp 1624635492
transform 1 0 13984 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_144
timestamp 1624635492
transform 1 0 14352 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_148
timestamp 1624635492
transform 1 0 14720 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_153
timestamp 1624635492
transform 1 0 15180 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_149
timestamp 1624635492
transform 1 0 14812 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__A1
timestamp 1624635492
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 14812 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1624635492
transform 1 0 14812 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_158
timestamp 1624635492
transform 1 0 15640 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_156
timestamp 1624635492
transform 1 0 15456 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1624635492
transform -1 0 16652 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_4_
timestamp 1624635492
transform -1 0 16468 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_176
timestamp 1624635492
transform 1 0 17296 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_173
timestamp 1624635492
transform 1 0 17020 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_169
timestamp 1624635492
transform 1 0 16652 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_176
timestamp 1624635492
transform 1 0 17296 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_172
timestamp 1624635492
transform 1 0 16928 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_167
timestamp 1624635492
transform 1 0 16468 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 17112 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1624635492
transform -1 0 17296 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1624635492
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_184
timestamp 1624635492
transform 1 0 18032 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_180
timestamp 1624635492
transform 1 0 17664 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_185
timestamp 1624635492
transform 1 0 18124 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_180
timestamp 1624635492
transform 1 0 17664 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 17480 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1624635492
transform -1 0 17664 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1624635492
transform -1 0 18032 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1624635492
transform -1 0 18400 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1624635492
transform -1 0 18124 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1624635492
transform 1 0 18308 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_193
timestamp 1624635492
transform 1 0 18860 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_188
timestamp 1624635492
transform 1 0 18400 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_196
timestamp 1624635492
transform 1 0 19136 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 19320 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_201
timestamp 1624635492
transform 1 0 19596 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_198
timestamp 1624635492
transform 1 0 19320 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_207
timestamp 1624635492
transform 1 0 20148 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1624635492
transform 1 0 19504 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1624635492
transform 1 0 19320 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1624635492
transform 1 0 19780 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_212
timestamp 1624635492
transform 1 0 20608 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1624635492
transform 1 0 20516 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_216
timestamp 1624635492
transform 1 0 20976 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_215
timestamp 1624635492
transform 1 0 20884 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1624635492
transform -1 0 21436 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1624635492
transform -1 0 21436 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1624635492
transform 1 0 21436 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_221
timestamp 1624635492
transform 1 0 21436 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1624635492
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1624635492
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1624635492
transform -1 0 3036 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1624635492
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output102
timestamp 1624635492
transform -1 0 1932 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1624635492
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_9
timestamp 1624635492
transform 1 0 1932 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1624635492
transform 1 0 3220 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp 1624635492
transform 1 0 3680 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1624635492
transform 1 0 4140 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_21
timestamp 1624635492
transform 1 0 3036 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_26
timestamp 1624635492
transform 1 0 3496 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_31
timestamp 1624635492
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1624635492
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1624635492
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_42
timestamp 1624635492
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_53
timestamp 1624635492
transform 1 0 5980 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_58
timestamp 1624635492
transform 1 0 6440 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1624635492
transform 1 0 7084 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1624635492
transform 1 0 8280 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_64
timestamp 1624635492
transform 1 0 6992 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_74
timestamp 1624635492
transform 1 0 7912 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9292 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 10672 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_87
timestamp 1624635492
transform 1 0 9108 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_98
timestamp 1624635492
transform 1 0 10120 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1624635492
transform -1 0 12696 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1624635492
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_106
timestamp 1624635492
transform 1 0 10856 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_112
timestamp 1624635492
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_115
timestamp 1624635492
transform 1 0 11684 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1624635492
transform -1 0 14444 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_126
timestamp 1624635492
transform 1 0 12696 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_134
timestamp 1624635492
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_145
timestamp 1624635492
transform 1 0 14444 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 16468 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A1
timestamp 1624635492
transform 1 0 14628 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1624635492
transform 1 0 14812 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_161
timestamp 1624635492
transform 1 0 15916 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1624635492
transform -1 0 18676 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1624635492
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A1
timestamp 1624635492
transform 1 0 17480 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_167
timestamp 1624635492
transform 1 0 16468 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_172
timestamp 1624635492
transform 1 0 16928 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_180
timestamp 1624635492
transform 1 0 17664 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1624635492
transform -1 0 20424 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1624635492
transform 1 0 18860 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_191
timestamp 1624635492
transform 1 0 18676 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_202
timestamp 1624635492
transform 1 0 19688 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_206
timestamp 1624635492
transform 1 0 20056 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1624635492
transform -1 0 20884 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1624635492
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output111
timestamp 1624635492
transform 1 0 21068 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_210
timestamp 1624635492
transform 1 0 20424 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_215
timestamp 1624635492
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_221
timestamp 1624635492
transform 1 0 21436 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1624635492
transform -1 0 3220 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1624635492
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output103
timestamp 1624635492
transform -1 0 1932 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1624635492
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_9
timestamp 1624635492
transform 1 0 1932 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_13
timestamp 1624635492
transform 1 0 2300 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1624635492
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1624635492
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__A1
timestamp 1624635492
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_23
timestamp 1624635492
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1624635492
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_30
timestamp 1624635492
transform 1 0 3864 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_41
timestamp 1624635492
transform 1 0 4876 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1624635492
transform 1 0 6716 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1624635492
transform 1 0 5704 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_22_49
timestamp 1624635492
transform 1 0 5612 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_59
timestamp 1624635492
transform 1 0 6532 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 7728 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 8188 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_70
timestamp 1624635492
transform 1 0 7544 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_75
timestamp 1624635492
transform 1 0 8004 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_79
timestamp 1624635492
transform 1 0 8372 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9292 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1624635492
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_85
timestamp 1624635492
transform 1 0 8924 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_87
timestamp 1624635492
transform 1 0 9108 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 11776 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_22_105
timestamp 1624635492
transform 1 0 10764 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_113
timestamp 1624635492
transform 1 0 11500 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1624635492
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 13616 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_132
timestamp 1624635492
transform 1 0 13248 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_139
timestamp 1624635492
transform 1 0 13892 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_144
timestamp 1624635492
transform 1 0 14352 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 15548 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1624635492
transform -1 0 15364 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_155
timestamp 1624635492
transform 1 0 15364 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 17204 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_173
timestamp 1624635492
transform 1 0 17020 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1624635492
transform -1 0 19320 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_6_
timestamp 1624635492
transform 1 0 19780 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1624635492
transform 1 0 19504 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_191
timestamp 1624635492
transform 1 0 18676 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_198
timestamp 1624635492
transform 1 0 19320 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_201
timestamp 1624635492
transform 1 0 19596 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1624635492
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output122
timestamp 1624635492
transform 1 0 21068 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_212
timestamp 1624635492
transform 1 0 20608 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_216
timestamp 1624635492
transform 1 0 20976 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1624635492
transform 1 0 21436 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 3864 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1624635492
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output104
timestamp 1624635492
transform -1 0 1932 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1624635492
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_9
timestamp 1624635492
transform 1 0 1932 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_13
timestamp 1624635492
transform 1 0 2300 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__A0
timestamp 1624635492
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_30
timestamp 1624635492
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_34
timestamp 1624635492
transform 1 0 4232 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 8096 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1624635492
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_46
timestamp 1624635492
transform 1 0 5336 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_54
timestamp 1624635492
transform 1 0 6072 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_58
timestamp 1624635492
transform 1 0 6440 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 8280 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_76
timestamp 1624635492
transform 1 0 8096 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 11408 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_94
timestamp 1624635492
transform 1 0 9752 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1624635492
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_112
timestamp 1624635492
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_115
timestamp 1624635492
transform 1 0 11684 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 13064 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_23_127
timestamp 1624635492
transform 1 0 12788 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1624635492
transform 1 0 15732 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1624635492
transform 1 0 14720 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_146
timestamp 1624635492
transform 1 0 14536 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_157
timestamp 1624635492
transform 1 0 15548 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_162
timestamp 1624635492
transform 1 0 16008 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1624635492
transform -1 0 18584 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1624635492
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_170
timestamp 1624635492
transform 1 0 16744 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_172
timestamp 1624635492
transform 1 0 16928 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_180
timestamp 1624635492
transform 1 0 17664 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1624635492
transform 1 0 18768 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1624635492
transform 1 0 19780 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_190
timestamp 1624635492
transform 1 0 18584 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_201
timestamp 1624635492
transform 1 0 19596 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1624635492
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output123
timestamp 1624635492
transform 1 0 21068 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_212
timestamp 1624635492
transform 1 0 20608 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_216
timestamp 1624635492
transform 1 0 20976 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_221
timestamp 1624635492
transform 1 0 21436 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1624635492
transform -1 0 3496 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1624635492
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output105
timestamp 1624635492
transform -1 0 1932 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output106
timestamp 1624635492
transform -1 0 2484 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1624635492
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_9
timestamp 1624635492
transform 1 0 1932 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_15
timestamp 1624635492
transform 1 0 2484 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 5520 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1624635492
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_26
timestamp 1624635492
transform 1 0 3496 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_30
timestamp 1624635492
transform 1 0 3864 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 8004 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_24_48
timestamp 1624635492
transform 1 0 5520 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_56
timestamp 1624635492
transform 1 0 6256 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_75
timestamp 1624635492
transform 1 0 8004 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_83
timestamp 1624635492
transform 1 0 8740 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1624635492
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 9568 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_87
timestamp 1624635492
transform 1 0 9108 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_92
timestamp 1624635492
transform 1 0 9568 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_104
timestamp 1624635492
transform 1 0 10672 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 12696 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1624635492
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_126
timestamp 1624635492
transform 1 0 12696 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_138
timestamp 1624635492
transform 1 0 13800 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_142
timestamp 1624635492
transform 1 0 14168 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_144
timestamp 1624635492
transform 1 0 14352 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 15548 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1624635492
transform -1 0 15364 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_155
timestamp 1624635492
transform 1 0 15364 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 17664 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_24_173
timestamp 1624635492
transform 1 0 17020 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_179
timestamp 1624635492
transform 1 0 17572 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1624635492
transform -1 0 20332 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1624635492
transform 1 0 19504 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A0
timestamp 1624635492
transform 1 0 19596 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_196
timestamp 1624635492
transform 1 0 19136 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_203
timestamp 1624635492
transform 1 0 19780 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1624635492
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output124
timestamp 1624635492
transform 1 0 21068 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output126
timestamp 1624635492
transform 1 0 20516 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_209
timestamp 1624635492
transform 1 0 20332 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1624635492
transform 1 0 20884 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1624635492
transform 1 0 21436 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp 1624635492
transform 1 0 2116 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _063_
timestamp 1624635492
transform 1 0 2576 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1624635492
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output107
timestamp 1624635492
transform -1 0 1932 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1624635492
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_9
timestamp 1624635492
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_14
timestamp 1624635492
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_19
timestamp 1624635492
transform 1 0 2852 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _064_
timestamp 1624635492
transform 1 0 3036 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4324 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3496 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1624635492
transform -1 0 4140 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_24
timestamp 1624635492
transform 1 0 3312 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_29
timestamp 1624635492
transform 1 0 3772 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_33
timestamp 1624635492
transform 1 0 4140 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1624635492
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A1
timestamp 1624635492
transform -1 0 6992 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A0
timestamp 1624635492
transform -1 0 6624 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_51
timestamp 1624635492
transform 1 0 5796 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_60
timestamp 1624635492
transform 1 0 6624 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 10028 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1624635492
transform -1 0 8004 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_64
timestamp 1624635492
transform 1 0 6992 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_75
timestamp 1624635492
transform 1 0 8004 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_97
timestamp 1624635492
transform 1 0 10028 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1624635492
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_109
timestamp 1624635492
transform 1 0 11132 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp 1624635492
transform 1 0 11500 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_117
timestamp 1624635492
transform 1 0 11868 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 13064 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_129
timestamp 1624635492
transform 1 0 12972 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_132
timestamp 1624635492
transform 1 0 13248 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_144
timestamp 1624635492
transform 1 0 14352 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_156
timestamp 1624635492
transform 1 0 15456 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1624635492
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_168
timestamp 1624635492
transform 1 0 16560 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_172
timestamp 1624635492
transform 1 0 16928 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_175
timestamp 1624635492
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_179
timestamp 1624635492
transform 1 0 17572 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_187
timestamp 1624635492
transform 1 0 18308 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1624635492
transform -1 0 20424 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1624635492
transform -1 0 19964 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 19504 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1624635492
transform -1 0 19044 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1624635492
transform -1 0 18676 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_191
timestamp 1624635492
transform 1 0 18676 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_195
timestamp 1624635492
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_200
timestamp 1624635492
transform 1 0 19504 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_205
timestamp 1624635492
transform 1 0 19964 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1624635492
transform -1 0 20884 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1624635492
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output125
timestamp 1624635492
transform 1 0 21068 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_210
timestamp 1624635492
transform 1 0 20424 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_215
timestamp 1624635492
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_221
timestamp 1624635492
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1624635492
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1624635492
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1624635492
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1624635492
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_9
timestamp 1624635492
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_9
timestamp 1624635492
transform 1 0 1932 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output109
timestamp 1624635492
transform -1 0 1932 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output108
timestamp 1624635492
transform -1 0 1932 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_14
timestamp 1624635492
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_14
timestamp 1624635492
transform 1 0 2392 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp 1624635492
transform 1 0 2116 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp 1624635492
transform 1 0 2116 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_19
timestamp 1624635492
transform 1 0 2852 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_19
timestamp 1624635492
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1624635492
transform 1 0 2576 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1624635492
transform 1 0 2576 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_30
timestamp 1624635492
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_28
timestamp 1624635492
transform 1 0 3680 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1624635492
transform 1 0 3312 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1624635492
transform -1 0 4048 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1624635492
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3036 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1624635492
transform -1 0 3864 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_27_39
timestamp 1624635492
transform 1 0 4692 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_35
timestamp 1624635492
transform 1 0 4324 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_40
timestamp 1624635492
transform 1 0 4784 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_36
timestamp 1624635492
transform 1 0 4416 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_32
timestamp 1624635492
transform 1 0 4048 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1624635492
transform -1 0 4692 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1624635492
transform 1 0 4600 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A
timestamp 1624635492
transform 1 0 4232 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1624635492
transform 1 0 4048 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_51
timestamp 1624635492
transform 1 0 5796 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_46
timestamp 1624635492
transform 1 0 5336 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1624635492
transform 1 0 4968 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1624635492
transform 1 0 5428 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_58
timestamp 1624635492
transform 1 0 6440 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_60
timestamp 1624635492
transform 1 0 6624 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_56
timestamp 1624635492
transform 1 0 6256 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 6440 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1624635492
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_62
timestamp 1624635492
transform 1 0 6808 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1624635492
transform 1 0 6900 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1624635492
transform -1 0 8648 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_26_64
timestamp 1624635492
transform 1 0 6992 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_72
timestamp 1624635492
transform 1 0 7728 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_82
timestamp 1624635492
transform 1 0 8648 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_72
timestamp 1624635492
transform 1 0 7728 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_84
timestamp 1624635492
transform 1 0 8832 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1624635492
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1624635492
transform 1 0 9108 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_27_100
timestamp 1624635492
transform 1 0 10304 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_96
timestamp 1624635492
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_99
timestamp 1624635492
transform 1 0 10212 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 10580 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1624635492
transform -1 0 11408 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_26_87
timestamp 1624635492
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1624635492
transform -1 0 11776 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1624635492
transform -1 0 12696 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1624635492
transform 1 0 11960 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1624635492
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_105
timestamp 1624635492
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_116
timestamp 1624635492
transform 1 0 11776 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_112
timestamp 1624635492
transform 1 0 11408 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_115
timestamp 1624635492
transform 1 0 11684 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_131
timestamp 1624635492
transform 1 0 13156 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_126
timestamp 1624635492
transform 1 0 12696 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_131
timestamp 1624635492
transform 1 0 13156 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_127
timestamp 1624635492
transform 1 0 12788 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1624635492
transform -1 0 14076 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1624635492
transform 1 0 13432 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1624635492
transform 1 0 12880 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_143
timestamp 1624635492
transform 1 0 14260 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_144
timestamp 1624635492
transform 1 0 14352 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1624635492
transform 1 0 14076 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1624635492
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1624635492
transform -1 0 14628 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1624635492
transform 1 0 16192 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1624635492
transform 1 0 15364 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1624635492
transform -1 0 15364 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 14812 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_155
timestamp 1624635492
transform 1 0 15364 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_163
timestamp 1624635492
transform 1 0 16100 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_147
timestamp 1624635492
transform 1 0 14628 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_151
timestamp 1624635492
transform 1 0 14996 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_164
timestamp 1624635492
transform 1 0 16192 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_172
timestamp 1624635492
transform 1 0 16928 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1624635492
transform 1 0 16652 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_173
timestamp 1624635492
transform 1 0 17020 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 16652 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1624635492
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1624635492
transform -1 0 17940 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1624635492
transform 1 0 17204 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_183
timestamp 1624635492
transform 1 0 17940 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_184
timestamp 1624635492
transform 1 0 18032 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 19596 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_26_192
timestamp 1624635492
transform 1 0 18768 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 19320 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_198
timestamp 1624635492
transform 1 0 19320 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_201
timestamp 1624635492
transform 1 0 19596 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_201
timestamp 1624635492
transform 1 0 19596 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1624635492
transform 1 0 19504 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_205
timestamp 1624635492
transform 1 0 19964 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_205
timestamp 1624635492
transform 1 0 19964 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1624635492
transform -1 0 19964 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1624635492
transform 1 0 19780 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1624635492
transform -1 0 20424 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1624635492
transform -1 0 20424 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_210
timestamp 1624635492
transform 1 0 20424 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_210
timestamp 1624635492
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1624635492
transform -1 0 20884 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1624635492
transform -1 0 20884 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_215
timestamp 1624635492
transform 1 0 20884 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_215
timestamp 1624635492
transform 1 0 20884 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output128
timestamp 1624635492
transform 1 0 21068 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output127
timestamp 1624635492
transform 1 0 21068 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_221
timestamp 1624635492
transform 1 0 21436 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_221
timestamp 1624635492
transform 1 0 21436 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1624635492
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1624635492
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1624635492
transform 1 0 2116 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1624635492
transform -1 0 3588 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1624635492
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output110
timestamp 1624635492
transform -1 0 1932 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1624635492
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_9
timestamp 1624635492
transform 1 0 1932 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_14
timestamp 1624635492
transform 1 0 2392 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1624635492
transform 1 0 4324 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1624635492
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1624635492
transform 1 0 3864 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1624635492
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_32
timestamp 1624635492
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 5612 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_28_44
timestamp 1624635492
transform 1 0 5152 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_48
timestamp 1624635492
transform 1 0 5520 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 7820 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 8280 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_65
timestamp 1624635492
transform 1 0 7084 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_76
timestamp 1624635492
transform 1 0 8096 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_80
timestamp 1624635492
transform 1 0 8464 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 9292 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1624635492
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_87
timestamp 1624635492
transform 1 0 9108 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 10948 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_105
timestamp 1624635492
transform 1 0 10764 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_123
timestamp 1624635492
transform 1 0 12420 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1624635492
transform -1 0 13984 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1624635492
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_129
timestamp 1624635492
transform 1 0 12972 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_140
timestamp 1624635492
transform 1 0 13984 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_144
timestamp 1624635492
transform 1 0 14352 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1624635492
transform 1 0 14812 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1624635492
transform -1 0 16652 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_147
timestamp 1624635492
transform 1 0 14628 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_158
timestamp 1624635492
transform 1 0 15640 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 18860 0 -1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_28_169
timestamp 1624635492
transform 1 0 16652 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_175
timestamp 1624635492
transform 1 0 17204 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1624635492
transform -1 0 20332 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 19320 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1624635492
transform 1 0 19504 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1624635492
transform -1 0 19872 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_193
timestamp 1624635492
transform 1 0 18860 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_198
timestamp 1624635492
transform 1 0 19320 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_201
timestamp 1624635492
transform 1 0 19596 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_204
timestamp 1624635492
transform 1 0 19872 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1624635492
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output129
timestamp 1624635492
transform 1 0 21068 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output130
timestamp 1624635492
transform 1 0 20516 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_209
timestamp 1624635492
transform 1 0 20332 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_215
timestamp 1624635492
transform 1 0 20884 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1624635492
transform 1 0 21436 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1624635492
transform 1 0 2668 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1624635492
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output92
timestamp 1624635492
transform -1 0 1932 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output93
timestamp 1624635492
transform -1 0 2484 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1624635492
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_9
timestamp 1624635492
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_15
timestamp 1624635492
transform 1 0 2484 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_20
timestamp 1624635492
transform 1 0 2944 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1624635492
transform -1 0 3956 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1624635492
transform 1 0 4140 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_31
timestamp 1624635492
transform 1 0 3956 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1624635492
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A1
timestamp 1624635492
transform -1 0 5336 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_42
timestamp 1624635492
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_46
timestamp 1624635492
transform 1 0 5336 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_54
timestamp 1624635492
transform 1 0 6072 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_58
timestamp 1624635492
transform 1 0 6440 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1624635492
transform 1 0 8464 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1624635492
transform 1 0 7452 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_29_66
timestamp 1624635492
transform 1 0 7176 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_78
timestamp 1624635492
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 9660 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_89
timestamp 1624635492
transform 1 0 9292 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1624635492
transform 1 0 9660 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1624635492
transform -1 0 12696 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1624635492
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_105
timestamp 1624635492
transform 1 0 10764 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_113
timestamp 1624635492
transform 1 0 11500 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_115
timestamp 1624635492
transform 1 0 11684 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1624635492
transform -1 0 15180 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_29_126
timestamp 1624635492
transform 1 0 12696 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_138
timestamp 1624635492
transform 1 0 13800 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1624635492
transform 1 0 15364 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_153
timestamp 1624635492
transform 1 0 15180 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_158
timestamp 1624635492
transform 1 0 15640 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1624635492
transform 1 0 17112 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1624635492
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1624635492
transform -1 0 18308 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_170
timestamp 1624635492
transform 1 0 16744 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_172
timestamp 1624635492
transform 1 0 16928 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_183
timestamp 1624635492
transform 1 0 17940 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_187
timestamp 1624635492
transform 1 0 18308 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1624635492
transform -1 0 20424 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 19964 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1624635492
transform -1 0 19504 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1624635492
transform -1 0 19136 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_193
timestamp 1624635492
transform 1 0 18860 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_196
timestamp 1624635492
transform 1 0 19136 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_200
timestamp 1624635492
transform 1 0 19504 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_205
timestamp 1624635492
transform 1 0 19964 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1624635492
transform -1 0 20884 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1624635492
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output112
timestamp 1624635492
transform 1 0 21068 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_210
timestamp 1624635492
transform 1 0 20424 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_215
timestamp 1624635492
transform 1 0 20884 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1624635492
transform 1 0 21436 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1624635492
transform 1 0 2116 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1624635492
transform 1 0 2576 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1624635492
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output94
timestamp 1624635492
transform -1 0 1932 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1624635492
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_9
timestamp 1624635492
transform 1 0 1932 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_14
timestamp 1624635492
transform 1 0 2392 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_19
timestamp 1624635492
transform 1 0 2852 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1624635492
transform 1 0 3312 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3036 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_28
timestamp 1624635492
transform 1 0 3680 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1624635492
transform 1 0 3864 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1624635492
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_32
timestamp 1624635492
transform 1 0 4048 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1624635492
transform 1 0 4232 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_40
timestamp 1624635492
transform 1 0 4784 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_36
timestamp 1624635492
transform 1 0 4416 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1624635492
transform 1 0 4600 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4968 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_30_58
timestamp 1624635492
transform 1 0 6440 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 7268 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_30_66
timestamp 1624635492
transform 1 0 7176 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_83
timestamp 1624635492
transform 1 0 8740 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1624635492
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_87
timestamp 1624635492
transform 1 0 9108 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_99
timestamp 1624635492
transform 1 0 10212 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 11960 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_30_111
timestamp 1624635492
transform 1 0 11316 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_117
timestamp 1624635492
transform 1 0 11868 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1624635492
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_134
timestamp 1624635492
transform 1 0 13432 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_142
timestamp 1624635492
transform 1 0 14168 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_144
timestamp 1624635492
transform 1 0 14352 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 14628 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_30_163
timestamp 1624635492
transform 1 0 16100 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_175
timestamp 1624635492
transform 1 0 17204 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_187
timestamp 1624635492
transform 1 0 18308 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1624635492
transform -1 0 20424 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 19320 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1624635492
transform 1 0 19504 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1624635492
transform 1 0 19780 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1624635492
transform 1 0 18676 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_193
timestamp 1624635492
transform 1 0 18860 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_198
timestamp 1624635492
transform 1 0 19320 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_201
timestamp 1624635492
transform 1 0 19596 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_205
timestamp 1624635492
transform 1 0 19964 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1624635492
transform -1 0 20884 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1624635492
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output113
timestamp 1624635492
transform 1 0 21068 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_210
timestamp 1624635492
transform 1 0 20424 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_215
timestamp 1624635492
transform 1 0 20884 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1624635492
transform 1 0 21436 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1624635492
transform 1 0 2116 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1624635492
transform 1 0 2576 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1624635492
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output95
timestamp 1624635492
transform -1 0 1932 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1624635492
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_9
timestamp 1624635492
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_14
timestamp 1624635492
transform 1 0 2392 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_19
timestamp 1624635492
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 4508 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1624635492
transform -1 0 4876 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_37
timestamp 1624635492
transform 1 0 4508 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_41
timestamp 1624635492
transform 1 0 4876 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1624635492
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1624635492
transform 1 0 5060 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_45
timestamp 1624635492
transform 1 0 5244 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_58
timestamp 1624635492
transform 1 0 6440 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 8280 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1624635492
transform 1 0 7268 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_31_66
timestamp 1624635492
transform 1 0 7176 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_76
timestamp 1624635492
transform 1 0 8096 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_94
timestamp 1624635492
transform 1 0 9752 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1624635492
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_106
timestamp 1624635492
transform 1 0 10856 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_115
timestamp 1624635492
transform 1 0 11684 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 13248 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_31_127
timestamp 1624635492
transform 1 0 12788 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_131
timestamp 1624635492
transform 1 0 13156 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_148
timestamp 1624635492
transform 1 0 14720 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_160
timestamp 1624635492
transform 1 0 15824 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1624635492
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1624635492
transform -1 0 18308 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_168
timestamp 1624635492
transform 1 0 16560 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_172
timestamp 1624635492
transform 1 0 16928 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_184
timestamp 1624635492
transform 1 0 18032 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_187
timestamp 1624635492
transform 1 0 18308 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1624635492
transform 1 0 20148 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1624635492
transform 1 0 19688 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1624635492
transform -1 0 19504 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1624635492
transform -1 0 19044 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1624635492
transform -1 0 18676 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_191
timestamp 1624635492
transform 1 0 18676 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_195
timestamp 1624635492
transform 1 0 19044 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_200
timestamp 1624635492
transform 1 0 19504 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_205
timestamp 1624635492
transform 1 0 19964 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1624635492
transform 1 0 20608 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1624635492
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output114
timestamp 1624635492
transform 1 0 21068 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_210
timestamp 1624635492
transform 1 0 20424 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_215
timestamp 1624635492
transform 1 0 20884 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_221
timestamp 1624635492
transform 1 0 21436 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1624635492
transform 1 0 2300 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1624635492
transform -1 0 3036 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1624635492
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output96
timestamp 1624635492
transform -1 0 1932 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1624635492
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_9
timestamp 1624635492
transform 1 0 1932 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_16
timestamp 1624635492
transform 1 0 2576 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1624635492
transform -1 0 3496 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 4048 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1624635492
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_21
timestamp 1624635492
transform 1 0 3036 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_26
timestamp 1624635492
transform 1 0 3496 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_30
timestamp 1624635492
transform 1 0 3864 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1624635492
transform 1 0 5704 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_48
timestamp 1624635492
transform 1 0 5520 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_52
timestamp 1624635492
transform 1 0 5888 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1624635492
transform 1 0 7728 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_32_64
timestamp 1624635492
transform 1 0 6992 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_81
timestamp 1624635492
transform 1 0 8556 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 10304 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1624635492
transform 1 0 9016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_85
timestamp 1624635492
transform 1 0 8924 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_87
timestamp 1624635492
transform 1 0 9108 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_99
timestamp 1624635492
transform 1 0 10212 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_116
timestamp 1624635492
transform 1 0 11776 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1624635492
transform 1 0 14260 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_128
timestamp 1624635492
transform 1 0 12880 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_140
timestamp 1624635492
transform 1 0 13984 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_144
timestamp 1624635492
transform 1 0 14352 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_156
timestamp 1624635492
transform 1 0 15456 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_168
timestamp 1624635492
transform 1 0 16560 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_180
timestamp 1624635492
transform 1 0 17664 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1624635492
transform 1 0 20056 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1624635492
transform 1 0 19504 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1624635492
transform -1 0 19872 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1624635492
transform 1 0 19136 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1624635492
transform 1 0 18768 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_198
timestamp 1624635492
transform 1 0 19320 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_201
timestamp 1624635492
transform 1 0 19596 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_204
timestamp 1624635492
transform 1 0 19872 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1624635492
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output115
timestamp 1624635492
transform 1 0 21068 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output121
timestamp 1624635492
transform 1 0 20516 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp 1624635492
transform 1 0 20332 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1624635492
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1624635492
transform 1 0 21436 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1624635492
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output97
timestamp 1624635492
transform -1 0 1932 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output98
timestamp 1624635492
transform -1 0 2484 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output99
timestamp 1624635492
transform -1 0 3036 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1624635492
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_9
timestamp 1624635492
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_15
timestamp 1624635492
transform 1 0 2484 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1624635492
transform 1 0 3772 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input79
timestamp 1624635492
transform -1 0 4876 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output100
timestamp 1624635492
transform -1 0 3588 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output101
timestamp 1624635492
transform -1 0 4416 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_21
timestamp 1624635492
transform 1 0 3036 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_27
timestamp 1624635492
transform 1 0 3588 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_30
timestamp 1624635492
transform 1 0 3864 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_36
timestamp 1624635492
transform 1 0 4416 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_41
timestamp 1624635492
transform 1 0 4876 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1624635492
transform 1 0 6440 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1624635492
transform -1 0 5980 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1624635492
transform -1 0 6716 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1624635492
transform -1 0 5244 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_45
timestamp 1624635492
transform 1 0 5244 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_49
timestamp 1624635492
transform 1 0 5612 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_53
timestamp 1624635492
transform 1 0 5980 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_57
timestamp 1624635492
transform 1 0 6348 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_61
timestamp 1624635492
transform 1 0 6716 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1624635492
transform 1 0 8096 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_73
timestamp 1624635492
transform 1 0 7820 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_79
timestamp 1624635492
transform 1 0 8372 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1624635492
transform 1 0 9108 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_88
timestamp 1624635492
transform 1 0 9200 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_100
timestamp 1624635492
transform 1 0 10304 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1624635492
transform 1 0 11776 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_112
timestamp 1624635492
transform 1 0 11408 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_117
timestamp 1624635492
transform 1 0 11868 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1624635492
transform 1 0 14444 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_129
timestamp 1624635492
transform 1 0 12972 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_141
timestamp 1624635492
transform 1 0 14076 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_146
timestamp 1624635492
transform 1 0 14536 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_158
timestamp 1624635492
transform 1 0 15640 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1624635492
transform 1 0 17112 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output90
timestamp 1624635492
transform -1 0 17756 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output120
timestamp 1624635492
transform 1 0 18124 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_170
timestamp 1624635492
transform 1 0 16744 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_175
timestamp 1624635492
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_181
timestamp 1624635492
transform 1 0 17756 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1624635492
transform 1 0 19780 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input88
timestamp 1624635492
transform -1 0 20332 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output118
timestamp 1624635492
transform 1 0 19228 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output119
timestamp 1624635492
transform 1 0 18676 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_189
timestamp 1624635492
transform 1 0 18492 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_195
timestamp 1624635492
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_201
timestamp 1624635492
transform 1 0 19596 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_204
timestamp 1624635492
transform 1 0 19872 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1624635492
transform -1 0 21896 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output116
timestamp 1624635492
transform 1 0 21068 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output117
timestamp 1624635492
transform 1 0 20516 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_209
timestamp 1624635492
transform 1 0 20332 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_215
timestamp 1624635492
transform 1 0 20884 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_221
timestamp 1624635492
transform 1 0 21436 0 1 20128
box -38 -48 222 592
<< labels >>
rlabel metal2 s 21822 0 21878 800 6 SC_IN_BOT
port 0 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 SC_OUT_BOT
port 1 nsew signal tristate
rlabel metal2 s 202 0 258 800 6 bottom_left_grid_pin_42_
port 2 nsew signal input
rlabel metal2 s 570 0 626 800 6 bottom_left_grid_pin_43_
port 3 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 bottom_left_grid_pin_44_
port 4 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 bottom_left_grid_pin_45_
port 5 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 bottom_left_grid_pin_46_
port 6 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 bottom_left_grid_pin_47_
port 7 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 bottom_left_grid_pin_48_
port 8 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 bottom_left_grid_pin_49_
port 9 nsew signal input
rlabel metal2 s 5722 22200 5778 23000 6 ccff_head
port 10 nsew signal input
rlabel metal2 s 17222 22200 17278 23000 6 ccff_tail
port 11 nsew signal tristate
rlabel metal3 s 0 3816 800 3936 6 chanx_left_in[0]
port 12 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 chanx_left_in[10]
port 13 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[11]
port 14 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[12]
port 15 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 chanx_left_in[13]
port 16 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[14]
port 17 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[15]
port 18 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[16]
port 19 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 chanx_left_in[17]
port 20 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[18]
port 21 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 chanx_left_in[19]
port 22 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 chanx_left_in[1]
port 23 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[2]
port 24 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 chanx_left_in[3]
port 25 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 chanx_left_in[4]
port 26 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 chanx_left_in[5]
port 27 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 chanx_left_in[6]
port 28 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 chanx_left_in[7]
port 29 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 chanx_left_in[8]
port 30 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[9]
port 31 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 chanx_left_out[0]
port 32 nsew signal tristate
rlabel metal3 s 0 17960 800 18080 6 chanx_left_out[10]
port 33 nsew signal tristate
rlabel metal3 s 0 18368 800 18488 6 chanx_left_out[11]
port 34 nsew signal tristate
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[12]
port 35 nsew signal tristate
rlabel metal3 s 0 19320 800 19440 6 chanx_left_out[13]
port 36 nsew signal tristate
rlabel metal3 s 0 19728 800 19848 6 chanx_left_out[14]
port 37 nsew signal tristate
rlabel metal3 s 0 20272 800 20392 6 chanx_left_out[15]
port 38 nsew signal tristate
rlabel metal3 s 0 20680 800 20800 6 chanx_left_out[16]
port 39 nsew signal tristate
rlabel metal3 s 0 21224 800 21344 6 chanx_left_out[17]
port 40 nsew signal tristate
rlabel metal3 s 0 21632 800 21752 6 chanx_left_out[18]
port 41 nsew signal tristate
rlabel metal3 s 0 22176 800 22296 6 chanx_left_out[19]
port 42 nsew signal tristate
rlabel metal3 s 0 13744 800 13864 6 chanx_left_out[1]
port 43 nsew signal tristate
rlabel metal3 s 0 14152 800 14272 6 chanx_left_out[2]
port 44 nsew signal tristate
rlabel metal3 s 0 14560 800 14680 6 chanx_left_out[3]
port 45 nsew signal tristate
rlabel metal3 s 0 15104 800 15224 6 chanx_left_out[4]
port 46 nsew signal tristate
rlabel metal3 s 0 15512 800 15632 6 chanx_left_out[5]
port 47 nsew signal tristate
rlabel metal3 s 0 16056 800 16176 6 chanx_left_out[6]
port 48 nsew signal tristate
rlabel metal3 s 0 16464 800 16584 6 chanx_left_out[7]
port 49 nsew signal tristate
rlabel metal3 s 0 17008 800 17128 6 chanx_left_out[8]
port 50 nsew signal tristate
rlabel metal3 s 0 17416 800 17536 6 chanx_left_out[9]
port 51 nsew signal tristate
rlabel metal3 s 22200 3816 23000 3936 6 chanx_right_in[0]
port 52 nsew signal input
rlabel metal3 s 22200 8576 23000 8696 6 chanx_right_in[10]
port 53 nsew signal input
rlabel metal3 s 22200 8984 23000 9104 6 chanx_right_in[11]
port 54 nsew signal input
rlabel metal3 s 22200 9392 23000 9512 6 chanx_right_in[12]
port 55 nsew signal input
rlabel metal3 s 22200 9936 23000 10056 6 chanx_right_in[13]
port 56 nsew signal input
rlabel metal3 s 22200 10344 23000 10464 6 chanx_right_in[14]
port 57 nsew signal input
rlabel metal3 s 22200 10888 23000 11008 6 chanx_right_in[15]
port 58 nsew signal input
rlabel metal3 s 22200 11296 23000 11416 6 chanx_right_in[16]
port 59 nsew signal input
rlabel metal3 s 22200 11840 23000 11960 6 chanx_right_in[17]
port 60 nsew signal input
rlabel metal3 s 22200 12248 23000 12368 6 chanx_right_in[18]
port 61 nsew signal input
rlabel metal3 s 22200 12792 23000 12912 6 chanx_right_in[19]
port 62 nsew signal input
rlabel metal3 s 22200 4360 23000 4480 6 chanx_right_in[1]
port 63 nsew signal input
rlabel metal3 s 22200 4768 23000 4888 6 chanx_right_in[2]
port 64 nsew signal input
rlabel metal3 s 22200 5176 23000 5296 6 chanx_right_in[3]
port 65 nsew signal input
rlabel metal3 s 22200 5720 23000 5840 6 chanx_right_in[4]
port 66 nsew signal input
rlabel metal3 s 22200 6128 23000 6248 6 chanx_right_in[5]
port 67 nsew signal input
rlabel metal3 s 22200 6672 23000 6792 6 chanx_right_in[6]
port 68 nsew signal input
rlabel metal3 s 22200 7080 23000 7200 6 chanx_right_in[7]
port 69 nsew signal input
rlabel metal3 s 22200 7624 23000 7744 6 chanx_right_in[8]
port 70 nsew signal input
rlabel metal3 s 22200 8032 23000 8152 6 chanx_right_in[9]
port 71 nsew signal input
rlabel metal3 s 22200 13200 23000 13320 6 chanx_right_out[0]
port 72 nsew signal tristate
rlabel metal3 s 22200 17960 23000 18080 6 chanx_right_out[10]
port 73 nsew signal tristate
rlabel metal3 s 22200 18368 23000 18488 6 chanx_right_out[11]
port 74 nsew signal tristate
rlabel metal3 s 22200 18776 23000 18896 6 chanx_right_out[12]
port 75 nsew signal tristate
rlabel metal3 s 22200 19320 23000 19440 6 chanx_right_out[13]
port 76 nsew signal tristate
rlabel metal3 s 22200 19728 23000 19848 6 chanx_right_out[14]
port 77 nsew signal tristate
rlabel metal3 s 22200 20272 23000 20392 6 chanx_right_out[15]
port 78 nsew signal tristate
rlabel metal3 s 22200 20680 23000 20800 6 chanx_right_out[16]
port 79 nsew signal tristate
rlabel metal3 s 22200 21224 23000 21344 6 chanx_right_out[17]
port 80 nsew signal tristate
rlabel metal3 s 22200 21632 23000 21752 6 chanx_right_out[18]
port 81 nsew signal tristate
rlabel metal3 s 22200 22176 23000 22296 6 chanx_right_out[19]
port 82 nsew signal tristate
rlabel metal3 s 22200 13744 23000 13864 6 chanx_right_out[1]
port 83 nsew signal tristate
rlabel metal3 s 22200 14152 23000 14272 6 chanx_right_out[2]
port 84 nsew signal tristate
rlabel metal3 s 22200 14560 23000 14680 6 chanx_right_out[3]
port 85 nsew signal tristate
rlabel metal3 s 22200 15104 23000 15224 6 chanx_right_out[4]
port 86 nsew signal tristate
rlabel metal3 s 22200 15512 23000 15632 6 chanx_right_out[5]
port 87 nsew signal tristate
rlabel metal3 s 22200 16056 23000 16176 6 chanx_right_out[6]
port 88 nsew signal tristate
rlabel metal3 s 22200 16464 23000 16584 6 chanx_right_out[7]
port 89 nsew signal tristate
rlabel metal3 s 22200 17008 23000 17128 6 chanx_right_out[8]
port 90 nsew signal tristate
rlabel metal3 s 22200 17416 23000 17536 6 chanx_right_out[9]
port 91 nsew signal tristate
rlabel metal2 s 3790 0 3846 800 6 chany_bottom_in[0]
port 92 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 chany_bottom_in[10]
port 93 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 chany_bottom_in[11]
port 94 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 chany_bottom_in[12]
port 95 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 chany_bottom_in[13]
port 96 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 chany_bottom_in[14]
port 97 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 chany_bottom_in[15]
port 98 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 chany_bottom_in[16]
port 99 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 chany_bottom_in[17]
port 100 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 chany_bottom_in[18]
port 101 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 chany_bottom_in[19]
port 102 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 chany_bottom_in[1]
port 103 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 chany_bottom_in[2]
port 104 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 chany_bottom_in[3]
port 105 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 chany_bottom_in[4]
port 106 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 chany_bottom_in[5]
port 107 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 chany_bottom_in[6]
port 108 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 chany_bottom_in[7]
port 109 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 chany_bottom_in[8]
port 110 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 chany_bottom_in[9]
port 111 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 chany_bottom_out[0]
port 112 nsew signal tristate
rlabel metal2 s 17314 0 17370 800 6 chany_bottom_out[10]
port 113 nsew signal tristate
rlabel metal2 s 17774 0 17830 800 6 chany_bottom_out[11]
port 114 nsew signal tristate
rlabel metal2 s 18234 0 18290 800 6 chany_bottom_out[12]
port 115 nsew signal tristate
rlabel metal2 s 18602 0 18658 800 6 chany_bottom_out[13]
port 116 nsew signal tristate
rlabel metal2 s 19062 0 19118 800 6 chany_bottom_out[14]
port 117 nsew signal tristate
rlabel metal2 s 19522 0 19578 800 6 chany_bottom_out[15]
port 118 nsew signal tristate
rlabel metal2 s 19982 0 20038 800 6 chany_bottom_out[16]
port 119 nsew signal tristate
rlabel metal2 s 20442 0 20498 800 6 chany_bottom_out[17]
port 120 nsew signal tristate
rlabel metal2 s 20902 0 20958 800 6 chany_bottom_out[18]
port 121 nsew signal tristate
rlabel metal2 s 21362 0 21418 800 6 chany_bottom_out[19]
port 122 nsew signal tristate
rlabel metal2 s 13266 0 13322 800 6 chany_bottom_out[1]
port 123 nsew signal tristate
rlabel metal2 s 13726 0 13782 800 6 chany_bottom_out[2]
port 124 nsew signal tristate
rlabel metal2 s 14094 0 14150 800 6 chany_bottom_out[3]
port 125 nsew signal tristate
rlabel metal2 s 14554 0 14610 800 6 chany_bottom_out[4]
port 126 nsew signal tristate
rlabel metal2 s 15014 0 15070 800 6 chany_bottom_out[5]
port 127 nsew signal tristate
rlabel metal2 s 15474 0 15530 800 6 chany_bottom_out[6]
port 128 nsew signal tristate
rlabel metal2 s 15934 0 15990 800 6 chany_bottom_out[7]
port 129 nsew signal tristate
rlabel metal2 s 16394 0 16450 800 6 chany_bottom_out[8]
port 130 nsew signal tristate
rlabel metal2 s 16854 0 16910 800 6 chany_bottom_out[9]
port 131 nsew signal tristate
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_34_
port 132 nsew signal input
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_35_
port 133 nsew signal input
rlabel metal3 s 0 960 800 1080 6 left_bottom_grid_pin_36_
port 134 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 left_bottom_grid_pin_37_
port 135 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 left_bottom_grid_pin_38_
port 136 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_39_
port 137 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 left_bottom_grid_pin_40_
port 138 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 left_bottom_grid_pin_41_
port 139 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 left_top_grid_pin_1_
port 140 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 prog_clk_0_S_in
port 141 nsew signal input
rlabel metal3 s 22200 144 23000 264 6 right_bottom_grid_pin_34_
port 142 nsew signal input
rlabel metal3 s 22200 552 23000 672 6 right_bottom_grid_pin_35_
port 143 nsew signal input
rlabel metal3 s 22200 960 23000 1080 6 right_bottom_grid_pin_36_
port 144 nsew signal input
rlabel metal3 s 22200 1504 23000 1624 6 right_bottom_grid_pin_37_
port 145 nsew signal input
rlabel metal3 s 22200 1912 23000 2032 6 right_bottom_grid_pin_38_
port 146 nsew signal input
rlabel metal3 s 22200 2456 23000 2576 6 right_bottom_grid_pin_39_
port 147 nsew signal input
rlabel metal3 s 22200 2864 23000 2984 6 right_bottom_grid_pin_40_
port 148 nsew signal input
rlabel metal3 s 22200 3408 23000 3528 6 right_bottom_grid_pin_41_
port 149 nsew signal input
rlabel metal3 s 22200 22584 23000 22704 6 right_top_grid_pin_1_
port 150 nsew signal input
rlabel metal4 s 18271 2128 18591 20720 6 VPWR
port 151 nsew power bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VPWR
port 152 nsew power bidirectional
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 153 nsew power bidirectional
rlabel metal4 s 14805 2128 15125 20720 6 VGND
port 154 nsew ground bidirectional
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 155 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
