magic
tech sky130A
magscale 1 2
timestamp 1679358067
<< obsli1 >>
rect 368 2159 494592 540753
<< obsm1 >>
rect 368 1980 494592 540784
<< metal2 >>
rect 3974 542200 4030 543000
rect 8482 542200 8538 543000
rect 12990 542200 13046 543000
rect 17498 542200 17554 543000
rect 22006 542200 22062 543000
rect 26514 542200 26570 543000
rect 31022 542200 31078 543000
rect 35530 542200 35586 543000
rect 40038 542200 40094 543000
rect 44546 542200 44602 543000
rect 49054 542200 49110 543000
rect 53562 542200 53618 543000
rect 58070 542200 58126 543000
rect 62578 542200 62634 543000
rect 67086 542200 67142 543000
rect 71594 542200 71650 543000
rect 76102 542200 76158 543000
rect 80610 542200 80666 543000
rect 85118 542200 85174 543000
rect 89626 542200 89682 543000
rect 94134 542200 94190 543000
rect 98642 542200 98698 543000
rect 103150 542200 103206 543000
rect 107658 542200 107714 543000
rect 112166 542200 112222 543000
rect 116674 542200 116730 543000
rect 121182 542200 121238 543000
rect 125690 542200 125746 543000
rect 130198 542200 130254 543000
rect 134706 542200 134762 543000
rect 139214 542200 139270 543000
rect 143722 542200 143778 543000
rect 148230 542200 148286 543000
rect 152738 542200 152794 543000
rect 157246 542200 157302 543000
rect 161754 542200 161810 543000
rect 166262 542200 166318 543000
rect 170770 542200 170826 543000
rect 175278 542200 175334 543000
rect 179786 542200 179842 543000
rect 184294 542200 184350 543000
rect 188802 542200 188858 543000
rect 193310 542200 193366 543000
rect 197818 542200 197874 543000
rect 202326 542200 202382 543000
rect 206834 542200 206890 543000
rect 211342 542200 211398 543000
rect 215850 542200 215906 543000
rect 220358 542200 220414 543000
rect 224866 542200 224922 543000
rect 229374 542200 229430 543000
rect 233882 542200 233938 543000
rect 238390 542200 238446 543000
rect 242898 542200 242954 543000
rect 247406 542200 247462 543000
rect 251914 542200 251970 543000
rect 256422 542200 256478 543000
rect 260930 542200 260986 543000
rect 265438 542200 265494 543000
rect 269946 542200 270002 543000
rect 274454 542200 274510 543000
rect 278962 542200 279018 543000
rect 283470 542200 283526 543000
rect 287978 542200 288034 543000
rect 292486 542200 292542 543000
rect 296994 542200 297050 543000
rect 301502 542200 301558 543000
rect 306010 542200 306066 543000
rect 310518 542200 310574 543000
rect 315026 542200 315082 543000
rect 319534 542200 319590 543000
rect 324042 542200 324098 543000
rect 328550 542200 328606 543000
rect 333058 542200 333114 543000
rect 337566 542200 337622 543000
rect 342074 542200 342130 543000
rect 346582 542200 346638 543000
rect 351090 542200 351146 543000
rect 355598 542200 355654 543000
rect 360106 542200 360162 543000
rect 364614 542200 364670 543000
rect 369122 542200 369178 543000
rect 373630 542200 373686 543000
rect 378138 542200 378194 543000
rect 382646 542200 382702 543000
rect 387154 542200 387210 543000
rect 391662 542200 391718 543000
rect 396170 542200 396226 543000
rect 400678 542200 400734 543000
rect 405186 542200 405242 543000
rect 409694 542200 409750 543000
rect 414202 542200 414258 543000
rect 418710 542200 418766 543000
rect 423218 542200 423274 543000
rect 427726 542200 427782 543000
rect 432234 542200 432290 543000
rect 436742 542200 436798 543000
rect 441250 542200 441306 543000
rect 445758 542200 445814 543000
rect 450266 542200 450322 543000
rect 454774 542200 454830 543000
rect 459282 542200 459338 543000
rect 463790 542200 463846 543000
rect 468298 542200 468354 543000
rect 472806 542200 472862 543000
rect 477314 542200 477370 543000
rect 481822 542200 481878 543000
rect 486330 542200 486386 543000
rect 490838 542200 490894 543000
rect 3974 0 4030 800
rect 9770 0 9826 800
rect 15566 0 15622 800
rect 21362 0 21418 800
rect 27158 0 27214 800
rect 32954 0 33010 800
rect 38750 0 38806 800
rect 44546 0 44602 800
rect 50342 0 50398 800
rect 56138 0 56194 800
rect 61934 0 61990 800
rect 67730 0 67786 800
rect 73526 0 73582 800
rect 79322 0 79378 800
rect 85118 0 85174 800
rect 90914 0 90970 800
rect 96710 0 96766 800
rect 102506 0 102562 800
rect 108302 0 108358 800
rect 114098 0 114154 800
rect 119894 0 119950 800
rect 125690 0 125746 800
rect 131486 0 131542 800
rect 137282 0 137338 800
rect 143078 0 143134 800
rect 148874 0 148930 800
rect 154670 0 154726 800
rect 160466 0 160522 800
rect 166262 0 166318 800
rect 172058 0 172114 800
rect 177854 0 177910 800
rect 183650 0 183706 800
rect 189446 0 189502 800
rect 195242 0 195298 800
rect 201038 0 201094 800
rect 206834 0 206890 800
rect 212630 0 212686 800
rect 218426 0 218482 800
rect 224222 0 224278 800
rect 230018 0 230074 800
rect 235814 0 235870 800
rect 241610 0 241666 800
rect 247406 0 247462 800
rect 253202 0 253258 800
rect 258998 0 259054 800
rect 264794 0 264850 800
rect 270590 0 270646 800
rect 276386 0 276442 800
rect 282182 0 282238 800
rect 287978 0 288034 800
rect 293774 0 293830 800
rect 299570 0 299626 800
rect 305366 0 305422 800
rect 311162 0 311218 800
rect 316958 0 317014 800
rect 322754 0 322810 800
rect 328550 0 328606 800
rect 334346 0 334402 800
rect 340142 0 340198 800
rect 345938 0 345994 800
rect 351734 0 351790 800
rect 357530 0 357586 800
rect 363326 0 363382 800
rect 369122 0 369178 800
rect 374918 0 374974 800
rect 380714 0 380770 800
rect 386510 0 386566 800
rect 392306 0 392362 800
rect 398102 0 398158 800
rect 403898 0 403954 800
rect 409694 0 409750 800
rect 415490 0 415546 800
rect 421286 0 421342 800
rect 427082 0 427138 800
rect 432878 0 432934 800
rect 438674 0 438730 800
rect 444470 0 444526 800
rect 450266 0 450322 800
rect 456062 0 456118 800
rect 461858 0 461914 800
rect 467654 0 467710 800
rect 473450 0 473506 800
rect 479246 0 479302 800
rect 485042 0 485098 800
rect 490838 0 490894 800
<< obsm2 >>
rect 754 542144 3918 542314
rect 4086 542144 8426 542314
rect 8594 542144 12934 542314
rect 13102 542144 17442 542314
rect 17610 542144 21950 542314
rect 22118 542144 26458 542314
rect 26626 542144 30966 542314
rect 31134 542144 35474 542314
rect 35642 542144 39982 542314
rect 40150 542144 44490 542314
rect 44658 542144 48998 542314
rect 49166 542144 53506 542314
rect 53674 542144 58014 542314
rect 58182 542144 62522 542314
rect 62690 542144 67030 542314
rect 67198 542144 71538 542314
rect 71706 542144 76046 542314
rect 76214 542144 80554 542314
rect 80722 542144 85062 542314
rect 85230 542144 89570 542314
rect 89738 542144 94078 542314
rect 94246 542144 98586 542314
rect 98754 542144 103094 542314
rect 103262 542144 107602 542314
rect 107770 542144 112110 542314
rect 112278 542144 116618 542314
rect 116786 542144 121126 542314
rect 121294 542144 125634 542314
rect 125802 542144 130142 542314
rect 130310 542144 134650 542314
rect 134818 542144 139158 542314
rect 139326 542144 143666 542314
rect 143834 542144 148174 542314
rect 148342 542144 152682 542314
rect 152850 542144 157190 542314
rect 157358 542144 161698 542314
rect 161866 542144 166206 542314
rect 166374 542144 170714 542314
rect 170882 542144 175222 542314
rect 175390 542144 179730 542314
rect 179898 542144 184238 542314
rect 184406 542144 188746 542314
rect 188914 542144 193254 542314
rect 193422 542144 197762 542314
rect 197930 542144 202270 542314
rect 202438 542144 206778 542314
rect 206946 542144 211286 542314
rect 211454 542144 215794 542314
rect 215962 542144 220302 542314
rect 220470 542144 224810 542314
rect 224978 542144 229318 542314
rect 229486 542144 233826 542314
rect 233994 542144 238334 542314
rect 238502 542144 242842 542314
rect 243010 542144 247350 542314
rect 247518 542144 251858 542314
rect 252026 542144 256366 542314
rect 256534 542144 260874 542314
rect 261042 542144 265382 542314
rect 265550 542144 269890 542314
rect 270058 542144 274398 542314
rect 274566 542144 278906 542314
rect 279074 542144 283414 542314
rect 283582 542144 287922 542314
rect 288090 542144 292430 542314
rect 292598 542144 296938 542314
rect 297106 542144 301446 542314
rect 301614 542144 305954 542314
rect 306122 542144 310462 542314
rect 310630 542144 314970 542314
rect 315138 542144 319478 542314
rect 319646 542144 323986 542314
rect 324154 542144 328494 542314
rect 328662 542144 333002 542314
rect 333170 542144 337510 542314
rect 337678 542144 342018 542314
rect 342186 542144 346526 542314
rect 346694 542144 351034 542314
rect 351202 542144 355542 542314
rect 355710 542144 360050 542314
rect 360218 542144 364558 542314
rect 364726 542144 369066 542314
rect 369234 542144 373574 542314
rect 373742 542144 378082 542314
rect 378250 542144 382590 542314
rect 382758 542144 387098 542314
rect 387266 542144 391606 542314
rect 391774 542144 396114 542314
rect 396282 542144 400622 542314
rect 400790 542144 405130 542314
rect 405298 542144 409638 542314
rect 409806 542144 414146 542314
rect 414314 542144 418654 542314
rect 418822 542144 423162 542314
rect 423330 542144 427670 542314
rect 427838 542144 432178 542314
rect 432346 542144 436686 542314
rect 436854 542144 441194 542314
rect 441362 542144 445702 542314
rect 445870 542144 450210 542314
rect 450378 542144 454718 542314
rect 454886 542144 459226 542314
rect 459394 542144 463734 542314
rect 463902 542144 468242 542314
rect 468410 542144 472750 542314
rect 472918 542144 477258 542314
rect 477426 542144 481766 542314
rect 481934 542144 486274 542314
rect 486442 542144 490782 542314
rect 490950 542144 494204 542314
rect 754 856 494204 542144
rect 754 734 3918 856
rect 4086 734 9714 856
rect 9882 734 15510 856
rect 15678 734 21306 856
rect 21474 734 27102 856
rect 27270 734 32898 856
rect 33066 734 38694 856
rect 38862 734 44490 856
rect 44658 734 50286 856
rect 50454 734 56082 856
rect 56250 734 61878 856
rect 62046 734 67674 856
rect 67842 734 73470 856
rect 73638 734 79266 856
rect 79434 734 85062 856
rect 85230 734 90858 856
rect 91026 734 96654 856
rect 96822 734 102450 856
rect 102618 734 108246 856
rect 108414 734 114042 856
rect 114210 734 119838 856
rect 120006 734 125634 856
rect 125802 734 131430 856
rect 131598 734 137226 856
rect 137394 734 143022 856
rect 143190 734 148818 856
rect 148986 734 154614 856
rect 154782 734 160410 856
rect 160578 734 166206 856
rect 166374 734 172002 856
rect 172170 734 177798 856
rect 177966 734 183594 856
rect 183762 734 189390 856
rect 189558 734 195186 856
rect 195354 734 200982 856
rect 201150 734 206778 856
rect 206946 734 212574 856
rect 212742 734 218370 856
rect 218538 734 224166 856
rect 224334 734 229962 856
rect 230130 734 235758 856
rect 235926 734 241554 856
rect 241722 734 247350 856
rect 247518 734 253146 856
rect 253314 734 258942 856
rect 259110 734 264738 856
rect 264906 734 270534 856
rect 270702 734 276330 856
rect 276498 734 282126 856
rect 282294 734 287922 856
rect 288090 734 293718 856
rect 293886 734 299514 856
rect 299682 734 305310 856
rect 305478 734 311106 856
rect 311274 734 316902 856
rect 317070 734 322698 856
rect 322866 734 328494 856
rect 328662 734 334290 856
rect 334458 734 340086 856
rect 340254 734 345882 856
rect 346050 734 351678 856
rect 351846 734 357474 856
rect 357642 734 363270 856
rect 363438 734 369066 856
rect 369234 734 374862 856
rect 375030 734 380658 856
rect 380826 734 386454 856
rect 386622 734 392250 856
rect 392418 734 398046 856
rect 398214 734 403842 856
rect 404010 734 409638 856
rect 409806 734 415434 856
rect 415602 734 421230 856
rect 421398 734 427026 856
rect 427194 734 432822 856
rect 432990 734 438618 856
rect 438786 734 444414 856
rect 444582 734 450210 856
rect 450378 734 456006 856
rect 456174 734 461802 856
rect 461970 734 467598 856
rect 467766 734 473394 856
rect 473562 734 479190 856
rect 479358 734 484986 856
rect 485154 734 490782 856
rect 490950 734 494204 856
<< metal3 >>
rect 0 537888 800 538008
rect 494200 536528 495000 536648
rect 0 532448 800 532568
rect 494200 531224 495000 531344
rect 0 527008 800 527128
rect 494200 525920 495000 526040
rect 0 521568 800 521688
rect 494200 520616 495000 520736
rect 0 516128 800 516248
rect 494200 515312 495000 515432
rect 0 510688 800 510808
rect 494200 510008 495000 510128
rect 0 505248 800 505368
rect 494200 504704 495000 504824
rect 0 499808 800 499928
rect 494200 499400 495000 499520
rect 0 494368 800 494488
rect 494200 494096 495000 494216
rect 0 488928 800 489048
rect 494200 488792 495000 488912
rect 0 483488 800 483608
rect 494200 483488 495000 483608
rect 0 478048 800 478168
rect 494200 478184 495000 478304
rect 494200 472880 495000 473000
rect 0 472608 800 472728
rect 494200 467576 495000 467696
rect 0 467168 800 467288
rect 494200 462272 495000 462392
rect 0 461728 800 461848
rect 494200 456968 495000 457088
rect 0 456288 800 456408
rect 494200 451664 495000 451784
rect 0 450848 800 450968
rect 494200 446360 495000 446480
rect 0 445408 800 445528
rect 494200 441056 495000 441176
rect 0 439968 800 440088
rect 494200 435752 495000 435872
rect 0 434528 800 434648
rect 494200 430448 495000 430568
rect 0 429088 800 429208
rect 494200 425144 495000 425264
rect 0 423648 800 423768
rect 494200 419840 495000 419960
rect 0 418208 800 418328
rect 494200 414536 495000 414656
rect 0 412768 800 412888
rect 494200 409232 495000 409352
rect 0 407328 800 407448
rect 494200 403928 495000 404048
rect 0 401888 800 402008
rect 494200 398624 495000 398744
rect 0 396448 800 396568
rect 494200 393320 495000 393440
rect 0 391008 800 391128
rect 494200 388016 495000 388136
rect 0 385568 800 385688
rect 494200 382712 495000 382832
rect 0 380128 800 380248
rect 494200 377408 495000 377528
rect 0 374688 800 374808
rect 494200 372104 495000 372224
rect 0 369248 800 369368
rect 494200 366800 495000 366920
rect 0 363808 800 363928
rect 494200 361496 495000 361616
rect 0 358368 800 358488
rect 494200 356192 495000 356312
rect 0 352928 800 353048
rect 494200 350888 495000 351008
rect 0 347488 800 347608
rect 494200 345584 495000 345704
rect 0 342048 800 342168
rect 494200 340280 495000 340400
rect 0 336608 800 336728
rect 494200 334976 495000 335096
rect 0 331168 800 331288
rect 494200 329672 495000 329792
rect 0 325728 800 325848
rect 494200 324368 495000 324488
rect 0 320288 800 320408
rect 494200 319064 495000 319184
rect 0 314848 800 314968
rect 494200 313760 495000 313880
rect 0 309408 800 309528
rect 494200 308456 495000 308576
rect 0 303968 800 304088
rect 494200 303152 495000 303272
rect 0 298528 800 298648
rect 494200 297848 495000 297968
rect 0 293088 800 293208
rect 494200 292544 495000 292664
rect 0 287648 800 287768
rect 494200 287240 495000 287360
rect 0 282208 800 282328
rect 494200 281936 495000 282056
rect 0 276768 800 276888
rect 494200 276632 495000 276752
rect 0 271328 800 271448
rect 494200 271328 495000 271448
rect 0 265888 800 266008
rect 494200 266024 495000 266144
rect 494200 260720 495000 260840
rect 0 260448 800 260568
rect 494200 255416 495000 255536
rect 0 255008 800 255128
rect 494200 250112 495000 250232
rect 0 249568 800 249688
rect 494200 244808 495000 244928
rect 0 244128 800 244248
rect 494200 239504 495000 239624
rect 0 238688 800 238808
rect 494200 234200 495000 234320
rect 0 233248 800 233368
rect 494200 228896 495000 229016
rect 0 227808 800 227928
rect 494200 223592 495000 223712
rect 0 222368 800 222488
rect 494200 218288 495000 218408
rect 0 216928 800 217048
rect 494200 212984 495000 213104
rect 0 211488 800 211608
rect 494200 207680 495000 207800
rect 0 206048 800 206168
rect 494200 202376 495000 202496
rect 0 200608 800 200728
rect 494200 197072 495000 197192
rect 0 195168 800 195288
rect 494200 191768 495000 191888
rect 0 189728 800 189848
rect 494200 186464 495000 186584
rect 0 184288 800 184408
rect 494200 181160 495000 181280
rect 0 178848 800 178968
rect 494200 175856 495000 175976
rect 0 173408 800 173528
rect 494200 170552 495000 170672
rect 0 167968 800 168088
rect 494200 165248 495000 165368
rect 0 162528 800 162648
rect 494200 159944 495000 160064
rect 0 157088 800 157208
rect 494200 154640 495000 154760
rect 0 151648 800 151768
rect 494200 149336 495000 149456
rect 0 146208 800 146328
rect 494200 144032 495000 144152
rect 0 140768 800 140888
rect 494200 138728 495000 138848
rect 0 135328 800 135448
rect 494200 133424 495000 133544
rect 0 129888 800 130008
rect 494200 128120 495000 128240
rect 0 124448 800 124568
rect 494200 122816 495000 122936
rect 0 119008 800 119128
rect 494200 117512 495000 117632
rect 0 113568 800 113688
rect 494200 112208 495000 112328
rect 0 108128 800 108248
rect 494200 106904 495000 107024
rect 0 102688 800 102808
rect 494200 101600 495000 101720
rect 0 97248 800 97368
rect 494200 96296 495000 96416
rect 0 91808 800 91928
rect 494200 90992 495000 91112
rect 0 86368 800 86488
rect 494200 85688 495000 85808
rect 0 80928 800 81048
rect 494200 80384 495000 80504
rect 0 75488 800 75608
rect 494200 75080 495000 75200
rect 0 70048 800 70168
rect 494200 69776 495000 69896
rect 0 64608 800 64728
rect 494200 64472 495000 64592
rect 0 59168 800 59288
rect 494200 59168 495000 59288
rect 0 53728 800 53848
rect 494200 53864 495000 53984
rect 494200 48560 495000 48680
rect 0 48288 800 48408
rect 494200 43256 495000 43376
rect 0 42848 800 42968
rect 494200 37952 495000 38072
rect 0 37408 800 37528
rect 494200 32648 495000 32768
rect 0 31968 800 32088
rect 494200 27344 495000 27464
rect 0 26528 800 26648
rect 494200 22040 495000 22160
rect 0 21088 800 21208
rect 494200 16736 495000 16856
rect 0 15648 800 15768
rect 494200 11432 495000 11552
rect 0 10208 800 10328
rect 494200 6128 495000 6248
rect 0 4768 800 4888
<< obsm3 >>
rect 749 538088 494200 540769
rect 880 537808 494200 538088
rect 749 536728 494200 537808
rect 749 536448 494120 536728
rect 749 532648 494200 536448
rect 880 532368 494200 532648
rect 749 531424 494200 532368
rect 749 531144 494120 531424
rect 749 527208 494200 531144
rect 880 526928 494200 527208
rect 749 526120 494200 526928
rect 749 525840 494120 526120
rect 749 521768 494200 525840
rect 880 521488 494200 521768
rect 749 520816 494200 521488
rect 749 520536 494120 520816
rect 749 516328 494200 520536
rect 880 516048 494200 516328
rect 749 515512 494200 516048
rect 749 515232 494120 515512
rect 749 510888 494200 515232
rect 880 510608 494200 510888
rect 749 510208 494200 510608
rect 749 509928 494120 510208
rect 749 505448 494200 509928
rect 880 505168 494200 505448
rect 749 504904 494200 505168
rect 749 504624 494120 504904
rect 749 500008 494200 504624
rect 880 499728 494200 500008
rect 749 499600 494200 499728
rect 749 499320 494120 499600
rect 749 494568 494200 499320
rect 880 494296 494200 494568
rect 880 494288 494120 494296
rect 749 494016 494120 494288
rect 749 489128 494200 494016
rect 880 488992 494200 489128
rect 880 488848 494120 488992
rect 749 488712 494120 488848
rect 749 483688 494200 488712
rect 880 483408 494120 483688
rect 749 478384 494200 483408
rect 749 478248 494120 478384
rect 880 478104 494120 478248
rect 880 477968 494200 478104
rect 749 473080 494200 477968
rect 749 472808 494120 473080
rect 880 472800 494120 472808
rect 880 472528 494200 472800
rect 749 467776 494200 472528
rect 749 467496 494120 467776
rect 749 467368 494200 467496
rect 880 467088 494200 467368
rect 749 462472 494200 467088
rect 749 462192 494120 462472
rect 749 461928 494200 462192
rect 880 461648 494200 461928
rect 749 457168 494200 461648
rect 749 456888 494120 457168
rect 749 456488 494200 456888
rect 880 456208 494200 456488
rect 749 451864 494200 456208
rect 749 451584 494120 451864
rect 749 451048 494200 451584
rect 880 450768 494200 451048
rect 749 446560 494200 450768
rect 749 446280 494120 446560
rect 749 445608 494200 446280
rect 880 445328 494200 445608
rect 749 441256 494200 445328
rect 749 440976 494120 441256
rect 749 440168 494200 440976
rect 880 439888 494200 440168
rect 749 435952 494200 439888
rect 749 435672 494120 435952
rect 749 434728 494200 435672
rect 880 434448 494200 434728
rect 749 430648 494200 434448
rect 749 430368 494120 430648
rect 749 429288 494200 430368
rect 880 429008 494200 429288
rect 749 425344 494200 429008
rect 749 425064 494120 425344
rect 749 423848 494200 425064
rect 880 423568 494200 423848
rect 749 420040 494200 423568
rect 749 419760 494120 420040
rect 749 418408 494200 419760
rect 880 418128 494200 418408
rect 749 414736 494200 418128
rect 749 414456 494120 414736
rect 749 412968 494200 414456
rect 880 412688 494200 412968
rect 749 409432 494200 412688
rect 749 409152 494120 409432
rect 749 407528 494200 409152
rect 880 407248 494200 407528
rect 749 404128 494200 407248
rect 749 403848 494120 404128
rect 749 402088 494200 403848
rect 880 401808 494200 402088
rect 749 398824 494200 401808
rect 749 398544 494120 398824
rect 749 396648 494200 398544
rect 880 396368 494200 396648
rect 749 393520 494200 396368
rect 749 393240 494120 393520
rect 749 391208 494200 393240
rect 880 390928 494200 391208
rect 749 388216 494200 390928
rect 749 387936 494120 388216
rect 749 385768 494200 387936
rect 880 385488 494200 385768
rect 749 382912 494200 385488
rect 749 382632 494120 382912
rect 749 380328 494200 382632
rect 880 380048 494200 380328
rect 749 377608 494200 380048
rect 749 377328 494120 377608
rect 749 374888 494200 377328
rect 880 374608 494200 374888
rect 749 372304 494200 374608
rect 749 372024 494120 372304
rect 749 369448 494200 372024
rect 880 369168 494200 369448
rect 749 367000 494200 369168
rect 749 366720 494120 367000
rect 749 364008 494200 366720
rect 880 363728 494200 364008
rect 749 361696 494200 363728
rect 749 361416 494120 361696
rect 749 358568 494200 361416
rect 880 358288 494200 358568
rect 749 356392 494200 358288
rect 749 356112 494120 356392
rect 749 353128 494200 356112
rect 880 352848 494200 353128
rect 749 351088 494200 352848
rect 749 350808 494120 351088
rect 749 347688 494200 350808
rect 880 347408 494200 347688
rect 749 345784 494200 347408
rect 749 345504 494120 345784
rect 749 342248 494200 345504
rect 880 341968 494200 342248
rect 749 340480 494200 341968
rect 749 340200 494120 340480
rect 749 336808 494200 340200
rect 880 336528 494200 336808
rect 749 335176 494200 336528
rect 749 334896 494120 335176
rect 749 331368 494200 334896
rect 880 331088 494200 331368
rect 749 329872 494200 331088
rect 749 329592 494120 329872
rect 749 325928 494200 329592
rect 880 325648 494200 325928
rect 749 324568 494200 325648
rect 749 324288 494120 324568
rect 749 320488 494200 324288
rect 880 320208 494200 320488
rect 749 319264 494200 320208
rect 749 318984 494120 319264
rect 749 315048 494200 318984
rect 880 314768 494200 315048
rect 749 313960 494200 314768
rect 749 313680 494120 313960
rect 749 309608 494200 313680
rect 880 309328 494200 309608
rect 749 308656 494200 309328
rect 749 308376 494120 308656
rect 749 304168 494200 308376
rect 880 303888 494200 304168
rect 749 303352 494200 303888
rect 749 303072 494120 303352
rect 749 298728 494200 303072
rect 880 298448 494200 298728
rect 749 298048 494200 298448
rect 749 297768 494120 298048
rect 749 293288 494200 297768
rect 880 293008 494200 293288
rect 749 292744 494200 293008
rect 749 292464 494120 292744
rect 749 287848 494200 292464
rect 880 287568 494200 287848
rect 749 287440 494200 287568
rect 749 287160 494120 287440
rect 749 282408 494200 287160
rect 880 282136 494200 282408
rect 880 282128 494120 282136
rect 749 281856 494120 282128
rect 749 276968 494200 281856
rect 880 276832 494200 276968
rect 880 276688 494120 276832
rect 749 276552 494120 276688
rect 749 271528 494200 276552
rect 880 271248 494120 271528
rect 749 266224 494200 271248
rect 749 266088 494120 266224
rect 880 265944 494120 266088
rect 880 265808 494200 265944
rect 749 260920 494200 265808
rect 749 260648 494120 260920
rect 880 260640 494120 260648
rect 880 260368 494200 260640
rect 749 255616 494200 260368
rect 749 255336 494120 255616
rect 749 255208 494200 255336
rect 880 254928 494200 255208
rect 749 250312 494200 254928
rect 749 250032 494120 250312
rect 749 249768 494200 250032
rect 880 249488 494200 249768
rect 749 245008 494200 249488
rect 749 244728 494120 245008
rect 749 244328 494200 244728
rect 880 244048 494200 244328
rect 749 239704 494200 244048
rect 749 239424 494120 239704
rect 749 238888 494200 239424
rect 880 238608 494200 238888
rect 749 234400 494200 238608
rect 749 234120 494120 234400
rect 749 233448 494200 234120
rect 880 233168 494200 233448
rect 749 229096 494200 233168
rect 749 228816 494120 229096
rect 749 228008 494200 228816
rect 880 227728 494200 228008
rect 749 223792 494200 227728
rect 749 223512 494120 223792
rect 749 222568 494200 223512
rect 880 222288 494200 222568
rect 749 218488 494200 222288
rect 749 218208 494120 218488
rect 749 217128 494200 218208
rect 880 216848 494200 217128
rect 749 213184 494200 216848
rect 749 212904 494120 213184
rect 749 211688 494200 212904
rect 880 211408 494200 211688
rect 749 207880 494200 211408
rect 749 207600 494120 207880
rect 749 206248 494200 207600
rect 880 205968 494200 206248
rect 749 202576 494200 205968
rect 749 202296 494120 202576
rect 749 200808 494200 202296
rect 880 200528 494200 200808
rect 749 197272 494200 200528
rect 749 196992 494120 197272
rect 749 195368 494200 196992
rect 880 195088 494200 195368
rect 749 191968 494200 195088
rect 749 191688 494120 191968
rect 749 189928 494200 191688
rect 880 189648 494200 189928
rect 749 186664 494200 189648
rect 749 186384 494120 186664
rect 749 184488 494200 186384
rect 880 184208 494200 184488
rect 749 181360 494200 184208
rect 749 181080 494120 181360
rect 749 179048 494200 181080
rect 880 178768 494200 179048
rect 749 176056 494200 178768
rect 749 175776 494120 176056
rect 749 173608 494200 175776
rect 880 173328 494200 173608
rect 749 170752 494200 173328
rect 749 170472 494120 170752
rect 749 168168 494200 170472
rect 880 167888 494200 168168
rect 749 165448 494200 167888
rect 749 165168 494120 165448
rect 749 162728 494200 165168
rect 880 162448 494200 162728
rect 749 160144 494200 162448
rect 749 159864 494120 160144
rect 749 157288 494200 159864
rect 880 157008 494200 157288
rect 749 154840 494200 157008
rect 749 154560 494120 154840
rect 749 151848 494200 154560
rect 880 151568 494200 151848
rect 749 149536 494200 151568
rect 749 149256 494120 149536
rect 749 146408 494200 149256
rect 880 146128 494200 146408
rect 749 144232 494200 146128
rect 749 143952 494120 144232
rect 749 140968 494200 143952
rect 880 140688 494200 140968
rect 749 138928 494200 140688
rect 749 138648 494120 138928
rect 749 135528 494200 138648
rect 880 135248 494200 135528
rect 749 133624 494200 135248
rect 749 133344 494120 133624
rect 749 130088 494200 133344
rect 880 129808 494200 130088
rect 749 128320 494200 129808
rect 749 128040 494120 128320
rect 749 124648 494200 128040
rect 880 124368 494200 124648
rect 749 123016 494200 124368
rect 749 122736 494120 123016
rect 749 119208 494200 122736
rect 880 118928 494200 119208
rect 749 117712 494200 118928
rect 749 117432 494120 117712
rect 749 113768 494200 117432
rect 880 113488 494200 113768
rect 749 112408 494200 113488
rect 749 112128 494120 112408
rect 749 108328 494200 112128
rect 880 108048 494200 108328
rect 749 107104 494200 108048
rect 749 106824 494120 107104
rect 749 102888 494200 106824
rect 880 102608 494200 102888
rect 749 101800 494200 102608
rect 749 101520 494120 101800
rect 749 97448 494200 101520
rect 880 97168 494200 97448
rect 749 96496 494200 97168
rect 749 96216 494120 96496
rect 749 92008 494200 96216
rect 880 91728 494200 92008
rect 749 91192 494200 91728
rect 749 90912 494120 91192
rect 749 86568 494200 90912
rect 880 86288 494200 86568
rect 749 85888 494200 86288
rect 749 85608 494120 85888
rect 749 81128 494200 85608
rect 880 80848 494200 81128
rect 749 80584 494200 80848
rect 749 80304 494120 80584
rect 749 75688 494200 80304
rect 880 75408 494200 75688
rect 749 75280 494200 75408
rect 749 75000 494120 75280
rect 749 70248 494200 75000
rect 880 69976 494200 70248
rect 880 69968 494120 69976
rect 749 69696 494120 69968
rect 749 64808 494200 69696
rect 880 64672 494200 64808
rect 880 64528 494120 64672
rect 749 64392 494120 64528
rect 749 59368 494200 64392
rect 880 59088 494120 59368
rect 749 54064 494200 59088
rect 749 53928 494120 54064
rect 880 53784 494120 53928
rect 880 53648 494200 53784
rect 749 48760 494200 53648
rect 749 48488 494120 48760
rect 880 48480 494120 48488
rect 880 48208 494200 48480
rect 749 43456 494200 48208
rect 749 43176 494120 43456
rect 749 43048 494200 43176
rect 880 42768 494200 43048
rect 749 38152 494200 42768
rect 749 37872 494120 38152
rect 749 37608 494200 37872
rect 880 37328 494200 37608
rect 749 32848 494200 37328
rect 749 32568 494120 32848
rect 749 32168 494200 32568
rect 880 31888 494200 32168
rect 749 27544 494200 31888
rect 749 27264 494120 27544
rect 749 26728 494200 27264
rect 880 26448 494200 26728
rect 749 22240 494200 26448
rect 749 21960 494120 22240
rect 749 21288 494200 21960
rect 880 21008 494200 21288
rect 749 16936 494200 21008
rect 749 16656 494120 16936
rect 749 15848 494200 16656
rect 880 15568 494200 15848
rect 749 11632 494200 15568
rect 749 11352 494120 11632
rect 749 10408 494200 11352
rect 880 10128 494200 10408
rect 749 6328 494200 10128
rect 749 6048 494120 6328
rect 749 4968 494200 6048
rect 880 4688 494200 4968
rect 749 2143 494200 4688
<< metal4 >>
rect -2552 -744 -1592 543656
rect -1192 616 -232 542296
rect 1024 -744 1664 543656
rect 1984 -744 2624 543656
rect 12424 34273 13064 543656
rect 13384 536508 14024 543656
rect 23824 536508 24464 543656
rect 24784 523777 25424 543656
rect 13384 473508 14024 480068
rect 23824 473508 24464 480068
rect 24784 473017 25424 480423
rect 13384 410508 14024 417068
rect 23824 410508 24464 417068
rect 24784 410017 25424 417831
rect 13384 347508 14024 354068
rect 23824 347508 24464 354068
rect 24784 347017 25424 354831
rect 13384 284508 14024 291068
rect 23824 284508 24464 291068
rect 24784 284017 25424 291831
rect 13384 221508 14024 228068
rect 23824 221508 24464 228068
rect 24784 221017 25424 228831
rect 13384 158508 14024 165068
rect 23824 158508 24464 165068
rect 24784 158017 25424 165831
rect 13384 95508 14024 102068
rect 23824 95508 24464 102068
rect 24784 95017 25424 102831
rect 13384 34273 14024 39068
rect 23824 34273 24464 39068
rect 24784 34273 25424 39831
rect 12424 -744 13064 13495
rect 13384 -744 14024 6068
rect 23824 -744 24464 6068
rect 24784 -744 25424 13495
rect 35224 -744 35864 543656
rect 36184 -744 36824 543656
rect 46624 536508 47264 543656
rect 47584 531257 48224 543656
rect 58024 531257 58664 543656
rect 58984 531257 59624 543656
rect 69424 531257 70064 543656
rect 70384 531257 71024 543656
rect 80824 531257 81464 543656
rect 81784 536508 82424 543656
rect 46624 473508 47264 480068
rect 47584 468801 48224 484231
rect 58024 468801 58664 484231
rect 58984 468801 59624 484231
rect 69424 468801 70064 484231
rect 70384 468801 71024 484231
rect 80824 468801 81464 484231
rect 81784 473508 82424 480068
rect 46624 410508 47264 417068
rect 47584 405801 48224 422591
rect 58024 405801 58664 422591
rect 58984 405801 59624 422591
rect 69424 405801 70064 422591
rect 70384 405801 71024 422591
rect 80824 405801 81464 422591
rect 81784 410508 82424 417068
rect 46624 347508 47264 354068
rect 47584 342801 48224 359591
rect 58024 342801 58664 359591
rect 58984 342801 59624 359591
rect 69424 342801 70064 359591
rect 70384 342801 71024 359591
rect 80824 342801 81464 359591
rect 81784 347508 82424 354068
rect 46624 284508 47264 291068
rect 47584 279801 48224 296591
rect 58024 279801 58664 296591
rect 58984 279801 59624 296591
rect 69424 279801 70064 296591
rect 70384 279801 71024 296591
rect 80824 279801 81464 296591
rect 81784 284508 82424 291068
rect 46624 221508 47264 228068
rect 47584 216801 48224 233591
rect 58024 216801 58664 233591
rect 58984 216801 59624 233591
rect 69424 216801 70064 233591
rect 70384 216801 71024 233591
rect 80824 216801 81464 233591
rect 81784 221508 82424 228068
rect 46624 158508 47264 165068
rect 47584 153801 48224 170591
rect 58024 153801 58664 170591
rect 58984 153801 59624 170591
rect 69424 153801 70064 170591
rect 70384 153801 71024 170591
rect 80824 153801 81464 170591
rect 81784 158508 82424 165068
rect 46624 95508 47264 102068
rect 47584 90801 48224 107591
rect 58024 90801 58664 107591
rect 58984 90801 59624 107591
rect 69424 90801 70064 107591
rect 70384 90801 71024 107591
rect 80824 90801 81464 107591
rect 81784 95508 82424 102068
rect 46624 32588 47264 39068
rect 46624 -744 47264 6068
rect 47584 -744 48224 44591
rect 58024 33049 58664 44591
rect 58984 33049 59624 44591
rect 69424 33049 70064 44591
rect 70384 33049 71024 44591
rect 58024 -744 58664 13495
rect 58984 -744 59624 13495
rect 69424 -744 70064 13495
rect 70384 -744 71024 13495
rect 80824 -744 81464 44591
rect 81784 32588 82424 39068
rect 81784 -744 82424 6068
rect 92224 -744 92864 543656
rect 93184 -744 93824 543656
rect 103624 536508 104264 543656
rect 104584 531257 105224 543656
rect 115024 531257 115664 543656
rect 115984 531257 116624 543656
rect 126424 531257 127064 543656
rect 127384 531257 128024 543656
rect 137824 531257 138464 543656
rect 138784 536508 139424 543656
rect 103624 473508 104264 480068
rect 104584 468801 105224 484231
rect 115024 468801 115664 484231
rect 115984 468801 116624 484231
rect 126424 468801 127064 484231
rect 127384 468801 128024 484231
rect 137824 468801 138464 484231
rect 138784 473508 139424 480068
rect 103624 410508 104264 417068
rect 104584 405801 105224 422591
rect 115024 405801 115664 422591
rect 115984 405801 116624 422591
rect 126424 405801 127064 422591
rect 127384 405801 128024 422591
rect 137824 405801 138464 422591
rect 138784 410508 139424 417068
rect 103624 347508 104264 354068
rect 104584 342801 105224 359591
rect 115024 342801 115664 359591
rect 115984 342801 116624 359591
rect 126424 342801 127064 359591
rect 127384 342801 128024 359591
rect 137824 342801 138464 359591
rect 138784 347508 139424 354068
rect 103624 284508 104264 291068
rect 104584 279801 105224 296591
rect 115024 279801 115664 296591
rect 115984 279801 116624 296591
rect 126424 279801 127064 296591
rect 127384 279801 128024 296591
rect 137824 279801 138464 296591
rect 138784 284508 139424 291068
rect 103624 221508 104264 228068
rect 104584 216801 105224 233591
rect 115024 216801 115664 233591
rect 115984 216801 116624 233591
rect 126424 216801 127064 233591
rect 127384 216801 128024 233591
rect 137824 216801 138464 233591
rect 138784 221508 139424 228068
rect 103624 158508 104264 165068
rect 104584 153801 105224 170591
rect 115024 153801 115664 170591
rect 115984 153801 116624 170591
rect 126424 153801 127064 170591
rect 127384 153801 128024 170591
rect 137824 153801 138464 170591
rect 138784 158508 139424 165068
rect 103624 95508 104264 102068
rect 104584 90801 105224 107591
rect 115024 90801 115664 107591
rect 115984 90801 116624 107591
rect 126424 90801 127064 107591
rect 127384 90801 128024 107591
rect 137824 90801 138464 107591
rect 138784 95508 139424 102068
rect 103624 32588 104264 39068
rect 103624 -744 104264 6068
rect 104584 -744 105224 44591
rect 115024 33049 115664 44591
rect 115984 33049 116624 44591
rect 126424 33049 127064 44591
rect 127384 33049 128024 44591
rect 115024 -744 115664 13495
rect 115984 -744 116624 13495
rect 126424 -744 127064 13495
rect 127384 -744 128024 13495
rect 137824 -744 138464 44591
rect 138784 32588 139424 39068
rect 138784 -744 139424 6068
rect 149224 -744 149864 543656
rect 150184 -744 150824 543656
rect 160624 536508 161264 543656
rect 161584 531257 162224 543656
rect 172024 531257 172664 543656
rect 172984 531257 173624 543656
rect 183424 531257 184064 543656
rect 184384 531257 185024 543656
rect 194824 531257 195464 543656
rect 195784 536508 196424 543656
rect 160624 473508 161264 480068
rect 161584 468801 162224 484231
rect 172024 468801 172664 484231
rect 172984 468801 173624 484231
rect 183424 468801 184064 484231
rect 184384 468801 185024 484231
rect 194824 468801 195464 484231
rect 195784 473508 196424 480068
rect 160624 410508 161264 417068
rect 161584 405801 162224 422591
rect 172024 405801 172664 422591
rect 172984 405801 173624 422591
rect 183424 405801 184064 422591
rect 184384 405801 185024 422591
rect 194824 405801 195464 422591
rect 195784 410508 196424 417068
rect 160624 347508 161264 354068
rect 161584 342801 162224 359591
rect 172024 342801 172664 359591
rect 172984 342801 173624 359591
rect 183424 342801 184064 359591
rect 184384 342801 185024 359591
rect 194824 342801 195464 359591
rect 195784 347508 196424 354068
rect 160624 284508 161264 291068
rect 161584 279801 162224 296591
rect 172024 279801 172664 296591
rect 172984 279801 173624 296591
rect 183424 279801 184064 296591
rect 184384 279801 185024 296591
rect 194824 279801 195464 296591
rect 195784 284508 196424 291068
rect 160624 221508 161264 228068
rect 161584 216801 162224 233591
rect 172024 216801 172664 233591
rect 172984 216801 173624 233591
rect 183424 216801 184064 233591
rect 184384 216801 185024 233591
rect 194824 216801 195464 233591
rect 195784 221508 196424 228068
rect 160624 158508 161264 165068
rect 161584 153801 162224 170591
rect 172024 153801 172664 170591
rect 172984 153801 173624 170591
rect 183424 153801 184064 170591
rect 184384 153801 185024 170591
rect 194824 153801 195464 170591
rect 195784 158508 196424 165068
rect 160624 95508 161264 102068
rect 161584 90801 162224 107591
rect 172024 90801 172664 107591
rect 172984 90801 173624 107591
rect 183424 90801 184064 107591
rect 184384 90801 185024 107591
rect 194824 90801 195464 107591
rect 195784 95508 196424 102068
rect 160624 32588 161264 39068
rect 160624 -744 161264 6068
rect 161584 -744 162224 44591
rect 172024 33049 172664 44591
rect 172984 33049 173624 44591
rect 183424 33049 184064 44591
rect 184384 33049 185024 44591
rect 172024 -744 172664 13495
rect 172984 -744 173624 13495
rect 183424 -744 184064 13495
rect 184384 -744 185024 13495
rect 194824 -744 195464 44591
rect 195784 32588 196424 39068
rect 195784 -744 196424 6068
rect 206224 -744 206864 543656
rect 207184 -744 207824 543656
rect 217624 536508 218264 543656
rect 218584 531257 219224 543656
rect 229024 531257 229664 543656
rect 229984 531257 230624 543656
rect 240424 531257 241064 543656
rect 241384 531257 242024 543656
rect 251824 531257 252464 543656
rect 252784 536508 253424 543656
rect 217624 473508 218264 480068
rect 218584 468801 219224 484231
rect 229024 468801 229664 484231
rect 229984 468801 230624 484231
rect 240424 468801 241064 484231
rect 241384 468801 242024 484231
rect 251824 468801 252464 484231
rect 252784 473508 253424 480068
rect 217624 410508 218264 417068
rect 218584 405801 219224 422591
rect 229024 405801 229664 422591
rect 229984 405801 230624 422591
rect 240424 405801 241064 422591
rect 241384 405801 242024 422591
rect 251824 405801 252464 422591
rect 252784 410508 253424 417068
rect 217624 347508 218264 354068
rect 218584 342801 219224 359591
rect 229024 342801 229664 359591
rect 229984 342801 230624 359591
rect 240424 342801 241064 359591
rect 241384 342801 242024 359591
rect 251824 342801 252464 359591
rect 252784 347508 253424 354068
rect 217624 284508 218264 291068
rect 218584 279801 219224 296591
rect 229024 279801 229664 296591
rect 229984 279801 230624 296591
rect 240424 279801 241064 296591
rect 241384 279801 242024 296591
rect 251824 279801 252464 296591
rect 252784 284508 253424 291068
rect 217624 221508 218264 228068
rect 218584 216801 219224 233591
rect 229024 216801 229664 233591
rect 229984 216801 230624 233591
rect 240424 216801 241064 233591
rect 241384 216801 242024 233591
rect 251824 216801 252464 233591
rect 252784 221508 253424 228068
rect 217624 158508 218264 165068
rect 218584 153801 219224 170591
rect 229024 153801 229664 170591
rect 229984 153801 230624 170591
rect 240424 153801 241064 170591
rect 241384 153801 242024 170591
rect 251824 153801 252464 170591
rect 252784 158508 253424 165068
rect 217624 95508 218264 102068
rect 218584 90801 219224 107591
rect 229024 90801 229664 107591
rect 229984 90801 230624 107591
rect 240424 90801 241064 107591
rect 241384 90801 242024 107591
rect 251824 90801 252464 107591
rect 252784 95508 253424 102068
rect 217624 32588 218264 39068
rect 217624 -744 218264 6068
rect 218584 -744 219224 44591
rect 229024 33049 229664 44591
rect 229984 33049 230624 44591
rect 240424 33049 241064 44591
rect 241384 33049 242024 44591
rect 229024 -744 229664 13495
rect 229984 -744 230624 13495
rect 240424 -744 241064 13495
rect 241384 -744 242024 13495
rect 251824 -744 252464 44591
rect 252784 32588 253424 39068
rect 252784 -744 253424 6068
rect 263224 -744 263864 543656
rect 264184 -744 264824 543656
rect 274624 536508 275264 543656
rect 275584 531257 276224 543656
rect 286024 531257 286664 543656
rect 286984 531257 287624 543656
rect 297424 531257 298064 543656
rect 298384 531257 299024 543656
rect 308824 531257 309464 543656
rect 309784 536508 310424 543656
rect 274624 473508 275264 480068
rect 275584 468801 276224 484231
rect 286024 468801 286664 484231
rect 286984 468801 287624 484231
rect 297424 468801 298064 484231
rect 298384 468801 299024 484231
rect 308824 468801 309464 484231
rect 309784 473508 310424 480068
rect 274624 410508 275264 417068
rect 275584 405801 276224 422591
rect 286024 405801 286664 422591
rect 286984 405801 287624 422591
rect 297424 405801 298064 422591
rect 298384 405801 299024 422591
rect 308824 405801 309464 422591
rect 309784 410508 310424 417068
rect 274624 347508 275264 354068
rect 275584 342801 276224 359591
rect 286024 342801 286664 359591
rect 286984 342801 287624 359591
rect 297424 342801 298064 359591
rect 298384 342801 299024 359591
rect 308824 342801 309464 359591
rect 309784 347508 310424 354068
rect 274624 284508 275264 291068
rect 275584 279801 276224 296591
rect 286024 279801 286664 296591
rect 286984 279801 287624 296591
rect 297424 279801 298064 296591
rect 298384 279801 299024 296591
rect 308824 279801 309464 296591
rect 309784 284508 310424 291068
rect 274624 221508 275264 228068
rect 275584 216801 276224 233591
rect 286024 216801 286664 233591
rect 286984 216801 287624 233591
rect 297424 216801 298064 233591
rect 298384 216801 299024 233591
rect 308824 216801 309464 233591
rect 309784 221508 310424 228068
rect 274624 158508 275264 165068
rect 275584 153801 276224 170591
rect 286024 153801 286664 170591
rect 286984 153801 287624 170591
rect 297424 153801 298064 170591
rect 298384 153801 299024 170591
rect 308824 153801 309464 170591
rect 309784 158508 310424 165068
rect 274624 95508 275264 102068
rect 275584 90801 276224 107591
rect 286024 90801 286664 107591
rect 286984 90801 287624 107591
rect 297424 90801 298064 107591
rect 298384 90801 299024 107591
rect 308824 90801 309464 107591
rect 309784 95508 310424 102068
rect 274624 32588 275264 39068
rect 274624 -744 275264 6068
rect 275584 -744 276224 44591
rect 286024 33049 286664 44591
rect 286984 33049 287624 44591
rect 297424 33049 298064 44591
rect 298384 33049 299024 44591
rect 286024 -744 286664 13495
rect 286984 -744 287624 13495
rect 297424 -744 298064 13495
rect 298384 -744 299024 13495
rect 308824 -744 309464 44591
rect 309784 32588 310424 39068
rect 309784 -744 310424 6068
rect 320224 -744 320864 543656
rect 321184 -744 321824 543656
rect 331624 536508 332264 543656
rect 332584 531257 333224 543656
rect 343024 531257 343664 543656
rect 343984 531257 344624 543656
rect 354424 531257 355064 543656
rect 355384 531257 356024 543656
rect 365824 531257 366464 543656
rect 366784 536508 367424 543656
rect 331624 473508 332264 480068
rect 332584 468801 333224 484231
rect 343024 468801 343664 484231
rect 343984 468801 344624 484231
rect 354424 468801 355064 484231
rect 355384 468801 356024 484231
rect 365824 468801 366464 484231
rect 366784 473508 367424 480068
rect 331624 410508 332264 417068
rect 332584 405801 333224 422591
rect 343024 405801 343664 422591
rect 343984 405801 344624 422591
rect 354424 405801 355064 422591
rect 355384 405801 356024 422591
rect 365824 405801 366464 422591
rect 366784 410508 367424 417068
rect 331624 347508 332264 354068
rect 332584 342801 333224 359591
rect 343024 342801 343664 359591
rect 343984 342801 344624 359591
rect 354424 342801 355064 359591
rect 355384 342801 356024 359591
rect 365824 342801 366464 359591
rect 366784 347508 367424 354068
rect 331624 284508 332264 291068
rect 332584 279801 333224 296591
rect 343024 279801 343664 296591
rect 343984 279801 344624 296591
rect 354424 279801 355064 296591
rect 355384 279801 356024 296591
rect 365824 279801 366464 296591
rect 366784 284508 367424 291068
rect 331624 221508 332264 228068
rect 332584 216801 333224 233591
rect 343024 216801 343664 233591
rect 343984 216801 344624 233591
rect 354424 216801 355064 233591
rect 355384 216801 356024 233591
rect 365824 216801 366464 233591
rect 366784 221508 367424 228068
rect 331624 158508 332264 165068
rect 332584 153801 333224 170591
rect 343024 153801 343664 170591
rect 343984 153801 344624 170591
rect 354424 153801 355064 170591
rect 355384 153801 356024 170591
rect 365824 153801 366464 170591
rect 366784 158508 367424 165068
rect 331624 95508 332264 102068
rect 332584 90801 333224 107591
rect 343024 90801 343664 107591
rect 343984 90801 344624 107591
rect 354424 90801 355064 107591
rect 355384 90801 356024 107591
rect 365824 90801 366464 107591
rect 366784 95508 367424 102068
rect 331624 32588 332264 39068
rect 331624 -744 332264 6068
rect 332584 -744 333224 44591
rect 343024 33049 343664 44591
rect 343984 33049 344624 44591
rect 354424 33049 355064 44591
rect 355384 33049 356024 44591
rect 343024 -744 343664 13495
rect 343984 -744 344624 13495
rect 354424 -744 355064 13495
rect 355384 -744 356024 13495
rect 365824 -744 366464 44591
rect 366784 32588 367424 39068
rect 366784 -744 367424 6068
rect 377224 -744 377864 543656
rect 378184 -744 378824 543656
rect 388624 536508 389264 543656
rect 389584 531257 390224 543656
rect 400024 531257 400664 543656
rect 400984 531257 401624 543656
rect 411424 531257 412064 543656
rect 412384 531257 413024 543656
rect 422824 531257 423464 543656
rect 423784 536508 424424 543656
rect 388624 473508 389264 480068
rect 389584 468801 390224 484231
rect 400024 468801 400664 484231
rect 400984 468801 401624 484231
rect 411424 468801 412064 484231
rect 412384 468801 413024 484231
rect 422824 468801 423464 484231
rect 423784 473508 424424 480068
rect 388624 410508 389264 417068
rect 389584 405801 390224 422591
rect 400024 405801 400664 422591
rect 400984 405801 401624 422591
rect 411424 405801 412064 422591
rect 412384 405801 413024 422591
rect 422824 405801 423464 422591
rect 423784 410508 424424 417068
rect 388624 347508 389264 354068
rect 389584 342801 390224 359591
rect 400024 342801 400664 359591
rect 400984 342801 401624 359591
rect 411424 342801 412064 359591
rect 412384 342801 413024 359591
rect 422824 342801 423464 359591
rect 423784 347508 424424 354068
rect 388624 284508 389264 291068
rect 389584 279801 390224 296591
rect 400024 279801 400664 296591
rect 400984 279801 401624 296591
rect 411424 279801 412064 296591
rect 412384 279801 413024 296591
rect 422824 279801 423464 296591
rect 423784 284508 424424 291068
rect 388624 221508 389264 228068
rect 389584 216801 390224 233591
rect 400024 216801 400664 233591
rect 400984 216801 401624 233591
rect 411424 216801 412064 233591
rect 412384 216801 413024 233591
rect 422824 216801 423464 233591
rect 423784 221508 424424 228068
rect 388624 158508 389264 165068
rect 389584 153801 390224 170591
rect 400024 153801 400664 170591
rect 400984 153801 401624 170591
rect 411424 153801 412064 170591
rect 412384 153801 413024 170591
rect 422824 153801 423464 170591
rect 423784 158508 424424 165068
rect 388624 95508 389264 102068
rect 389584 90801 390224 107591
rect 400024 90801 400664 107591
rect 400984 90801 401624 107591
rect 411424 90801 412064 107591
rect 412384 90801 413024 107591
rect 422824 90801 423464 107591
rect 423784 95508 424424 102068
rect 388624 32588 389264 39068
rect 388624 -744 389264 6068
rect 389584 -744 390224 44591
rect 400024 33049 400664 44591
rect 400984 33049 401624 44591
rect 411424 33049 412064 44591
rect 412384 33049 413024 44591
rect 400024 -744 400664 13495
rect 400984 -744 401624 13495
rect 411424 -744 412064 13495
rect 412384 -744 413024 13495
rect 422824 -744 423464 44591
rect 423784 32588 424424 39068
rect 423784 -744 424424 6068
rect 434224 -744 434864 543656
rect 435184 -744 435824 543656
rect 445624 536508 446264 543656
rect 446584 536017 447224 543656
rect 457024 536017 457664 543656
rect 457984 536017 458624 543656
rect 468424 536017 469064 543656
rect 469384 536017 470024 543656
rect 479824 536017 480464 543656
rect 480784 536508 481424 543656
rect 445624 473508 446264 480068
rect 446584 473017 447224 481375
rect 457024 473017 457664 481375
rect 457984 473017 458624 481375
rect 468424 473017 469064 481375
rect 469384 473017 470024 481375
rect 479824 473017 480464 481375
rect 480784 473508 481424 480068
rect 445624 410508 446264 417068
rect 446584 410017 447224 417287
rect 457024 410017 457664 417287
rect 457984 410017 458624 417287
rect 468424 410017 469064 417287
rect 469384 410017 470024 417287
rect 479824 410017 480464 417287
rect 480784 410508 481424 417068
rect 445624 347508 446264 354068
rect 446584 347017 447224 354287
rect 457024 347017 457664 354287
rect 457984 347017 458624 354287
rect 468424 347017 469064 354287
rect 469384 347017 470024 354287
rect 479824 347017 480464 354287
rect 480784 347508 481424 354068
rect 445624 284508 446264 291068
rect 446584 284017 447224 291287
rect 457024 284017 457664 291287
rect 457984 284017 458624 291287
rect 468424 284017 469064 291287
rect 469384 284017 470024 291287
rect 479824 284017 480464 291287
rect 480784 284508 481424 291068
rect 445624 221508 446264 228068
rect 446584 221017 447224 228287
rect 457024 221017 457664 228287
rect 457984 221017 458624 228287
rect 468424 221017 469064 228287
rect 469384 221017 470024 228287
rect 479824 221017 480464 228287
rect 480784 221508 481424 228068
rect 445624 158508 446264 165068
rect 446584 158017 447224 165287
rect 457024 158017 457664 165287
rect 457984 158017 458624 165287
rect 468424 158017 469064 165287
rect 469384 158017 470024 165287
rect 479824 158017 480464 165287
rect 480784 158508 481424 165068
rect 445624 95508 446264 102068
rect 446584 95017 447224 102287
rect 457024 95017 457664 102287
rect 457984 95017 458624 102287
rect 468424 95017 469064 102287
rect 469384 95017 470024 102287
rect 479824 95017 480464 102287
rect 480784 95508 481424 102068
rect 445624 32588 446264 39068
rect 446584 32233 447224 39287
rect 457024 32233 457664 39287
rect 457984 32233 458624 39287
rect 445624 -744 446264 6068
rect 446584 -744 447224 12135
rect 457024 -744 457664 12135
rect 457984 -744 458624 12135
rect 468424 -744 469064 39287
rect 469384 -744 470024 39287
rect 479824 -744 480464 39287
rect 480784 32588 481424 39068
rect 480784 -744 481424 6068
rect 491224 -744 491864 543656
rect 492184 -744 492824 543656
rect 495192 616 496152 542296
rect 496552 -744 497512 543656
<< obsm4 >>
rect 8944 34193 12344 534448
rect 13144 523697 24704 534448
rect 25504 523697 35144 534448
rect 13144 480503 35144 523697
rect 13144 480148 24704 480503
rect 13144 473428 13304 480148
rect 14104 473428 23744 480148
rect 24544 473428 24704 480148
rect 13144 472937 24704 473428
rect 25504 472937 35144 480503
rect 13144 417911 35144 472937
rect 13144 417148 24704 417911
rect 13144 410428 13304 417148
rect 14104 410428 23744 417148
rect 24544 410428 24704 417148
rect 13144 409937 24704 410428
rect 25504 409937 35144 417911
rect 13144 354911 35144 409937
rect 13144 354148 24704 354911
rect 13144 347428 13304 354148
rect 14104 347428 23744 354148
rect 24544 347428 24704 354148
rect 13144 346937 24704 347428
rect 25504 346937 35144 354911
rect 13144 291911 35144 346937
rect 13144 291148 24704 291911
rect 13144 284428 13304 291148
rect 14104 284428 23744 291148
rect 24544 284428 24704 291148
rect 13144 283937 24704 284428
rect 25504 283937 35144 291911
rect 13144 228911 35144 283937
rect 13144 228148 24704 228911
rect 13144 221428 13304 228148
rect 14104 221428 23744 228148
rect 24544 221428 24704 228148
rect 13144 220937 24704 221428
rect 25504 220937 35144 228911
rect 13144 165911 35144 220937
rect 13144 165148 24704 165911
rect 13144 158428 13304 165148
rect 14104 158428 23744 165148
rect 24544 158428 24704 165148
rect 13144 157937 24704 158428
rect 25504 157937 35144 165911
rect 13144 102911 35144 157937
rect 13144 102148 24704 102911
rect 13144 95428 13304 102148
rect 14104 95428 23744 102148
rect 24544 95428 24704 102148
rect 13144 94937 24704 95428
rect 25504 94937 35144 102911
rect 13144 39911 35144 94937
rect 13144 39148 24704 39911
rect 13144 34193 13304 39148
rect 14104 34193 23744 39148
rect 24544 34193 24704 39148
rect 25504 34193 35144 39911
rect 8944 13575 35144 34193
rect 8944 8128 12344 13575
rect 13144 8128 24704 13575
rect 25504 8128 35144 13575
rect 35944 8128 36104 534448
rect 36904 531177 47504 534448
rect 48304 531177 57944 534448
rect 58744 531177 58904 534448
rect 59704 531177 69344 534448
rect 70144 531177 70304 534448
rect 71104 531177 80744 534448
rect 81544 531177 92144 534448
rect 36904 484311 92144 531177
rect 36904 480148 47504 484311
rect 36904 473428 46544 480148
rect 47344 473428 47504 480148
rect 36904 468721 47504 473428
rect 48304 468721 57944 484311
rect 58744 468721 58904 484311
rect 59704 468721 69344 484311
rect 70144 468721 70304 484311
rect 71104 468721 80744 484311
rect 81544 480148 92144 484311
rect 81544 473428 81704 480148
rect 82504 473428 92144 480148
rect 81544 468721 92144 473428
rect 36904 422671 92144 468721
rect 36904 417148 47504 422671
rect 36904 410428 46544 417148
rect 47344 410428 47504 417148
rect 36904 405721 47504 410428
rect 48304 405721 57944 422671
rect 58744 405721 58904 422671
rect 59704 405721 69344 422671
rect 70144 405721 70304 422671
rect 71104 405721 80744 422671
rect 81544 417148 92144 422671
rect 81544 410428 81704 417148
rect 82504 410428 92144 417148
rect 81544 405721 92144 410428
rect 36904 359671 92144 405721
rect 36904 354148 47504 359671
rect 36904 347428 46544 354148
rect 47344 347428 47504 354148
rect 36904 342721 47504 347428
rect 48304 342721 57944 359671
rect 58744 342721 58904 359671
rect 59704 342721 69344 359671
rect 70144 342721 70304 359671
rect 71104 342721 80744 359671
rect 81544 354148 92144 359671
rect 81544 347428 81704 354148
rect 82504 347428 92144 354148
rect 81544 342721 92144 347428
rect 36904 296671 92144 342721
rect 36904 291148 47504 296671
rect 36904 284428 46544 291148
rect 47344 284428 47504 291148
rect 36904 279721 47504 284428
rect 48304 279721 57944 296671
rect 58744 279721 58904 296671
rect 59704 279721 69344 296671
rect 70144 279721 70304 296671
rect 71104 279721 80744 296671
rect 81544 291148 92144 296671
rect 81544 284428 81704 291148
rect 82504 284428 92144 291148
rect 81544 279721 92144 284428
rect 36904 233671 92144 279721
rect 36904 228148 47504 233671
rect 36904 221428 46544 228148
rect 47344 221428 47504 228148
rect 36904 216721 47504 221428
rect 48304 216721 57944 233671
rect 58744 216721 58904 233671
rect 59704 216721 69344 233671
rect 70144 216721 70304 233671
rect 71104 216721 80744 233671
rect 81544 228148 92144 233671
rect 81544 221428 81704 228148
rect 82504 221428 92144 228148
rect 81544 216721 92144 221428
rect 36904 170671 92144 216721
rect 36904 165148 47504 170671
rect 36904 158428 46544 165148
rect 47344 158428 47504 165148
rect 36904 153721 47504 158428
rect 48304 153721 57944 170671
rect 58744 153721 58904 170671
rect 59704 153721 69344 170671
rect 70144 153721 70304 170671
rect 71104 153721 80744 170671
rect 81544 165148 92144 170671
rect 81544 158428 81704 165148
rect 82504 158428 92144 165148
rect 81544 153721 92144 158428
rect 36904 107671 92144 153721
rect 36904 102148 47504 107671
rect 36904 95428 46544 102148
rect 47344 95428 47504 102148
rect 36904 90721 47504 95428
rect 48304 90721 57944 107671
rect 58744 90721 58904 107671
rect 59704 90721 69344 107671
rect 70144 90721 70304 107671
rect 71104 90721 80744 107671
rect 81544 102148 92144 107671
rect 81544 95428 81704 102148
rect 82504 95428 92144 102148
rect 81544 90721 92144 95428
rect 36904 44671 92144 90721
rect 36904 39148 47504 44671
rect 36904 32508 46544 39148
rect 47344 32508 47504 39148
rect 36904 8128 47504 32508
rect 48304 32969 57944 44671
rect 58744 32969 58904 44671
rect 59704 32969 69344 44671
rect 70144 32969 70304 44671
rect 71104 32969 80744 44671
rect 48304 13575 80744 32969
rect 48304 8128 57944 13575
rect 58744 8128 58904 13575
rect 59704 8128 69344 13575
rect 70144 8128 70304 13575
rect 71104 8128 80744 13575
rect 81544 39148 92144 44671
rect 81544 32508 81704 39148
rect 82504 32508 92144 39148
rect 81544 8128 92144 32508
rect 92944 8128 93104 534448
rect 93904 531177 104504 534448
rect 105304 531177 114944 534448
rect 115744 531177 115904 534448
rect 116704 531177 126344 534448
rect 127144 531177 127304 534448
rect 128104 531177 137744 534448
rect 138544 531177 149144 534448
rect 93904 484311 149144 531177
rect 93904 480148 104504 484311
rect 93904 473428 103544 480148
rect 104344 473428 104504 480148
rect 93904 468721 104504 473428
rect 105304 468721 114944 484311
rect 115744 468721 115904 484311
rect 116704 468721 126344 484311
rect 127144 468721 127304 484311
rect 128104 468721 137744 484311
rect 138544 480148 149144 484311
rect 138544 473428 138704 480148
rect 139504 473428 149144 480148
rect 138544 468721 149144 473428
rect 93904 422671 149144 468721
rect 93904 417148 104504 422671
rect 93904 410428 103544 417148
rect 104344 410428 104504 417148
rect 93904 405721 104504 410428
rect 105304 405721 114944 422671
rect 115744 405721 115904 422671
rect 116704 405721 126344 422671
rect 127144 405721 127304 422671
rect 128104 405721 137744 422671
rect 138544 417148 149144 422671
rect 138544 410428 138704 417148
rect 139504 410428 149144 417148
rect 138544 405721 149144 410428
rect 93904 359671 149144 405721
rect 93904 354148 104504 359671
rect 93904 347428 103544 354148
rect 104344 347428 104504 354148
rect 93904 342721 104504 347428
rect 105304 342721 114944 359671
rect 115744 342721 115904 359671
rect 116704 342721 126344 359671
rect 127144 342721 127304 359671
rect 128104 342721 137744 359671
rect 138544 354148 149144 359671
rect 138544 347428 138704 354148
rect 139504 347428 149144 354148
rect 138544 342721 149144 347428
rect 93904 296671 149144 342721
rect 93904 291148 104504 296671
rect 93904 284428 103544 291148
rect 104344 284428 104504 291148
rect 93904 279721 104504 284428
rect 105304 279721 114944 296671
rect 115744 279721 115904 296671
rect 116704 279721 126344 296671
rect 127144 279721 127304 296671
rect 128104 279721 137744 296671
rect 138544 291148 149144 296671
rect 138544 284428 138704 291148
rect 139504 284428 149144 291148
rect 138544 279721 149144 284428
rect 93904 233671 149144 279721
rect 93904 228148 104504 233671
rect 93904 221428 103544 228148
rect 104344 221428 104504 228148
rect 93904 216721 104504 221428
rect 105304 216721 114944 233671
rect 115744 216721 115904 233671
rect 116704 216721 126344 233671
rect 127144 216721 127304 233671
rect 128104 216721 137744 233671
rect 138544 228148 149144 233671
rect 138544 221428 138704 228148
rect 139504 221428 149144 228148
rect 138544 216721 149144 221428
rect 93904 170671 149144 216721
rect 93904 165148 104504 170671
rect 93904 158428 103544 165148
rect 104344 158428 104504 165148
rect 93904 153721 104504 158428
rect 105304 153721 114944 170671
rect 115744 153721 115904 170671
rect 116704 153721 126344 170671
rect 127144 153721 127304 170671
rect 128104 153721 137744 170671
rect 138544 165148 149144 170671
rect 138544 158428 138704 165148
rect 139504 158428 149144 165148
rect 138544 153721 149144 158428
rect 93904 107671 149144 153721
rect 93904 102148 104504 107671
rect 93904 95428 103544 102148
rect 104344 95428 104504 102148
rect 93904 90721 104504 95428
rect 105304 90721 114944 107671
rect 115744 90721 115904 107671
rect 116704 90721 126344 107671
rect 127144 90721 127304 107671
rect 128104 90721 137744 107671
rect 138544 102148 149144 107671
rect 138544 95428 138704 102148
rect 139504 95428 149144 102148
rect 138544 90721 149144 95428
rect 93904 44671 149144 90721
rect 93904 39148 104504 44671
rect 93904 32508 103544 39148
rect 104344 32508 104504 39148
rect 93904 8128 104504 32508
rect 105304 32969 114944 44671
rect 115744 32969 115904 44671
rect 116704 32969 126344 44671
rect 127144 32969 127304 44671
rect 128104 32969 137744 44671
rect 105304 13575 137744 32969
rect 105304 8128 114944 13575
rect 115744 8128 115904 13575
rect 116704 8128 126344 13575
rect 127144 8128 127304 13575
rect 128104 8128 137744 13575
rect 138544 39148 149144 44671
rect 138544 32508 138704 39148
rect 139504 32508 149144 39148
rect 138544 8128 149144 32508
rect 149944 8128 150104 534448
rect 150904 531177 161504 534448
rect 162304 531177 171944 534448
rect 172744 531177 172904 534448
rect 173704 531177 183344 534448
rect 184144 531177 184304 534448
rect 185104 531177 194744 534448
rect 195544 531177 206144 534448
rect 150904 484311 206144 531177
rect 150904 480148 161504 484311
rect 150904 473428 160544 480148
rect 161344 473428 161504 480148
rect 150904 468721 161504 473428
rect 162304 468721 171944 484311
rect 172744 468721 172904 484311
rect 173704 468721 183344 484311
rect 184144 468721 184304 484311
rect 185104 468721 194744 484311
rect 195544 480148 206144 484311
rect 195544 473428 195704 480148
rect 196504 473428 206144 480148
rect 195544 468721 206144 473428
rect 150904 422671 206144 468721
rect 150904 417148 161504 422671
rect 150904 410428 160544 417148
rect 161344 410428 161504 417148
rect 150904 405721 161504 410428
rect 162304 405721 171944 422671
rect 172744 405721 172904 422671
rect 173704 405721 183344 422671
rect 184144 405721 184304 422671
rect 185104 405721 194744 422671
rect 195544 417148 206144 422671
rect 195544 410428 195704 417148
rect 196504 410428 206144 417148
rect 195544 405721 206144 410428
rect 150904 359671 206144 405721
rect 150904 354148 161504 359671
rect 150904 347428 160544 354148
rect 161344 347428 161504 354148
rect 150904 342721 161504 347428
rect 162304 342721 171944 359671
rect 172744 342721 172904 359671
rect 173704 342721 183344 359671
rect 184144 342721 184304 359671
rect 185104 342721 194744 359671
rect 195544 354148 206144 359671
rect 195544 347428 195704 354148
rect 196504 347428 206144 354148
rect 195544 342721 206144 347428
rect 150904 296671 206144 342721
rect 150904 291148 161504 296671
rect 150904 284428 160544 291148
rect 161344 284428 161504 291148
rect 150904 279721 161504 284428
rect 162304 279721 171944 296671
rect 172744 279721 172904 296671
rect 173704 279721 183344 296671
rect 184144 279721 184304 296671
rect 185104 279721 194744 296671
rect 195544 291148 206144 296671
rect 195544 284428 195704 291148
rect 196504 284428 206144 291148
rect 195544 279721 206144 284428
rect 150904 233671 206144 279721
rect 150904 228148 161504 233671
rect 150904 221428 160544 228148
rect 161344 221428 161504 228148
rect 150904 216721 161504 221428
rect 162304 216721 171944 233671
rect 172744 216721 172904 233671
rect 173704 216721 183344 233671
rect 184144 216721 184304 233671
rect 185104 216721 194744 233671
rect 195544 228148 206144 233671
rect 195544 221428 195704 228148
rect 196504 221428 206144 228148
rect 195544 216721 206144 221428
rect 150904 170671 206144 216721
rect 150904 165148 161504 170671
rect 150904 158428 160544 165148
rect 161344 158428 161504 165148
rect 150904 153721 161504 158428
rect 162304 153721 171944 170671
rect 172744 153721 172904 170671
rect 173704 153721 183344 170671
rect 184144 153721 184304 170671
rect 185104 153721 194744 170671
rect 195544 165148 206144 170671
rect 195544 158428 195704 165148
rect 196504 158428 206144 165148
rect 195544 153721 206144 158428
rect 150904 107671 206144 153721
rect 150904 102148 161504 107671
rect 150904 95428 160544 102148
rect 161344 95428 161504 102148
rect 150904 90721 161504 95428
rect 162304 90721 171944 107671
rect 172744 90721 172904 107671
rect 173704 90721 183344 107671
rect 184144 90721 184304 107671
rect 185104 90721 194744 107671
rect 195544 102148 206144 107671
rect 195544 95428 195704 102148
rect 196504 95428 206144 102148
rect 195544 90721 206144 95428
rect 150904 44671 206144 90721
rect 150904 39148 161504 44671
rect 150904 32508 160544 39148
rect 161344 32508 161504 39148
rect 150904 8128 161504 32508
rect 162304 32969 171944 44671
rect 172744 32969 172904 44671
rect 173704 32969 183344 44671
rect 184144 32969 184304 44671
rect 185104 32969 194744 44671
rect 162304 13575 194744 32969
rect 162304 8128 171944 13575
rect 172744 8128 172904 13575
rect 173704 8128 183344 13575
rect 184144 8128 184304 13575
rect 185104 8128 194744 13575
rect 195544 39148 206144 44671
rect 195544 32508 195704 39148
rect 196504 32508 206144 39148
rect 195544 8128 206144 32508
rect 206944 8128 207104 534448
rect 207904 531177 218504 534448
rect 219304 531177 228944 534448
rect 229744 531177 229904 534448
rect 230704 531177 240344 534448
rect 241144 531177 241304 534448
rect 242104 531177 251744 534448
rect 252544 531177 263144 534448
rect 207904 484311 263144 531177
rect 207904 480148 218504 484311
rect 207904 473428 217544 480148
rect 218344 473428 218504 480148
rect 207904 468721 218504 473428
rect 219304 468721 228944 484311
rect 229744 468721 229904 484311
rect 230704 468721 240344 484311
rect 241144 468721 241304 484311
rect 242104 468721 251744 484311
rect 252544 480148 263144 484311
rect 252544 473428 252704 480148
rect 253504 473428 263144 480148
rect 252544 468721 263144 473428
rect 207904 422671 263144 468721
rect 207904 417148 218504 422671
rect 207904 410428 217544 417148
rect 218344 410428 218504 417148
rect 207904 405721 218504 410428
rect 219304 405721 228944 422671
rect 229744 405721 229904 422671
rect 230704 405721 240344 422671
rect 241144 405721 241304 422671
rect 242104 405721 251744 422671
rect 252544 417148 263144 422671
rect 252544 410428 252704 417148
rect 253504 410428 263144 417148
rect 252544 405721 263144 410428
rect 207904 359671 263144 405721
rect 207904 354148 218504 359671
rect 207904 347428 217544 354148
rect 218344 347428 218504 354148
rect 207904 342721 218504 347428
rect 219304 342721 228944 359671
rect 229744 342721 229904 359671
rect 230704 342721 240344 359671
rect 241144 342721 241304 359671
rect 242104 342721 251744 359671
rect 252544 354148 263144 359671
rect 252544 347428 252704 354148
rect 253504 347428 263144 354148
rect 252544 342721 263144 347428
rect 207904 296671 263144 342721
rect 207904 291148 218504 296671
rect 207904 284428 217544 291148
rect 218344 284428 218504 291148
rect 207904 279721 218504 284428
rect 219304 279721 228944 296671
rect 229744 279721 229904 296671
rect 230704 279721 240344 296671
rect 241144 279721 241304 296671
rect 242104 279721 251744 296671
rect 252544 291148 263144 296671
rect 252544 284428 252704 291148
rect 253504 284428 263144 291148
rect 252544 279721 263144 284428
rect 207904 233671 263144 279721
rect 207904 228148 218504 233671
rect 207904 221428 217544 228148
rect 218344 221428 218504 228148
rect 207904 216721 218504 221428
rect 219304 216721 228944 233671
rect 229744 216721 229904 233671
rect 230704 216721 240344 233671
rect 241144 216721 241304 233671
rect 242104 216721 251744 233671
rect 252544 228148 263144 233671
rect 252544 221428 252704 228148
rect 253504 221428 263144 228148
rect 252544 216721 263144 221428
rect 207904 170671 263144 216721
rect 207904 165148 218504 170671
rect 207904 158428 217544 165148
rect 218344 158428 218504 165148
rect 207904 153721 218504 158428
rect 219304 153721 228944 170671
rect 229744 153721 229904 170671
rect 230704 153721 240344 170671
rect 241144 153721 241304 170671
rect 242104 153721 251744 170671
rect 252544 165148 263144 170671
rect 252544 158428 252704 165148
rect 253504 158428 263144 165148
rect 252544 153721 263144 158428
rect 207904 107671 263144 153721
rect 207904 102148 218504 107671
rect 207904 95428 217544 102148
rect 218344 95428 218504 102148
rect 207904 90721 218504 95428
rect 219304 90721 228944 107671
rect 229744 90721 229904 107671
rect 230704 90721 240344 107671
rect 241144 90721 241304 107671
rect 242104 90721 251744 107671
rect 252544 102148 263144 107671
rect 252544 95428 252704 102148
rect 253504 95428 263144 102148
rect 252544 90721 263144 95428
rect 207904 44671 263144 90721
rect 207904 39148 218504 44671
rect 207904 32508 217544 39148
rect 218344 32508 218504 39148
rect 207904 8128 218504 32508
rect 219304 32969 228944 44671
rect 229744 32969 229904 44671
rect 230704 32969 240344 44671
rect 241144 32969 241304 44671
rect 242104 32969 251744 44671
rect 219304 13575 251744 32969
rect 219304 8128 228944 13575
rect 229744 8128 229904 13575
rect 230704 8128 240344 13575
rect 241144 8128 241304 13575
rect 242104 8128 251744 13575
rect 252544 39148 263144 44671
rect 252544 32508 252704 39148
rect 253504 32508 263144 39148
rect 252544 8128 263144 32508
rect 263944 8128 264104 534448
rect 264904 531177 275504 534448
rect 276304 531177 285944 534448
rect 286744 531177 286904 534448
rect 287704 531177 297344 534448
rect 298144 531177 298304 534448
rect 299104 531177 308744 534448
rect 309544 531177 320144 534448
rect 264904 484311 320144 531177
rect 264904 480148 275504 484311
rect 264904 473428 274544 480148
rect 275344 473428 275504 480148
rect 264904 468721 275504 473428
rect 276304 468721 285944 484311
rect 286744 468721 286904 484311
rect 287704 468721 297344 484311
rect 298144 468721 298304 484311
rect 299104 468721 308744 484311
rect 309544 480148 320144 484311
rect 309544 473428 309704 480148
rect 310504 473428 320144 480148
rect 309544 468721 320144 473428
rect 264904 422671 320144 468721
rect 264904 417148 275504 422671
rect 264904 410428 274544 417148
rect 275344 410428 275504 417148
rect 264904 405721 275504 410428
rect 276304 405721 285944 422671
rect 286744 405721 286904 422671
rect 287704 405721 297344 422671
rect 298144 405721 298304 422671
rect 299104 405721 308744 422671
rect 309544 417148 320144 422671
rect 309544 410428 309704 417148
rect 310504 410428 320144 417148
rect 309544 405721 320144 410428
rect 264904 359671 320144 405721
rect 264904 354148 275504 359671
rect 264904 347428 274544 354148
rect 275344 347428 275504 354148
rect 264904 342721 275504 347428
rect 276304 342721 285944 359671
rect 286744 342721 286904 359671
rect 287704 342721 297344 359671
rect 298144 342721 298304 359671
rect 299104 342721 308744 359671
rect 309544 354148 320144 359671
rect 309544 347428 309704 354148
rect 310504 347428 320144 354148
rect 309544 342721 320144 347428
rect 264904 296671 320144 342721
rect 264904 291148 275504 296671
rect 264904 284428 274544 291148
rect 275344 284428 275504 291148
rect 264904 279721 275504 284428
rect 276304 279721 285944 296671
rect 286744 279721 286904 296671
rect 287704 279721 297344 296671
rect 298144 279721 298304 296671
rect 299104 279721 308744 296671
rect 309544 291148 320144 296671
rect 309544 284428 309704 291148
rect 310504 284428 320144 291148
rect 309544 279721 320144 284428
rect 264904 233671 320144 279721
rect 264904 228148 275504 233671
rect 264904 221428 274544 228148
rect 275344 221428 275504 228148
rect 264904 216721 275504 221428
rect 276304 216721 285944 233671
rect 286744 216721 286904 233671
rect 287704 216721 297344 233671
rect 298144 216721 298304 233671
rect 299104 216721 308744 233671
rect 309544 228148 320144 233671
rect 309544 221428 309704 228148
rect 310504 221428 320144 228148
rect 309544 216721 320144 221428
rect 264904 170671 320144 216721
rect 264904 165148 275504 170671
rect 264904 158428 274544 165148
rect 275344 158428 275504 165148
rect 264904 153721 275504 158428
rect 276304 153721 285944 170671
rect 286744 153721 286904 170671
rect 287704 153721 297344 170671
rect 298144 153721 298304 170671
rect 299104 153721 308744 170671
rect 309544 165148 320144 170671
rect 309544 158428 309704 165148
rect 310504 158428 320144 165148
rect 309544 153721 320144 158428
rect 264904 107671 320144 153721
rect 264904 102148 275504 107671
rect 264904 95428 274544 102148
rect 275344 95428 275504 102148
rect 264904 90721 275504 95428
rect 276304 90721 285944 107671
rect 286744 90721 286904 107671
rect 287704 90721 297344 107671
rect 298144 90721 298304 107671
rect 299104 90721 308744 107671
rect 309544 102148 320144 107671
rect 309544 95428 309704 102148
rect 310504 95428 320144 102148
rect 309544 90721 320144 95428
rect 264904 44671 320144 90721
rect 264904 39148 275504 44671
rect 264904 32508 274544 39148
rect 275344 32508 275504 39148
rect 264904 8128 275504 32508
rect 276304 32969 285944 44671
rect 286744 32969 286904 44671
rect 287704 32969 297344 44671
rect 298144 32969 298304 44671
rect 299104 32969 308744 44671
rect 276304 13575 308744 32969
rect 276304 8128 285944 13575
rect 286744 8128 286904 13575
rect 287704 8128 297344 13575
rect 298144 8128 298304 13575
rect 299104 8128 308744 13575
rect 309544 39148 320144 44671
rect 309544 32508 309704 39148
rect 310504 32508 320144 39148
rect 309544 8128 320144 32508
rect 320944 8128 321104 534448
rect 321904 531177 332504 534448
rect 333304 531177 342944 534448
rect 343744 531177 343904 534448
rect 344704 531177 354344 534448
rect 355144 531177 355304 534448
rect 356104 531177 365744 534448
rect 366544 531177 377144 534448
rect 321904 484311 377144 531177
rect 321904 480148 332504 484311
rect 321904 473428 331544 480148
rect 332344 473428 332504 480148
rect 321904 468721 332504 473428
rect 333304 468721 342944 484311
rect 343744 468721 343904 484311
rect 344704 468721 354344 484311
rect 355144 468721 355304 484311
rect 356104 468721 365744 484311
rect 366544 480148 377144 484311
rect 366544 473428 366704 480148
rect 367504 473428 377144 480148
rect 366544 468721 377144 473428
rect 321904 422671 377144 468721
rect 321904 417148 332504 422671
rect 321904 410428 331544 417148
rect 332344 410428 332504 417148
rect 321904 405721 332504 410428
rect 333304 405721 342944 422671
rect 343744 405721 343904 422671
rect 344704 405721 354344 422671
rect 355144 405721 355304 422671
rect 356104 405721 365744 422671
rect 366544 417148 377144 422671
rect 366544 410428 366704 417148
rect 367504 410428 377144 417148
rect 366544 405721 377144 410428
rect 321904 359671 377144 405721
rect 321904 354148 332504 359671
rect 321904 347428 331544 354148
rect 332344 347428 332504 354148
rect 321904 342721 332504 347428
rect 333304 342721 342944 359671
rect 343744 342721 343904 359671
rect 344704 342721 354344 359671
rect 355144 342721 355304 359671
rect 356104 342721 365744 359671
rect 366544 354148 377144 359671
rect 366544 347428 366704 354148
rect 367504 347428 377144 354148
rect 366544 342721 377144 347428
rect 321904 296671 377144 342721
rect 321904 291148 332504 296671
rect 321904 284428 331544 291148
rect 332344 284428 332504 291148
rect 321904 279721 332504 284428
rect 333304 279721 342944 296671
rect 343744 279721 343904 296671
rect 344704 279721 354344 296671
rect 355144 279721 355304 296671
rect 356104 279721 365744 296671
rect 366544 291148 377144 296671
rect 366544 284428 366704 291148
rect 367504 284428 377144 291148
rect 366544 279721 377144 284428
rect 321904 233671 377144 279721
rect 321904 228148 332504 233671
rect 321904 221428 331544 228148
rect 332344 221428 332504 228148
rect 321904 216721 332504 221428
rect 333304 216721 342944 233671
rect 343744 216721 343904 233671
rect 344704 216721 354344 233671
rect 355144 216721 355304 233671
rect 356104 216721 365744 233671
rect 366544 228148 377144 233671
rect 366544 221428 366704 228148
rect 367504 221428 377144 228148
rect 366544 216721 377144 221428
rect 321904 170671 377144 216721
rect 321904 165148 332504 170671
rect 321904 158428 331544 165148
rect 332344 158428 332504 165148
rect 321904 153721 332504 158428
rect 333304 153721 342944 170671
rect 343744 153721 343904 170671
rect 344704 153721 354344 170671
rect 355144 153721 355304 170671
rect 356104 153721 365744 170671
rect 366544 165148 377144 170671
rect 366544 158428 366704 165148
rect 367504 158428 377144 165148
rect 366544 153721 377144 158428
rect 321904 107671 377144 153721
rect 321904 102148 332504 107671
rect 321904 95428 331544 102148
rect 332344 95428 332504 102148
rect 321904 90721 332504 95428
rect 333304 90721 342944 107671
rect 343744 90721 343904 107671
rect 344704 90721 354344 107671
rect 355144 90721 355304 107671
rect 356104 90721 365744 107671
rect 366544 102148 377144 107671
rect 366544 95428 366704 102148
rect 367504 95428 377144 102148
rect 366544 90721 377144 95428
rect 321904 44671 377144 90721
rect 321904 39148 332504 44671
rect 321904 32508 331544 39148
rect 332344 32508 332504 39148
rect 321904 8128 332504 32508
rect 333304 32969 342944 44671
rect 343744 32969 343904 44671
rect 344704 32969 354344 44671
rect 355144 32969 355304 44671
rect 356104 32969 365744 44671
rect 333304 13575 365744 32969
rect 333304 8128 342944 13575
rect 343744 8128 343904 13575
rect 344704 8128 354344 13575
rect 355144 8128 355304 13575
rect 356104 8128 365744 13575
rect 366544 39148 377144 44671
rect 366544 32508 366704 39148
rect 367504 32508 377144 39148
rect 366544 8128 377144 32508
rect 377944 8128 378104 534448
rect 378904 531177 389504 534448
rect 390304 531177 399944 534448
rect 400744 531177 400904 534448
rect 401704 531177 411344 534448
rect 412144 531177 412304 534448
rect 413104 531177 422744 534448
rect 423544 531177 434144 534448
rect 378904 484311 434144 531177
rect 378904 480148 389504 484311
rect 378904 473428 388544 480148
rect 389344 473428 389504 480148
rect 378904 468721 389504 473428
rect 390304 468721 399944 484311
rect 400744 468721 400904 484311
rect 401704 468721 411344 484311
rect 412144 468721 412304 484311
rect 413104 468721 422744 484311
rect 423544 480148 434144 484311
rect 423544 473428 423704 480148
rect 424504 473428 434144 480148
rect 423544 468721 434144 473428
rect 378904 422671 434144 468721
rect 378904 417148 389504 422671
rect 378904 410428 388544 417148
rect 389344 410428 389504 417148
rect 378904 405721 389504 410428
rect 390304 405721 399944 422671
rect 400744 405721 400904 422671
rect 401704 405721 411344 422671
rect 412144 405721 412304 422671
rect 413104 405721 422744 422671
rect 423544 417148 434144 422671
rect 423544 410428 423704 417148
rect 424504 410428 434144 417148
rect 423544 405721 434144 410428
rect 378904 359671 434144 405721
rect 378904 354148 389504 359671
rect 378904 347428 388544 354148
rect 389344 347428 389504 354148
rect 378904 342721 389504 347428
rect 390304 342721 399944 359671
rect 400744 342721 400904 359671
rect 401704 342721 411344 359671
rect 412144 342721 412304 359671
rect 413104 342721 422744 359671
rect 423544 354148 434144 359671
rect 423544 347428 423704 354148
rect 424504 347428 434144 354148
rect 423544 342721 434144 347428
rect 378904 296671 434144 342721
rect 378904 291148 389504 296671
rect 378904 284428 388544 291148
rect 389344 284428 389504 291148
rect 378904 279721 389504 284428
rect 390304 279721 399944 296671
rect 400744 279721 400904 296671
rect 401704 279721 411344 296671
rect 412144 279721 412304 296671
rect 413104 279721 422744 296671
rect 423544 291148 434144 296671
rect 423544 284428 423704 291148
rect 424504 284428 434144 291148
rect 423544 279721 434144 284428
rect 378904 233671 434144 279721
rect 378904 228148 389504 233671
rect 378904 221428 388544 228148
rect 389344 221428 389504 228148
rect 378904 216721 389504 221428
rect 390304 216721 399944 233671
rect 400744 216721 400904 233671
rect 401704 216721 411344 233671
rect 412144 216721 412304 233671
rect 413104 216721 422744 233671
rect 423544 228148 434144 233671
rect 423544 221428 423704 228148
rect 424504 221428 434144 228148
rect 423544 216721 434144 221428
rect 378904 170671 434144 216721
rect 378904 165148 389504 170671
rect 378904 158428 388544 165148
rect 389344 158428 389504 165148
rect 378904 153721 389504 158428
rect 390304 153721 399944 170671
rect 400744 153721 400904 170671
rect 401704 153721 411344 170671
rect 412144 153721 412304 170671
rect 413104 153721 422744 170671
rect 423544 165148 434144 170671
rect 423544 158428 423704 165148
rect 424504 158428 434144 165148
rect 423544 153721 434144 158428
rect 378904 107671 434144 153721
rect 378904 102148 389504 107671
rect 378904 95428 388544 102148
rect 389344 95428 389504 102148
rect 378904 90721 389504 95428
rect 390304 90721 399944 107671
rect 400744 90721 400904 107671
rect 401704 90721 411344 107671
rect 412144 90721 412304 107671
rect 413104 90721 422744 107671
rect 423544 102148 434144 107671
rect 423544 95428 423704 102148
rect 424504 95428 434144 102148
rect 423544 90721 434144 95428
rect 378904 44671 434144 90721
rect 378904 39148 389504 44671
rect 378904 32508 388544 39148
rect 389344 32508 389504 39148
rect 378904 8128 389504 32508
rect 390304 32969 399944 44671
rect 400744 32969 400904 44671
rect 401704 32969 411344 44671
rect 412144 32969 412304 44671
rect 413104 32969 422744 44671
rect 390304 13575 422744 32969
rect 390304 8128 399944 13575
rect 400744 8128 400904 13575
rect 401704 8128 411344 13575
rect 412144 8128 412304 13575
rect 413104 8128 422744 13575
rect 423544 39148 434144 44671
rect 423544 32508 423704 39148
rect 424504 32508 434144 39148
rect 423544 8128 434144 32508
rect 434944 8128 435104 534448
rect 435904 481455 486264 534448
rect 435904 480148 446504 481455
rect 435904 473428 445544 480148
rect 446344 473428 446504 480148
rect 435904 472937 446504 473428
rect 447304 472937 456944 481455
rect 457744 472937 457904 481455
rect 458704 472937 468344 481455
rect 469144 472937 469304 481455
rect 470104 472937 479744 481455
rect 480544 480148 486264 481455
rect 480544 473428 480704 480148
rect 481504 473428 486264 480148
rect 480544 472937 486264 473428
rect 435904 417367 486264 472937
rect 435904 417148 446504 417367
rect 435904 410428 445544 417148
rect 446344 410428 446504 417148
rect 435904 409937 446504 410428
rect 447304 409937 456944 417367
rect 457744 409937 457904 417367
rect 458704 409937 468344 417367
rect 469144 409937 469304 417367
rect 470104 409937 479744 417367
rect 480544 417148 486264 417367
rect 480544 410428 480704 417148
rect 481504 410428 486264 417148
rect 480544 409937 486264 410428
rect 435904 354367 486264 409937
rect 435904 354148 446504 354367
rect 435904 347428 445544 354148
rect 446344 347428 446504 354148
rect 435904 346937 446504 347428
rect 447304 346937 456944 354367
rect 457744 346937 457904 354367
rect 458704 346937 468344 354367
rect 469144 346937 469304 354367
rect 470104 346937 479744 354367
rect 480544 354148 486264 354367
rect 480544 347428 480704 354148
rect 481504 347428 486264 354148
rect 480544 346937 486264 347428
rect 435904 291367 486264 346937
rect 435904 291148 446504 291367
rect 435904 284428 445544 291148
rect 446344 284428 446504 291148
rect 435904 283937 446504 284428
rect 447304 283937 456944 291367
rect 457744 283937 457904 291367
rect 458704 283937 468344 291367
rect 469144 283937 469304 291367
rect 470104 283937 479744 291367
rect 480544 291148 486264 291367
rect 480544 284428 480704 291148
rect 481504 284428 486264 291148
rect 480544 283937 486264 284428
rect 435904 228367 486264 283937
rect 435904 228148 446504 228367
rect 435904 221428 445544 228148
rect 446344 221428 446504 228148
rect 435904 220937 446504 221428
rect 447304 220937 456944 228367
rect 457744 220937 457904 228367
rect 458704 220937 468344 228367
rect 469144 220937 469304 228367
rect 470104 220937 479744 228367
rect 480544 228148 486264 228367
rect 480544 221428 480704 228148
rect 481504 221428 486264 228148
rect 480544 220937 486264 221428
rect 435904 165367 486264 220937
rect 435904 165148 446504 165367
rect 435904 158428 445544 165148
rect 446344 158428 446504 165148
rect 435904 157937 446504 158428
rect 447304 157937 456944 165367
rect 457744 157937 457904 165367
rect 458704 157937 468344 165367
rect 469144 157937 469304 165367
rect 470104 157937 479744 165367
rect 480544 165148 486264 165367
rect 480544 158428 480704 165148
rect 481504 158428 486264 165148
rect 480544 157937 486264 158428
rect 435904 102367 486264 157937
rect 435904 102148 446504 102367
rect 435904 95428 445544 102148
rect 446344 95428 446504 102148
rect 435904 94937 446504 95428
rect 447304 94937 456944 102367
rect 457744 94937 457904 102367
rect 458704 94937 468344 102367
rect 469144 94937 469304 102367
rect 470104 94937 479744 102367
rect 480544 102148 486264 102367
rect 480544 95428 480704 102148
rect 481504 95428 486264 102148
rect 480544 94937 486264 95428
rect 435904 39367 486264 94937
rect 435904 39148 446504 39367
rect 435904 32508 445544 39148
rect 446344 32508 446504 39148
rect 435904 32153 446504 32508
rect 447304 32153 456944 39367
rect 457744 32153 457904 39367
rect 458704 32153 468344 39367
rect 435904 12215 468344 32153
rect 435904 8128 446504 12215
rect 447304 8128 456944 12215
rect 457744 8128 457904 12215
rect 458704 8128 468344 12215
rect 469144 8128 469304 39367
rect 470104 8128 479744 39367
rect 480544 39148 486264 39367
rect 480544 32508 480704 39148
rect 481504 32508 486264 39148
rect 480544 8128 486264 32508
<< metal5 >>
rect -2552 542696 497512 543656
rect -1192 541336 496152 542296
rect -2552 539356 497512 539996
rect -2552 530136 497512 530776
rect -2552 528856 497512 529496
rect -2552 519636 497512 520276
rect -2552 518356 497512 518996
rect -2552 509136 497512 509776
rect -2552 507856 497512 508496
rect -2552 498636 497512 499276
rect -2552 497356 497512 497996
rect -2552 488136 497512 488776
rect -2552 486856 497512 487496
rect -2552 477636 497512 478276
rect -2552 476356 497512 476996
rect -2552 467136 497512 467776
rect -2552 465856 497512 466496
rect -2552 456636 497512 457276
rect -2552 455356 497512 455996
rect -2552 446136 497512 446776
rect -2552 444856 497512 445496
rect -2552 435636 497512 436276
rect -2552 434356 497512 434996
rect -2552 425136 497512 425776
rect -2552 423856 497512 424496
rect -2552 414636 497512 415276
rect -2552 413356 497512 413996
rect -2552 404136 497512 404776
rect -2552 402856 497512 403496
rect -2552 393636 497512 394276
rect -2552 392356 497512 392996
rect -2552 383136 497512 383776
rect -2552 381856 497512 382496
rect -2552 372636 497512 373276
rect -2552 371356 497512 371996
rect -2552 362136 497512 362776
rect -2552 360856 497512 361496
rect -2552 351636 497512 352276
rect -2552 350356 497512 350996
rect -2552 341136 497512 341776
rect -2552 339856 497512 340496
rect -2552 330636 497512 331276
rect -2552 329356 497512 329996
rect -2552 320136 497512 320776
rect -2552 318856 497512 319496
rect -2552 309636 497512 310276
rect -2552 308356 497512 308996
rect -2552 299136 497512 299776
rect -2552 297856 497512 298496
rect -2552 288636 497512 289276
rect -2552 287356 497512 287996
rect -2552 278136 497512 278776
rect -2552 276856 497512 277496
rect -2552 267636 497512 268276
rect -2552 266356 497512 266996
rect -2552 257136 497512 257776
rect -2552 255856 497512 256496
rect -2552 246636 497512 247276
rect -2552 245356 497512 245996
rect -2552 236136 497512 236776
rect -2552 234856 497512 235496
rect -2552 225636 497512 226276
rect -2552 224356 497512 224996
rect -2552 215136 497512 215776
rect -2552 213856 497512 214496
rect -2552 204636 497512 205276
rect -2552 203356 497512 203996
rect -2552 194136 497512 194776
rect -2552 192856 497512 193496
rect -2552 183636 497512 184276
rect -2552 182356 497512 182996
rect -2552 173136 497512 173776
rect -2552 171856 497512 172496
rect -2552 162636 497512 163276
rect -2552 161356 497512 161996
rect -2552 152136 497512 152776
rect -2552 150856 497512 151496
rect -2552 141636 497512 142276
rect -2552 140356 497512 140996
rect -2552 131136 497512 131776
rect -2552 129856 497512 130496
rect -2552 120636 497512 121276
rect -2552 119356 497512 119996
rect -2552 110136 497512 110776
rect -2552 108856 497512 109496
rect -2552 99636 497512 100276
rect -2552 98356 497512 98996
rect -2552 89136 497512 89776
rect -2552 87856 497512 88496
rect -2552 78636 497512 79276
rect -2552 77356 497512 77996
rect -2552 68136 497512 68776
rect -2552 66856 497512 67496
rect -2552 57636 497512 58276
rect -2552 56356 497512 56996
rect -2552 47136 497512 47776
rect -2552 45856 497512 46496
rect -2552 36636 497512 37276
rect -2552 35356 497512 35996
rect -2552 26136 497512 26776
rect -2552 24856 497512 25496
rect -2552 15636 497512 16276
rect -2552 14356 497512 14996
rect -2552 5136 497512 5776
rect -2552 3856 497512 4496
rect -1192 616 496152 1576
rect -2552 -744 497512 216
<< labels >>
rlabel metal4 s -2552 -744 -1592 543656 4 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 -744 497512 216 8 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 542696 497512 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 496552 -744 497512 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1984 -744 2624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 -744 14024 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 34273 14024 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 95508 14024 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 158508 14024 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 221508 14024 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 284508 14024 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 347508 14024 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 410508 14024 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 473508 14024 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 536508 14024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 -744 25424 13495 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 34273 25424 39831 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 95017 25424 102831 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 158017 25424 165831 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 221017 25424 228831 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 284017 25424 291831 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 347017 25424 354831 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 410017 25424 417831 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 473017 25424 480423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 523777 25424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 36184 -744 36824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 -744 48224 44591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 90801 48224 107591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 153801 48224 170591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 216801 48224 233591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 279801 48224 296591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 342801 48224 359591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 405801 48224 422591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 468801 48224 484231 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 531257 48224 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 -744 59624 13495 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 33049 59624 44591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 90801 59624 107591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 153801 59624 170591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 216801 59624 233591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 279801 59624 296591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 342801 59624 359591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 405801 59624 422591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 468801 59624 484231 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 531257 59624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 -744 71024 13495 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 33049 71024 44591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 90801 71024 107591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 153801 71024 170591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 216801 71024 233591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 279801 71024 296591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 342801 71024 359591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 405801 71024 422591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 468801 71024 484231 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 531257 71024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 -744 82424 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 32588 82424 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 95508 82424 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 158508 82424 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 221508 82424 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 284508 82424 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 347508 82424 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 410508 82424 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 473508 82424 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 536508 82424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 93184 -744 93824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 -744 105224 44591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 90801 105224 107591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 153801 105224 170591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 216801 105224 233591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 279801 105224 296591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 342801 105224 359591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 405801 105224 422591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 468801 105224 484231 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 531257 105224 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 -744 116624 13495 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 33049 116624 44591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 90801 116624 107591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 153801 116624 170591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 216801 116624 233591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 279801 116624 296591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 342801 116624 359591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 405801 116624 422591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 468801 116624 484231 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 531257 116624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 -744 128024 13495 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 33049 128024 44591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 90801 128024 107591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 153801 128024 170591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 216801 128024 233591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 279801 128024 296591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 342801 128024 359591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 405801 128024 422591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 468801 128024 484231 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 531257 128024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 -744 139424 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 32588 139424 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 95508 139424 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 158508 139424 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 221508 139424 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 284508 139424 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 347508 139424 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 410508 139424 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 473508 139424 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 536508 139424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 150184 -744 150824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 -744 162224 44591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 90801 162224 107591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 153801 162224 170591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 216801 162224 233591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 279801 162224 296591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 342801 162224 359591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 405801 162224 422591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 468801 162224 484231 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 531257 162224 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 -744 173624 13495 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 33049 173624 44591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 90801 173624 107591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 153801 173624 170591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 216801 173624 233591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 279801 173624 296591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 342801 173624 359591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 405801 173624 422591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 468801 173624 484231 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 531257 173624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 -744 185024 13495 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 33049 185024 44591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 90801 185024 107591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 153801 185024 170591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 216801 185024 233591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 279801 185024 296591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 342801 185024 359591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 405801 185024 422591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 468801 185024 484231 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 531257 185024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 -744 196424 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 32588 196424 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 95508 196424 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 158508 196424 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 221508 196424 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 284508 196424 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 347508 196424 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 410508 196424 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 473508 196424 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 536508 196424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 207184 -744 207824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 -744 219224 44591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 90801 219224 107591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 153801 219224 170591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 216801 219224 233591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 279801 219224 296591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 342801 219224 359591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 405801 219224 422591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 468801 219224 484231 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 531257 219224 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 -744 230624 13495 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 33049 230624 44591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 90801 230624 107591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 153801 230624 170591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 216801 230624 233591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 279801 230624 296591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 342801 230624 359591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 405801 230624 422591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 468801 230624 484231 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 531257 230624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 -744 242024 13495 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 33049 242024 44591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 90801 242024 107591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 153801 242024 170591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 216801 242024 233591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 279801 242024 296591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 342801 242024 359591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 405801 242024 422591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 468801 242024 484231 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 531257 242024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 -744 253424 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 32588 253424 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 95508 253424 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 158508 253424 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 221508 253424 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 284508 253424 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 347508 253424 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 410508 253424 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 473508 253424 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 536508 253424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 264184 -744 264824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 -744 276224 44591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 90801 276224 107591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 153801 276224 170591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 216801 276224 233591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 279801 276224 296591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 342801 276224 359591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 405801 276224 422591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 468801 276224 484231 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 531257 276224 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 -744 287624 13495 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 33049 287624 44591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 90801 287624 107591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 153801 287624 170591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 216801 287624 233591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 279801 287624 296591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 342801 287624 359591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 405801 287624 422591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 468801 287624 484231 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 531257 287624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 -744 299024 13495 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 33049 299024 44591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 90801 299024 107591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 153801 299024 170591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 216801 299024 233591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 279801 299024 296591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 342801 299024 359591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 405801 299024 422591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 468801 299024 484231 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 531257 299024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 -744 310424 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 32588 310424 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 95508 310424 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 158508 310424 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 221508 310424 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 284508 310424 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 347508 310424 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 410508 310424 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 473508 310424 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 536508 310424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 321184 -744 321824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 -744 333224 44591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 90801 333224 107591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 153801 333224 170591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 216801 333224 233591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 279801 333224 296591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 342801 333224 359591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 405801 333224 422591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 468801 333224 484231 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 531257 333224 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 -744 344624 13495 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 33049 344624 44591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 90801 344624 107591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 153801 344624 170591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 216801 344624 233591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 279801 344624 296591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 342801 344624 359591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 405801 344624 422591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 468801 344624 484231 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 531257 344624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 -744 356024 13495 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 33049 356024 44591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 90801 356024 107591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 153801 356024 170591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 216801 356024 233591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 279801 356024 296591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 342801 356024 359591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 405801 356024 422591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 468801 356024 484231 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 531257 356024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 -744 367424 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 32588 367424 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 95508 367424 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 158508 367424 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 221508 367424 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 284508 367424 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 347508 367424 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 410508 367424 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 473508 367424 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 536508 367424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 378184 -744 378824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 -744 390224 44591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 90801 390224 107591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 153801 390224 170591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 216801 390224 233591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 279801 390224 296591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 342801 390224 359591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 405801 390224 422591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 468801 390224 484231 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 531257 390224 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 -744 401624 13495 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 33049 401624 44591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 90801 401624 107591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 153801 401624 170591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 216801 401624 233591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 279801 401624 296591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 342801 401624 359591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 405801 401624 422591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 468801 401624 484231 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 531257 401624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 -744 413024 13495 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 33049 413024 44591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 90801 413024 107591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 153801 413024 170591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 216801 413024 233591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 279801 413024 296591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 342801 413024 359591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 405801 413024 422591 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 468801 413024 484231 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 531257 413024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 -744 424424 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 32588 424424 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 95508 424424 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 158508 424424 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 221508 424424 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 284508 424424 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 347508 424424 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 410508 424424 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 473508 424424 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 536508 424424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 435184 -744 435824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 -744 447224 12135 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 32233 447224 39287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 95017 447224 102287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 158017 447224 165287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 221017 447224 228287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 284017 447224 291287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 347017 447224 354287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 410017 447224 417287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 473017 447224 481375 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 536017 447224 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 -744 458624 12135 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 32233 458624 39287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 95017 458624 102287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 158017 458624 165287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 221017 458624 228287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 284017 458624 291287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 347017 458624 354287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 410017 458624 417287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 473017 458624 481375 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 536017 458624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 -744 470024 39287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 95017 470024 102287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 158017 470024 165287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 221017 470024 228287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 284017 470024 291287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 347017 470024 354287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 410017 470024 417287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 473017 470024 481375 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 536017 470024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 -744 481424 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 32588 481424 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 95508 481424 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 158508 481424 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 221508 481424 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 284508 481424 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 347508 481424 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 410508 481424 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 473508 481424 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 536508 481424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 492184 -744 492824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 5136 497512 5776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 15636 497512 16276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 26136 497512 26776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 36636 497512 37276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 47136 497512 47776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 57636 497512 58276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 68136 497512 68776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 78636 497512 79276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 89136 497512 89776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 99636 497512 100276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 110136 497512 110776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 120636 497512 121276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 131136 497512 131776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 141636 497512 142276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 152136 497512 152776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 162636 497512 163276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 173136 497512 173776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 183636 497512 184276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 194136 497512 194776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 204636 497512 205276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 215136 497512 215776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 225636 497512 226276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 236136 497512 236776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 246636 497512 247276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 257136 497512 257776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 267636 497512 268276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 278136 497512 278776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 288636 497512 289276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 299136 497512 299776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 309636 497512 310276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 320136 497512 320776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 330636 497512 331276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 341136 497512 341776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 351636 497512 352276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 362136 497512 362776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 372636 497512 373276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 383136 497512 383776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 393636 497512 394276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 404136 497512 404776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 414636 497512 415276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 425136 497512 425776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 435636 497512 436276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 446136 497512 446776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 456636 497512 457276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 467136 497512 467776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 477636 497512 478276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 488136 497512 488776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 498636 497512 499276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 509136 497512 509776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 519636 497512 520276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 530136 497512 530776 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s -1192 616 -232 542296 4 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -1192 616 496152 1576 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -1192 541336 496152 542296 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 495192 616 496152 542296 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 1024 -744 1664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12424 -744 13064 13495 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12424 34273 13064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 -744 24464 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 34273 24464 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 95508 24464 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 158508 24464 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 221508 24464 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 284508 24464 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 347508 24464 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 410508 24464 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 473508 24464 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 536508 24464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 35224 -744 35864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 -744 47264 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 32588 47264 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 95508 47264 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 158508 47264 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 221508 47264 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 284508 47264 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 347508 47264 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 410508 47264 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 473508 47264 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 536508 47264 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 -744 58664 13495 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 33049 58664 44591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 90801 58664 107591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 153801 58664 170591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 216801 58664 233591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 279801 58664 296591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 342801 58664 359591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 405801 58664 422591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 468801 58664 484231 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 531257 58664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 -744 70064 13495 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 33049 70064 44591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 90801 70064 107591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 153801 70064 170591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 216801 70064 233591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 279801 70064 296591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 342801 70064 359591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 405801 70064 422591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 468801 70064 484231 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 531257 70064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 -744 81464 44591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 90801 81464 107591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 153801 81464 170591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 216801 81464 233591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 279801 81464 296591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 342801 81464 359591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 405801 81464 422591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 468801 81464 484231 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 531257 81464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 92224 -744 92864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 -744 104264 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 32588 104264 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 95508 104264 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 158508 104264 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 221508 104264 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 284508 104264 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 347508 104264 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 410508 104264 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 473508 104264 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 536508 104264 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 -744 115664 13495 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 33049 115664 44591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 90801 115664 107591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 153801 115664 170591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 216801 115664 233591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 279801 115664 296591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 342801 115664 359591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 405801 115664 422591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 468801 115664 484231 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 531257 115664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 -744 127064 13495 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 33049 127064 44591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 90801 127064 107591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 153801 127064 170591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 216801 127064 233591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 279801 127064 296591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 342801 127064 359591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 405801 127064 422591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 468801 127064 484231 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 531257 127064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 -744 138464 44591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 90801 138464 107591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 153801 138464 170591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 216801 138464 233591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 279801 138464 296591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 342801 138464 359591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 405801 138464 422591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 468801 138464 484231 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 531257 138464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 149224 -744 149864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 -744 161264 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 32588 161264 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 95508 161264 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 158508 161264 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 221508 161264 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 284508 161264 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 347508 161264 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 410508 161264 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 473508 161264 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 536508 161264 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 -744 172664 13495 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 33049 172664 44591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 90801 172664 107591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 153801 172664 170591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 216801 172664 233591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 279801 172664 296591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 342801 172664 359591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 405801 172664 422591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 468801 172664 484231 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 531257 172664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 -744 184064 13495 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 33049 184064 44591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 90801 184064 107591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 153801 184064 170591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 216801 184064 233591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 279801 184064 296591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 342801 184064 359591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 405801 184064 422591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 468801 184064 484231 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 531257 184064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 -744 195464 44591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 90801 195464 107591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 153801 195464 170591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 216801 195464 233591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 279801 195464 296591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 342801 195464 359591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 405801 195464 422591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 468801 195464 484231 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 531257 195464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 206224 -744 206864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 -744 218264 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 32588 218264 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 95508 218264 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 158508 218264 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 221508 218264 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 284508 218264 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 347508 218264 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 410508 218264 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 473508 218264 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 536508 218264 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 -744 229664 13495 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 33049 229664 44591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 90801 229664 107591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 153801 229664 170591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 216801 229664 233591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 279801 229664 296591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 342801 229664 359591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 405801 229664 422591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 468801 229664 484231 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 531257 229664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 -744 241064 13495 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 33049 241064 44591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 90801 241064 107591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 153801 241064 170591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 216801 241064 233591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 279801 241064 296591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 342801 241064 359591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 405801 241064 422591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 468801 241064 484231 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 531257 241064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 -744 252464 44591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 90801 252464 107591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 153801 252464 170591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 216801 252464 233591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 279801 252464 296591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 342801 252464 359591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 405801 252464 422591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 468801 252464 484231 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 531257 252464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 263224 -744 263864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 -744 275264 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 32588 275264 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 95508 275264 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 158508 275264 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 221508 275264 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 284508 275264 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 347508 275264 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 410508 275264 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 473508 275264 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 536508 275264 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 -744 286664 13495 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 33049 286664 44591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 90801 286664 107591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 153801 286664 170591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 216801 286664 233591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 279801 286664 296591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 342801 286664 359591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 405801 286664 422591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 468801 286664 484231 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 531257 286664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 -744 298064 13495 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 33049 298064 44591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 90801 298064 107591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 153801 298064 170591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 216801 298064 233591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 279801 298064 296591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 342801 298064 359591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 405801 298064 422591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 468801 298064 484231 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 531257 298064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 -744 309464 44591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 90801 309464 107591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 153801 309464 170591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 216801 309464 233591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 279801 309464 296591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 342801 309464 359591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 405801 309464 422591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 468801 309464 484231 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 531257 309464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 320224 -744 320864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 -744 332264 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 32588 332264 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 95508 332264 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 158508 332264 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 221508 332264 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 284508 332264 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 347508 332264 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 410508 332264 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 473508 332264 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 536508 332264 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 -744 343664 13495 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 33049 343664 44591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 90801 343664 107591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 153801 343664 170591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 216801 343664 233591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 279801 343664 296591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 342801 343664 359591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 405801 343664 422591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 468801 343664 484231 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 531257 343664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 -744 355064 13495 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 33049 355064 44591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 90801 355064 107591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 153801 355064 170591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 216801 355064 233591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 279801 355064 296591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 342801 355064 359591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 405801 355064 422591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 468801 355064 484231 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 531257 355064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 -744 366464 44591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 90801 366464 107591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 153801 366464 170591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 216801 366464 233591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 279801 366464 296591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 342801 366464 359591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 405801 366464 422591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 468801 366464 484231 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 531257 366464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 377224 -744 377864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 -744 389264 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 32588 389264 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 95508 389264 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 158508 389264 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 221508 389264 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 284508 389264 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 347508 389264 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 410508 389264 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 473508 389264 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 536508 389264 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 -744 400664 13495 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 33049 400664 44591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 90801 400664 107591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 153801 400664 170591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 216801 400664 233591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 279801 400664 296591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 342801 400664 359591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 405801 400664 422591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 468801 400664 484231 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 531257 400664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 -744 412064 13495 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 33049 412064 44591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 90801 412064 107591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 153801 412064 170591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 216801 412064 233591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 279801 412064 296591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 342801 412064 359591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 405801 412064 422591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 468801 412064 484231 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 531257 412064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 -744 423464 44591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 90801 423464 107591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 153801 423464 170591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 216801 423464 233591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 279801 423464 296591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 342801 423464 359591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 405801 423464 422591 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 468801 423464 484231 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 531257 423464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 434224 -744 434864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 -744 446264 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 32588 446264 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 95508 446264 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 158508 446264 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 221508 446264 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 284508 446264 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 347508 446264 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 410508 446264 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 473508 446264 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 536508 446264 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 -744 457664 12135 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 32233 457664 39287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 95017 457664 102287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 158017 457664 165287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 221017 457664 228287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 284017 457664 291287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 347017 457664 354287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 410017 457664 417287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 473017 457664 481375 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 536017 457664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 -744 469064 39287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 95017 469064 102287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 158017 469064 165287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 221017 469064 228287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 284017 469064 291287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 347017 469064 354287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 410017 469064 417287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 473017 469064 481375 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 536017 469064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 -744 480464 39287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 95017 480464 102287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 158017 480464 165287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 221017 480464 228287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 284017 480464 291287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 347017 480464 354287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 410017 480464 417287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 473017 480464 481375 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 536017 480464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 491224 -744 491864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 3856 497512 4496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 14356 497512 14996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 24856 497512 25496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 35356 497512 35996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 45856 497512 46496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 56356 497512 56996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 66856 497512 67496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 77356 497512 77996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 87856 497512 88496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 98356 497512 98996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 108856 497512 109496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 119356 497512 119996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 129856 497512 130496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 140356 497512 140996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 150856 497512 151496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 161356 497512 161996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 171856 497512 172496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 182356 497512 182996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 192856 497512 193496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 203356 497512 203996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 213856 497512 214496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 224356 497512 224996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 234856 497512 235496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 245356 497512 245996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 255856 497512 256496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 266356 497512 266996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 276856 497512 277496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 287356 497512 287996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 297856 497512 298496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 308356 497512 308996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 318856 497512 319496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 329356 497512 329996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 339856 497512 340496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 350356 497512 350996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 360856 497512 361496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 371356 497512 371996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 381856 497512 382496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 392356 497512 392996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 402856 497512 403496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 413356 497512 413996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 423856 497512 424496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 434356 497512 434996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 444856 497512 445496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 455356 497512 455996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 465856 497512 466496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 476356 497512 476996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 486856 497512 487496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 497356 497512 497996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 507856 497512 508496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 518356 497512 518996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 528856 497512 529496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 539356 497512 539996 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 73526 0 73582 800 6 ccff_head
port 3 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 ccff_tail
port 4 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 clk
port 5 nsew signal input
rlabel metal2 s 12990 542200 13046 543000 6 gfpga_pad_io_soc_dir[0]
port 6 nsew signal output
rlabel metal3 s 0 97248 800 97368 6 gfpga_pad_io_soc_dir[100]
port 7 nsew signal output
rlabel metal3 s 0 113568 800 113688 6 gfpga_pad_io_soc_dir[101]
port 8 nsew signal output
rlabel metal3 s 0 129888 800 130008 6 gfpga_pad_io_soc_dir[102]
port 9 nsew signal output
rlabel metal3 s 0 146208 800 146328 6 gfpga_pad_io_soc_dir[103]
port 10 nsew signal output
rlabel metal3 s 0 162528 800 162648 6 gfpga_pad_io_soc_dir[104]
port 11 nsew signal output
rlabel metal3 s 0 178848 800 178968 6 gfpga_pad_io_soc_dir[105]
port 12 nsew signal output
rlabel metal3 s 0 195168 800 195288 6 gfpga_pad_io_soc_dir[106]
port 13 nsew signal output
rlabel metal3 s 0 211488 800 211608 6 gfpga_pad_io_soc_dir[107]
port 14 nsew signal output
rlabel metal3 s 0 227808 800 227928 6 gfpga_pad_io_soc_dir[108]
port 15 nsew signal output
rlabel metal3 s 0 244128 800 244248 6 gfpga_pad_io_soc_dir[109]
port 16 nsew signal output
rlabel metal2 s 152738 542200 152794 543000 6 gfpga_pad_io_soc_dir[10]
port 17 nsew signal output
rlabel metal3 s 0 260448 800 260568 6 gfpga_pad_io_soc_dir[110]
port 18 nsew signal output
rlabel metal3 s 0 276768 800 276888 6 gfpga_pad_io_soc_dir[111]
port 19 nsew signal output
rlabel metal3 s 0 293088 800 293208 6 gfpga_pad_io_soc_dir[112]
port 20 nsew signal output
rlabel metal3 s 0 309408 800 309528 6 gfpga_pad_io_soc_dir[113]
port 21 nsew signal output
rlabel metal3 s 0 325728 800 325848 6 gfpga_pad_io_soc_dir[114]
port 22 nsew signal output
rlabel metal3 s 0 342048 800 342168 6 gfpga_pad_io_soc_dir[115]
port 23 nsew signal output
rlabel metal3 s 0 358368 800 358488 6 gfpga_pad_io_soc_dir[116]
port 24 nsew signal output
rlabel metal3 s 0 374688 800 374808 6 gfpga_pad_io_soc_dir[117]
port 25 nsew signal output
rlabel metal3 s 0 391008 800 391128 6 gfpga_pad_io_soc_dir[118]
port 26 nsew signal output
rlabel metal3 s 0 407328 800 407448 6 gfpga_pad_io_soc_dir[119]
port 27 nsew signal output
rlabel metal2 s 166262 542200 166318 543000 6 gfpga_pad_io_soc_dir[11]
port 28 nsew signal output
rlabel metal3 s 0 423648 800 423768 6 gfpga_pad_io_soc_dir[120]
port 29 nsew signal output
rlabel metal3 s 0 439968 800 440088 6 gfpga_pad_io_soc_dir[121]
port 30 nsew signal output
rlabel metal3 s 0 456288 800 456408 6 gfpga_pad_io_soc_dir[122]
port 31 nsew signal output
rlabel metal3 s 0 472608 800 472728 6 gfpga_pad_io_soc_dir[123]
port 32 nsew signal output
rlabel metal3 s 0 488928 800 489048 6 gfpga_pad_io_soc_dir[124]
port 33 nsew signal output
rlabel metal3 s 0 505248 800 505368 6 gfpga_pad_io_soc_dir[125]
port 34 nsew signal output
rlabel metal3 s 0 521568 800 521688 6 gfpga_pad_io_soc_dir[126]
port 35 nsew signal output
rlabel metal3 s 0 537888 800 538008 6 gfpga_pad_io_soc_dir[127]
port 36 nsew signal output
rlabel metal2 s 179786 542200 179842 543000 6 gfpga_pad_io_soc_dir[12]
port 37 nsew signal output
rlabel metal2 s 193310 542200 193366 543000 6 gfpga_pad_io_soc_dir[13]
port 38 nsew signal output
rlabel metal2 s 206834 542200 206890 543000 6 gfpga_pad_io_soc_dir[14]
port 39 nsew signal output
rlabel metal2 s 220358 542200 220414 543000 6 gfpga_pad_io_soc_dir[15]
port 40 nsew signal output
rlabel metal2 s 233882 542200 233938 543000 6 gfpga_pad_io_soc_dir[16]
port 41 nsew signal output
rlabel metal2 s 247406 542200 247462 543000 6 gfpga_pad_io_soc_dir[17]
port 42 nsew signal output
rlabel metal2 s 260930 542200 260986 543000 6 gfpga_pad_io_soc_dir[18]
port 43 nsew signal output
rlabel metal2 s 274454 542200 274510 543000 6 gfpga_pad_io_soc_dir[19]
port 44 nsew signal output
rlabel metal2 s 26514 542200 26570 543000 6 gfpga_pad_io_soc_dir[1]
port 45 nsew signal output
rlabel metal2 s 287978 542200 288034 543000 6 gfpga_pad_io_soc_dir[20]
port 46 nsew signal output
rlabel metal2 s 301502 542200 301558 543000 6 gfpga_pad_io_soc_dir[21]
port 47 nsew signal output
rlabel metal2 s 315026 542200 315082 543000 6 gfpga_pad_io_soc_dir[22]
port 48 nsew signal output
rlabel metal2 s 328550 542200 328606 543000 6 gfpga_pad_io_soc_dir[23]
port 49 nsew signal output
rlabel metal2 s 342074 542200 342130 543000 6 gfpga_pad_io_soc_dir[24]
port 50 nsew signal output
rlabel metal2 s 355598 542200 355654 543000 6 gfpga_pad_io_soc_dir[25]
port 51 nsew signal output
rlabel metal2 s 369122 542200 369178 543000 6 gfpga_pad_io_soc_dir[26]
port 52 nsew signal output
rlabel metal2 s 382646 542200 382702 543000 6 gfpga_pad_io_soc_dir[27]
port 53 nsew signal output
rlabel metal2 s 396170 542200 396226 543000 6 gfpga_pad_io_soc_dir[28]
port 54 nsew signal output
rlabel metal2 s 409694 542200 409750 543000 6 gfpga_pad_io_soc_dir[29]
port 55 nsew signal output
rlabel metal2 s 40038 542200 40094 543000 6 gfpga_pad_io_soc_dir[2]
port 56 nsew signal output
rlabel metal2 s 423218 542200 423274 543000 6 gfpga_pad_io_soc_dir[30]
port 57 nsew signal output
rlabel metal2 s 436742 542200 436798 543000 6 gfpga_pad_io_soc_dir[31]
port 58 nsew signal output
rlabel metal2 s 450266 542200 450322 543000 6 gfpga_pad_io_soc_dir[32]
port 59 nsew signal output
rlabel metal2 s 463790 542200 463846 543000 6 gfpga_pad_io_soc_dir[33]
port 60 nsew signal output
rlabel metal2 s 477314 542200 477370 543000 6 gfpga_pad_io_soc_dir[34]
port 61 nsew signal output
rlabel metal2 s 490838 542200 490894 543000 6 gfpga_pad_io_soc_dir[35]
port 62 nsew signal output
rlabel metal3 s 494200 520616 495000 520736 6 gfpga_pad_io_soc_dir[36]
port 63 nsew signal output
rlabel metal3 s 494200 504704 495000 504824 6 gfpga_pad_io_soc_dir[37]
port 64 nsew signal output
rlabel metal3 s 494200 488792 495000 488912 6 gfpga_pad_io_soc_dir[38]
port 65 nsew signal output
rlabel metal3 s 494200 472880 495000 473000 6 gfpga_pad_io_soc_dir[39]
port 66 nsew signal output
rlabel metal2 s 53562 542200 53618 543000 6 gfpga_pad_io_soc_dir[3]
port 67 nsew signal output
rlabel metal3 s 494200 456968 495000 457088 6 gfpga_pad_io_soc_dir[40]
port 68 nsew signal output
rlabel metal3 s 494200 441056 495000 441176 6 gfpga_pad_io_soc_dir[41]
port 69 nsew signal output
rlabel metal3 s 494200 425144 495000 425264 6 gfpga_pad_io_soc_dir[42]
port 70 nsew signal output
rlabel metal3 s 494200 409232 495000 409352 6 gfpga_pad_io_soc_dir[43]
port 71 nsew signal output
rlabel metal3 s 494200 393320 495000 393440 6 gfpga_pad_io_soc_dir[44]
port 72 nsew signal output
rlabel metal3 s 494200 377408 495000 377528 6 gfpga_pad_io_soc_dir[45]
port 73 nsew signal output
rlabel metal3 s 494200 361496 495000 361616 6 gfpga_pad_io_soc_dir[46]
port 74 nsew signal output
rlabel metal3 s 494200 345584 495000 345704 6 gfpga_pad_io_soc_dir[47]
port 75 nsew signal output
rlabel metal3 s 494200 329672 495000 329792 6 gfpga_pad_io_soc_dir[48]
port 76 nsew signal output
rlabel metal3 s 494200 313760 495000 313880 6 gfpga_pad_io_soc_dir[49]
port 77 nsew signal output
rlabel metal2 s 71594 542200 71650 543000 6 gfpga_pad_io_soc_dir[4]
port 78 nsew signal output
rlabel metal3 s 494200 297848 495000 297968 6 gfpga_pad_io_soc_dir[50]
port 79 nsew signal output
rlabel metal3 s 494200 281936 495000 282056 6 gfpga_pad_io_soc_dir[51]
port 80 nsew signal output
rlabel metal3 s 494200 266024 495000 266144 6 gfpga_pad_io_soc_dir[52]
port 81 nsew signal output
rlabel metal3 s 494200 250112 495000 250232 6 gfpga_pad_io_soc_dir[53]
port 82 nsew signal output
rlabel metal3 s 494200 234200 495000 234320 6 gfpga_pad_io_soc_dir[54]
port 83 nsew signal output
rlabel metal3 s 494200 218288 495000 218408 6 gfpga_pad_io_soc_dir[55]
port 84 nsew signal output
rlabel metal3 s 494200 202376 495000 202496 6 gfpga_pad_io_soc_dir[56]
port 85 nsew signal output
rlabel metal3 s 494200 186464 495000 186584 6 gfpga_pad_io_soc_dir[57]
port 86 nsew signal output
rlabel metal3 s 494200 170552 495000 170672 6 gfpga_pad_io_soc_dir[58]
port 87 nsew signal output
rlabel metal3 s 494200 154640 495000 154760 6 gfpga_pad_io_soc_dir[59]
port 88 nsew signal output
rlabel metal2 s 85118 542200 85174 543000 6 gfpga_pad_io_soc_dir[5]
port 89 nsew signal output
rlabel metal3 s 494200 138728 495000 138848 6 gfpga_pad_io_soc_dir[60]
port 90 nsew signal output
rlabel metal3 s 494200 122816 495000 122936 6 gfpga_pad_io_soc_dir[61]
port 91 nsew signal output
rlabel metal3 s 494200 106904 495000 107024 6 gfpga_pad_io_soc_dir[62]
port 92 nsew signal output
rlabel metal3 s 494200 90992 495000 91112 6 gfpga_pad_io_soc_dir[63]
port 93 nsew signal output
rlabel metal3 s 494200 75080 495000 75200 6 gfpga_pad_io_soc_dir[64]
port 94 nsew signal output
rlabel metal3 s 494200 59168 495000 59288 6 gfpga_pad_io_soc_dir[65]
port 95 nsew signal output
rlabel metal3 s 494200 43256 495000 43376 6 gfpga_pad_io_soc_dir[66]
port 96 nsew signal output
rlabel metal3 s 494200 27344 495000 27464 6 gfpga_pad_io_soc_dir[67]
port 97 nsew signal output
rlabel metal2 s 479246 0 479302 800 6 gfpga_pad_io_soc_dir[68]
port 98 nsew signal output
rlabel metal2 s 461858 0 461914 800 6 gfpga_pad_io_soc_dir[69]
port 99 nsew signal output
rlabel metal2 s 98642 542200 98698 543000 6 gfpga_pad_io_soc_dir[6]
port 100 nsew signal output
rlabel metal2 s 444470 0 444526 800 6 gfpga_pad_io_soc_dir[70]
port 101 nsew signal output
rlabel metal2 s 427082 0 427138 800 6 gfpga_pad_io_soc_dir[71]
port 102 nsew signal output
rlabel metal2 s 409694 0 409750 800 6 gfpga_pad_io_soc_dir[72]
port 103 nsew signal output
rlabel metal2 s 392306 0 392362 800 6 gfpga_pad_io_soc_dir[73]
port 104 nsew signal output
rlabel metal2 s 374918 0 374974 800 6 gfpga_pad_io_soc_dir[74]
port 105 nsew signal output
rlabel metal2 s 357530 0 357586 800 6 gfpga_pad_io_soc_dir[75]
port 106 nsew signal output
rlabel metal2 s 340142 0 340198 800 6 gfpga_pad_io_soc_dir[76]
port 107 nsew signal output
rlabel metal2 s 322754 0 322810 800 6 gfpga_pad_io_soc_dir[77]
port 108 nsew signal output
rlabel metal2 s 305366 0 305422 800 6 gfpga_pad_io_soc_dir[78]
port 109 nsew signal output
rlabel metal2 s 287978 0 288034 800 6 gfpga_pad_io_soc_dir[79]
port 110 nsew signal output
rlabel metal2 s 112166 542200 112222 543000 6 gfpga_pad_io_soc_dir[7]
port 111 nsew signal output
rlabel metal2 s 270590 0 270646 800 6 gfpga_pad_io_soc_dir[80]
port 112 nsew signal output
rlabel metal2 s 253202 0 253258 800 6 gfpga_pad_io_soc_dir[81]
port 113 nsew signal output
rlabel metal2 s 235814 0 235870 800 6 gfpga_pad_io_soc_dir[82]
port 114 nsew signal output
rlabel metal2 s 218426 0 218482 800 6 gfpga_pad_io_soc_dir[83]
port 115 nsew signal output
rlabel metal2 s 201038 0 201094 800 6 gfpga_pad_io_soc_dir[84]
port 116 nsew signal output
rlabel metal2 s 183650 0 183706 800 6 gfpga_pad_io_soc_dir[85]
port 117 nsew signal output
rlabel metal2 s 166262 0 166318 800 6 gfpga_pad_io_soc_dir[86]
port 118 nsew signal output
rlabel metal2 s 148874 0 148930 800 6 gfpga_pad_io_soc_dir[87]
port 119 nsew signal output
rlabel metal2 s 131486 0 131542 800 6 gfpga_pad_io_soc_dir[88]
port 120 nsew signal output
rlabel metal2 s 114098 0 114154 800 6 gfpga_pad_io_soc_dir[89]
port 121 nsew signal output
rlabel metal2 s 125690 542200 125746 543000 6 gfpga_pad_io_soc_dir[8]
port 122 nsew signal output
rlabel metal2 s 96710 0 96766 800 6 gfpga_pad_io_soc_dir[90]
port 123 nsew signal output
rlabel metal2 s 79322 0 79378 800 6 gfpga_pad_io_soc_dir[91]
port 124 nsew signal output
rlabel metal2 s 56138 0 56194 800 6 gfpga_pad_io_soc_dir[92]
port 125 nsew signal output
rlabel metal2 s 38750 0 38806 800 6 gfpga_pad_io_soc_dir[93]
port 126 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 gfpga_pad_io_soc_dir[94]
port 127 nsew signal output
rlabel metal2 s 3974 0 4030 800 6 gfpga_pad_io_soc_dir[95]
port 128 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 gfpga_pad_io_soc_dir[96]
port 129 nsew signal output
rlabel metal3 s 0 48288 800 48408 6 gfpga_pad_io_soc_dir[97]
port 130 nsew signal output
rlabel metal3 s 0 64608 800 64728 6 gfpga_pad_io_soc_dir[98]
port 131 nsew signal output
rlabel metal3 s 0 80928 800 81048 6 gfpga_pad_io_soc_dir[99]
port 132 nsew signal output
rlabel metal2 s 139214 542200 139270 543000 6 gfpga_pad_io_soc_dir[9]
port 133 nsew signal output
rlabel metal2 s 3974 542200 4030 543000 6 gfpga_pad_io_soc_in[0]
port 134 nsew signal input
rlabel metal3 s 0 86368 800 86488 6 gfpga_pad_io_soc_in[100]
port 135 nsew signal input
rlabel metal3 s 0 102688 800 102808 6 gfpga_pad_io_soc_in[101]
port 136 nsew signal input
rlabel metal3 s 0 119008 800 119128 6 gfpga_pad_io_soc_in[102]
port 137 nsew signal input
rlabel metal3 s 0 135328 800 135448 6 gfpga_pad_io_soc_in[103]
port 138 nsew signal input
rlabel metal3 s 0 151648 800 151768 6 gfpga_pad_io_soc_in[104]
port 139 nsew signal input
rlabel metal3 s 0 167968 800 168088 6 gfpga_pad_io_soc_in[105]
port 140 nsew signal input
rlabel metal3 s 0 184288 800 184408 6 gfpga_pad_io_soc_in[106]
port 141 nsew signal input
rlabel metal3 s 0 200608 800 200728 6 gfpga_pad_io_soc_in[107]
port 142 nsew signal input
rlabel metal3 s 0 216928 800 217048 6 gfpga_pad_io_soc_in[108]
port 143 nsew signal input
rlabel metal3 s 0 233248 800 233368 6 gfpga_pad_io_soc_in[109]
port 144 nsew signal input
rlabel metal2 s 143722 542200 143778 543000 6 gfpga_pad_io_soc_in[10]
port 145 nsew signal input
rlabel metal3 s 0 249568 800 249688 6 gfpga_pad_io_soc_in[110]
port 146 nsew signal input
rlabel metal3 s 0 265888 800 266008 6 gfpga_pad_io_soc_in[111]
port 147 nsew signal input
rlabel metal3 s 0 282208 800 282328 6 gfpga_pad_io_soc_in[112]
port 148 nsew signal input
rlabel metal3 s 0 298528 800 298648 6 gfpga_pad_io_soc_in[113]
port 149 nsew signal input
rlabel metal3 s 0 314848 800 314968 6 gfpga_pad_io_soc_in[114]
port 150 nsew signal input
rlabel metal3 s 0 331168 800 331288 6 gfpga_pad_io_soc_in[115]
port 151 nsew signal input
rlabel metal3 s 0 347488 800 347608 6 gfpga_pad_io_soc_in[116]
port 152 nsew signal input
rlabel metal3 s 0 363808 800 363928 6 gfpga_pad_io_soc_in[117]
port 153 nsew signal input
rlabel metal3 s 0 380128 800 380248 6 gfpga_pad_io_soc_in[118]
port 154 nsew signal input
rlabel metal3 s 0 396448 800 396568 6 gfpga_pad_io_soc_in[119]
port 155 nsew signal input
rlabel metal2 s 157246 542200 157302 543000 6 gfpga_pad_io_soc_in[11]
port 156 nsew signal input
rlabel metal3 s 0 412768 800 412888 6 gfpga_pad_io_soc_in[120]
port 157 nsew signal input
rlabel metal3 s 0 429088 800 429208 6 gfpga_pad_io_soc_in[121]
port 158 nsew signal input
rlabel metal3 s 0 445408 800 445528 6 gfpga_pad_io_soc_in[122]
port 159 nsew signal input
rlabel metal3 s 0 461728 800 461848 6 gfpga_pad_io_soc_in[123]
port 160 nsew signal input
rlabel metal3 s 0 478048 800 478168 6 gfpga_pad_io_soc_in[124]
port 161 nsew signal input
rlabel metal3 s 0 494368 800 494488 6 gfpga_pad_io_soc_in[125]
port 162 nsew signal input
rlabel metal3 s 0 510688 800 510808 6 gfpga_pad_io_soc_in[126]
port 163 nsew signal input
rlabel metal3 s 0 527008 800 527128 6 gfpga_pad_io_soc_in[127]
port 164 nsew signal input
rlabel metal2 s 170770 542200 170826 543000 6 gfpga_pad_io_soc_in[12]
port 165 nsew signal input
rlabel metal2 s 184294 542200 184350 543000 6 gfpga_pad_io_soc_in[13]
port 166 nsew signal input
rlabel metal2 s 197818 542200 197874 543000 6 gfpga_pad_io_soc_in[14]
port 167 nsew signal input
rlabel metal2 s 211342 542200 211398 543000 6 gfpga_pad_io_soc_in[15]
port 168 nsew signal input
rlabel metal2 s 224866 542200 224922 543000 6 gfpga_pad_io_soc_in[16]
port 169 nsew signal input
rlabel metal2 s 238390 542200 238446 543000 6 gfpga_pad_io_soc_in[17]
port 170 nsew signal input
rlabel metal2 s 251914 542200 251970 543000 6 gfpga_pad_io_soc_in[18]
port 171 nsew signal input
rlabel metal2 s 265438 542200 265494 543000 6 gfpga_pad_io_soc_in[19]
port 172 nsew signal input
rlabel metal2 s 17498 542200 17554 543000 6 gfpga_pad_io_soc_in[1]
port 173 nsew signal input
rlabel metal2 s 278962 542200 279018 543000 6 gfpga_pad_io_soc_in[20]
port 174 nsew signal input
rlabel metal2 s 292486 542200 292542 543000 6 gfpga_pad_io_soc_in[21]
port 175 nsew signal input
rlabel metal2 s 306010 542200 306066 543000 6 gfpga_pad_io_soc_in[22]
port 176 nsew signal input
rlabel metal2 s 319534 542200 319590 543000 6 gfpga_pad_io_soc_in[23]
port 177 nsew signal input
rlabel metal2 s 333058 542200 333114 543000 6 gfpga_pad_io_soc_in[24]
port 178 nsew signal input
rlabel metal2 s 346582 542200 346638 543000 6 gfpga_pad_io_soc_in[25]
port 179 nsew signal input
rlabel metal2 s 360106 542200 360162 543000 6 gfpga_pad_io_soc_in[26]
port 180 nsew signal input
rlabel metal2 s 373630 542200 373686 543000 6 gfpga_pad_io_soc_in[27]
port 181 nsew signal input
rlabel metal2 s 387154 542200 387210 543000 6 gfpga_pad_io_soc_in[28]
port 182 nsew signal input
rlabel metal2 s 400678 542200 400734 543000 6 gfpga_pad_io_soc_in[29]
port 183 nsew signal input
rlabel metal2 s 31022 542200 31078 543000 6 gfpga_pad_io_soc_in[2]
port 184 nsew signal input
rlabel metal2 s 414202 542200 414258 543000 6 gfpga_pad_io_soc_in[30]
port 185 nsew signal input
rlabel metal2 s 427726 542200 427782 543000 6 gfpga_pad_io_soc_in[31]
port 186 nsew signal input
rlabel metal2 s 441250 542200 441306 543000 6 gfpga_pad_io_soc_in[32]
port 187 nsew signal input
rlabel metal2 s 454774 542200 454830 543000 6 gfpga_pad_io_soc_in[33]
port 188 nsew signal input
rlabel metal2 s 468298 542200 468354 543000 6 gfpga_pad_io_soc_in[34]
port 189 nsew signal input
rlabel metal2 s 481822 542200 481878 543000 6 gfpga_pad_io_soc_in[35]
port 190 nsew signal input
rlabel metal3 s 494200 531224 495000 531344 6 gfpga_pad_io_soc_in[36]
port 191 nsew signal input
rlabel metal3 s 494200 515312 495000 515432 6 gfpga_pad_io_soc_in[37]
port 192 nsew signal input
rlabel metal3 s 494200 499400 495000 499520 6 gfpga_pad_io_soc_in[38]
port 193 nsew signal input
rlabel metal3 s 494200 483488 495000 483608 6 gfpga_pad_io_soc_in[39]
port 194 nsew signal input
rlabel metal2 s 44546 542200 44602 543000 6 gfpga_pad_io_soc_in[3]
port 195 nsew signal input
rlabel metal3 s 494200 467576 495000 467696 6 gfpga_pad_io_soc_in[40]
port 196 nsew signal input
rlabel metal3 s 494200 451664 495000 451784 6 gfpga_pad_io_soc_in[41]
port 197 nsew signal input
rlabel metal3 s 494200 435752 495000 435872 6 gfpga_pad_io_soc_in[42]
port 198 nsew signal input
rlabel metal3 s 494200 419840 495000 419960 6 gfpga_pad_io_soc_in[43]
port 199 nsew signal input
rlabel metal3 s 494200 403928 495000 404048 6 gfpga_pad_io_soc_in[44]
port 200 nsew signal input
rlabel metal3 s 494200 388016 495000 388136 6 gfpga_pad_io_soc_in[45]
port 201 nsew signal input
rlabel metal3 s 494200 372104 495000 372224 6 gfpga_pad_io_soc_in[46]
port 202 nsew signal input
rlabel metal3 s 494200 356192 495000 356312 6 gfpga_pad_io_soc_in[47]
port 203 nsew signal input
rlabel metal3 s 494200 340280 495000 340400 6 gfpga_pad_io_soc_in[48]
port 204 nsew signal input
rlabel metal3 s 494200 324368 495000 324488 6 gfpga_pad_io_soc_in[49]
port 205 nsew signal input
rlabel metal2 s 62578 542200 62634 543000 6 gfpga_pad_io_soc_in[4]
port 206 nsew signal input
rlabel metal3 s 494200 308456 495000 308576 6 gfpga_pad_io_soc_in[50]
port 207 nsew signal input
rlabel metal3 s 494200 292544 495000 292664 6 gfpga_pad_io_soc_in[51]
port 208 nsew signal input
rlabel metal3 s 494200 276632 495000 276752 6 gfpga_pad_io_soc_in[52]
port 209 nsew signal input
rlabel metal3 s 494200 260720 495000 260840 6 gfpga_pad_io_soc_in[53]
port 210 nsew signal input
rlabel metal3 s 494200 244808 495000 244928 6 gfpga_pad_io_soc_in[54]
port 211 nsew signal input
rlabel metal3 s 494200 228896 495000 229016 6 gfpga_pad_io_soc_in[55]
port 212 nsew signal input
rlabel metal3 s 494200 212984 495000 213104 6 gfpga_pad_io_soc_in[56]
port 213 nsew signal input
rlabel metal3 s 494200 197072 495000 197192 6 gfpga_pad_io_soc_in[57]
port 214 nsew signal input
rlabel metal3 s 494200 181160 495000 181280 6 gfpga_pad_io_soc_in[58]
port 215 nsew signal input
rlabel metal3 s 494200 165248 495000 165368 6 gfpga_pad_io_soc_in[59]
port 216 nsew signal input
rlabel metal2 s 76102 542200 76158 543000 6 gfpga_pad_io_soc_in[5]
port 217 nsew signal input
rlabel metal3 s 494200 149336 495000 149456 6 gfpga_pad_io_soc_in[60]
port 218 nsew signal input
rlabel metal3 s 494200 133424 495000 133544 6 gfpga_pad_io_soc_in[61]
port 219 nsew signal input
rlabel metal3 s 494200 117512 495000 117632 6 gfpga_pad_io_soc_in[62]
port 220 nsew signal input
rlabel metal3 s 494200 101600 495000 101720 6 gfpga_pad_io_soc_in[63]
port 221 nsew signal input
rlabel metal3 s 494200 85688 495000 85808 6 gfpga_pad_io_soc_in[64]
port 222 nsew signal input
rlabel metal3 s 494200 69776 495000 69896 6 gfpga_pad_io_soc_in[65]
port 223 nsew signal input
rlabel metal3 s 494200 53864 495000 53984 6 gfpga_pad_io_soc_in[66]
port 224 nsew signal input
rlabel metal3 s 494200 37952 495000 38072 6 gfpga_pad_io_soc_in[67]
port 225 nsew signal input
rlabel metal2 s 490838 0 490894 800 6 gfpga_pad_io_soc_in[68]
port 226 nsew signal input
rlabel metal2 s 473450 0 473506 800 6 gfpga_pad_io_soc_in[69]
port 227 nsew signal input
rlabel metal2 s 89626 542200 89682 543000 6 gfpga_pad_io_soc_in[6]
port 228 nsew signal input
rlabel metal2 s 456062 0 456118 800 6 gfpga_pad_io_soc_in[70]
port 229 nsew signal input
rlabel metal2 s 438674 0 438730 800 6 gfpga_pad_io_soc_in[71]
port 230 nsew signal input
rlabel metal2 s 421286 0 421342 800 6 gfpga_pad_io_soc_in[72]
port 231 nsew signal input
rlabel metal2 s 403898 0 403954 800 6 gfpga_pad_io_soc_in[73]
port 232 nsew signal input
rlabel metal2 s 386510 0 386566 800 6 gfpga_pad_io_soc_in[74]
port 233 nsew signal input
rlabel metal2 s 369122 0 369178 800 6 gfpga_pad_io_soc_in[75]
port 234 nsew signal input
rlabel metal2 s 351734 0 351790 800 6 gfpga_pad_io_soc_in[76]
port 235 nsew signal input
rlabel metal2 s 334346 0 334402 800 6 gfpga_pad_io_soc_in[77]
port 236 nsew signal input
rlabel metal2 s 316958 0 317014 800 6 gfpga_pad_io_soc_in[78]
port 237 nsew signal input
rlabel metal2 s 299570 0 299626 800 6 gfpga_pad_io_soc_in[79]
port 238 nsew signal input
rlabel metal2 s 103150 542200 103206 543000 6 gfpga_pad_io_soc_in[7]
port 239 nsew signal input
rlabel metal2 s 282182 0 282238 800 6 gfpga_pad_io_soc_in[80]
port 240 nsew signal input
rlabel metal2 s 264794 0 264850 800 6 gfpga_pad_io_soc_in[81]
port 241 nsew signal input
rlabel metal2 s 247406 0 247462 800 6 gfpga_pad_io_soc_in[82]
port 242 nsew signal input
rlabel metal2 s 230018 0 230074 800 6 gfpga_pad_io_soc_in[83]
port 243 nsew signal input
rlabel metal2 s 212630 0 212686 800 6 gfpga_pad_io_soc_in[84]
port 244 nsew signal input
rlabel metal2 s 195242 0 195298 800 6 gfpga_pad_io_soc_in[85]
port 245 nsew signal input
rlabel metal2 s 177854 0 177910 800 6 gfpga_pad_io_soc_in[86]
port 246 nsew signal input
rlabel metal2 s 160466 0 160522 800 6 gfpga_pad_io_soc_in[87]
port 247 nsew signal input
rlabel metal2 s 143078 0 143134 800 6 gfpga_pad_io_soc_in[88]
port 248 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 gfpga_pad_io_soc_in[89]
port 249 nsew signal input
rlabel metal2 s 116674 542200 116730 543000 6 gfpga_pad_io_soc_in[8]
port 250 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 gfpga_pad_io_soc_in[90]
port 251 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 gfpga_pad_io_soc_in[91]
port 252 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 gfpga_pad_io_soc_in[92]
port 253 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 gfpga_pad_io_soc_in[93]
port 254 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 gfpga_pad_io_soc_in[94]
port 255 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 gfpga_pad_io_soc_in[95]
port 256 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 gfpga_pad_io_soc_in[96]
port 257 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 gfpga_pad_io_soc_in[97]
port 258 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 gfpga_pad_io_soc_in[98]
port 259 nsew signal input
rlabel metal3 s 0 70048 800 70168 6 gfpga_pad_io_soc_in[99]
port 260 nsew signal input
rlabel metal2 s 130198 542200 130254 543000 6 gfpga_pad_io_soc_in[9]
port 261 nsew signal input
rlabel metal2 s 8482 542200 8538 543000 6 gfpga_pad_io_soc_out[0]
port 262 nsew signal output
rlabel metal3 s 0 91808 800 91928 6 gfpga_pad_io_soc_out[100]
port 263 nsew signal output
rlabel metal3 s 0 108128 800 108248 6 gfpga_pad_io_soc_out[101]
port 264 nsew signal output
rlabel metal3 s 0 124448 800 124568 6 gfpga_pad_io_soc_out[102]
port 265 nsew signal output
rlabel metal3 s 0 140768 800 140888 6 gfpga_pad_io_soc_out[103]
port 266 nsew signal output
rlabel metal3 s 0 157088 800 157208 6 gfpga_pad_io_soc_out[104]
port 267 nsew signal output
rlabel metal3 s 0 173408 800 173528 6 gfpga_pad_io_soc_out[105]
port 268 nsew signal output
rlabel metal3 s 0 189728 800 189848 6 gfpga_pad_io_soc_out[106]
port 269 nsew signal output
rlabel metal3 s 0 206048 800 206168 6 gfpga_pad_io_soc_out[107]
port 270 nsew signal output
rlabel metal3 s 0 222368 800 222488 6 gfpga_pad_io_soc_out[108]
port 271 nsew signal output
rlabel metal3 s 0 238688 800 238808 6 gfpga_pad_io_soc_out[109]
port 272 nsew signal output
rlabel metal2 s 148230 542200 148286 543000 6 gfpga_pad_io_soc_out[10]
port 273 nsew signal output
rlabel metal3 s 0 255008 800 255128 6 gfpga_pad_io_soc_out[110]
port 274 nsew signal output
rlabel metal3 s 0 271328 800 271448 6 gfpga_pad_io_soc_out[111]
port 275 nsew signal output
rlabel metal3 s 0 287648 800 287768 6 gfpga_pad_io_soc_out[112]
port 276 nsew signal output
rlabel metal3 s 0 303968 800 304088 6 gfpga_pad_io_soc_out[113]
port 277 nsew signal output
rlabel metal3 s 0 320288 800 320408 6 gfpga_pad_io_soc_out[114]
port 278 nsew signal output
rlabel metal3 s 0 336608 800 336728 6 gfpga_pad_io_soc_out[115]
port 279 nsew signal output
rlabel metal3 s 0 352928 800 353048 6 gfpga_pad_io_soc_out[116]
port 280 nsew signal output
rlabel metal3 s 0 369248 800 369368 6 gfpga_pad_io_soc_out[117]
port 281 nsew signal output
rlabel metal3 s 0 385568 800 385688 6 gfpga_pad_io_soc_out[118]
port 282 nsew signal output
rlabel metal3 s 0 401888 800 402008 6 gfpga_pad_io_soc_out[119]
port 283 nsew signal output
rlabel metal2 s 161754 542200 161810 543000 6 gfpga_pad_io_soc_out[11]
port 284 nsew signal output
rlabel metal3 s 0 418208 800 418328 6 gfpga_pad_io_soc_out[120]
port 285 nsew signal output
rlabel metal3 s 0 434528 800 434648 6 gfpga_pad_io_soc_out[121]
port 286 nsew signal output
rlabel metal3 s 0 450848 800 450968 6 gfpga_pad_io_soc_out[122]
port 287 nsew signal output
rlabel metal3 s 0 467168 800 467288 6 gfpga_pad_io_soc_out[123]
port 288 nsew signal output
rlabel metal3 s 0 483488 800 483608 6 gfpga_pad_io_soc_out[124]
port 289 nsew signal output
rlabel metal3 s 0 499808 800 499928 6 gfpga_pad_io_soc_out[125]
port 290 nsew signal output
rlabel metal3 s 0 516128 800 516248 6 gfpga_pad_io_soc_out[126]
port 291 nsew signal output
rlabel metal3 s 0 532448 800 532568 6 gfpga_pad_io_soc_out[127]
port 292 nsew signal output
rlabel metal2 s 175278 542200 175334 543000 6 gfpga_pad_io_soc_out[12]
port 293 nsew signal output
rlabel metal2 s 188802 542200 188858 543000 6 gfpga_pad_io_soc_out[13]
port 294 nsew signal output
rlabel metal2 s 202326 542200 202382 543000 6 gfpga_pad_io_soc_out[14]
port 295 nsew signal output
rlabel metal2 s 215850 542200 215906 543000 6 gfpga_pad_io_soc_out[15]
port 296 nsew signal output
rlabel metal2 s 229374 542200 229430 543000 6 gfpga_pad_io_soc_out[16]
port 297 nsew signal output
rlabel metal2 s 242898 542200 242954 543000 6 gfpga_pad_io_soc_out[17]
port 298 nsew signal output
rlabel metal2 s 256422 542200 256478 543000 6 gfpga_pad_io_soc_out[18]
port 299 nsew signal output
rlabel metal2 s 269946 542200 270002 543000 6 gfpga_pad_io_soc_out[19]
port 300 nsew signal output
rlabel metal2 s 22006 542200 22062 543000 6 gfpga_pad_io_soc_out[1]
port 301 nsew signal output
rlabel metal2 s 283470 542200 283526 543000 6 gfpga_pad_io_soc_out[20]
port 302 nsew signal output
rlabel metal2 s 296994 542200 297050 543000 6 gfpga_pad_io_soc_out[21]
port 303 nsew signal output
rlabel metal2 s 310518 542200 310574 543000 6 gfpga_pad_io_soc_out[22]
port 304 nsew signal output
rlabel metal2 s 324042 542200 324098 543000 6 gfpga_pad_io_soc_out[23]
port 305 nsew signal output
rlabel metal2 s 337566 542200 337622 543000 6 gfpga_pad_io_soc_out[24]
port 306 nsew signal output
rlabel metal2 s 351090 542200 351146 543000 6 gfpga_pad_io_soc_out[25]
port 307 nsew signal output
rlabel metal2 s 364614 542200 364670 543000 6 gfpga_pad_io_soc_out[26]
port 308 nsew signal output
rlabel metal2 s 378138 542200 378194 543000 6 gfpga_pad_io_soc_out[27]
port 309 nsew signal output
rlabel metal2 s 391662 542200 391718 543000 6 gfpga_pad_io_soc_out[28]
port 310 nsew signal output
rlabel metal2 s 405186 542200 405242 543000 6 gfpga_pad_io_soc_out[29]
port 311 nsew signal output
rlabel metal2 s 35530 542200 35586 543000 6 gfpga_pad_io_soc_out[2]
port 312 nsew signal output
rlabel metal2 s 418710 542200 418766 543000 6 gfpga_pad_io_soc_out[30]
port 313 nsew signal output
rlabel metal2 s 432234 542200 432290 543000 6 gfpga_pad_io_soc_out[31]
port 314 nsew signal output
rlabel metal2 s 445758 542200 445814 543000 6 gfpga_pad_io_soc_out[32]
port 315 nsew signal output
rlabel metal2 s 459282 542200 459338 543000 6 gfpga_pad_io_soc_out[33]
port 316 nsew signal output
rlabel metal2 s 472806 542200 472862 543000 6 gfpga_pad_io_soc_out[34]
port 317 nsew signal output
rlabel metal2 s 486330 542200 486386 543000 6 gfpga_pad_io_soc_out[35]
port 318 nsew signal output
rlabel metal3 s 494200 525920 495000 526040 6 gfpga_pad_io_soc_out[36]
port 319 nsew signal output
rlabel metal3 s 494200 510008 495000 510128 6 gfpga_pad_io_soc_out[37]
port 320 nsew signal output
rlabel metal3 s 494200 494096 495000 494216 6 gfpga_pad_io_soc_out[38]
port 321 nsew signal output
rlabel metal3 s 494200 478184 495000 478304 6 gfpga_pad_io_soc_out[39]
port 322 nsew signal output
rlabel metal2 s 49054 542200 49110 543000 6 gfpga_pad_io_soc_out[3]
port 323 nsew signal output
rlabel metal3 s 494200 462272 495000 462392 6 gfpga_pad_io_soc_out[40]
port 324 nsew signal output
rlabel metal3 s 494200 446360 495000 446480 6 gfpga_pad_io_soc_out[41]
port 325 nsew signal output
rlabel metal3 s 494200 430448 495000 430568 6 gfpga_pad_io_soc_out[42]
port 326 nsew signal output
rlabel metal3 s 494200 414536 495000 414656 6 gfpga_pad_io_soc_out[43]
port 327 nsew signal output
rlabel metal3 s 494200 398624 495000 398744 6 gfpga_pad_io_soc_out[44]
port 328 nsew signal output
rlabel metal3 s 494200 382712 495000 382832 6 gfpga_pad_io_soc_out[45]
port 329 nsew signal output
rlabel metal3 s 494200 366800 495000 366920 6 gfpga_pad_io_soc_out[46]
port 330 nsew signal output
rlabel metal3 s 494200 350888 495000 351008 6 gfpga_pad_io_soc_out[47]
port 331 nsew signal output
rlabel metal3 s 494200 334976 495000 335096 6 gfpga_pad_io_soc_out[48]
port 332 nsew signal output
rlabel metal3 s 494200 319064 495000 319184 6 gfpga_pad_io_soc_out[49]
port 333 nsew signal output
rlabel metal2 s 67086 542200 67142 543000 6 gfpga_pad_io_soc_out[4]
port 334 nsew signal output
rlabel metal3 s 494200 303152 495000 303272 6 gfpga_pad_io_soc_out[50]
port 335 nsew signal output
rlabel metal3 s 494200 287240 495000 287360 6 gfpga_pad_io_soc_out[51]
port 336 nsew signal output
rlabel metal3 s 494200 271328 495000 271448 6 gfpga_pad_io_soc_out[52]
port 337 nsew signal output
rlabel metal3 s 494200 255416 495000 255536 6 gfpga_pad_io_soc_out[53]
port 338 nsew signal output
rlabel metal3 s 494200 239504 495000 239624 6 gfpga_pad_io_soc_out[54]
port 339 nsew signal output
rlabel metal3 s 494200 223592 495000 223712 6 gfpga_pad_io_soc_out[55]
port 340 nsew signal output
rlabel metal3 s 494200 207680 495000 207800 6 gfpga_pad_io_soc_out[56]
port 341 nsew signal output
rlabel metal3 s 494200 191768 495000 191888 6 gfpga_pad_io_soc_out[57]
port 342 nsew signal output
rlabel metal3 s 494200 175856 495000 175976 6 gfpga_pad_io_soc_out[58]
port 343 nsew signal output
rlabel metal3 s 494200 159944 495000 160064 6 gfpga_pad_io_soc_out[59]
port 344 nsew signal output
rlabel metal2 s 80610 542200 80666 543000 6 gfpga_pad_io_soc_out[5]
port 345 nsew signal output
rlabel metal3 s 494200 144032 495000 144152 6 gfpga_pad_io_soc_out[60]
port 346 nsew signal output
rlabel metal3 s 494200 128120 495000 128240 6 gfpga_pad_io_soc_out[61]
port 347 nsew signal output
rlabel metal3 s 494200 112208 495000 112328 6 gfpga_pad_io_soc_out[62]
port 348 nsew signal output
rlabel metal3 s 494200 96296 495000 96416 6 gfpga_pad_io_soc_out[63]
port 349 nsew signal output
rlabel metal3 s 494200 80384 495000 80504 6 gfpga_pad_io_soc_out[64]
port 350 nsew signal output
rlabel metal3 s 494200 64472 495000 64592 6 gfpga_pad_io_soc_out[65]
port 351 nsew signal output
rlabel metal3 s 494200 48560 495000 48680 6 gfpga_pad_io_soc_out[66]
port 352 nsew signal output
rlabel metal3 s 494200 32648 495000 32768 6 gfpga_pad_io_soc_out[67]
port 353 nsew signal output
rlabel metal2 s 485042 0 485098 800 6 gfpga_pad_io_soc_out[68]
port 354 nsew signal output
rlabel metal2 s 467654 0 467710 800 6 gfpga_pad_io_soc_out[69]
port 355 nsew signal output
rlabel metal2 s 94134 542200 94190 543000 6 gfpga_pad_io_soc_out[6]
port 356 nsew signal output
rlabel metal2 s 450266 0 450322 800 6 gfpga_pad_io_soc_out[70]
port 357 nsew signal output
rlabel metal2 s 432878 0 432934 800 6 gfpga_pad_io_soc_out[71]
port 358 nsew signal output
rlabel metal2 s 415490 0 415546 800 6 gfpga_pad_io_soc_out[72]
port 359 nsew signal output
rlabel metal2 s 398102 0 398158 800 6 gfpga_pad_io_soc_out[73]
port 360 nsew signal output
rlabel metal2 s 380714 0 380770 800 6 gfpga_pad_io_soc_out[74]
port 361 nsew signal output
rlabel metal2 s 363326 0 363382 800 6 gfpga_pad_io_soc_out[75]
port 362 nsew signal output
rlabel metal2 s 345938 0 345994 800 6 gfpga_pad_io_soc_out[76]
port 363 nsew signal output
rlabel metal2 s 328550 0 328606 800 6 gfpga_pad_io_soc_out[77]
port 364 nsew signal output
rlabel metal2 s 311162 0 311218 800 6 gfpga_pad_io_soc_out[78]
port 365 nsew signal output
rlabel metal2 s 293774 0 293830 800 6 gfpga_pad_io_soc_out[79]
port 366 nsew signal output
rlabel metal2 s 107658 542200 107714 543000 6 gfpga_pad_io_soc_out[7]
port 367 nsew signal output
rlabel metal2 s 276386 0 276442 800 6 gfpga_pad_io_soc_out[80]
port 368 nsew signal output
rlabel metal2 s 258998 0 259054 800 6 gfpga_pad_io_soc_out[81]
port 369 nsew signal output
rlabel metal2 s 241610 0 241666 800 6 gfpga_pad_io_soc_out[82]
port 370 nsew signal output
rlabel metal2 s 224222 0 224278 800 6 gfpga_pad_io_soc_out[83]
port 371 nsew signal output
rlabel metal2 s 206834 0 206890 800 6 gfpga_pad_io_soc_out[84]
port 372 nsew signal output
rlabel metal2 s 189446 0 189502 800 6 gfpga_pad_io_soc_out[85]
port 373 nsew signal output
rlabel metal2 s 172058 0 172114 800 6 gfpga_pad_io_soc_out[86]
port 374 nsew signal output
rlabel metal2 s 154670 0 154726 800 6 gfpga_pad_io_soc_out[87]
port 375 nsew signal output
rlabel metal2 s 137282 0 137338 800 6 gfpga_pad_io_soc_out[88]
port 376 nsew signal output
rlabel metal2 s 119894 0 119950 800 6 gfpga_pad_io_soc_out[89]
port 377 nsew signal output
rlabel metal2 s 121182 542200 121238 543000 6 gfpga_pad_io_soc_out[8]
port 378 nsew signal output
rlabel metal2 s 102506 0 102562 800 6 gfpga_pad_io_soc_out[90]
port 379 nsew signal output
rlabel metal2 s 85118 0 85174 800 6 gfpga_pad_io_soc_out[91]
port 380 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 gfpga_pad_io_soc_out[92]
port 381 nsew signal output
rlabel metal2 s 44546 0 44602 800 6 gfpga_pad_io_soc_out[93]
port 382 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 gfpga_pad_io_soc_out[94]
port 383 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 gfpga_pad_io_soc_out[95]
port 384 nsew signal output
rlabel metal3 s 0 26528 800 26648 6 gfpga_pad_io_soc_out[96]
port 385 nsew signal output
rlabel metal3 s 0 42848 800 42968 6 gfpga_pad_io_soc_out[97]
port 386 nsew signal output
rlabel metal3 s 0 59168 800 59288 6 gfpga_pad_io_soc_out[98]
port 387 nsew signal output
rlabel metal3 s 0 75488 800 75608 6 gfpga_pad_io_soc_out[99]
port 388 nsew signal output
rlabel metal2 s 134706 542200 134762 543000 6 gfpga_pad_io_soc_out[9]
port 389 nsew signal output
rlabel metal3 s 494200 11432 495000 11552 6 isol_n
port 390 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 prog_clk
port 391 nsew signal input
rlabel metal3 s 494200 16736 495000 16856 6 prog_reset
port 392 nsew signal input
rlabel metal3 s 494200 22040 495000 22160 6 reset
port 393 nsew signal input
rlabel metal2 s 58070 542200 58126 543000 6 sc_head
port 394 nsew signal input
rlabel metal3 s 494200 536528 495000 536648 6 sc_tail
port 395 nsew signal output
rlabel metal3 s 494200 6128 495000 6248 6 test_enable
port 396 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 495000 543000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 82835136
string GDS_FILE /home/hosni/OpenFPGA/clear/openlane/fpga_core/runs/23_03_20_17_16/results/signoff/fpga_core.magic.gds
string GDS_START 36294118
<< end >>

