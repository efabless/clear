magic
tech sky130A
magscale 1 2
timestamp 1625783076
<< locali >>
rect 6285 16031 6319 16201
rect 9137 15351 9171 15521
rect 16129 14535 16163 15113
rect 9505 13243 9539 13413
rect 9597 10455 9631 10557
rect 9597 8347 9631 8585
rect 6653 6171 6687 6273
<< viali >>
rect 1869 17289 1903 17323
rect 4445 17289 4479 17323
rect 7573 17289 7607 17323
rect 7941 17289 7975 17323
rect 13277 17289 13311 17323
rect 14013 17289 14047 17323
rect 15025 17289 15059 17323
rect 1409 17221 1443 17255
rect 2145 17221 2179 17255
rect 2881 17221 2915 17255
rect 4629 17221 4663 17255
rect 5089 17221 5123 17255
rect 5457 17221 5491 17255
rect 5917 17221 5951 17255
rect 6561 17221 6595 17255
rect 6929 17221 6963 17255
rect 8309 17221 8343 17255
rect 13553 17221 13587 17255
rect 14565 17221 14599 17255
rect 2513 17153 2547 17187
rect 3709 17153 3743 17187
rect 7389 17153 7423 17187
rect 13001 17153 13035 17187
rect 15577 17153 15611 17187
rect 3985 17085 4019 17119
rect 4169 17085 4203 17119
rect 8493 17085 8527 17119
rect 8953 17085 8987 17119
rect 9229 17085 9263 17119
rect 9413 17085 9447 17119
rect 9680 17085 9714 17119
rect 11345 17085 11379 17119
rect 13737 17085 13771 17119
rect 14289 17085 14323 17119
rect 14933 17085 14967 17119
rect 1593 17017 1627 17051
rect 1961 17017 1995 17051
rect 2329 17017 2363 17051
rect 2697 17017 2731 17051
rect 3065 17017 3099 17051
rect 3525 17017 3559 17051
rect 4353 17017 4387 17051
rect 4813 17017 4847 17051
rect 5273 17017 5307 17051
rect 5641 17017 5675 17051
rect 6101 17017 6135 17051
rect 6745 17017 6779 17051
rect 7113 17017 7147 17051
rect 7665 17017 7699 17051
rect 8033 17017 8067 17051
rect 10977 17017 11011 17051
rect 11621 17017 11655 17051
rect 12173 17017 12207 17051
rect 13369 17017 13403 17051
rect 14105 17017 14139 17051
rect 14749 17017 14783 17051
rect 6377 16949 6411 16983
rect 8677 16949 8711 16983
rect 10793 16949 10827 16983
rect 11529 16949 11563 16983
rect 12081 16949 12115 16983
rect 12357 16949 12391 16983
rect 12725 16949 12759 16983
rect 12817 16949 12851 16983
rect 15393 16949 15427 16983
rect 1869 16745 1903 16779
rect 2145 16745 2179 16779
rect 4629 16745 4663 16779
rect 5089 16745 5123 16779
rect 8493 16745 8527 16779
rect 8769 16745 8803 16779
rect 11437 16745 11471 16779
rect 12725 16745 12759 16779
rect 14473 16745 14507 16779
rect 15669 16745 15703 16779
rect 1409 16677 1443 16711
rect 2605 16677 2639 16711
rect 3065 16677 3099 16711
rect 3433 16677 3467 16711
rect 3893 16677 3927 16711
rect 4261 16677 4295 16711
rect 4445 16677 4479 16711
rect 5610 16677 5644 16711
rect 7082 16677 7116 16711
rect 11529 16677 11563 16711
rect 12357 16677 12391 16711
rect 1593 16609 1627 16643
rect 1961 16609 1995 16643
rect 2329 16609 2363 16643
rect 2789 16609 2823 16643
rect 3249 16609 3283 16643
rect 3617 16609 3651 16643
rect 4077 16609 4111 16643
rect 4813 16609 4847 16643
rect 4997 16609 5031 16643
rect 5273 16609 5307 16643
rect 8585 16609 8619 16643
rect 8953 16609 8987 16643
rect 9393 16609 9427 16643
rect 10609 16609 10643 16643
rect 12265 16609 12299 16643
rect 13838 16609 13872 16643
rect 14565 16609 14599 16643
rect 14749 16609 14783 16643
rect 14933 16609 14967 16643
rect 15485 16609 15519 16643
rect 5365 16541 5399 16575
rect 6837 16541 6871 16575
rect 9137 16541 9171 16575
rect 11621 16541 11655 16575
rect 12449 16541 12483 16575
rect 14105 16541 14139 16575
rect 6745 16473 6779 16507
rect 8217 16473 8251 16507
rect 2421 16405 2455 16439
rect 10517 16405 10551 16439
rect 10793 16405 10827 16439
rect 11069 16405 11103 16439
rect 11897 16405 11931 16439
rect 15209 16405 15243 16439
rect 2421 16201 2455 16235
rect 2881 16201 2915 16235
rect 3157 16201 3191 16235
rect 3617 16201 3651 16235
rect 3893 16201 3927 16235
rect 4077 16201 4111 16235
rect 4721 16201 4755 16235
rect 5641 16201 5675 16235
rect 6009 16201 6043 16235
rect 6285 16201 6319 16235
rect 7297 16201 7331 16235
rect 7573 16201 7607 16235
rect 7849 16201 7883 16235
rect 8493 16201 8527 16235
rect 9597 16201 9631 16235
rect 13645 16201 13679 16235
rect 1409 16133 1443 16167
rect 5917 16133 5951 16167
rect 4353 16065 4387 16099
rect 8217 16133 8251 16167
rect 7021 16065 7055 16099
rect 8861 16065 8895 16099
rect 9873 16065 9907 16099
rect 10149 16065 10183 16099
rect 10885 16065 10919 16099
rect 11069 16065 11103 16099
rect 1961 15997 1995 16031
rect 2237 15997 2271 16031
rect 2513 15997 2547 16031
rect 3065 15997 3099 16031
rect 3341 15997 3375 16031
rect 3433 15997 3467 16031
rect 3709 15997 3743 16031
rect 4537 15997 4571 16031
rect 4905 15997 4939 16031
rect 5457 15997 5491 16031
rect 5733 15997 5767 16031
rect 6193 15997 6227 16031
rect 6285 15997 6319 16031
rect 7481 15997 7515 16031
rect 7757 15997 7791 16031
rect 8033 15997 8067 16031
rect 8309 15997 8343 16031
rect 11161 15997 11195 16031
rect 11897 15997 11931 16031
rect 12173 15997 12207 16031
rect 13829 15997 13863 16031
rect 14085 15997 14119 16031
rect 15485 15997 15519 16031
rect 1593 15929 1627 15963
rect 6837 15929 6871 15963
rect 8953 15929 8987 15963
rect 10241 15929 10275 15963
rect 12440 15929 12474 15963
rect 15301 15929 15335 15963
rect 1777 15861 1811 15895
rect 2145 15861 2179 15895
rect 2697 15861 2731 15895
rect 4261 15861 4295 15895
rect 5089 15861 5123 15895
rect 5365 15861 5399 15895
rect 6469 15861 6503 15895
rect 6929 15861 6963 15895
rect 9045 15861 9079 15895
rect 9413 15861 9447 15895
rect 10333 15861 10367 15895
rect 10701 15861 10735 15895
rect 11529 15861 11563 15895
rect 11805 15861 11839 15895
rect 13553 15861 13587 15895
rect 15209 15861 15243 15895
rect 1501 15657 1535 15691
rect 1777 15657 1811 15691
rect 2329 15657 2363 15691
rect 7205 15657 7239 15691
rect 7297 15657 7331 15691
rect 8125 15657 8159 15691
rect 9505 15657 9539 15691
rect 9965 15657 9999 15691
rect 10333 15657 10367 15691
rect 10793 15657 10827 15691
rect 11161 15657 11195 15691
rect 11529 15657 11563 15691
rect 12909 15657 12943 15691
rect 13369 15657 13403 15691
rect 14657 15657 14691 15691
rect 1593 15589 1627 15623
rect 3341 15589 3375 15623
rect 11621 15589 11655 15623
rect 15485 15589 15519 15623
rect 1961 15521 1995 15555
rect 2237 15521 2271 15555
rect 2513 15521 2547 15555
rect 2605 15521 2639 15555
rect 2881 15521 2915 15555
rect 5937 15521 5971 15555
rect 6193 15521 6227 15555
rect 6377 15521 6411 15555
rect 6837 15521 6871 15555
rect 7665 15521 7699 15555
rect 8769 15521 8803 15555
rect 9137 15521 9171 15555
rect 9597 15521 9631 15555
rect 10701 15521 10735 15555
rect 12541 15521 12575 15555
rect 14013 15521 14047 15555
rect 14749 15521 14783 15555
rect 3157 15453 3191 15487
rect 6561 15453 6595 15487
rect 6745 15453 6779 15487
rect 7757 15453 7791 15487
rect 7849 15453 7883 15487
rect 8493 15453 8527 15487
rect 2053 15385 2087 15419
rect 4721 15385 4755 15419
rect 9413 15453 9447 15487
rect 10885 15453 10919 15487
rect 11713 15453 11747 15487
rect 12357 15453 12391 15487
rect 12449 15453 12483 15487
rect 13461 15453 13495 15487
rect 13645 15453 13679 15487
rect 14473 15453 14507 15487
rect 15301 15453 15335 15487
rect 13001 15385 13035 15419
rect 2789 15317 2823 15351
rect 3065 15317 3099 15351
rect 3617 15317 3651 15351
rect 4813 15317 4847 15351
rect 8585 15317 8619 15351
rect 9137 15317 9171 15351
rect 10241 15317 10275 15351
rect 12081 15317 12115 15351
rect 13921 15317 13955 15351
rect 15117 15317 15151 15351
rect 1961 15113 1995 15147
rect 6745 15113 6779 15147
rect 7757 15113 7791 15147
rect 8585 15113 8619 15147
rect 9873 15113 9907 15147
rect 11345 15113 11379 15147
rect 12909 15113 12943 15147
rect 13001 15113 13035 15147
rect 14013 15113 14047 15147
rect 14933 15113 14967 15147
rect 16129 15113 16163 15147
rect 3341 15045 3375 15079
rect 5825 15045 5859 15079
rect 7665 15045 7699 15079
rect 11529 15045 11563 15079
rect 2789 14977 2823 15011
rect 3157 14977 3191 15011
rect 3893 14977 3927 15011
rect 4445 14977 4479 15011
rect 7297 14977 7331 15011
rect 8309 14977 8343 15011
rect 9137 14977 9171 15011
rect 9965 14977 9999 15011
rect 12357 14977 12391 15011
rect 13553 14977 13587 15011
rect 14197 14977 14231 15011
rect 14381 14977 14415 15011
rect 15393 14977 15427 15011
rect 15485 14977 15519 15011
rect 1777 14909 1811 14943
rect 6285 14909 6319 14943
rect 7113 14909 7147 14943
rect 8125 14909 8159 14943
rect 8953 14909 8987 14943
rect 9045 14909 9079 14943
rect 9689 14909 9723 14943
rect 10232 14909 10266 14943
rect 11897 14909 11931 14943
rect 12541 14909 12575 14943
rect 13461 14909 13495 14943
rect 1593 14841 1627 14875
rect 2513 14841 2547 14875
rect 4690 14841 4724 14875
rect 6101 14841 6135 14875
rect 15301 14841 15335 14875
rect 1501 14773 1535 14807
rect 2145 14773 2179 14807
rect 2605 14773 2639 14807
rect 3065 14773 3099 14807
rect 3709 14773 3743 14807
rect 3801 14773 3835 14807
rect 6561 14773 6595 14807
rect 7205 14773 7239 14807
rect 8217 14773 8251 14807
rect 9505 14773 9539 14807
rect 11805 14773 11839 14807
rect 12449 14773 12483 14807
rect 13369 14773 13403 14807
rect 14473 14773 14507 14807
rect 14841 14773 14875 14807
rect 1593 14569 1627 14603
rect 1961 14569 1995 14603
rect 5365 14569 5399 14603
rect 6377 14569 6411 14603
rect 6837 14569 6871 14603
rect 7297 14569 7331 14603
rect 7665 14569 7699 14603
rect 8033 14569 8067 14603
rect 8769 14569 8803 14603
rect 10057 14569 10091 14603
rect 10425 14569 10459 14603
rect 14197 14569 14231 14603
rect 14565 14569 14599 14603
rect 4138 14501 4172 14535
rect 5825 14501 5859 14535
rect 6469 14501 6503 14535
rect 11244 14501 11278 14535
rect 12633 14501 12667 14535
rect 14841 14501 14875 14535
rect 15117 14501 15151 14535
rect 15301 14501 15335 14535
rect 16129 14501 16163 14535
rect 1501 14433 1535 14467
rect 1777 14433 1811 14467
rect 3085 14433 3119 14467
rect 5733 14433 5767 14467
rect 6193 14433 6227 14467
rect 7205 14433 7239 14467
rect 9597 14433 9631 14467
rect 10701 14433 10735 14467
rect 10977 14433 11011 14467
rect 12817 14433 12851 14467
rect 13084 14433 13118 14467
rect 15577 14433 15611 14467
rect 3341 14365 3375 14399
rect 3893 14365 3927 14399
rect 5917 14365 5951 14399
rect 6653 14365 6687 14399
rect 7389 14365 7423 14399
rect 8125 14365 8159 14399
rect 8309 14365 8343 14399
rect 8953 14365 8987 14399
rect 9689 14365 9723 14399
rect 9873 14365 9907 14399
rect 10333 14365 10367 14399
rect 14473 14365 14507 14399
rect 5273 14297 5307 14331
rect 9229 14297 9263 14331
rect 12357 14297 12391 14331
rect 15393 14297 15427 14331
rect 8493 14229 8527 14263
rect 10885 14229 10919 14263
rect 12541 14229 12575 14263
rect 1777 14025 1811 14059
rect 2145 14025 2179 14059
rect 4077 14025 4111 14059
rect 5273 14025 5307 14059
rect 7021 14025 7055 14059
rect 9965 14025 9999 14059
rect 11713 14025 11747 14059
rect 13369 14025 13403 14059
rect 14289 14025 14323 14059
rect 5365 13957 5399 13991
rect 9873 13957 9907 13991
rect 11437 13957 11471 13991
rect 13461 13957 13495 13991
rect 2789 13889 2823 13923
rect 3617 13889 3651 13923
rect 4721 13889 4755 13923
rect 5917 13889 5951 13923
rect 12265 13889 12299 13923
rect 12817 13889 12851 13923
rect 14013 13889 14047 13923
rect 14565 13889 14599 13923
rect 1409 13821 1443 13855
rect 1961 13821 1995 13855
rect 5733 13821 5767 13855
rect 6561 13821 6595 13855
rect 8145 13821 8179 13855
rect 8401 13821 8435 13855
rect 8493 13821 8527 13855
rect 8760 13821 8794 13855
rect 11078 13821 11112 13855
rect 11345 13821 11379 13855
rect 12173 13821 12207 13855
rect 13829 13821 13863 13855
rect 1593 13753 1627 13787
rect 2513 13753 2547 13787
rect 3341 13753 3375 13787
rect 4445 13753 4479 13787
rect 5089 13753 5123 13787
rect 12909 13753 12943 13787
rect 13921 13753 13955 13787
rect 15485 13753 15519 13787
rect 15577 13753 15611 13787
rect 2605 13685 2639 13719
rect 2973 13685 3007 13719
rect 3433 13685 3467 13719
rect 3893 13685 3927 13719
rect 4537 13685 4571 13719
rect 5825 13685 5859 13719
rect 6745 13685 6779 13719
rect 12081 13685 12115 13719
rect 13001 13685 13035 13719
rect 2697 13481 2731 13515
rect 3065 13481 3099 13515
rect 3985 13481 4019 13515
rect 5457 13481 5491 13515
rect 7665 13481 7699 13515
rect 8677 13481 8711 13515
rect 8953 13481 8987 13515
rect 9597 13481 9631 13515
rect 10425 13481 10459 13515
rect 12173 13481 12207 13515
rect 13553 13481 13587 13515
rect 13921 13481 13955 13515
rect 14657 13481 14691 13515
rect 15071 13481 15105 13515
rect 15393 13481 15427 13515
rect 15485 13481 15519 13515
rect 3525 13413 3559 13447
rect 5917 13413 5951 13447
rect 7849 13413 7883 13447
rect 9505 13413 9539 13447
rect 9965 13413 9999 13447
rect 11538 13413 11572 13447
rect 12633 13413 12667 13447
rect 14105 13413 14139 13447
rect 14381 13413 14415 13447
rect 1685 13345 1719 13379
rect 5825 13345 5859 13379
rect 6541 13345 6575 13379
rect 3157 13277 3191 13311
rect 3341 13277 3375 13311
rect 6101 13277 6135 13311
rect 6285 13277 6319 13311
rect 12541 13345 12575 13379
rect 15000 13345 15034 13379
rect 15669 13345 15703 13379
rect 10057 13277 10091 13311
rect 10241 13277 10275 13311
rect 11805 13277 11839 13311
rect 12725 13277 12759 13311
rect 13001 13277 13035 13311
rect 13185 13277 13219 13311
rect 13461 13277 13495 13311
rect 5181 13209 5215 13243
rect 9505 13209 9539 13243
rect 1501 13141 1535 13175
rect 7941 13141 7975 13175
rect 11989 13141 12023 13175
rect 13829 13141 13863 13175
rect 14749 13141 14783 13175
rect 1777 12937 1811 12971
rect 3249 12937 3283 12971
rect 4721 12937 4755 12971
rect 6469 12937 6503 12971
rect 8401 12937 8435 12971
rect 9781 12937 9815 12971
rect 11713 12937 11747 12971
rect 14381 12937 14415 12971
rect 15669 12937 15703 12971
rect 1409 12869 1443 12903
rect 8125 12869 8159 12903
rect 12541 12869 12575 12903
rect 14197 12869 14231 12903
rect 2697 12801 2731 12835
rect 5457 12801 5491 12835
rect 6009 12801 6043 12835
rect 6193 12801 6227 12835
rect 7021 12801 7055 12835
rect 7849 12801 7883 12835
rect 10425 12801 10459 12835
rect 10885 12801 10919 12835
rect 12265 12801 12299 12835
rect 13093 12801 13127 12835
rect 13369 12801 13403 12835
rect 15301 12801 15335 12835
rect 1593 12733 1627 12767
rect 1961 12733 1995 12767
rect 3341 12733 3375 12767
rect 5917 12733 5951 12767
rect 8309 12733 8343 12767
rect 9505 12733 9539 12767
rect 10977 12733 11011 12767
rect 12081 12733 12115 12767
rect 13645 12733 13679 12767
rect 14933 12733 14967 12767
rect 15025 12733 15059 12767
rect 3586 12665 3620 12699
rect 6837 12665 6871 12699
rect 7757 12665 7791 12699
rect 8585 12665 8619 12699
rect 12909 12665 12943 12699
rect 13829 12665 13863 12699
rect 14105 12665 14139 12699
rect 2789 12597 2823 12631
rect 2881 12597 2915 12631
rect 5549 12597 5583 12631
rect 6929 12597 6963 12631
rect 7297 12597 7331 12631
rect 7665 12597 7699 12631
rect 9689 12597 9723 12631
rect 10149 12597 10183 12631
rect 10241 12597 10275 12631
rect 11069 12597 11103 12631
rect 11437 12597 11471 12631
rect 12173 12597 12207 12631
rect 13001 12597 13035 12631
rect 1777 12393 1811 12427
rect 3433 12393 3467 12427
rect 3985 12393 4019 12427
rect 4813 12393 4847 12427
rect 4905 12393 4939 12427
rect 5365 12393 5399 12427
rect 5825 12393 5859 12427
rect 6745 12393 6779 12427
rect 8953 12393 8987 12427
rect 10609 12393 10643 12427
rect 12633 12393 12667 12427
rect 1593 12325 1627 12359
rect 7542 12325 7576 12359
rect 1961 12257 1995 12291
rect 2053 12257 2087 12291
rect 2320 12257 2354 12291
rect 5733 12257 5767 12291
rect 6837 12257 6871 12291
rect 8769 12257 8803 12291
rect 9393 12257 9427 12291
rect 11520 12257 11554 12291
rect 12909 12257 12943 12291
rect 13829 12257 13863 12291
rect 4721 12189 4755 12223
rect 6009 12189 6043 12223
rect 6653 12189 6687 12223
rect 7297 12189 7331 12223
rect 9137 12189 9171 12223
rect 11253 12189 11287 12223
rect 13185 12189 13219 12223
rect 10517 12121 10551 12155
rect 1501 12053 1535 12087
rect 3617 12053 3651 12087
rect 5273 12053 5307 12087
rect 6285 12053 6319 12087
rect 7205 12053 7239 12087
rect 8677 12053 8711 12087
rect 10885 12053 10919 12087
rect 11069 12053 11103 12087
rect 3801 11849 3835 11883
rect 4721 11849 4755 11883
rect 9781 11849 9815 11883
rect 9965 11849 9999 11883
rect 5549 11781 5583 11815
rect 10793 11781 10827 11815
rect 11897 11781 11931 11815
rect 4445 11713 4479 11747
rect 5181 11713 5215 11747
rect 5365 11713 5399 11747
rect 6469 11713 6503 11747
rect 8493 11713 8527 11747
rect 10425 11713 10459 11747
rect 10609 11713 10643 11747
rect 11345 11713 11379 11747
rect 2533 11645 2567 11679
rect 2789 11645 2823 11679
rect 5733 11645 5767 11679
rect 8401 11645 8435 11679
rect 11713 11645 11747 11679
rect 6714 11577 6748 11611
rect 11253 11577 11287 11611
rect 11989 11577 12023 11611
rect 1409 11509 1443 11543
rect 3525 11509 3559 11543
rect 3893 11509 3927 11543
rect 4261 11509 4295 11543
rect 4353 11509 4387 11543
rect 5089 11509 5123 11543
rect 7849 11509 7883 11543
rect 7941 11509 7975 11543
rect 8309 11509 8343 11543
rect 8769 11509 8803 11543
rect 9597 11509 9631 11543
rect 10333 11509 10367 11543
rect 11161 11509 11195 11543
rect 12173 11509 12207 11543
rect 12449 11509 12483 11543
rect 1869 11305 1903 11339
rect 2237 11305 2271 11339
rect 5365 11305 5399 11339
rect 6745 11305 6779 11339
rect 7113 11305 7147 11339
rect 7205 11305 7239 11339
rect 7665 11305 7699 11339
rect 9781 11305 9815 11339
rect 10241 11305 10275 11339
rect 3249 11237 3283 11271
rect 5028 11237 5062 11271
rect 1593 11169 1627 11203
rect 5273 11169 5307 11203
rect 5733 11169 5767 11203
rect 8309 11169 8343 11203
rect 9321 11169 9355 11203
rect 12745 11169 12779 11203
rect 2329 11101 2363 11135
rect 2421 11101 2455 11135
rect 3341 11101 3375 11135
rect 3525 11101 3559 11135
rect 5825 11101 5859 11135
rect 6009 11101 6043 11135
rect 6285 11101 6319 11135
rect 7389 11101 7423 11135
rect 8401 11101 8435 11135
rect 8585 11101 8619 11135
rect 9505 11101 9539 11135
rect 9689 11101 9723 11135
rect 13001 11101 13035 11135
rect 1409 11033 1443 11067
rect 3893 11033 3927 11067
rect 8861 11033 8895 11067
rect 10149 11033 10183 11067
rect 2881 10965 2915 10999
rect 7941 10965 7975 10999
rect 11621 10965 11655 10999
rect 1501 10761 1535 10795
rect 2053 10761 2087 10795
rect 3985 10761 4019 10795
rect 5457 10761 5491 10795
rect 7665 10761 7699 10795
rect 10701 10761 10735 10795
rect 14197 10761 14231 10795
rect 2697 10625 2731 10659
rect 3525 10625 3559 10659
rect 6009 10625 6043 10659
rect 7113 10625 7147 10659
rect 9137 10625 9171 10659
rect 9781 10625 9815 10659
rect 10333 10625 10367 10659
rect 10517 10625 10551 10659
rect 11253 10625 11287 10659
rect 12265 10625 12299 10659
rect 12817 10625 12851 10659
rect 1685 10557 1719 10591
rect 2421 10557 2455 10591
rect 5365 10557 5399 10591
rect 7297 10557 7331 10591
rect 8870 10557 8904 10591
rect 9229 10557 9263 10591
rect 9505 10557 9539 10591
rect 9597 10557 9631 10591
rect 3249 10489 3283 10523
rect 3709 10489 3743 10523
rect 5120 10489 5154 10523
rect 5917 10489 5951 10523
rect 11161 10489 11195 10523
rect 12081 10489 12115 10523
rect 13084 10489 13118 10523
rect 2513 10421 2547 10455
rect 2881 10421 2915 10455
rect 3341 10421 3375 10455
rect 5825 10421 5859 10455
rect 6561 10421 6595 10455
rect 7205 10421 7239 10455
rect 7757 10421 7791 10455
rect 9597 10421 9631 10455
rect 9873 10421 9907 10455
rect 10241 10421 10275 10455
rect 11069 10421 11103 10455
rect 11713 10421 11747 10455
rect 12173 10421 12207 10455
rect 12633 10421 12667 10455
rect 14473 10421 14507 10455
rect 14657 10421 14691 10455
rect 1777 10217 1811 10251
rect 3893 10217 3927 10251
rect 5457 10217 5491 10251
rect 7941 10217 7975 10251
rect 8401 10217 8435 10251
rect 8769 10217 8803 10251
rect 9505 10217 9539 10251
rect 14749 10217 14783 10251
rect 15209 10217 15243 10251
rect 1593 10149 1627 10183
rect 11170 10149 11204 10183
rect 12642 10149 12676 10183
rect 13645 10149 13679 10183
rect 15485 10149 15519 10183
rect 1961 10081 1995 10115
rect 4261 10081 4295 10115
rect 5825 10081 5859 10115
rect 6092 10081 6126 10115
rect 8309 10081 8343 10115
rect 9597 10081 9631 10115
rect 11437 10081 11471 10115
rect 12909 10081 12943 10115
rect 13737 10081 13771 10115
rect 4353 10013 4387 10047
rect 4537 10013 4571 10047
rect 8585 10013 8619 10047
rect 9413 10013 9447 10047
rect 13461 10013 13495 10047
rect 14841 10013 14875 10047
rect 14933 10013 14967 10047
rect 1409 9945 1443 9979
rect 4813 9945 4847 9979
rect 7205 9945 7239 9979
rect 9965 9945 9999 9979
rect 11529 9945 11563 9979
rect 15669 9945 15703 9979
rect 4997 9877 5031 9911
rect 10057 9877 10091 9911
rect 13001 9877 13035 9911
rect 14105 9877 14139 9911
rect 14381 9877 14415 9911
rect 6469 9673 6503 9707
rect 8493 9605 8527 9639
rect 9965 9605 9999 9639
rect 13001 9605 13035 9639
rect 4261 9537 4295 9571
rect 5181 9537 5215 9571
rect 5917 9537 5951 9571
rect 10517 9537 10551 9571
rect 12357 9537 12391 9571
rect 13645 9537 13679 9571
rect 14289 9537 14323 9571
rect 14381 9537 14415 9571
rect 4997 9469 5031 9503
rect 5825 9469 5859 9503
rect 7849 9469 7883 9503
rect 9781 9469 9815 9503
rect 14197 9469 14231 9503
rect 4077 9401 4111 9435
rect 7582 9401 7616 9435
rect 10793 9401 10827 9435
rect 12541 9401 12575 9435
rect 13369 9401 13403 9435
rect 3709 9333 3743 9367
rect 4169 9333 4203 9367
rect 4537 9333 4571 9367
rect 4905 9333 4939 9367
rect 5365 9333 5399 9367
rect 5733 9333 5767 9367
rect 6193 9333 6227 9367
rect 10333 9333 10367 9367
rect 10425 9333 10459 9367
rect 10977 9333 11011 9367
rect 11253 9333 11287 9367
rect 12449 9333 12483 9367
rect 12909 9333 12943 9367
rect 13461 9333 13495 9367
rect 13829 9333 13863 9367
rect 3341 9129 3375 9163
rect 5273 9129 5307 9163
rect 7205 9129 7239 9163
rect 9505 9129 9539 9163
rect 9965 9129 9999 9163
rect 10333 9129 10367 9163
rect 10425 9129 10459 9163
rect 1409 9061 1443 9095
rect 5610 9061 5644 9095
rect 1593 8993 1627 9027
rect 4160 8993 4194 9027
rect 8217 8993 8251 9027
rect 8953 8993 8987 9027
rect 9597 8993 9631 9027
rect 11060 8993 11094 9027
rect 12909 8993 12943 9027
rect 13369 8993 13403 9027
rect 3433 8925 3467 8959
rect 3617 8925 3651 8959
rect 3893 8925 3927 8959
rect 5365 8925 5399 8959
rect 6929 8925 6963 8959
rect 7113 8925 7147 8959
rect 7941 8925 7975 8959
rect 8125 8925 8159 8959
rect 8769 8925 8803 8959
rect 9689 8925 9723 8959
rect 10517 8925 10551 8959
rect 10793 8925 10827 8959
rect 12633 8925 12667 8959
rect 12817 8925 12851 8959
rect 6745 8857 6779 8891
rect 8585 8857 8619 8891
rect 2973 8789 3007 8823
rect 7573 8789 7607 8823
rect 7757 8789 7791 8823
rect 9137 8789 9171 8823
rect 12173 8789 12207 8823
rect 12449 8789 12483 8823
rect 13277 8789 13311 8823
rect 1593 8585 1627 8619
rect 3985 8585 4019 8619
rect 8493 8585 8527 8619
rect 9597 8585 9631 8619
rect 11345 8585 11379 8619
rect 11897 8585 11931 8619
rect 14289 8585 14323 8619
rect 5089 8517 5123 8551
rect 6285 8517 6319 8551
rect 4445 8449 4479 8483
rect 4537 8449 4571 8483
rect 5641 8449 5675 8483
rect 5917 8449 5951 8483
rect 6469 8449 6503 8483
rect 9137 8449 9171 8483
rect 1777 8381 1811 8415
rect 2513 8381 2547 8415
rect 2780 8381 2814 8415
rect 6736 8381 6770 8415
rect 7941 8381 7975 8415
rect 8125 8381 8159 8415
rect 8309 8381 8343 8415
rect 8861 8381 8895 8415
rect 12173 8449 12207 8483
rect 9689 8381 9723 8415
rect 9965 8381 9999 8415
rect 12357 8381 12391 8415
rect 12909 8381 12943 8415
rect 13165 8381 13199 8415
rect 5457 8313 5491 8347
rect 8953 8313 8987 8347
rect 9597 8313 9631 8347
rect 10232 8313 10266 8347
rect 12449 8313 12483 8347
rect 3893 8245 3927 8279
rect 4353 8245 4387 8279
rect 4997 8245 5031 8279
rect 5549 8245 5583 8279
rect 7849 8245 7883 8279
rect 9505 8245 9539 8279
rect 9873 8245 9907 8279
rect 11805 8245 11839 8279
rect 12817 8245 12851 8279
rect 1501 8041 1535 8075
rect 1777 8041 1811 8075
rect 4077 8041 4111 8075
rect 4445 8041 4479 8075
rect 5181 8041 5215 8075
rect 7297 8041 7331 8075
rect 7757 8041 7791 8075
rect 8585 8041 8619 8075
rect 9137 8041 9171 8075
rect 9505 8041 9539 8075
rect 10885 8041 10919 8075
rect 11437 8041 11471 8075
rect 12541 8041 12575 8075
rect 13001 8041 13035 8075
rect 13369 8041 13403 8075
rect 13737 8041 13771 8075
rect 1593 7973 1627 8007
rect 7389 7973 7423 8007
rect 8493 7973 8527 8007
rect 11345 7973 11379 8007
rect 12909 7973 12943 8007
rect 1961 7905 1995 7939
rect 3709 7905 3743 7939
rect 3985 7905 4019 7939
rect 4905 7905 4939 7939
rect 6478 7905 6512 7939
rect 6745 7905 6779 7939
rect 8033 7905 8067 7939
rect 10517 7905 10551 7939
rect 12173 7905 12207 7939
rect 4537 7837 4571 7871
rect 4629 7837 4663 7871
rect 7205 7837 7239 7871
rect 8309 7837 8343 7871
rect 9597 7837 9631 7871
rect 9689 7837 9723 7871
rect 10241 7837 10275 7871
rect 10425 7837 10459 7871
rect 11529 7837 11563 7871
rect 11989 7837 12023 7871
rect 12081 7837 12115 7871
rect 12817 7837 12851 7871
rect 5089 7769 5123 7803
rect 5365 7769 5399 7803
rect 10977 7769 11011 7803
rect 3525 7701 3559 7735
rect 6837 7701 6871 7735
rect 7849 7701 7883 7735
rect 8953 7701 8987 7735
rect 10057 7701 10091 7735
rect 13461 7701 13495 7735
rect 2145 7497 2179 7531
rect 2881 7497 2915 7531
rect 4445 7497 4479 7531
rect 5549 7497 5583 7531
rect 6653 7497 6687 7531
rect 6929 7497 6963 7531
rect 8401 7497 8435 7531
rect 11437 7497 11471 7531
rect 4353 7429 4387 7463
rect 8493 7429 8527 7463
rect 9321 7429 9355 7463
rect 9505 7429 9539 7463
rect 5089 7361 5123 7395
rect 6193 7361 6227 7395
rect 7021 7361 7055 7395
rect 9045 7361 9079 7395
rect 9689 7361 9723 7395
rect 11897 7361 11931 7395
rect 12081 7361 12115 7395
rect 1961 7293 1995 7327
rect 2973 7293 3007 7327
rect 4905 7293 4939 7327
rect 5365 7293 5399 7327
rect 8861 7293 8895 7327
rect 8953 7293 8987 7327
rect 11253 7293 11287 7327
rect 12173 7293 12207 7327
rect 1593 7225 1627 7259
rect 3240 7225 3274 7259
rect 4813 7225 4847 7259
rect 7266 7225 7300 7259
rect 9956 7225 9990 7259
rect 1501 7157 1535 7191
rect 1777 7157 1811 7191
rect 2329 7157 2363 7191
rect 5917 7157 5951 7191
rect 6009 7157 6043 7191
rect 6469 7157 6503 7191
rect 11069 7157 11103 7191
rect 12541 7157 12575 7191
rect 12633 7157 12667 7191
rect 13001 7157 13035 7191
rect 8953 6953 8987 6987
rect 10609 6953 10643 6987
rect 13553 6953 13587 6987
rect 3433 6885 3467 6919
rect 4353 6885 4387 6919
rect 4537 6885 4571 6919
rect 5917 6885 5951 6919
rect 9382 6885 9416 6919
rect 10977 6885 11011 6919
rect 1593 6817 1627 6851
rect 2125 6817 2159 6851
rect 4997 6817 5031 6851
rect 5457 6817 5491 6851
rect 6009 6817 6043 6851
rect 6561 6817 6595 6851
rect 7840 6817 7874 6851
rect 9137 6817 9171 6851
rect 11877 6817 11911 6851
rect 13461 6817 13495 6851
rect 1869 6749 1903 6783
rect 6193 6749 6227 6783
rect 7481 6749 7515 6783
rect 7573 6749 7607 6783
rect 11069 6749 11103 6783
rect 11253 6749 11287 6783
rect 11621 6749 11655 6783
rect 13645 6749 13679 6783
rect 3893 6681 3927 6715
rect 4813 6681 4847 6715
rect 5549 6681 5583 6715
rect 6377 6681 6411 6715
rect 6745 6681 6779 6715
rect 10517 6681 10551 6715
rect 13001 6681 13035 6715
rect 13093 6681 13127 6715
rect 1501 6613 1535 6647
rect 3249 6613 3283 6647
rect 3709 6613 3743 6647
rect 4261 6613 4295 6647
rect 5273 6613 5307 6647
rect 6929 6613 6963 6647
rect 7021 6613 7055 6647
rect 11437 6613 11471 6647
rect 3249 6409 3283 6443
rect 3617 6409 3651 6443
rect 8769 6409 8803 6443
rect 9137 6409 9171 6443
rect 9321 6409 9355 6443
rect 10609 6409 10643 6443
rect 12541 6409 12575 6443
rect 13093 6409 13127 6443
rect 14289 6409 14323 6443
rect 15209 6409 15243 6443
rect 3801 6341 3835 6375
rect 13185 6341 13219 6375
rect 4353 6273 4387 6307
rect 5181 6273 5215 6307
rect 5365 6273 5399 6307
rect 6101 6273 6135 6307
rect 6561 6273 6595 6307
rect 6653 6273 6687 6307
rect 8309 6273 8343 6307
rect 9965 6273 9999 6307
rect 11253 6273 11287 6307
rect 11897 6273 11931 6307
rect 13369 6273 13403 6307
rect 2973 6205 3007 6239
rect 5089 6205 5123 6239
rect 6009 6205 6043 6239
rect 9413 6205 9447 6239
rect 10149 6205 10183 6239
rect 11069 6205 11103 6239
rect 1501 6137 1535 6171
rect 2706 6137 2740 6171
rect 4169 6137 4203 6171
rect 6653 6137 6687 6171
rect 6745 6137 6779 6171
rect 8042 6137 8076 6171
rect 12173 6137 12207 6171
rect 1593 6069 1627 6103
rect 3065 6069 3099 6103
rect 3433 6069 3467 6103
rect 4261 6069 4295 6103
rect 4721 6069 4755 6103
rect 5549 6069 5583 6103
rect 5917 6069 5951 6103
rect 6929 6069 6963 6103
rect 8401 6069 8435 6103
rect 8677 6069 8711 6103
rect 9597 6069 9631 6103
rect 10057 6069 10091 6103
rect 10517 6069 10551 6103
rect 10977 6069 11011 6103
rect 11437 6069 11471 6103
rect 12081 6069 12115 6103
rect 12633 6069 12667 6103
rect 12817 6069 12851 6103
rect 15393 6069 15427 6103
rect 1777 5865 1811 5899
rect 2513 5865 2547 5899
rect 2973 5865 3007 5899
rect 3433 5865 3467 5899
rect 3893 5865 3927 5899
rect 4261 5865 4295 5899
rect 5181 5865 5215 5899
rect 8125 5865 8159 5899
rect 9781 5865 9815 5899
rect 11437 5865 11471 5899
rect 11805 5865 11839 5899
rect 12633 5865 12667 5899
rect 14933 5865 14967 5899
rect 6408 5797 6442 5831
rect 10241 5797 10275 5831
rect 11161 5797 11195 5831
rect 11529 5797 11563 5831
rect 14381 5797 14415 5831
rect 15669 5797 15703 5831
rect 1685 5729 1719 5763
rect 1961 5729 1995 5763
rect 3341 5729 3375 5763
rect 4905 5729 4939 5763
rect 6653 5729 6687 5763
rect 7297 5729 7331 5763
rect 8217 5729 8251 5763
rect 8769 5729 8803 5763
rect 10149 5729 10183 5763
rect 12081 5729 12115 5763
rect 13369 5729 13403 5763
rect 14749 5729 14783 5763
rect 15485 5729 15519 5763
rect 2237 5661 2271 5695
rect 2421 5661 2455 5695
rect 3617 5661 3651 5695
rect 4353 5661 4387 5695
rect 4445 5661 4479 5695
rect 7389 5661 7423 5695
rect 7573 5661 7607 5695
rect 8309 5661 8343 5695
rect 10333 5661 10367 5695
rect 12449 5661 12483 5695
rect 13093 5661 13127 5695
rect 13277 5661 13311 5695
rect 15117 5661 15151 5695
rect 8585 5593 8619 5627
rect 9137 5593 9171 5627
rect 13737 5593 13771 5627
rect 1501 5525 1535 5559
rect 2881 5525 2915 5559
rect 4721 5525 4755 5559
rect 5273 5525 5307 5559
rect 6745 5525 6779 5559
rect 6929 5525 6963 5559
rect 7757 5525 7791 5559
rect 8953 5525 8987 5559
rect 9321 5525 9355 5559
rect 9597 5525 9631 5559
rect 10609 5525 10643 5559
rect 10885 5525 10919 5559
rect 11069 5525 11103 5559
rect 11989 5525 12023 5559
rect 12817 5525 12851 5559
rect 13829 5525 13863 5559
rect 14013 5525 14047 5559
rect 15209 5525 15243 5559
rect 2513 5321 2547 5355
rect 5273 5321 5307 5355
rect 6469 5321 6503 5355
rect 11069 5321 11103 5355
rect 13369 5321 13403 5355
rect 15393 5321 15427 5355
rect 1409 5253 1443 5287
rect 2605 5253 2639 5287
rect 7297 5253 7331 5287
rect 8309 5253 8343 5287
rect 10057 5253 10091 5287
rect 14841 5253 14875 5287
rect 1961 5185 1995 5219
rect 3065 5185 3099 5219
rect 3249 5185 3283 5219
rect 6009 5185 6043 5219
rect 6101 5185 6135 5219
rect 6929 5185 6963 5219
rect 7113 5185 7147 5219
rect 7849 5185 7883 5219
rect 9689 5185 9723 5219
rect 10701 5185 10735 5219
rect 11989 5185 12023 5219
rect 1593 5117 1627 5151
rect 2973 5117 3007 5151
rect 3617 5117 3651 5151
rect 3893 5117 3927 5151
rect 4160 5117 4194 5151
rect 6837 5117 6871 5151
rect 9965 5117 9999 5151
rect 10517 5117 10551 5151
rect 10885 5117 10919 5151
rect 13461 5117 13495 5151
rect 13717 5117 13751 5151
rect 15209 5117 15243 5151
rect 3709 5049 3743 5083
rect 5917 5049 5951 5083
rect 9422 5049 9456 5083
rect 11253 5049 11287 5083
rect 12256 5049 12290 5083
rect 2053 4981 2087 5015
rect 2145 4981 2179 5015
rect 3433 4981 3467 5015
rect 5365 4981 5399 5015
rect 5549 4981 5583 5015
rect 7665 4981 7699 5015
rect 7757 4981 7791 5015
rect 8125 4981 8159 5015
rect 9781 4981 9815 5015
rect 10425 4981 10459 5015
rect 11345 4981 11379 5015
rect 11713 4981 11747 5015
rect 14933 4981 14967 5015
rect 15485 4981 15519 5015
rect 2053 4777 2087 4811
rect 2881 4777 2915 4811
rect 3893 4777 3927 4811
rect 6009 4777 6043 4811
rect 6745 4777 6779 4811
rect 7205 4777 7239 4811
rect 7389 4777 7423 4811
rect 7757 4777 7791 4811
rect 7849 4777 7883 4811
rect 9965 4777 9999 4811
rect 13185 4777 13219 4811
rect 13829 4777 13863 4811
rect 15485 4777 15519 4811
rect 2513 4709 2547 4743
rect 3341 4709 3375 4743
rect 7021 4709 7055 4743
rect 9321 4709 9355 4743
rect 11468 4709 11502 4743
rect 13737 4709 13771 4743
rect 14749 4709 14783 4743
rect 1685 4641 1719 4675
rect 1961 4641 1995 4675
rect 2421 4641 2455 4675
rect 3249 4641 3283 4675
rect 4261 4641 4295 4675
rect 4353 4641 4387 4675
rect 4905 4641 4939 4675
rect 5181 4641 5215 4675
rect 5457 4641 5491 4675
rect 5549 4641 5583 4675
rect 5825 4641 5859 4675
rect 6377 4641 6411 4675
rect 6561 4641 6595 4675
rect 8585 4641 8619 4675
rect 9873 4641 9907 4675
rect 11713 4641 11747 4675
rect 12072 4641 12106 4675
rect 14841 4641 14875 4675
rect 15577 4641 15611 4675
rect 2697 4573 2731 4607
rect 3525 4573 3559 4607
rect 4445 4573 4479 4607
rect 8033 4573 8067 4607
rect 8677 4573 8711 4607
rect 8861 4573 8895 4607
rect 10149 4573 10183 4607
rect 11805 4573 11839 4607
rect 13553 4573 13587 4607
rect 14933 4573 14967 4607
rect 5273 4505 5307 4539
rect 5733 4505 5767 4539
rect 6837 4505 6871 4539
rect 9137 4505 9171 4539
rect 13277 4505 13311 4539
rect 1501 4437 1535 4471
rect 1777 4437 1811 4471
rect 4721 4437 4755 4471
rect 4997 4437 5031 4471
rect 6193 4437 6227 4471
rect 8217 4437 8251 4471
rect 9505 4437 9539 4471
rect 10333 4437 10367 4471
rect 14197 4437 14231 4471
rect 14381 4437 14415 4471
rect 15209 4437 15243 4471
rect 3065 4233 3099 4267
rect 5089 4233 5123 4267
rect 7941 4233 7975 4267
rect 11069 4233 11103 4267
rect 15117 4233 15151 4267
rect 4905 4165 4939 4199
rect 1409 4097 1443 4131
rect 4445 4097 4479 4131
rect 5641 4097 5675 4131
rect 6469 4097 6503 4131
rect 8401 4097 8435 4131
rect 8585 4097 8619 4131
rect 9505 4097 9539 4131
rect 9597 4097 9631 4131
rect 10701 4097 10735 4131
rect 12173 4097 12207 4131
rect 13001 4097 13035 4131
rect 14197 4097 14231 4131
rect 14565 4097 14599 4131
rect 15393 4097 15427 4131
rect 1593 4029 1627 4063
rect 1961 4029 1995 4063
rect 2237 4029 2271 4063
rect 2421 4029 2455 4063
rect 2789 4029 2823 4063
rect 4721 4029 4755 4063
rect 6101 4029 6135 4063
rect 6725 4029 6759 4063
rect 8769 4029 8803 4063
rect 9137 4029 9171 4063
rect 10609 4029 10643 4063
rect 11161 4029 11195 4063
rect 11345 4029 11379 4063
rect 11897 4029 11931 4063
rect 14013 4029 14047 4063
rect 14105 4029 14139 4063
rect 15577 4029 15611 4063
rect 2973 3961 3007 3995
rect 4178 3961 4212 3995
rect 5457 3961 5491 3995
rect 8953 3961 8987 3995
rect 9689 3961 9723 3995
rect 12265 3961 12299 3995
rect 13185 3961 13219 3995
rect 14749 3961 14783 3995
rect 14933 3961 14967 3995
rect 15209 3961 15243 3995
rect 1777 3893 1811 3927
rect 2053 3893 2087 3927
rect 2605 3893 2639 3927
rect 4629 3893 4663 3927
rect 5549 3893 5583 3927
rect 6193 3893 6227 3927
rect 7849 3893 7883 3927
rect 8309 3893 8343 3927
rect 10057 3893 10091 3927
rect 10149 3893 10183 3927
rect 10517 3893 10551 3927
rect 11713 3893 11747 3927
rect 12357 3893 12391 3927
rect 12725 3893 12759 3927
rect 13093 3893 13127 3927
rect 13553 3893 13587 3927
rect 13645 3893 13679 3927
rect 3525 3689 3559 3723
rect 4353 3689 4387 3723
rect 5825 3689 5859 3723
rect 8953 3689 8987 3723
rect 9781 3689 9815 3723
rect 9873 3689 9907 3723
rect 11345 3689 11379 3723
rect 12173 3689 12207 3723
rect 12909 3689 12943 3723
rect 14933 3689 14967 3723
rect 15393 3689 15427 3723
rect 1593 3621 1627 3655
rect 1961 3621 1995 3655
rect 4077 3621 4111 3655
rect 6193 3621 6227 3655
rect 10333 3621 10367 3655
rect 11897 3621 11931 3655
rect 14473 3621 14507 3655
rect 14657 3621 14691 3655
rect 15025 3621 15059 3655
rect 15485 3621 15519 3655
rect 2412 3553 2446 3587
rect 5477 3553 5511 3587
rect 6009 3553 6043 3587
rect 6837 3553 6871 3587
rect 6929 3553 6963 3587
rect 7481 3553 7515 3587
rect 7573 3553 7607 3587
rect 7840 3553 7874 3587
rect 9321 3553 9355 3587
rect 11253 3553 11287 3587
rect 12265 3553 12299 3587
rect 12817 3553 12851 3587
rect 13369 3553 13403 3587
rect 13553 3553 13587 3587
rect 13737 3553 13771 3587
rect 13921 3553 13955 3587
rect 2145 3485 2179 3519
rect 3709 3485 3743 3519
rect 5733 3485 5767 3519
rect 6377 3485 6411 3519
rect 7113 3485 7147 3519
rect 9965 3485 9999 3519
rect 11437 3485 11471 3519
rect 12633 3485 12667 3519
rect 3893 3417 3927 3451
rect 1501 3349 1535 3383
rect 1869 3349 1903 3383
rect 6469 3349 6503 3383
rect 7297 3349 7331 3383
rect 9137 3349 9171 3383
rect 9413 3349 9447 3383
rect 10609 3349 10643 3383
rect 10885 3349 10919 3383
rect 11805 3349 11839 3383
rect 13277 3349 13311 3383
rect 14105 3349 14139 3383
rect 4353 3145 4387 3179
rect 5549 3145 5583 3179
rect 8309 3145 8343 3179
rect 14289 3145 14323 3179
rect 14473 3145 14507 3179
rect 2145 3077 2179 3111
rect 2881 3077 2915 3111
rect 6561 3077 6595 3111
rect 11437 3077 11471 3111
rect 11989 3077 12023 3111
rect 2513 3009 2547 3043
rect 3249 3009 3283 3043
rect 3801 3009 3835 3043
rect 5089 3009 5123 3043
rect 6009 3009 6043 3043
rect 6193 3009 6227 3043
rect 7941 3009 7975 3043
rect 9689 3009 9723 3043
rect 11161 3009 11195 3043
rect 12265 3009 12299 3043
rect 12909 3009 12943 3043
rect 15577 3009 15611 3043
rect 1593 2941 1627 2975
rect 2329 2941 2363 2975
rect 3065 2941 3099 2975
rect 3433 2941 3467 2975
rect 3985 2941 4019 2975
rect 4905 2941 4939 2975
rect 7685 2941 7719 2975
rect 8217 2941 8251 2975
rect 11253 2941 11287 2975
rect 11805 2941 11839 2975
rect 12449 2941 12483 2975
rect 14565 2941 14599 2975
rect 15025 2941 15059 2975
rect 1409 2873 1443 2907
rect 1961 2873 1995 2907
rect 2697 2873 2731 2907
rect 3893 2873 3927 2907
rect 9444 2873 9478 2907
rect 10894 2873 10928 2907
rect 13154 2873 13188 2907
rect 15301 2873 15335 2907
rect 1869 2805 1903 2839
rect 4445 2805 4479 2839
rect 4813 2805 4847 2839
rect 5273 2805 5307 2839
rect 5917 2805 5951 2839
rect 8033 2805 8067 2839
rect 9781 2805 9815 2839
rect 12357 2805 12391 2839
rect 12817 2805 12851 2839
rect 14749 2805 14783 2839
rect 1777 2601 1811 2635
rect 3525 2601 3559 2635
rect 3893 2601 3927 2635
rect 4537 2601 4571 2635
rect 4905 2601 4939 2635
rect 5549 2601 5583 2635
rect 6009 2601 6043 2635
rect 9229 2601 9263 2635
rect 9597 2601 9631 2635
rect 10057 2601 10091 2635
rect 10425 2601 10459 2635
rect 10885 2601 10919 2635
rect 11253 2601 11287 2635
rect 12449 2601 12483 2635
rect 13277 2601 13311 2635
rect 13369 2601 13403 2635
rect 14197 2601 14231 2635
rect 1593 2533 1627 2567
rect 2320 2533 2354 2567
rect 5457 2533 5491 2567
rect 5917 2533 5951 2567
rect 7113 2533 7147 2567
rect 7849 2533 7883 2567
rect 9689 2533 9723 2567
rect 11897 2533 11931 2567
rect 14289 2533 14323 2567
rect 1961 2465 1995 2499
rect 3709 2465 3743 2499
rect 4077 2465 4111 2499
rect 4353 2465 4387 2499
rect 6745 2465 6779 2499
rect 7481 2465 7515 2499
rect 8401 2465 8435 2499
rect 8953 2465 8987 2499
rect 10517 2465 10551 2499
rect 12541 2465 12575 2499
rect 13921 2465 13955 2499
rect 14841 2465 14875 2499
rect 15485 2465 15519 2499
rect 2053 2397 2087 2431
rect 4997 2397 5031 2431
rect 5181 2397 5215 2431
rect 6193 2397 6227 2431
rect 7665 2397 7699 2431
rect 9781 2397 9815 2431
rect 10609 2397 10643 2431
rect 11345 2397 11379 2431
rect 11437 2397 11471 2431
rect 12633 2397 12667 2431
rect 13553 2397 13587 2431
rect 14565 2397 14599 2431
rect 1409 2329 1443 2363
rect 7297 2329 7331 2363
rect 12081 2329 12115 2363
rect 12909 2329 12943 2363
rect 3433 2261 3467 2295
rect 4261 2261 4295 2295
rect 6653 2261 6687 2295
rect 7021 2261 7055 2295
rect 8125 2261 8159 2295
rect 8861 2261 8895 2295
rect 13829 2261 13863 2295
rect 15669 2261 15703 2295
<< metal1 >>
rect 3970 17552 3976 17604
rect 4028 17592 4034 17604
rect 7742 17592 7748 17604
rect 4028 17564 7748 17592
rect 4028 17552 4034 17564
rect 7742 17552 7748 17564
rect 7800 17552 7806 17604
rect 4338 17484 4344 17536
rect 4396 17524 4402 17536
rect 7466 17524 7472 17536
rect 4396 17496 7472 17524
rect 4396 17484 4402 17496
rect 7466 17484 7472 17496
rect 7524 17484 7530 17536
rect 1104 17434 16008 17456
rect 1104 17382 3480 17434
rect 3532 17382 3544 17434
rect 3596 17382 3608 17434
rect 3660 17382 3672 17434
rect 3724 17382 8478 17434
rect 8530 17382 8542 17434
rect 8594 17382 8606 17434
rect 8658 17382 8670 17434
rect 8722 17382 13475 17434
rect 13527 17382 13539 17434
rect 13591 17382 13603 17434
rect 13655 17382 13667 17434
rect 13719 17382 16008 17434
rect 1104 17360 16008 17382
rect 934 17280 940 17332
rect 992 17320 998 17332
rect 1857 17323 1915 17329
rect 1857 17320 1869 17323
rect 992 17292 1869 17320
rect 992 17280 998 17292
rect 1857 17289 1869 17292
rect 1903 17289 1915 17323
rect 1857 17283 1915 17289
rect 4433 17323 4491 17329
rect 4433 17289 4445 17323
rect 4479 17320 4491 17323
rect 7098 17320 7104 17332
rect 4479 17292 7104 17320
rect 4479 17289 4491 17292
rect 4433 17283 4491 17289
rect 7098 17280 7104 17292
rect 7156 17280 7162 17332
rect 7374 17280 7380 17332
rect 7432 17320 7438 17332
rect 7561 17323 7619 17329
rect 7561 17320 7573 17323
rect 7432 17292 7573 17320
rect 7432 17280 7438 17292
rect 7561 17289 7573 17292
rect 7607 17289 7619 17323
rect 7561 17283 7619 17289
rect 7929 17323 7987 17329
rect 7929 17289 7941 17323
rect 7975 17320 7987 17323
rect 12618 17320 12624 17332
rect 7975 17292 12624 17320
rect 7975 17289 7987 17292
rect 7929 17283 7987 17289
rect 12618 17280 12624 17292
rect 12676 17280 12682 17332
rect 13265 17323 13323 17329
rect 13265 17289 13277 17323
rect 13311 17320 13323 17323
rect 13906 17320 13912 17332
rect 13311 17292 13912 17320
rect 13311 17289 13323 17292
rect 13265 17283 13323 17289
rect 13906 17280 13912 17292
rect 13964 17280 13970 17332
rect 14001 17323 14059 17329
rect 14001 17289 14013 17323
rect 14047 17320 14059 17323
rect 14826 17320 14832 17332
rect 14047 17292 14832 17320
rect 14047 17289 14059 17292
rect 14001 17283 14059 17289
rect 14826 17280 14832 17292
rect 14884 17280 14890 17332
rect 15010 17320 15016 17332
rect 14971 17292 15016 17320
rect 15010 17280 15016 17292
rect 15068 17280 15074 17332
rect 566 17212 572 17264
rect 624 17252 630 17264
rect 1397 17255 1455 17261
rect 1397 17252 1409 17255
rect 624 17224 1409 17252
rect 624 17212 630 17224
rect 1397 17221 1409 17224
rect 1443 17221 1455 17255
rect 1397 17215 1455 17221
rect 1486 17212 1492 17264
rect 1544 17252 1550 17264
rect 2133 17255 2191 17261
rect 2133 17252 2145 17255
rect 1544 17224 2145 17252
rect 1544 17212 1550 17224
rect 2133 17221 2145 17224
rect 2179 17221 2191 17255
rect 2133 17215 2191 17221
rect 2222 17212 2228 17264
rect 2280 17252 2286 17264
rect 2869 17255 2927 17261
rect 2869 17252 2881 17255
rect 2280 17224 2881 17252
rect 2280 17212 2286 17224
rect 2869 17221 2881 17224
rect 2915 17221 2927 17255
rect 4614 17252 4620 17264
rect 4575 17224 4620 17252
rect 2869 17215 2927 17221
rect 4614 17212 4620 17224
rect 4672 17212 4678 17264
rect 5074 17252 5080 17264
rect 5035 17224 5080 17252
rect 5074 17212 5080 17224
rect 5132 17212 5138 17264
rect 5442 17252 5448 17264
rect 5403 17224 5448 17252
rect 5442 17212 5448 17224
rect 5500 17212 5506 17264
rect 5902 17252 5908 17264
rect 5863 17224 5908 17252
rect 5902 17212 5908 17224
rect 5960 17212 5966 17264
rect 6270 17212 6276 17264
rect 6328 17252 6334 17264
rect 6549 17255 6607 17261
rect 6549 17252 6561 17255
rect 6328 17224 6561 17252
rect 6328 17212 6334 17224
rect 6549 17221 6561 17224
rect 6595 17221 6607 17255
rect 6549 17215 6607 17221
rect 6730 17212 6736 17264
rect 6788 17252 6794 17264
rect 6917 17255 6975 17261
rect 6917 17252 6929 17255
rect 6788 17224 6929 17252
rect 6788 17212 6794 17224
rect 6917 17221 6929 17224
rect 6963 17221 6975 17255
rect 7834 17252 7840 17264
rect 6917 17215 6975 17221
rect 7024 17224 7840 17252
rect 1762 17144 1768 17196
rect 1820 17184 1826 17196
rect 2501 17187 2559 17193
rect 2501 17184 2513 17187
rect 1820 17156 2513 17184
rect 1820 17144 1826 17156
rect 2501 17153 2513 17156
rect 2547 17153 2559 17187
rect 2501 17147 2559 17153
rect 3697 17187 3755 17193
rect 3697 17153 3709 17187
rect 3743 17184 3755 17187
rect 7024 17184 7052 17224
rect 7834 17212 7840 17224
rect 7892 17212 7898 17264
rect 8297 17255 8355 17261
rect 8297 17221 8309 17255
rect 8343 17252 8355 17255
rect 9214 17252 9220 17264
rect 8343 17224 9220 17252
rect 8343 17221 8355 17224
rect 8297 17215 8355 17221
rect 9214 17212 9220 17224
rect 9272 17212 9278 17264
rect 12158 17212 12164 17264
rect 12216 17252 12222 17264
rect 13541 17255 13599 17261
rect 13541 17252 13553 17255
rect 12216 17224 13553 17252
rect 12216 17212 12222 17224
rect 13541 17221 13553 17224
rect 13587 17221 13599 17255
rect 13541 17215 13599 17221
rect 14274 17212 14280 17264
rect 14332 17252 14338 17264
rect 14553 17255 14611 17261
rect 14553 17252 14565 17255
rect 14332 17224 14565 17252
rect 14332 17212 14338 17224
rect 14553 17221 14565 17224
rect 14599 17221 14611 17255
rect 14553 17215 14611 17221
rect 3743 17156 7052 17184
rect 7377 17187 7435 17193
rect 3743 17153 3755 17156
rect 3697 17147 3755 17153
rect 7377 17153 7389 17187
rect 7423 17184 7435 17187
rect 9122 17184 9128 17196
rect 7423 17156 9128 17184
rect 7423 17153 7435 17156
rect 7377 17147 7435 17153
rect 3970 17116 3976 17128
rect 3931 17088 3976 17116
rect 3970 17076 3976 17088
rect 4028 17076 4034 17128
rect 4157 17119 4215 17125
rect 4157 17085 4169 17119
rect 4203 17116 4215 17119
rect 7558 17116 7564 17128
rect 4203 17088 7564 17116
rect 4203 17085 4215 17088
rect 4157 17079 4215 17085
rect 7558 17076 7564 17088
rect 7616 17076 7622 17128
rect 8496 17125 8524 17156
rect 9122 17144 9128 17156
rect 9180 17144 9186 17196
rect 11054 17144 11060 17196
rect 11112 17184 11118 17196
rect 12989 17187 13047 17193
rect 11112 17156 12388 17184
rect 11112 17144 11118 17156
rect 8481 17119 8539 17125
rect 8481 17085 8493 17119
rect 8527 17085 8539 17119
rect 8481 17079 8539 17085
rect 8846 17076 8852 17128
rect 8904 17116 8910 17128
rect 8941 17119 8999 17125
rect 8941 17116 8953 17119
rect 8904 17088 8953 17116
rect 8904 17076 8910 17088
rect 8941 17085 8953 17088
rect 8987 17116 8999 17119
rect 9217 17119 9275 17125
rect 9217 17116 9229 17119
rect 8987 17088 9229 17116
rect 8987 17085 8999 17088
rect 8941 17079 8999 17085
rect 9217 17085 9229 17088
rect 9263 17085 9275 17119
rect 9217 17079 9275 17085
rect 9401 17119 9459 17125
rect 9401 17085 9413 17119
rect 9447 17085 9459 17119
rect 9401 17079 9459 17085
rect 9668 17119 9726 17125
rect 9668 17085 9680 17119
rect 9714 17116 9726 17119
rect 10502 17116 10508 17128
rect 9714 17088 10508 17116
rect 9714 17085 9726 17088
rect 9668 17079 9726 17085
rect 1581 17051 1639 17057
rect 1581 17017 1593 17051
rect 1627 17048 1639 17051
rect 1670 17048 1676 17060
rect 1627 17020 1676 17048
rect 1627 17017 1639 17020
rect 1581 17011 1639 17017
rect 1670 17008 1676 17020
rect 1728 17008 1734 17060
rect 1949 17051 2007 17057
rect 1949 17017 1961 17051
rect 1995 17048 2007 17051
rect 2130 17048 2136 17060
rect 1995 17020 2136 17048
rect 1995 17017 2007 17020
rect 1949 17011 2007 17017
rect 2130 17008 2136 17020
rect 2188 17008 2194 17060
rect 2222 17008 2228 17060
rect 2280 17048 2286 17060
rect 2317 17051 2375 17057
rect 2317 17048 2329 17051
rect 2280 17020 2329 17048
rect 2280 17008 2286 17020
rect 2317 17017 2329 17020
rect 2363 17017 2375 17051
rect 2682 17048 2688 17060
rect 2643 17020 2688 17048
rect 2317 17011 2375 17017
rect 2682 17008 2688 17020
rect 2740 17008 2746 17060
rect 2866 17008 2872 17060
rect 2924 17048 2930 17060
rect 3053 17051 3111 17057
rect 3053 17048 3065 17051
rect 2924 17020 3065 17048
rect 2924 17008 2930 17020
rect 3053 17017 3065 17020
rect 3099 17017 3111 17051
rect 3053 17011 3111 17017
rect 3513 17051 3571 17057
rect 3513 17017 3525 17051
rect 3559 17017 3571 17051
rect 4338 17048 4344 17060
rect 4299 17020 4344 17048
rect 3513 17011 3571 17017
rect 3528 16980 3556 17011
rect 4338 17008 4344 17020
rect 4396 17008 4402 17060
rect 4798 17048 4804 17060
rect 4759 17020 4804 17048
rect 4798 17008 4804 17020
rect 4856 17008 4862 17060
rect 5074 17008 5080 17060
rect 5132 17048 5138 17060
rect 5261 17051 5319 17057
rect 5261 17048 5273 17051
rect 5132 17020 5273 17048
rect 5132 17008 5138 17020
rect 5261 17017 5273 17020
rect 5307 17017 5319 17051
rect 5626 17048 5632 17060
rect 5587 17020 5632 17048
rect 5261 17011 5319 17017
rect 5626 17008 5632 17020
rect 5684 17008 5690 17060
rect 5810 17008 5816 17060
rect 5868 17048 5874 17060
rect 6089 17051 6147 17057
rect 6089 17048 6101 17051
rect 5868 17020 6101 17048
rect 5868 17008 5874 17020
rect 6089 17017 6101 17020
rect 6135 17017 6147 17051
rect 6730 17048 6736 17060
rect 6691 17020 6736 17048
rect 6089 17011 6147 17017
rect 6730 17008 6736 17020
rect 6788 17008 6794 17060
rect 7098 17048 7104 17060
rect 7059 17020 7104 17048
rect 7098 17008 7104 17020
rect 7156 17008 7162 17060
rect 7650 17048 7656 17060
rect 7392 17020 7656 17048
rect 5442 16980 5448 16992
rect 3528 16952 5448 16980
rect 5442 16940 5448 16952
rect 5500 16940 5506 16992
rect 6365 16983 6423 16989
rect 6365 16949 6377 16983
rect 6411 16980 6423 16983
rect 7392 16980 7420 17020
rect 7650 17008 7656 17020
rect 7708 17008 7714 17060
rect 8018 17048 8024 17060
rect 7979 17020 8024 17048
rect 8018 17008 8024 17020
rect 8076 17008 8082 17060
rect 8110 17008 8116 17060
rect 8168 17048 8174 17060
rect 8168 17020 8800 17048
rect 8168 17008 8174 17020
rect 6411 16952 7420 16980
rect 6411 16949 6423 16952
rect 6365 16943 6423 16949
rect 8202 16940 8208 16992
rect 8260 16980 8266 16992
rect 8665 16983 8723 16989
rect 8665 16980 8677 16983
rect 8260 16952 8677 16980
rect 8260 16940 8266 16952
rect 8665 16949 8677 16952
rect 8711 16949 8723 16983
rect 8772 16980 8800 17020
rect 9122 17008 9128 17060
rect 9180 17048 9186 17060
rect 9416 17048 9444 17079
rect 10502 17076 10508 17088
rect 10560 17076 10566 17128
rect 11333 17119 11391 17125
rect 11333 17085 11345 17119
rect 11379 17116 11391 17119
rect 12250 17116 12256 17128
rect 11379 17088 12256 17116
rect 11379 17085 11391 17088
rect 11333 17079 11391 17085
rect 12250 17076 12256 17088
rect 12308 17076 12314 17128
rect 9180 17020 9444 17048
rect 9180 17008 9186 17020
rect 9766 17008 9772 17060
rect 9824 17048 9830 17060
rect 10965 17051 11023 17057
rect 10965 17048 10977 17051
rect 9824 17020 10977 17048
rect 9824 17008 9830 17020
rect 10965 17017 10977 17020
rect 11011 17017 11023 17051
rect 10965 17011 11023 17017
rect 11609 17051 11667 17057
rect 11609 17017 11621 17051
rect 11655 17048 11667 17051
rect 11790 17048 11796 17060
rect 11655 17020 11796 17048
rect 11655 17017 11667 17020
rect 11609 17011 11667 17017
rect 11790 17008 11796 17020
rect 11848 17008 11854 17060
rect 11974 17008 11980 17060
rect 12032 17048 12038 17060
rect 12161 17051 12219 17057
rect 12161 17048 12173 17051
rect 12032 17020 12173 17048
rect 12032 17008 12038 17020
rect 12161 17017 12173 17020
rect 12207 17017 12219 17051
rect 12161 17011 12219 17017
rect 9858 16980 9864 16992
rect 8772 16952 9864 16980
rect 8665 16943 8723 16949
rect 9858 16940 9864 16952
rect 9916 16940 9922 16992
rect 10778 16980 10784 16992
rect 10739 16952 10784 16980
rect 10778 16940 10784 16952
rect 10836 16940 10842 16992
rect 11514 16980 11520 16992
rect 11475 16952 11520 16980
rect 11514 16940 11520 16952
rect 11572 16940 11578 16992
rect 12069 16983 12127 16989
rect 12069 16949 12081 16983
rect 12115 16980 12127 16983
rect 12250 16980 12256 16992
rect 12115 16952 12256 16980
rect 12115 16949 12127 16952
rect 12069 16943 12127 16949
rect 12250 16940 12256 16952
rect 12308 16940 12314 16992
rect 12360 16989 12388 17156
rect 12989 17153 13001 17187
rect 13035 17184 13047 17187
rect 13906 17184 13912 17196
rect 13035 17156 13912 17184
rect 13035 17153 13047 17156
rect 12989 17147 13047 17153
rect 13906 17144 13912 17156
rect 13964 17144 13970 17196
rect 15565 17187 15623 17193
rect 15565 17184 15577 17187
rect 14476 17156 15577 17184
rect 13262 17076 13268 17128
rect 13320 17116 13326 17128
rect 13725 17119 13783 17125
rect 13725 17116 13737 17119
rect 13320 17088 13737 17116
rect 13320 17076 13326 17088
rect 13725 17085 13737 17088
rect 13771 17085 13783 17119
rect 14277 17119 14335 17125
rect 14277 17116 14289 17119
rect 13725 17079 13783 17085
rect 13832 17088 14289 17116
rect 12894 17008 12900 17060
rect 12952 17048 12958 17060
rect 13357 17051 13415 17057
rect 13357 17048 13369 17051
rect 12952 17020 13369 17048
rect 12952 17008 12958 17020
rect 13357 17017 13369 17020
rect 13403 17048 13415 17051
rect 13832 17048 13860 17088
rect 14277 17085 14289 17088
rect 14323 17085 14335 17119
rect 14277 17079 14335 17085
rect 14093 17051 14151 17057
rect 14093 17048 14105 17051
rect 13403 17020 13860 17048
rect 13924 17020 14105 17048
rect 13403 17017 13415 17020
rect 13357 17011 13415 17017
rect 12345 16983 12403 16989
rect 12345 16949 12357 16983
rect 12391 16949 12403 16983
rect 12710 16980 12716 16992
rect 12671 16952 12716 16980
rect 12345 16943 12403 16949
rect 12710 16940 12716 16952
rect 12768 16940 12774 16992
rect 12805 16983 12863 16989
rect 12805 16949 12817 16983
rect 12851 16980 12863 16983
rect 12986 16980 12992 16992
rect 12851 16952 12992 16980
rect 12851 16949 12863 16952
rect 12805 16943 12863 16949
rect 12986 16940 12992 16952
rect 13044 16940 13050 16992
rect 13814 16940 13820 16992
rect 13872 16980 13878 16992
rect 13924 16980 13952 17020
rect 14093 17017 14105 17020
rect 14139 17048 14151 17051
rect 14476 17048 14504 17156
rect 15565 17153 15577 17156
rect 15611 17153 15623 17187
rect 15565 17147 15623 17153
rect 14550 17076 14556 17128
rect 14608 17116 14614 17128
rect 14921 17119 14979 17125
rect 14921 17116 14933 17119
rect 14608 17088 14933 17116
rect 14608 17076 14614 17088
rect 14921 17085 14933 17088
rect 14967 17085 14979 17119
rect 14921 17079 14979 17085
rect 14737 17051 14795 17057
rect 14737 17048 14749 17051
rect 14139 17020 14504 17048
rect 14568 17020 14749 17048
rect 14139 17017 14151 17020
rect 14093 17011 14151 17017
rect 13872 16952 13952 16980
rect 13872 16940 13878 16952
rect 14182 16940 14188 16992
rect 14240 16980 14246 16992
rect 14568 16980 14596 17020
rect 14737 17017 14749 17020
rect 14783 17017 14795 17051
rect 14737 17011 14795 17017
rect 14240 16952 14596 16980
rect 14240 16940 14246 16952
rect 15286 16940 15292 16992
rect 15344 16980 15350 16992
rect 15381 16983 15439 16989
rect 15381 16980 15393 16983
rect 15344 16952 15393 16980
rect 15344 16940 15350 16952
rect 15381 16949 15393 16952
rect 15427 16949 15439 16983
rect 15381 16943 15439 16949
rect 1104 16890 16008 16912
rect 1104 16838 5979 16890
rect 6031 16838 6043 16890
rect 6095 16838 6107 16890
rect 6159 16838 6171 16890
rect 6223 16838 10976 16890
rect 11028 16838 11040 16890
rect 11092 16838 11104 16890
rect 11156 16838 11168 16890
rect 11220 16838 16008 16890
rect 1104 16816 16008 16838
rect 1854 16776 1860 16788
rect 1815 16748 1860 16776
rect 1854 16736 1860 16748
rect 1912 16736 1918 16788
rect 2130 16776 2136 16788
rect 2091 16748 2136 16776
rect 2130 16736 2136 16748
rect 2188 16736 2194 16788
rect 4617 16779 4675 16785
rect 4617 16776 4629 16779
rect 4448 16748 4629 16776
rect 1394 16708 1400 16720
rect 1355 16680 1400 16708
rect 1394 16668 1400 16680
rect 1452 16668 1458 16720
rect 2590 16668 2596 16720
rect 2648 16708 2654 16720
rect 3050 16708 3056 16720
rect 2648 16680 2693 16708
rect 3011 16680 3056 16708
rect 2648 16668 2654 16680
rect 3050 16668 3056 16680
rect 3108 16668 3114 16720
rect 3326 16668 3332 16720
rect 3384 16708 3390 16720
rect 3421 16711 3479 16717
rect 3421 16708 3433 16711
rect 3384 16680 3433 16708
rect 3384 16668 3390 16680
rect 3421 16677 3433 16680
rect 3467 16677 3479 16711
rect 3878 16708 3884 16720
rect 3839 16680 3884 16708
rect 3421 16671 3479 16677
rect 3878 16668 3884 16680
rect 3936 16668 3942 16720
rect 4246 16708 4252 16720
rect 4207 16680 4252 16708
rect 4246 16668 4252 16680
rect 4304 16668 4310 16720
rect 4448 16717 4476 16748
rect 4617 16745 4629 16748
rect 4663 16745 4675 16779
rect 5074 16776 5080 16788
rect 5035 16748 5080 16776
rect 4617 16739 4675 16745
rect 5074 16736 5080 16748
rect 5132 16736 5138 16788
rect 8110 16776 8116 16788
rect 5276 16748 8116 16776
rect 4433 16711 4491 16717
rect 4433 16677 4445 16711
rect 4479 16677 4491 16711
rect 4433 16671 4491 16677
rect 1578 16640 1584 16652
rect 1539 16612 1584 16640
rect 1578 16600 1584 16612
rect 1636 16600 1642 16652
rect 1946 16640 1952 16652
rect 1907 16612 1952 16640
rect 1946 16600 1952 16612
rect 2004 16600 2010 16652
rect 2317 16643 2375 16649
rect 2317 16609 2329 16643
rect 2363 16640 2375 16643
rect 2406 16640 2412 16652
rect 2363 16612 2412 16640
rect 2363 16609 2375 16612
rect 2317 16603 2375 16609
rect 2406 16600 2412 16612
rect 2464 16600 2470 16652
rect 2777 16643 2835 16649
rect 2777 16609 2789 16643
rect 2823 16609 2835 16643
rect 3234 16640 3240 16652
rect 3195 16612 3240 16640
rect 2777 16603 2835 16609
rect 2792 16516 2820 16603
rect 3234 16600 3240 16612
rect 3292 16600 3298 16652
rect 3605 16643 3663 16649
rect 3605 16609 3617 16643
rect 3651 16640 3663 16643
rect 3786 16640 3792 16652
rect 3651 16612 3792 16640
rect 3651 16609 3663 16612
rect 3605 16603 3663 16609
rect 3786 16600 3792 16612
rect 3844 16600 3850 16652
rect 3970 16600 3976 16652
rect 4028 16640 4034 16652
rect 4065 16643 4123 16649
rect 4065 16640 4077 16643
rect 4028 16612 4077 16640
rect 4028 16600 4034 16612
rect 4065 16609 4077 16612
rect 4111 16609 4123 16643
rect 4065 16603 4123 16609
rect 4801 16643 4859 16649
rect 4801 16609 4813 16643
rect 4847 16640 4859 16643
rect 4890 16640 4896 16652
rect 4847 16612 4896 16640
rect 4847 16609 4859 16612
rect 4801 16603 4859 16609
rect 4890 16600 4896 16612
rect 4948 16600 4954 16652
rect 5276 16649 5304 16748
rect 8110 16736 8116 16748
rect 8168 16736 8174 16788
rect 8294 16736 8300 16788
rect 8352 16776 8358 16788
rect 8481 16779 8539 16785
rect 8481 16776 8493 16779
rect 8352 16748 8493 16776
rect 8352 16736 8358 16748
rect 8481 16745 8493 16748
rect 8527 16745 8539 16779
rect 8481 16739 8539 16745
rect 8757 16779 8815 16785
rect 8757 16745 8769 16779
rect 8803 16745 8815 16779
rect 8757 16739 8815 16745
rect 11425 16779 11483 16785
rect 11425 16745 11437 16779
rect 11471 16776 11483 16779
rect 11882 16776 11888 16788
rect 11471 16748 11888 16776
rect 11471 16745 11483 16748
rect 11425 16739 11483 16745
rect 5534 16668 5540 16720
rect 5592 16717 5598 16720
rect 5592 16711 5656 16717
rect 5592 16677 5610 16711
rect 5644 16677 5656 16711
rect 5592 16671 5656 16677
rect 5592 16668 5598 16671
rect 6638 16668 6644 16720
rect 6696 16708 6702 16720
rect 7070 16711 7128 16717
rect 7070 16708 7082 16711
rect 6696 16680 7082 16708
rect 6696 16668 6702 16680
rect 7070 16677 7082 16680
rect 7116 16677 7128 16711
rect 8772 16708 8800 16739
rect 11882 16736 11888 16748
rect 11940 16736 11946 16788
rect 12713 16779 12771 16785
rect 12713 16745 12725 16779
rect 12759 16776 12771 16779
rect 13906 16776 13912 16788
rect 12759 16748 13912 16776
rect 12759 16745 12771 16748
rect 12713 16739 12771 16745
rect 13906 16736 13912 16748
rect 13964 16736 13970 16788
rect 14461 16779 14519 16785
rect 14461 16745 14473 16779
rect 14507 16776 14519 16779
rect 14642 16776 14648 16788
rect 14507 16748 14648 16776
rect 14507 16745 14519 16748
rect 14461 16739 14519 16745
rect 14642 16736 14648 16748
rect 14700 16736 14706 16788
rect 15657 16779 15715 16785
rect 15657 16745 15669 16779
rect 15703 16776 15715 16779
rect 16942 16776 16948 16788
rect 15703 16748 16948 16776
rect 15703 16745 15715 16748
rect 15657 16739 15715 16745
rect 16942 16736 16948 16748
rect 17000 16736 17006 16788
rect 7070 16671 7128 16677
rect 7208 16680 8800 16708
rect 11517 16711 11575 16717
rect 4985 16643 5043 16649
rect 4985 16609 4997 16643
rect 5031 16640 5043 16643
rect 5261 16643 5319 16649
rect 5261 16640 5273 16643
rect 5031 16612 5273 16640
rect 5031 16609 5043 16612
rect 4985 16603 5043 16609
rect 5261 16609 5273 16612
rect 5307 16609 5319 16643
rect 5261 16603 5319 16609
rect 5442 16600 5448 16652
rect 5500 16640 5506 16652
rect 7208 16640 7236 16680
rect 11517 16677 11529 16711
rect 11563 16708 11575 16711
rect 12158 16708 12164 16720
rect 11563 16680 12164 16708
rect 11563 16677 11575 16680
rect 11517 16671 11575 16677
rect 12158 16668 12164 16680
rect 12216 16668 12222 16720
rect 12345 16711 12403 16717
rect 12345 16677 12357 16711
rect 12391 16708 12403 16711
rect 12526 16708 12532 16720
rect 12391 16680 12532 16708
rect 12391 16677 12403 16680
rect 12345 16671 12403 16677
rect 12526 16668 12532 16680
rect 12584 16668 12590 16720
rect 5500 16612 7236 16640
rect 5500 16600 5506 16612
rect 8294 16600 8300 16652
rect 8352 16640 8358 16652
rect 8573 16643 8631 16649
rect 8573 16640 8585 16643
rect 8352 16612 8585 16640
rect 8352 16600 8358 16612
rect 8573 16609 8585 16612
rect 8619 16609 8631 16643
rect 8938 16640 8944 16652
rect 8899 16612 8944 16640
rect 8573 16603 8631 16609
rect 8938 16600 8944 16612
rect 8996 16600 9002 16652
rect 9381 16643 9439 16649
rect 9381 16640 9393 16643
rect 9048 16612 9393 16640
rect 5353 16575 5411 16581
rect 5353 16541 5365 16575
rect 5399 16541 5411 16575
rect 5353 16535 5411 16541
rect 6825 16575 6883 16581
rect 6825 16541 6837 16575
rect 6871 16541 6883 16575
rect 6825 16535 6883 16541
rect 2774 16464 2780 16516
rect 2832 16464 2838 16516
rect 2406 16436 2412 16448
rect 2367 16408 2412 16436
rect 2406 16396 2412 16408
rect 2464 16396 2470 16448
rect 5368 16436 5396 16535
rect 6638 16464 6644 16516
rect 6696 16504 6702 16516
rect 6733 16507 6791 16513
rect 6733 16504 6745 16507
rect 6696 16476 6745 16504
rect 6696 16464 6702 16476
rect 6733 16473 6745 16476
rect 6779 16473 6791 16507
rect 6733 16467 6791 16473
rect 6362 16436 6368 16448
rect 5368 16408 6368 16436
rect 6362 16396 6368 16408
rect 6420 16436 6426 16448
rect 6840 16436 6868 16535
rect 8205 16507 8263 16513
rect 8205 16473 8217 16507
rect 8251 16504 8263 16507
rect 8846 16504 8852 16516
rect 8251 16476 8852 16504
rect 8251 16473 8263 16476
rect 8205 16467 8263 16473
rect 8846 16464 8852 16476
rect 8904 16504 8910 16516
rect 9048 16504 9076 16612
rect 9381 16609 9393 16612
rect 9427 16609 9439 16643
rect 9381 16603 9439 16609
rect 9950 16600 9956 16652
rect 10008 16640 10014 16652
rect 10410 16640 10416 16652
rect 10008 16612 10416 16640
rect 10008 16600 10014 16612
rect 10410 16600 10416 16612
rect 10468 16640 10474 16652
rect 10597 16643 10655 16649
rect 10597 16640 10609 16643
rect 10468 16612 10609 16640
rect 10468 16600 10474 16612
rect 10597 16609 10609 16612
rect 10643 16609 10655 16643
rect 10597 16603 10655 16609
rect 11698 16600 11704 16652
rect 11756 16640 11762 16652
rect 12253 16643 12311 16649
rect 12253 16640 12265 16643
rect 11756 16612 12265 16640
rect 11756 16600 11762 16612
rect 12253 16609 12265 16612
rect 12299 16609 12311 16643
rect 12253 16603 12311 16609
rect 13814 16600 13820 16652
rect 13872 16649 13878 16652
rect 13872 16640 13884 16649
rect 13872 16612 13917 16640
rect 13872 16603 13884 16612
rect 13872 16600 13878 16603
rect 14458 16600 14464 16652
rect 14516 16640 14522 16652
rect 14553 16643 14611 16649
rect 14553 16640 14565 16643
rect 14516 16612 14565 16640
rect 14516 16600 14522 16612
rect 14553 16609 14565 16612
rect 14599 16609 14611 16643
rect 14734 16640 14740 16652
rect 14695 16612 14740 16640
rect 14553 16603 14611 16609
rect 14734 16600 14740 16612
rect 14792 16600 14798 16652
rect 14921 16643 14979 16649
rect 14921 16609 14933 16643
rect 14967 16640 14979 16643
rect 15286 16640 15292 16652
rect 14967 16612 15292 16640
rect 14967 16609 14979 16612
rect 14921 16603 14979 16609
rect 15286 16600 15292 16612
rect 15344 16600 15350 16652
rect 15470 16640 15476 16652
rect 15431 16612 15476 16640
rect 15470 16600 15476 16612
rect 15528 16600 15534 16652
rect 9122 16532 9128 16584
rect 9180 16572 9186 16584
rect 11609 16575 11667 16581
rect 9180 16544 9225 16572
rect 9180 16532 9186 16544
rect 11609 16541 11621 16575
rect 11655 16572 11667 16575
rect 12437 16575 12495 16581
rect 12437 16572 12449 16575
rect 11655 16544 12449 16572
rect 11655 16541 11667 16544
rect 11609 16535 11667 16541
rect 12437 16541 12449 16544
rect 12483 16541 12495 16575
rect 12437 16535 12495 16541
rect 14093 16575 14151 16581
rect 14093 16541 14105 16575
rect 14139 16572 14151 16575
rect 14182 16572 14188 16584
rect 14139 16544 14188 16572
rect 14139 16541 14151 16544
rect 14093 16535 14151 16541
rect 11624 16504 11652 16535
rect 14182 16532 14188 16544
rect 14240 16532 14246 16584
rect 16022 16504 16028 16516
rect 8904 16476 9076 16504
rect 10520 16476 11652 16504
rect 14200 16476 16028 16504
rect 8904 16464 8910 16476
rect 10520 16448 10548 16476
rect 6420 16408 6868 16436
rect 6420 16396 6426 16408
rect 7006 16396 7012 16448
rect 7064 16436 7070 16448
rect 10042 16436 10048 16448
rect 7064 16408 10048 16436
rect 7064 16396 7070 16408
rect 10042 16396 10048 16408
rect 10100 16396 10106 16448
rect 10502 16436 10508 16448
rect 10463 16408 10508 16436
rect 10502 16396 10508 16408
rect 10560 16396 10566 16448
rect 10686 16396 10692 16448
rect 10744 16436 10750 16448
rect 10781 16439 10839 16445
rect 10781 16436 10793 16439
rect 10744 16408 10793 16436
rect 10744 16396 10750 16408
rect 10781 16405 10793 16408
rect 10827 16405 10839 16439
rect 11054 16436 11060 16448
rect 11015 16408 11060 16436
rect 10781 16399 10839 16405
rect 11054 16396 11060 16408
rect 11112 16396 11118 16448
rect 11146 16396 11152 16448
rect 11204 16436 11210 16448
rect 11885 16439 11943 16445
rect 11885 16436 11897 16439
rect 11204 16408 11897 16436
rect 11204 16396 11210 16408
rect 11885 16405 11897 16408
rect 11931 16405 11943 16439
rect 11885 16399 11943 16405
rect 12066 16396 12072 16448
rect 12124 16436 12130 16448
rect 13170 16436 13176 16448
rect 12124 16408 13176 16436
rect 12124 16396 12130 16408
rect 13170 16396 13176 16408
rect 13228 16396 13234 16448
rect 13354 16396 13360 16448
rect 13412 16436 13418 16448
rect 14200 16436 14228 16476
rect 16022 16464 16028 16476
rect 16080 16464 16086 16516
rect 15194 16436 15200 16448
rect 13412 16408 14228 16436
rect 15155 16408 15200 16436
rect 13412 16396 13418 16408
rect 15194 16396 15200 16408
rect 15252 16396 15258 16448
rect 1104 16346 16008 16368
rect 1104 16294 3480 16346
rect 3532 16294 3544 16346
rect 3596 16294 3608 16346
rect 3660 16294 3672 16346
rect 3724 16294 8478 16346
rect 8530 16294 8542 16346
rect 8594 16294 8606 16346
rect 8658 16294 8670 16346
rect 8722 16294 13475 16346
rect 13527 16294 13539 16346
rect 13591 16294 13603 16346
rect 13655 16294 13667 16346
rect 13719 16294 16008 16346
rect 1104 16272 16008 16294
rect 2409 16235 2467 16241
rect 2409 16201 2421 16235
rect 2455 16232 2467 16235
rect 2682 16232 2688 16244
rect 2455 16204 2688 16232
rect 2455 16201 2467 16204
rect 2409 16195 2467 16201
rect 2682 16192 2688 16204
rect 2740 16192 2746 16244
rect 2774 16192 2780 16244
rect 2832 16232 2838 16244
rect 2869 16235 2927 16241
rect 2869 16232 2881 16235
rect 2832 16204 2881 16232
rect 2832 16192 2838 16204
rect 2869 16201 2881 16204
rect 2915 16201 2927 16235
rect 2869 16195 2927 16201
rect 3145 16235 3203 16241
rect 3145 16201 3157 16235
rect 3191 16232 3203 16235
rect 3234 16232 3240 16244
rect 3191 16204 3240 16232
rect 3191 16201 3203 16204
rect 3145 16195 3203 16201
rect 3234 16192 3240 16204
rect 3292 16192 3298 16244
rect 3605 16235 3663 16241
rect 3605 16201 3617 16235
rect 3651 16232 3663 16235
rect 3786 16232 3792 16244
rect 3651 16204 3792 16232
rect 3651 16201 3663 16204
rect 3605 16195 3663 16201
rect 3786 16192 3792 16204
rect 3844 16192 3850 16244
rect 3881 16235 3939 16241
rect 3881 16201 3893 16235
rect 3927 16232 3939 16235
rect 3970 16232 3976 16244
rect 3927 16204 3976 16232
rect 3927 16201 3939 16204
rect 3881 16195 3939 16201
rect 3970 16192 3976 16204
rect 4028 16192 4034 16244
rect 4065 16235 4123 16241
rect 4065 16201 4077 16235
rect 4111 16232 4123 16235
rect 4246 16232 4252 16244
rect 4111 16204 4252 16232
rect 4111 16201 4123 16204
rect 4065 16195 4123 16201
rect 4246 16192 4252 16204
rect 4304 16232 4310 16244
rect 4709 16235 4767 16241
rect 4304 16204 4660 16232
rect 4304 16192 4310 16204
rect 1397 16167 1455 16173
rect 1397 16133 1409 16167
rect 1443 16164 1455 16167
rect 2958 16164 2964 16176
rect 1443 16136 2964 16164
rect 1443 16133 1455 16136
rect 1397 16127 1455 16133
rect 2958 16124 2964 16136
rect 3016 16124 3022 16176
rect 4154 16164 4160 16176
rect 3068 16136 4160 16164
rect 1949 16031 2007 16037
rect 1949 15997 1961 16031
rect 1995 16028 2007 16031
rect 2038 16028 2044 16040
rect 1995 16000 2044 16028
rect 1995 15997 2007 16000
rect 1949 15991 2007 15997
rect 2038 15988 2044 16000
rect 2096 15988 2102 16040
rect 2225 16031 2283 16037
rect 2225 15997 2237 16031
rect 2271 15997 2283 16031
rect 2225 15991 2283 15997
rect 2501 16031 2559 16037
rect 2501 15997 2513 16031
rect 2547 16028 2559 16031
rect 2958 16028 2964 16040
rect 2547 16000 2964 16028
rect 2547 15997 2559 16000
rect 2501 15991 2559 15997
rect 1581 15963 1639 15969
rect 1581 15929 1593 15963
rect 1627 15929 1639 15963
rect 1581 15923 1639 15929
rect 1596 15892 1624 15923
rect 1765 15895 1823 15901
rect 1765 15892 1777 15895
rect 1596 15864 1777 15892
rect 1765 15861 1777 15864
rect 1811 15861 1823 15895
rect 1765 15855 1823 15861
rect 2133 15895 2191 15901
rect 2133 15861 2145 15895
rect 2179 15892 2191 15895
rect 2240 15892 2268 15991
rect 2958 15988 2964 16000
rect 3016 15988 3022 16040
rect 3068 16037 3096 16136
rect 4154 16124 4160 16136
rect 4212 16124 4218 16176
rect 4632 16164 4660 16204
rect 4709 16201 4721 16235
rect 4755 16232 4767 16235
rect 4798 16232 4804 16244
rect 4755 16204 4804 16232
rect 4755 16201 4767 16204
rect 4709 16195 4767 16201
rect 4798 16192 4804 16204
rect 4856 16192 4862 16244
rect 5626 16232 5632 16244
rect 5587 16204 5632 16232
rect 5626 16192 5632 16204
rect 5684 16192 5690 16244
rect 5810 16192 5816 16244
rect 5868 16232 5874 16244
rect 5997 16235 6055 16241
rect 5997 16232 6009 16235
rect 5868 16204 6009 16232
rect 5868 16192 5874 16204
rect 5997 16201 6009 16204
rect 6043 16201 6055 16235
rect 5997 16195 6055 16201
rect 6273 16235 6331 16241
rect 6273 16201 6285 16235
rect 6319 16232 6331 16235
rect 6454 16232 6460 16244
rect 6319 16204 6460 16232
rect 6319 16201 6331 16204
rect 6273 16195 6331 16201
rect 6454 16192 6460 16204
rect 6512 16232 6518 16244
rect 7006 16232 7012 16244
rect 6512 16204 7012 16232
rect 6512 16192 6518 16204
rect 7006 16192 7012 16204
rect 7064 16192 7070 16244
rect 7098 16192 7104 16244
rect 7156 16232 7162 16244
rect 7285 16235 7343 16241
rect 7285 16232 7297 16235
rect 7156 16204 7297 16232
rect 7156 16192 7162 16204
rect 7285 16201 7297 16204
rect 7331 16201 7343 16235
rect 7285 16195 7343 16201
rect 7466 16192 7472 16244
rect 7524 16232 7530 16244
rect 7561 16235 7619 16241
rect 7561 16232 7573 16235
rect 7524 16204 7573 16232
rect 7524 16192 7530 16204
rect 7561 16201 7573 16204
rect 7607 16201 7619 16235
rect 7561 16195 7619 16201
rect 7742 16192 7748 16244
rect 7800 16232 7806 16244
rect 7837 16235 7895 16241
rect 7837 16232 7849 16235
rect 7800 16204 7849 16232
rect 7800 16192 7806 16204
rect 7837 16201 7849 16204
rect 7883 16201 7895 16235
rect 7837 16195 7895 16201
rect 8294 16192 8300 16244
rect 8352 16232 8358 16244
rect 8481 16235 8539 16241
rect 8481 16232 8493 16235
rect 8352 16204 8493 16232
rect 8352 16192 8358 16204
rect 8481 16201 8493 16204
rect 8527 16201 8539 16235
rect 9582 16232 9588 16244
rect 9543 16204 9588 16232
rect 8481 16195 8539 16201
rect 9582 16192 9588 16204
rect 9640 16192 9646 16244
rect 10318 16232 10324 16244
rect 9692 16204 10324 16232
rect 5905 16167 5963 16173
rect 4632 16136 5856 16164
rect 3234 16056 3240 16108
rect 3292 16096 3298 16108
rect 3292 16068 3740 16096
rect 3292 16056 3298 16068
rect 3053 16031 3111 16037
rect 3053 15997 3065 16031
rect 3099 15997 3111 16031
rect 3053 15991 3111 15997
rect 3329 16031 3387 16037
rect 3329 15997 3341 16031
rect 3375 15997 3387 16031
rect 3329 15991 3387 15997
rect 3344 15960 3372 15991
rect 3418 15988 3424 16040
rect 3476 16028 3482 16040
rect 3712 16037 3740 16068
rect 3970 16056 3976 16108
rect 4028 16096 4034 16108
rect 4341 16099 4399 16105
rect 4341 16096 4353 16099
rect 4028 16068 4353 16096
rect 4028 16056 4034 16068
rect 4341 16065 4353 16068
rect 4387 16065 4399 16099
rect 4341 16059 4399 16065
rect 3697 16031 3755 16037
rect 3476 16000 3521 16028
rect 3476 15988 3482 16000
rect 3697 15997 3709 16031
rect 3743 16028 3755 16031
rect 4525 16031 4583 16037
rect 4525 16028 4537 16031
rect 3743 16000 4537 16028
rect 3743 15997 3755 16000
rect 3697 15991 3755 15997
rect 4525 15997 4537 16000
rect 4571 15997 4583 16031
rect 4525 15991 4583 15997
rect 4893 16031 4951 16037
rect 4893 15997 4905 16031
rect 4939 16028 4951 16031
rect 5445 16031 5503 16037
rect 4939 16000 5120 16028
rect 4939 15997 4951 16000
rect 4893 15991 4951 15997
rect 3344 15932 4292 15960
rect 2590 15892 2596 15904
rect 2179 15864 2596 15892
rect 2179 15861 2191 15864
rect 2133 15855 2191 15861
rect 2590 15852 2596 15864
rect 2648 15852 2654 15904
rect 2685 15895 2743 15901
rect 2685 15861 2697 15895
rect 2731 15892 2743 15895
rect 2866 15892 2872 15904
rect 2731 15864 2872 15892
rect 2731 15861 2743 15864
rect 2685 15855 2743 15861
rect 2866 15852 2872 15864
rect 2924 15852 2930 15904
rect 3418 15852 3424 15904
rect 3476 15892 3482 15904
rect 3970 15892 3976 15904
rect 3476 15864 3976 15892
rect 3476 15852 3482 15864
rect 3970 15852 3976 15864
rect 4028 15852 4034 15904
rect 4264 15901 4292 15932
rect 5092 15904 5120 16000
rect 5445 15997 5457 16031
rect 5491 15997 5503 16031
rect 5718 16028 5724 16040
rect 5679 16000 5724 16028
rect 5445 15991 5503 15997
rect 4249 15895 4307 15901
rect 4249 15861 4261 15895
rect 4295 15892 4307 15895
rect 4338 15892 4344 15904
rect 4295 15864 4344 15892
rect 4295 15861 4307 15864
rect 4249 15855 4307 15861
rect 4338 15852 4344 15864
rect 4396 15852 4402 15904
rect 5074 15892 5080 15904
rect 5035 15864 5080 15892
rect 5074 15852 5080 15864
rect 5132 15852 5138 15904
rect 5353 15895 5411 15901
rect 5353 15861 5365 15895
rect 5399 15892 5411 15895
rect 5460 15892 5488 15991
rect 5718 15988 5724 16000
rect 5776 15988 5782 16040
rect 5828 15960 5856 16136
rect 5905 16133 5917 16167
rect 5951 16164 5963 16167
rect 6730 16164 6736 16176
rect 5951 16136 6736 16164
rect 5951 16133 5963 16136
rect 5905 16127 5963 16133
rect 6730 16124 6736 16136
rect 6788 16124 6794 16176
rect 8018 16124 8024 16176
rect 8076 16164 8082 16176
rect 8205 16167 8263 16173
rect 8205 16164 8217 16167
rect 8076 16136 8217 16164
rect 8076 16124 8082 16136
rect 8205 16133 8217 16136
rect 8251 16164 8263 16167
rect 9692 16164 9720 16204
rect 10318 16192 10324 16204
rect 10376 16192 10382 16244
rect 10870 16192 10876 16244
rect 10928 16232 10934 16244
rect 10928 16204 11836 16232
rect 10928 16192 10934 16204
rect 11698 16164 11704 16176
rect 8251 16136 9720 16164
rect 9876 16136 11704 16164
rect 8251 16133 8263 16136
rect 8205 16127 8263 16133
rect 6638 16056 6644 16108
rect 6696 16096 6702 16108
rect 7009 16099 7067 16105
rect 7009 16096 7021 16099
rect 6696 16068 7021 16096
rect 6696 16056 6702 16068
rect 7009 16065 7021 16068
rect 7055 16065 7067 16099
rect 7009 16059 7067 16065
rect 7650 16056 7656 16108
rect 7708 16096 7714 16108
rect 8846 16096 8852 16108
rect 7708 16068 8432 16096
rect 8807 16068 8852 16096
rect 7708 16056 7714 16068
rect 6181 16031 6239 16037
rect 6181 15997 6193 16031
rect 6227 16028 6239 16031
rect 6273 16031 6331 16037
rect 6273 16028 6285 16031
rect 6227 16000 6285 16028
rect 6227 15997 6239 16000
rect 6181 15991 6239 15997
rect 6273 15997 6285 16000
rect 6319 15997 6331 16031
rect 6273 15991 6331 15997
rect 6380 16000 7420 16028
rect 6380 15960 6408 16000
rect 5828 15932 6408 15960
rect 6825 15963 6883 15969
rect 6825 15929 6837 15963
rect 6871 15960 6883 15963
rect 7282 15960 7288 15972
rect 6871 15932 7288 15960
rect 6871 15929 6883 15932
rect 6825 15923 6883 15929
rect 7282 15920 7288 15932
rect 7340 15920 7346 15972
rect 7392 15960 7420 16000
rect 7466 15988 7472 16040
rect 7524 16028 7530 16040
rect 7745 16031 7803 16037
rect 7524 16000 7569 16028
rect 7524 15988 7530 16000
rect 7745 15997 7757 16031
rect 7791 16028 7803 16031
rect 7834 16028 7840 16040
rect 7791 16000 7840 16028
rect 7791 15997 7803 16000
rect 7745 15991 7803 15997
rect 7834 15988 7840 16000
rect 7892 15988 7898 16040
rect 8021 16031 8079 16037
rect 8021 15997 8033 16031
rect 8067 15997 8079 16031
rect 8294 16028 8300 16040
rect 8255 16000 8300 16028
rect 8021 15991 8079 15997
rect 7926 15960 7932 15972
rect 7392 15932 7932 15960
rect 7926 15920 7932 15932
rect 7984 15920 7990 15972
rect 8036 15960 8064 15991
rect 8294 15988 8300 16000
rect 8352 15988 8358 16040
rect 8404 16028 8432 16068
rect 8846 16056 8852 16068
rect 8904 16056 8910 16108
rect 9876 16105 9904 16136
rect 11698 16124 11704 16136
rect 11756 16124 11762 16176
rect 9861 16099 9919 16105
rect 9861 16065 9873 16099
rect 9907 16065 9919 16099
rect 9861 16059 9919 16065
rect 10137 16099 10195 16105
rect 10137 16065 10149 16099
rect 10183 16096 10195 16099
rect 10226 16096 10232 16108
rect 10183 16068 10232 16096
rect 10183 16065 10195 16068
rect 10137 16059 10195 16065
rect 10226 16056 10232 16068
rect 10284 16096 10290 16108
rect 10778 16096 10784 16108
rect 10284 16068 10784 16096
rect 10284 16056 10290 16068
rect 10778 16056 10784 16068
rect 10836 16096 10842 16108
rect 10873 16099 10931 16105
rect 10873 16096 10885 16099
rect 10836 16068 10885 16096
rect 10836 16056 10842 16068
rect 10873 16065 10885 16068
rect 10919 16065 10931 16099
rect 11054 16096 11060 16108
rect 11015 16068 11060 16096
rect 10873 16059 10931 16065
rect 11054 16056 11060 16068
rect 11112 16056 11118 16108
rect 11146 16028 11152 16040
rect 8404 16000 10364 16028
rect 11107 16000 11152 16028
rect 8754 15960 8760 15972
rect 8036 15932 8760 15960
rect 8754 15920 8760 15932
rect 8812 15920 8818 15972
rect 8941 15963 8999 15969
rect 8941 15929 8953 15963
rect 8987 15960 8999 15963
rect 9766 15960 9772 15972
rect 8987 15932 9772 15960
rect 8987 15929 8999 15932
rect 8941 15923 8999 15929
rect 9766 15920 9772 15932
rect 9824 15920 9830 15972
rect 9950 15920 9956 15972
rect 10008 15960 10014 15972
rect 10229 15963 10287 15969
rect 10229 15960 10241 15963
rect 10008 15932 10241 15960
rect 10008 15920 10014 15932
rect 10229 15929 10241 15932
rect 10275 15929 10287 15963
rect 10336 15960 10364 16000
rect 11146 15988 11152 16000
rect 11204 15988 11210 16040
rect 11698 15988 11704 16040
rect 11756 15988 11762 16040
rect 11808 16028 11836 16204
rect 11974 16192 11980 16244
rect 12032 16232 12038 16244
rect 12032 16204 13216 16232
rect 12032 16192 12038 16204
rect 13188 16164 13216 16204
rect 13262 16192 13268 16244
rect 13320 16232 13326 16244
rect 13633 16235 13691 16241
rect 13633 16232 13645 16235
rect 13320 16204 13645 16232
rect 13320 16192 13326 16204
rect 13633 16201 13645 16204
rect 13679 16201 13691 16235
rect 15746 16232 15752 16244
rect 13633 16195 13691 16201
rect 13740 16204 15752 16232
rect 13740 16164 13768 16204
rect 15746 16192 15752 16204
rect 15804 16192 15810 16244
rect 13188 16136 13768 16164
rect 12084 16068 12296 16096
rect 11885 16031 11943 16037
rect 11885 16028 11897 16031
rect 11808 16000 11897 16028
rect 11885 15997 11897 16000
rect 11931 15997 11943 16031
rect 11885 15991 11943 15997
rect 11606 15960 11612 15972
rect 10336 15932 11612 15960
rect 10229 15923 10287 15929
rect 11606 15920 11612 15932
rect 11664 15920 11670 15972
rect 11716 15960 11744 15988
rect 12084 15960 12112 16068
rect 12161 16031 12219 16037
rect 12161 15997 12173 16031
rect 12207 15997 12219 16031
rect 12268 16028 12296 16068
rect 13354 16028 13360 16040
rect 12268 16000 13360 16028
rect 12161 15991 12219 15997
rect 11716 15932 12112 15960
rect 5626 15892 5632 15904
rect 5399 15864 5632 15892
rect 5399 15861 5411 15864
rect 5353 15855 5411 15861
rect 5626 15852 5632 15864
rect 5684 15852 5690 15904
rect 5810 15852 5816 15904
rect 5868 15892 5874 15904
rect 6457 15895 6515 15901
rect 6457 15892 6469 15895
rect 5868 15864 6469 15892
rect 5868 15852 5874 15864
rect 6457 15861 6469 15864
rect 6503 15861 6515 15895
rect 6457 15855 6515 15861
rect 6917 15895 6975 15901
rect 6917 15861 6929 15895
rect 6963 15892 6975 15895
rect 7190 15892 7196 15904
rect 6963 15864 7196 15892
rect 6963 15861 6975 15864
rect 6917 15855 6975 15861
rect 7190 15852 7196 15864
rect 7248 15852 7254 15904
rect 9033 15895 9091 15901
rect 9033 15861 9045 15895
rect 9079 15892 9091 15895
rect 9214 15892 9220 15904
rect 9079 15864 9220 15892
rect 9079 15861 9091 15864
rect 9033 15855 9091 15861
rect 9214 15852 9220 15864
rect 9272 15852 9278 15904
rect 9398 15892 9404 15904
rect 9359 15864 9404 15892
rect 9398 15852 9404 15864
rect 9456 15852 9462 15904
rect 10318 15892 10324 15904
rect 10279 15864 10324 15892
rect 10318 15852 10324 15864
rect 10376 15852 10382 15904
rect 10689 15895 10747 15901
rect 10689 15861 10701 15895
rect 10735 15892 10747 15895
rect 11330 15892 11336 15904
rect 10735 15864 11336 15892
rect 10735 15861 10747 15864
rect 10689 15855 10747 15861
rect 11330 15852 11336 15864
rect 11388 15852 11394 15904
rect 11517 15895 11575 15901
rect 11517 15861 11529 15895
rect 11563 15892 11575 15895
rect 11698 15892 11704 15904
rect 11563 15864 11704 15892
rect 11563 15861 11575 15864
rect 11517 15855 11575 15861
rect 11698 15852 11704 15864
rect 11756 15852 11762 15904
rect 11793 15895 11851 15901
rect 11793 15861 11805 15895
rect 11839 15892 11851 15895
rect 12066 15892 12072 15904
rect 11839 15864 12072 15892
rect 11839 15861 11851 15864
rect 11793 15855 11851 15861
rect 12066 15852 12072 15864
rect 12124 15852 12130 15904
rect 12176 15892 12204 15991
rect 13354 15988 13360 16000
rect 13412 15988 13418 16040
rect 13817 16031 13875 16037
rect 13817 15997 13829 16031
rect 13863 15997 13875 16031
rect 13817 15991 13875 15997
rect 12428 15963 12486 15969
rect 12428 15929 12440 15963
rect 12474 15960 12486 15963
rect 12526 15960 12532 15972
rect 12474 15932 12532 15960
rect 12474 15929 12486 15932
rect 12428 15923 12486 15929
rect 12526 15920 12532 15932
rect 12584 15920 12590 15972
rect 12802 15960 12808 15972
rect 12636 15932 12808 15960
rect 12636 15892 12664 15932
rect 12802 15920 12808 15932
rect 12860 15960 12866 15972
rect 13832 15960 13860 15991
rect 13906 15988 13912 16040
rect 13964 16028 13970 16040
rect 14073 16031 14131 16037
rect 14073 16028 14085 16031
rect 13964 16000 14085 16028
rect 13964 15988 13970 16000
rect 14073 15997 14085 16000
rect 14119 15997 14131 16031
rect 14073 15991 14131 15997
rect 14918 15988 14924 16040
rect 14976 16028 14982 16040
rect 15473 16031 15531 16037
rect 15473 16028 15485 16031
rect 14976 16000 15485 16028
rect 14976 15988 14982 16000
rect 15473 15997 15485 16000
rect 15519 15997 15531 16031
rect 15473 15991 15531 15997
rect 14182 15960 14188 15972
rect 12860 15932 14188 15960
rect 12860 15920 12866 15932
rect 14182 15920 14188 15932
rect 14240 15920 14246 15972
rect 15286 15960 15292 15972
rect 15247 15932 15292 15960
rect 15286 15920 15292 15932
rect 15344 15920 15350 15972
rect 12176 15864 12664 15892
rect 13541 15895 13599 15901
rect 13541 15861 13553 15895
rect 13587 15892 13599 15895
rect 13814 15892 13820 15904
rect 13587 15864 13820 15892
rect 13587 15861 13599 15864
rect 13541 15855 13599 15861
rect 13814 15852 13820 15864
rect 13872 15852 13878 15904
rect 14366 15852 14372 15904
rect 14424 15892 14430 15904
rect 15010 15892 15016 15904
rect 14424 15864 15016 15892
rect 14424 15852 14430 15864
rect 15010 15852 15016 15864
rect 15068 15892 15074 15904
rect 15197 15895 15255 15901
rect 15197 15892 15209 15895
rect 15068 15864 15209 15892
rect 15068 15852 15074 15864
rect 15197 15861 15209 15864
rect 15243 15861 15255 15895
rect 15197 15855 15255 15861
rect 1104 15802 16008 15824
rect 1104 15750 5979 15802
rect 6031 15750 6043 15802
rect 6095 15750 6107 15802
rect 6159 15750 6171 15802
rect 6223 15750 10976 15802
rect 11028 15750 11040 15802
rect 11092 15750 11104 15802
rect 11156 15750 11168 15802
rect 11220 15750 16008 15802
rect 1104 15728 16008 15750
rect 1486 15688 1492 15700
rect 1447 15660 1492 15688
rect 1486 15648 1492 15660
rect 1544 15648 1550 15700
rect 1765 15691 1823 15697
rect 1765 15688 1777 15691
rect 1596 15660 1777 15688
rect 1596 15629 1624 15660
rect 1765 15657 1777 15660
rect 1811 15657 1823 15691
rect 1765 15651 1823 15657
rect 1946 15648 1952 15700
rect 2004 15688 2010 15700
rect 2317 15691 2375 15697
rect 2317 15688 2329 15691
rect 2004 15660 2329 15688
rect 2004 15648 2010 15660
rect 2317 15657 2329 15660
rect 2363 15657 2375 15691
rect 2317 15651 2375 15657
rect 2746 15660 4936 15688
rect 1581 15623 1639 15629
rect 1581 15589 1593 15623
rect 1627 15589 1639 15623
rect 2746 15620 2774 15660
rect 1581 15583 1639 15589
rect 2240 15592 2774 15620
rect 1949 15555 2007 15561
rect 1949 15521 1961 15555
rect 1995 15552 2007 15555
rect 2130 15552 2136 15564
rect 1995 15524 2136 15552
rect 1995 15521 2007 15524
rect 1949 15515 2007 15521
rect 2130 15512 2136 15524
rect 2188 15512 2194 15564
rect 2240 15561 2268 15592
rect 3142 15580 3148 15632
rect 3200 15620 3206 15632
rect 3329 15623 3387 15629
rect 3329 15620 3341 15623
rect 3200 15592 3341 15620
rect 3200 15580 3206 15592
rect 3329 15589 3341 15592
rect 3375 15589 3387 15623
rect 4908 15620 4936 15660
rect 5074 15648 5080 15700
rect 5132 15688 5138 15700
rect 7006 15688 7012 15700
rect 5132 15660 7012 15688
rect 5132 15648 5138 15660
rect 7006 15648 7012 15660
rect 7064 15648 7070 15700
rect 7190 15688 7196 15700
rect 7151 15660 7196 15688
rect 7190 15648 7196 15660
rect 7248 15648 7254 15700
rect 7282 15648 7288 15700
rect 7340 15688 7346 15700
rect 7340 15660 7385 15688
rect 7340 15648 7346 15660
rect 7466 15648 7472 15700
rect 7524 15688 7530 15700
rect 8113 15691 8171 15697
rect 8113 15688 8125 15691
rect 7524 15660 8125 15688
rect 7524 15648 7530 15660
rect 8113 15657 8125 15660
rect 8159 15657 8171 15691
rect 8113 15651 8171 15657
rect 8294 15648 8300 15700
rect 8352 15688 8358 15700
rect 9030 15688 9036 15700
rect 8352 15660 9036 15688
rect 8352 15648 8358 15660
rect 9030 15648 9036 15660
rect 9088 15648 9094 15700
rect 9398 15648 9404 15700
rect 9456 15688 9462 15700
rect 9493 15691 9551 15697
rect 9493 15688 9505 15691
rect 9456 15660 9505 15688
rect 9456 15648 9462 15660
rect 9493 15657 9505 15660
rect 9539 15657 9551 15691
rect 9950 15688 9956 15700
rect 9911 15660 9956 15688
rect 9493 15651 9551 15657
rect 9950 15648 9956 15660
rect 10008 15648 10014 15700
rect 10318 15688 10324 15700
rect 10279 15660 10324 15688
rect 10318 15648 10324 15660
rect 10376 15648 10382 15700
rect 10686 15648 10692 15700
rect 10744 15688 10750 15700
rect 10781 15691 10839 15697
rect 10781 15688 10793 15691
rect 10744 15660 10793 15688
rect 10744 15648 10750 15660
rect 10781 15657 10793 15660
rect 10827 15657 10839 15691
rect 10781 15651 10839 15657
rect 11149 15691 11207 15697
rect 11149 15657 11161 15691
rect 11195 15657 11207 15691
rect 11149 15651 11207 15657
rect 11517 15691 11575 15697
rect 11517 15657 11529 15691
rect 11563 15688 11575 15691
rect 11698 15688 11704 15700
rect 11563 15660 11704 15688
rect 11563 15657 11575 15660
rect 11517 15651 11575 15657
rect 11164 15620 11192 15651
rect 11698 15648 11704 15660
rect 11756 15648 11762 15700
rect 12526 15688 12532 15700
rect 12406 15660 12532 15688
rect 4908 15592 11192 15620
rect 3329 15583 3387 15589
rect 11330 15580 11336 15632
rect 11388 15620 11394 15632
rect 11609 15623 11667 15629
rect 11609 15620 11621 15623
rect 11388 15592 11621 15620
rect 11388 15580 11394 15592
rect 11609 15589 11621 15592
rect 11655 15589 11667 15623
rect 12406 15620 12434 15660
rect 12526 15648 12532 15660
rect 12584 15648 12590 15700
rect 12897 15691 12955 15697
rect 12897 15657 12909 15691
rect 12943 15688 12955 15691
rect 13357 15691 13415 15697
rect 13357 15688 13369 15691
rect 12943 15660 13369 15688
rect 12943 15657 12955 15660
rect 12897 15651 12955 15657
rect 13357 15657 13369 15660
rect 13403 15657 13415 15691
rect 13357 15651 13415 15657
rect 13722 15648 13728 15700
rect 13780 15688 13786 15700
rect 13998 15688 14004 15700
rect 13780 15660 14004 15688
rect 13780 15648 13786 15660
rect 13998 15648 14004 15660
rect 14056 15688 14062 15700
rect 14645 15691 14703 15697
rect 14645 15688 14657 15691
rect 14056 15660 14657 15688
rect 14056 15648 14062 15660
rect 14645 15657 14657 15660
rect 14691 15657 14703 15691
rect 14645 15651 14703 15657
rect 13262 15620 13268 15632
rect 11609 15583 11667 15589
rect 12360 15592 13268 15620
rect 2225 15555 2283 15561
rect 2225 15521 2237 15555
rect 2271 15521 2283 15555
rect 2498 15552 2504 15564
rect 2459 15524 2504 15552
rect 2225 15515 2283 15521
rect 2498 15512 2504 15524
rect 2556 15512 2562 15564
rect 2593 15555 2651 15561
rect 2593 15521 2605 15555
rect 2639 15552 2651 15555
rect 2869 15555 2927 15561
rect 2639 15524 2673 15552
rect 2639 15521 2651 15524
rect 2593 15515 2651 15521
rect 2869 15521 2881 15555
rect 2915 15552 2927 15555
rect 3160 15552 3188 15580
rect 2915 15524 3188 15552
rect 5925 15555 5983 15561
rect 2915 15521 2927 15524
rect 2869 15515 2927 15521
rect 5925 15521 5937 15555
rect 5971 15552 5983 15555
rect 6086 15552 6092 15564
rect 5971 15524 6092 15552
rect 5971 15521 5983 15524
rect 5925 15515 5983 15521
rect 2608 15484 2636 15515
rect 6086 15512 6092 15524
rect 6144 15512 6150 15564
rect 6181 15555 6239 15561
rect 6181 15521 6193 15555
rect 6227 15552 6239 15555
rect 6270 15552 6276 15564
rect 6227 15524 6276 15552
rect 6227 15521 6239 15524
rect 6181 15515 6239 15521
rect 6270 15512 6276 15524
rect 6328 15512 6334 15564
rect 6365 15555 6423 15561
rect 6365 15521 6377 15555
rect 6411 15552 6423 15555
rect 6454 15552 6460 15564
rect 6411 15524 6460 15552
rect 6411 15521 6423 15524
rect 6365 15515 6423 15521
rect 6454 15512 6460 15524
rect 6512 15512 6518 15564
rect 6822 15552 6828 15564
rect 6783 15524 6828 15552
rect 6822 15512 6828 15524
rect 6880 15512 6886 15564
rect 7653 15555 7711 15561
rect 7653 15521 7665 15555
rect 7699 15552 7711 15555
rect 8294 15552 8300 15564
rect 7699 15524 8300 15552
rect 7699 15521 7711 15524
rect 7653 15515 7711 15521
rect 8294 15512 8300 15524
rect 8352 15512 8358 15564
rect 8754 15552 8760 15564
rect 8715 15524 8760 15552
rect 8754 15512 8760 15524
rect 8812 15552 8818 15564
rect 9125 15555 9183 15561
rect 9125 15552 9137 15555
rect 8812 15524 9137 15552
rect 8812 15512 8818 15524
rect 9125 15521 9137 15524
rect 9171 15521 9183 15555
rect 9125 15515 9183 15521
rect 9306 15512 9312 15564
rect 9364 15552 9370 15564
rect 9585 15555 9643 15561
rect 9585 15552 9597 15555
rect 9364 15524 9597 15552
rect 9364 15512 9370 15524
rect 9585 15521 9597 15524
rect 9631 15521 9643 15555
rect 9585 15515 9643 15521
rect 9858 15512 9864 15564
rect 9916 15552 9922 15564
rect 10689 15555 10747 15561
rect 10689 15552 10701 15555
rect 9916 15524 10701 15552
rect 9916 15512 9922 15524
rect 10689 15521 10701 15524
rect 10735 15552 10747 15555
rect 10778 15552 10784 15564
rect 10735 15524 10784 15552
rect 10735 15521 10747 15524
rect 10689 15515 10747 15521
rect 10778 15512 10784 15524
rect 10836 15512 10842 15564
rect 3145 15487 3203 15493
rect 3145 15484 3157 15487
rect 2424 15456 3157 15484
rect 1578 15376 1584 15428
rect 1636 15416 1642 15428
rect 2041 15419 2099 15425
rect 2041 15416 2053 15419
rect 1636 15388 2053 15416
rect 1636 15376 1642 15388
rect 2041 15385 2053 15388
rect 2087 15385 2099 15419
rect 2041 15379 2099 15385
rect 198 15308 204 15360
rect 256 15348 262 15360
rect 2424 15348 2452 15456
rect 3145 15453 3157 15456
rect 3191 15453 3203 15487
rect 6549 15487 6607 15493
rect 6549 15484 6561 15487
rect 3145 15447 3203 15453
rect 6196 15456 6561 15484
rect 4709 15419 4767 15425
rect 4709 15385 4721 15419
rect 4755 15416 4767 15419
rect 4890 15416 4896 15428
rect 4755 15388 4896 15416
rect 4755 15385 4767 15388
rect 4709 15379 4767 15385
rect 4890 15376 4896 15388
rect 4948 15376 4954 15428
rect 256 15320 2452 15348
rect 256 15308 262 15320
rect 2774 15308 2780 15360
rect 2832 15348 2838 15360
rect 3053 15351 3111 15357
rect 2832 15320 2877 15348
rect 2832 15308 2838 15320
rect 3053 15317 3065 15351
rect 3099 15348 3111 15351
rect 3326 15348 3332 15360
rect 3099 15320 3332 15348
rect 3099 15317 3111 15320
rect 3053 15311 3111 15317
rect 3326 15308 3332 15320
rect 3384 15308 3390 15360
rect 3605 15351 3663 15357
rect 3605 15317 3617 15351
rect 3651 15348 3663 15351
rect 4154 15348 4160 15360
rect 3651 15320 4160 15348
rect 3651 15317 3663 15320
rect 3605 15311 3663 15317
rect 4154 15308 4160 15320
rect 4212 15348 4218 15360
rect 4614 15348 4620 15360
rect 4212 15320 4620 15348
rect 4212 15308 4218 15320
rect 4614 15308 4620 15320
rect 4672 15308 4678 15360
rect 4801 15351 4859 15357
rect 4801 15317 4813 15351
rect 4847 15348 4859 15351
rect 5534 15348 5540 15360
rect 4847 15320 5540 15348
rect 4847 15317 4859 15320
rect 4801 15311 4859 15317
rect 5534 15308 5540 15320
rect 5592 15348 5598 15360
rect 6196 15348 6224 15456
rect 6549 15453 6561 15456
rect 6595 15453 6607 15487
rect 6730 15484 6736 15496
rect 6691 15456 6736 15484
rect 6549 15447 6607 15453
rect 6564 15416 6592 15447
rect 6730 15444 6736 15456
rect 6788 15444 6794 15496
rect 7742 15484 7748 15496
rect 7703 15456 7748 15484
rect 7742 15444 7748 15456
rect 7800 15444 7806 15496
rect 7837 15487 7895 15493
rect 7837 15453 7849 15487
rect 7883 15453 7895 15487
rect 7837 15447 7895 15453
rect 8481 15487 8539 15493
rect 8481 15453 8493 15487
rect 8527 15484 8539 15487
rect 8938 15484 8944 15496
rect 8527 15456 8944 15484
rect 8527 15453 8539 15456
rect 8481 15447 8539 15453
rect 7852 15416 7880 15447
rect 8938 15444 8944 15456
rect 8996 15444 9002 15496
rect 9401 15487 9459 15493
rect 9401 15453 9413 15487
rect 9447 15484 9459 15487
rect 10502 15484 10508 15496
rect 9447 15456 10508 15484
rect 9447 15453 9459 15456
rect 9401 15447 9459 15453
rect 10502 15444 10508 15456
rect 10560 15484 10566 15496
rect 10873 15487 10931 15493
rect 10873 15484 10885 15487
rect 10560 15456 10885 15484
rect 10560 15444 10566 15456
rect 10873 15453 10885 15456
rect 10919 15453 10931 15487
rect 10873 15447 10931 15453
rect 11698 15444 11704 15496
rect 11756 15484 11762 15496
rect 12360 15493 12388 15592
rect 13262 15580 13268 15592
rect 13320 15620 13326 15632
rect 15473 15623 15531 15629
rect 13320 15592 14412 15620
rect 13320 15580 13326 15592
rect 12529 15555 12587 15561
rect 12529 15521 12541 15555
rect 12575 15552 12587 15555
rect 12894 15552 12900 15564
rect 12575 15524 12900 15552
rect 12575 15521 12587 15524
rect 12529 15515 12587 15521
rect 12894 15512 12900 15524
rect 12952 15512 12958 15564
rect 13170 15512 13176 15564
rect 13228 15552 13234 15564
rect 13998 15552 14004 15564
rect 13228 15524 14004 15552
rect 13228 15512 13234 15524
rect 13998 15512 14004 15524
rect 14056 15512 14062 15564
rect 12345 15487 12403 15493
rect 11756 15456 11801 15484
rect 11756 15444 11762 15456
rect 12345 15453 12357 15487
rect 12391 15453 12403 15487
rect 12345 15447 12403 15453
rect 12434 15444 12440 15496
rect 12492 15484 12498 15496
rect 12492 15456 12537 15484
rect 12492 15444 12498 15456
rect 13078 15444 13084 15496
rect 13136 15484 13142 15496
rect 13449 15487 13507 15493
rect 13449 15484 13461 15487
rect 13136 15456 13461 15484
rect 13136 15444 13142 15456
rect 13449 15453 13461 15456
rect 13495 15453 13507 15487
rect 13449 15447 13507 15453
rect 13633 15487 13691 15493
rect 13633 15453 13645 15487
rect 13679 15484 13691 15487
rect 13814 15484 13820 15496
rect 13679 15456 13820 15484
rect 13679 15453 13691 15456
rect 13633 15447 13691 15453
rect 13814 15444 13820 15456
rect 13872 15484 13878 15496
rect 14274 15484 14280 15496
rect 13872 15456 14280 15484
rect 13872 15444 13878 15456
rect 14274 15444 14280 15456
rect 14332 15444 14338 15496
rect 14384 15484 14412 15592
rect 15473 15589 15485 15623
rect 15519 15620 15531 15623
rect 15654 15620 15660 15632
rect 15519 15592 15660 15620
rect 15519 15589 15531 15592
rect 15473 15583 15531 15589
rect 14737 15555 14795 15561
rect 14737 15521 14749 15555
rect 14783 15552 14795 15555
rect 15010 15552 15016 15564
rect 14783 15524 15016 15552
rect 14783 15521 14795 15524
rect 14737 15515 14795 15521
rect 15010 15512 15016 15524
rect 15068 15512 15074 15564
rect 14461 15487 14519 15493
rect 14461 15484 14473 15487
rect 14384 15456 14473 15484
rect 14461 15453 14473 15456
rect 14507 15453 14519 15487
rect 14461 15447 14519 15453
rect 15102 15444 15108 15496
rect 15160 15484 15166 15496
rect 15289 15487 15347 15493
rect 15289 15484 15301 15487
rect 15160 15456 15301 15484
rect 15160 15444 15166 15456
rect 15289 15453 15301 15456
rect 15335 15453 15347 15487
rect 15289 15447 15347 15453
rect 6564 15388 7880 15416
rect 7926 15376 7932 15428
rect 7984 15416 7990 15428
rect 10594 15416 10600 15428
rect 7984 15388 10600 15416
rect 7984 15376 7990 15388
rect 10594 15376 10600 15388
rect 10652 15376 10658 15428
rect 12986 15416 12992 15428
rect 12947 15388 12992 15416
rect 12986 15376 12992 15388
rect 13044 15376 13050 15428
rect 15488 15416 15516 15583
rect 15654 15580 15660 15592
rect 15712 15580 15718 15632
rect 13740 15388 15516 15416
rect 5592 15320 6224 15348
rect 5592 15308 5598 15320
rect 7834 15308 7840 15360
rect 7892 15348 7898 15360
rect 8573 15351 8631 15357
rect 8573 15348 8585 15351
rect 7892 15320 8585 15348
rect 7892 15308 7898 15320
rect 8573 15317 8585 15320
rect 8619 15317 8631 15351
rect 8573 15311 8631 15317
rect 9125 15351 9183 15357
rect 9125 15317 9137 15351
rect 9171 15348 9183 15351
rect 10134 15348 10140 15360
rect 9171 15320 10140 15348
rect 9171 15317 9183 15320
rect 9125 15311 9183 15317
rect 10134 15308 10140 15320
rect 10192 15308 10198 15360
rect 10229 15351 10287 15357
rect 10229 15317 10241 15351
rect 10275 15348 10287 15351
rect 11790 15348 11796 15360
rect 10275 15320 11796 15348
rect 10275 15317 10287 15320
rect 10229 15311 10287 15317
rect 11790 15308 11796 15320
rect 11848 15308 11854 15360
rect 12069 15351 12127 15357
rect 12069 15317 12081 15351
rect 12115 15348 12127 15351
rect 13740 15348 13768 15388
rect 13906 15348 13912 15360
rect 12115 15320 13768 15348
rect 13867 15320 13912 15348
rect 12115 15317 12127 15320
rect 12069 15311 12127 15317
rect 13906 15308 13912 15320
rect 13964 15308 13970 15360
rect 15105 15351 15163 15357
rect 15105 15317 15117 15351
rect 15151 15348 15163 15351
rect 15286 15348 15292 15360
rect 15151 15320 15292 15348
rect 15151 15317 15163 15320
rect 15105 15311 15163 15317
rect 15286 15308 15292 15320
rect 15344 15308 15350 15360
rect 1104 15258 16008 15280
rect 1104 15206 3480 15258
rect 3532 15206 3544 15258
rect 3596 15206 3608 15258
rect 3660 15206 3672 15258
rect 3724 15206 8478 15258
rect 8530 15206 8542 15258
rect 8594 15206 8606 15258
rect 8658 15206 8670 15258
rect 8722 15206 13475 15258
rect 13527 15206 13539 15258
rect 13591 15206 13603 15258
rect 13655 15206 13667 15258
rect 13719 15206 16008 15258
rect 1104 15184 16008 15206
rect 1949 15147 2007 15153
rect 1949 15113 1961 15147
rect 1995 15144 2007 15147
rect 2222 15144 2228 15156
rect 1995 15116 2228 15144
rect 1995 15113 2007 15116
rect 1949 15107 2007 15113
rect 2222 15104 2228 15116
rect 2280 15104 2286 15156
rect 2866 15104 2872 15156
rect 2924 15144 2930 15156
rect 4062 15144 4068 15156
rect 2924 15116 4068 15144
rect 2924 15104 2930 15116
rect 4062 15104 4068 15116
rect 4120 15104 4126 15156
rect 6362 15144 6368 15156
rect 4448 15116 6368 15144
rect 2958 15076 2964 15088
rect 1780 15048 2964 15076
rect 1780 14949 1808 15048
rect 2958 15036 2964 15048
rect 3016 15036 3022 15088
rect 3329 15079 3387 15085
rect 3329 15045 3341 15079
rect 3375 15045 3387 15079
rect 3329 15039 3387 15045
rect 2774 15008 2780 15020
rect 2735 14980 2780 15008
rect 2774 14968 2780 14980
rect 2832 14968 2838 15020
rect 3142 15008 3148 15020
rect 3103 14980 3148 15008
rect 3142 14968 3148 14980
rect 3200 14968 3206 15020
rect 1765 14943 1823 14949
rect 1765 14909 1777 14943
rect 1811 14909 1823 14943
rect 1765 14903 1823 14909
rect 1578 14872 1584 14884
rect 1539 14844 1584 14872
rect 1578 14832 1584 14844
rect 1636 14832 1642 14884
rect 2501 14875 2559 14881
rect 2501 14841 2513 14875
rect 2547 14872 2559 14875
rect 3344 14872 3372 15039
rect 3786 15036 3792 15088
rect 3844 15076 3850 15088
rect 4448 15076 4476 15116
rect 6362 15104 6368 15116
rect 6420 15104 6426 15156
rect 6733 15147 6791 15153
rect 6733 15113 6745 15147
rect 6779 15144 6791 15147
rect 6822 15144 6828 15156
rect 6779 15116 6828 15144
rect 6779 15113 6791 15116
rect 6733 15107 6791 15113
rect 6822 15104 6828 15116
rect 6880 15104 6886 15156
rect 7742 15144 7748 15156
rect 7703 15116 7748 15144
rect 7742 15104 7748 15116
rect 7800 15104 7806 15156
rect 8294 15104 8300 15156
rect 8352 15144 8358 15156
rect 8573 15147 8631 15153
rect 8573 15144 8585 15147
rect 8352 15116 8585 15144
rect 8352 15104 8358 15116
rect 8573 15113 8585 15116
rect 8619 15113 8631 15147
rect 8573 15107 8631 15113
rect 9122 15104 9128 15156
rect 9180 15144 9186 15156
rect 9861 15147 9919 15153
rect 9180 15116 9720 15144
rect 9180 15104 9186 15116
rect 9692 15088 9720 15116
rect 9861 15113 9873 15147
rect 9907 15144 9919 15147
rect 10870 15144 10876 15156
rect 9907 15116 10876 15144
rect 9907 15113 9919 15116
rect 9861 15107 9919 15113
rect 10870 15104 10876 15116
rect 10928 15104 10934 15156
rect 11333 15147 11391 15153
rect 11333 15113 11345 15147
rect 11379 15144 11391 15147
rect 11698 15144 11704 15156
rect 11379 15116 11704 15144
rect 11379 15113 11391 15116
rect 11333 15107 11391 15113
rect 11698 15104 11704 15116
rect 11756 15104 11762 15156
rect 12434 15104 12440 15156
rect 12492 15144 12498 15156
rect 12897 15147 12955 15153
rect 12897 15144 12909 15147
rect 12492 15116 12909 15144
rect 12492 15104 12498 15116
rect 12897 15113 12909 15116
rect 12943 15113 12955 15147
rect 12897 15107 12955 15113
rect 12989 15147 13047 15153
rect 12989 15113 13001 15147
rect 13035 15144 13047 15147
rect 13078 15144 13084 15156
rect 13035 15116 13084 15144
rect 13035 15113 13047 15116
rect 12989 15107 13047 15113
rect 13078 15104 13084 15116
rect 13136 15104 13142 15156
rect 14001 15147 14059 15153
rect 14001 15113 14013 15147
rect 14047 15144 14059 15147
rect 14090 15144 14096 15156
rect 14047 15116 14096 15144
rect 14047 15113 14059 15116
rect 14001 15107 14059 15113
rect 14090 15104 14096 15116
rect 14148 15104 14154 15156
rect 14921 15147 14979 15153
rect 14921 15144 14933 15147
rect 14200 15116 14933 15144
rect 3844 15048 4476 15076
rect 3844 15036 3850 15048
rect 3878 15008 3884 15020
rect 3839 14980 3884 15008
rect 3878 14968 3884 14980
rect 3936 14968 3942 15020
rect 4448 15017 4476 15048
rect 5813 15079 5871 15085
rect 5813 15045 5825 15079
rect 5859 15076 5871 15079
rect 6270 15076 6276 15088
rect 5859 15048 6276 15076
rect 5859 15045 5871 15048
rect 5813 15039 5871 15045
rect 6270 15036 6276 15048
rect 6328 15036 6334 15088
rect 7098 15036 7104 15088
rect 7156 15076 7162 15088
rect 7653 15079 7711 15085
rect 7653 15076 7665 15079
rect 7156 15048 7665 15076
rect 7156 15036 7162 15048
rect 7653 15045 7665 15048
rect 7699 15076 7711 15079
rect 9582 15076 9588 15088
rect 7699 15048 9588 15076
rect 7699 15045 7711 15048
rect 7653 15039 7711 15045
rect 9582 15036 9588 15048
rect 9640 15036 9646 15088
rect 9674 15036 9680 15088
rect 9732 15076 9738 15088
rect 11517 15079 11575 15085
rect 9732 15048 9996 15076
rect 9732 15036 9738 15048
rect 4433 15011 4491 15017
rect 4433 14977 4445 15011
rect 4479 14977 4491 15011
rect 4433 14971 4491 14977
rect 6086 14968 6092 15020
rect 6144 15008 6150 15020
rect 7282 15008 7288 15020
rect 6144 14980 7288 15008
rect 6144 14968 6150 14980
rect 7282 14968 7288 14980
rect 7340 15008 7346 15020
rect 9968 15017 9996 15048
rect 11517 15045 11529 15079
rect 11563 15076 11575 15079
rect 11974 15076 11980 15088
rect 11563 15048 11980 15076
rect 11563 15045 11575 15048
rect 11517 15039 11575 15045
rect 11974 15036 11980 15048
rect 12032 15036 12038 15088
rect 12710 15036 12716 15088
rect 12768 15076 12774 15088
rect 14200 15076 14228 15116
rect 14921 15113 14933 15116
rect 14967 15113 14979 15147
rect 16114 15144 16120 15156
rect 16075 15116 16120 15144
rect 14921 15107 14979 15113
rect 16114 15104 16120 15116
rect 16172 15104 16178 15156
rect 12768 15048 14228 15076
rect 12768 15036 12774 15048
rect 14274 15036 14280 15088
rect 14332 15076 14338 15088
rect 14332 15048 15516 15076
rect 14332 15036 14338 15048
rect 8297 15011 8355 15017
rect 8297 15008 8309 15011
rect 7340 14980 8309 15008
rect 7340 14968 7346 14980
rect 8297 14977 8309 14980
rect 8343 15008 8355 15011
rect 9125 15011 9183 15017
rect 9125 15008 9137 15011
rect 8343 14980 9137 15008
rect 8343 14977 8355 14980
rect 8297 14971 8355 14977
rect 9125 14977 9137 14980
rect 9171 14977 9183 15011
rect 9125 14971 9183 14977
rect 9953 15011 10011 15017
rect 9953 14977 9965 15011
rect 9999 14977 10011 15011
rect 9953 14971 10011 14977
rect 12345 15011 12403 15017
rect 12345 14977 12357 15011
rect 12391 15008 12403 15011
rect 13078 15008 13084 15020
rect 12391 14980 13084 15008
rect 12391 14977 12403 14980
rect 12345 14971 12403 14977
rect 13078 14968 13084 14980
rect 13136 14968 13142 15020
rect 13262 14968 13268 15020
rect 13320 15008 13326 15020
rect 13541 15011 13599 15017
rect 13541 15008 13553 15011
rect 13320 14980 13553 15008
rect 13320 14968 13326 14980
rect 13541 14977 13553 14980
rect 13587 15008 13599 15011
rect 13722 15008 13728 15020
rect 13587 14980 13728 15008
rect 13587 14977 13599 14980
rect 13541 14971 13599 14977
rect 13722 14968 13728 14980
rect 13780 15008 13786 15020
rect 14185 15011 14243 15017
rect 14185 15008 14197 15011
rect 13780 14980 14197 15008
rect 13780 14968 13786 14980
rect 14185 14977 14197 14980
rect 14231 14977 14243 15011
rect 14185 14971 14243 14977
rect 14369 15011 14427 15017
rect 14369 14977 14381 15011
rect 14415 15008 14427 15011
rect 14734 15008 14740 15020
rect 14415 14980 14740 15008
rect 14415 14977 14427 14980
rect 14369 14971 14427 14977
rect 14734 14968 14740 14980
rect 14792 15008 14798 15020
rect 15102 15008 15108 15020
rect 14792 14980 15108 15008
rect 14792 14968 14798 14980
rect 15102 14968 15108 14980
rect 15160 14968 15166 15020
rect 15286 14968 15292 15020
rect 15344 15008 15350 15020
rect 15488 15017 15516 15048
rect 15381 15011 15439 15017
rect 15381 15008 15393 15011
rect 15344 14980 15393 15008
rect 15344 14968 15350 14980
rect 15381 14977 15393 14980
rect 15427 14977 15439 15011
rect 15381 14971 15439 14977
rect 15473 15011 15531 15017
rect 15473 14977 15485 15011
rect 15519 14977 15531 15011
rect 15473 14971 15531 14977
rect 6273 14943 6331 14949
rect 6273 14909 6285 14943
rect 6319 14940 6331 14943
rect 6822 14940 6828 14952
rect 6319 14912 6828 14940
rect 6319 14909 6331 14912
rect 6273 14903 6331 14909
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 7098 14940 7104 14952
rect 7059 14912 7104 14940
rect 7098 14900 7104 14912
rect 7156 14900 7162 14952
rect 8113 14943 8171 14949
rect 8113 14909 8125 14943
rect 8159 14940 8171 14943
rect 8754 14940 8760 14952
rect 8159 14912 8760 14940
rect 8159 14909 8171 14912
rect 8113 14903 8171 14909
rect 8754 14900 8760 14912
rect 8812 14900 8818 14952
rect 8938 14940 8944 14952
rect 8899 14912 8944 14940
rect 8938 14900 8944 14912
rect 8996 14900 9002 14952
rect 9033 14943 9091 14949
rect 9033 14909 9045 14943
rect 9079 14940 9091 14943
rect 9306 14940 9312 14952
rect 9079 14912 9312 14940
rect 9079 14909 9091 14912
rect 9033 14903 9091 14909
rect 9306 14900 9312 14912
rect 9364 14940 9370 14952
rect 9582 14940 9588 14952
rect 9364 14912 9588 14940
rect 9364 14900 9370 14912
rect 9582 14900 9588 14912
rect 9640 14900 9646 14952
rect 9677 14943 9735 14949
rect 9677 14909 9689 14943
rect 9723 14940 9735 14943
rect 9766 14940 9772 14952
rect 9723 14912 9772 14940
rect 9723 14909 9735 14912
rect 9677 14903 9735 14909
rect 9766 14900 9772 14912
rect 9824 14900 9830 14952
rect 10226 14949 10232 14952
rect 10220 14903 10232 14949
rect 10284 14940 10290 14952
rect 10284 14912 10320 14940
rect 10226 14900 10232 14903
rect 10284 14900 10290 14912
rect 11422 14900 11428 14952
rect 11480 14940 11486 14952
rect 11885 14943 11943 14949
rect 11885 14940 11897 14943
rect 11480 14912 11897 14940
rect 11480 14900 11486 14912
rect 11885 14909 11897 14912
rect 11931 14909 11943 14943
rect 11885 14903 11943 14909
rect 12529 14943 12587 14949
rect 12529 14909 12541 14943
rect 12575 14940 12587 14943
rect 12710 14940 12716 14952
rect 12575 14912 12716 14940
rect 12575 14909 12587 14912
rect 12529 14903 12587 14909
rect 12710 14900 12716 14912
rect 12768 14900 12774 14952
rect 13354 14900 13360 14952
rect 13412 14940 13418 14952
rect 13449 14943 13507 14949
rect 13449 14940 13461 14943
rect 13412 14912 13461 14940
rect 13412 14900 13418 14912
rect 13449 14909 13461 14912
rect 13495 14909 13507 14943
rect 13449 14903 13507 14909
rect 2547 14844 3372 14872
rect 3528 14844 4200 14872
rect 2547 14841 2559 14844
rect 2501 14835 2559 14841
rect 1486 14804 1492 14816
rect 1447 14776 1492 14804
rect 1486 14764 1492 14776
rect 1544 14764 1550 14816
rect 2130 14804 2136 14816
rect 2091 14776 2136 14804
rect 2130 14764 2136 14776
rect 2188 14764 2194 14816
rect 2590 14804 2596 14816
rect 2551 14776 2596 14804
rect 2590 14764 2596 14776
rect 2648 14764 2654 14816
rect 2958 14764 2964 14816
rect 3016 14804 3022 14816
rect 3053 14807 3111 14813
rect 3053 14804 3065 14807
rect 3016 14776 3065 14804
rect 3016 14764 3022 14776
rect 3053 14773 3065 14776
rect 3099 14804 3111 14807
rect 3528 14804 3556 14844
rect 3694 14804 3700 14816
rect 3099 14776 3556 14804
rect 3655 14776 3700 14804
rect 3099 14773 3111 14776
rect 3053 14767 3111 14773
rect 3694 14764 3700 14776
rect 3752 14764 3758 14816
rect 3789 14807 3847 14813
rect 3789 14773 3801 14807
rect 3835 14804 3847 14807
rect 4062 14804 4068 14816
rect 3835 14776 4068 14804
rect 3835 14773 3847 14776
rect 3789 14767 3847 14773
rect 4062 14764 4068 14776
rect 4120 14764 4126 14816
rect 4172 14804 4200 14844
rect 4522 14832 4528 14884
rect 4580 14872 4586 14884
rect 4678 14875 4736 14881
rect 4678 14872 4690 14875
rect 4580 14844 4690 14872
rect 4580 14832 4586 14844
rect 4678 14841 4690 14844
rect 4724 14872 4736 14875
rect 5258 14872 5264 14884
rect 4724 14844 5264 14872
rect 4724 14841 4736 14844
rect 4678 14835 4736 14841
rect 5258 14832 5264 14844
rect 5316 14832 5322 14884
rect 5718 14832 5724 14884
rect 5776 14872 5782 14884
rect 6089 14875 6147 14881
rect 6089 14872 6101 14875
rect 5776 14844 6101 14872
rect 5776 14832 5782 14844
rect 6089 14841 6101 14844
rect 6135 14872 6147 14875
rect 6454 14872 6460 14884
rect 6135 14844 6460 14872
rect 6135 14841 6147 14844
rect 6089 14835 6147 14841
rect 6454 14832 6460 14844
rect 6512 14832 6518 14884
rect 6638 14832 6644 14884
rect 6696 14872 6702 14884
rect 10134 14872 10140 14884
rect 6696 14844 10140 14872
rect 6696 14832 6702 14844
rect 10134 14832 10140 14844
rect 10192 14832 10198 14884
rect 15289 14875 15347 14881
rect 15289 14872 15301 14875
rect 14844 14844 15301 14872
rect 4982 14804 4988 14816
rect 4172 14776 4988 14804
rect 4982 14764 4988 14776
rect 5040 14764 5046 14816
rect 5810 14764 5816 14816
rect 5868 14804 5874 14816
rect 6549 14807 6607 14813
rect 6549 14804 6561 14807
rect 5868 14776 6561 14804
rect 5868 14764 5874 14776
rect 6549 14773 6561 14776
rect 6595 14773 6607 14807
rect 6549 14767 6607 14773
rect 6822 14764 6828 14816
rect 6880 14804 6886 14816
rect 7193 14807 7251 14813
rect 7193 14804 7205 14807
rect 6880 14776 7205 14804
rect 6880 14764 6886 14776
rect 7193 14773 7205 14776
rect 7239 14804 7251 14807
rect 7558 14804 7564 14816
rect 7239 14776 7564 14804
rect 7239 14773 7251 14776
rect 7193 14767 7251 14773
rect 7558 14764 7564 14776
rect 7616 14764 7622 14816
rect 8205 14807 8263 14813
rect 8205 14773 8217 14807
rect 8251 14804 8263 14807
rect 8938 14804 8944 14816
rect 8251 14776 8944 14804
rect 8251 14773 8263 14776
rect 8205 14767 8263 14773
rect 8938 14764 8944 14776
rect 8996 14764 9002 14816
rect 9490 14804 9496 14816
rect 9451 14776 9496 14804
rect 9490 14764 9496 14776
rect 9548 14764 9554 14816
rect 9582 14764 9588 14816
rect 9640 14804 9646 14816
rect 11606 14804 11612 14816
rect 9640 14776 11612 14804
rect 9640 14764 9646 14776
rect 11606 14764 11612 14776
rect 11664 14764 11670 14816
rect 11790 14804 11796 14816
rect 11751 14776 11796 14804
rect 11790 14764 11796 14776
rect 11848 14764 11854 14816
rect 11974 14764 11980 14816
rect 12032 14804 12038 14816
rect 12158 14804 12164 14816
rect 12032 14776 12164 14804
rect 12032 14764 12038 14776
rect 12158 14764 12164 14776
rect 12216 14764 12222 14816
rect 12434 14764 12440 14816
rect 12492 14804 12498 14816
rect 12492 14776 12537 14804
rect 12492 14764 12498 14776
rect 13262 14764 13268 14816
rect 13320 14804 13326 14816
rect 13357 14807 13415 14813
rect 13357 14804 13369 14807
rect 13320 14776 13369 14804
rect 13320 14764 13326 14776
rect 13357 14773 13369 14776
rect 13403 14773 13415 14807
rect 13357 14767 13415 14773
rect 14461 14807 14519 14813
rect 14461 14773 14473 14807
rect 14507 14804 14519 14807
rect 14550 14804 14556 14816
rect 14507 14776 14556 14804
rect 14507 14773 14519 14776
rect 14461 14767 14519 14773
rect 14550 14764 14556 14776
rect 14608 14764 14614 14816
rect 14844 14813 14872 14844
rect 15289 14841 15301 14844
rect 15335 14841 15347 14875
rect 15289 14835 15347 14841
rect 14829 14807 14887 14813
rect 14829 14773 14841 14807
rect 14875 14773 14887 14807
rect 14829 14767 14887 14773
rect 1104 14714 16008 14736
rect 1104 14662 5979 14714
rect 6031 14662 6043 14714
rect 6095 14662 6107 14714
rect 6159 14662 6171 14714
rect 6223 14662 10976 14714
rect 11028 14662 11040 14714
rect 11092 14662 11104 14714
rect 11156 14662 11168 14714
rect 11220 14662 16008 14714
rect 1104 14640 16008 14662
rect 1581 14603 1639 14609
rect 1581 14569 1593 14603
rect 1627 14600 1639 14603
rect 1670 14600 1676 14612
rect 1627 14572 1676 14600
rect 1627 14569 1639 14572
rect 1581 14563 1639 14569
rect 1670 14560 1676 14572
rect 1728 14560 1734 14612
rect 1949 14603 2007 14609
rect 1949 14569 1961 14603
rect 1995 14600 2007 14603
rect 2774 14600 2780 14612
rect 1995 14572 2780 14600
rect 1995 14569 2007 14572
rect 1949 14563 2007 14569
rect 2774 14560 2780 14572
rect 2832 14560 2838 14612
rect 3694 14560 3700 14612
rect 3752 14600 3758 14612
rect 5353 14603 5411 14609
rect 5353 14600 5365 14603
rect 3752 14572 5365 14600
rect 3752 14560 3758 14572
rect 5353 14569 5365 14572
rect 5399 14569 5411 14603
rect 6362 14600 6368 14612
rect 6323 14572 6368 14600
rect 5353 14563 5411 14569
rect 6362 14560 6368 14572
rect 6420 14600 6426 14612
rect 6546 14600 6552 14612
rect 6420 14572 6552 14600
rect 6420 14560 6426 14572
rect 6546 14560 6552 14572
rect 6604 14560 6610 14612
rect 6730 14560 6736 14612
rect 6788 14600 6794 14612
rect 6825 14603 6883 14609
rect 6825 14600 6837 14603
rect 6788 14572 6837 14600
rect 6788 14560 6794 14572
rect 6825 14569 6837 14572
rect 6871 14569 6883 14603
rect 6825 14563 6883 14569
rect 7285 14603 7343 14609
rect 7285 14569 7297 14603
rect 7331 14600 7343 14603
rect 7653 14603 7711 14609
rect 7653 14600 7665 14603
rect 7331 14572 7665 14600
rect 7331 14569 7343 14572
rect 7285 14563 7343 14569
rect 7653 14569 7665 14572
rect 7699 14569 7711 14603
rect 7653 14563 7711 14569
rect 8021 14603 8079 14609
rect 8021 14569 8033 14603
rect 8067 14600 8079 14603
rect 8202 14600 8208 14612
rect 8067 14572 8208 14600
rect 8067 14569 8079 14572
rect 8021 14563 8079 14569
rect 8202 14560 8208 14572
rect 8260 14560 8266 14612
rect 8754 14600 8760 14612
rect 8667 14572 8760 14600
rect 8754 14560 8760 14572
rect 8812 14600 8818 14612
rect 9398 14600 9404 14612
rect 8812 14572 9404 14600
rect 8812 14560 8818 14572
rect 9398 14560 9404 14572
rect 9456 14560 9462 14612
rect 9858 14600 9864 14612
rect 9508 14572 9864 14600
rect 2792 14532 2820 14560
rect 3878 14532 3884 14544
rect 2792 14504 3884 14532
rect 3878 14492 3884 14504
rect 3936 14532 3942 14544
rect 4126 14535 4184 14541
rect 4126 14532 4138 14535
rect 3936 14504 4138 14532
rect 3936 14492 3942 14504
rect 4126 14501 4138 14504
rect 4172 14501 4184 14535
rect 4126 14495 4184 14501
rect 5813 14535 5871 14541
rect 5813 14501 5825 14535
rect 5859 14532 5871 14535
rect 6457 14535 6515 14541
rect 6457 14532 6469 14535
rect 5859 14504 6469 14532
rect 5859 14501 5871 14504
rect 5813 14495 5871 14501
rect 6457 14501 6469 14504
rect 6503 14532 6515 14535
rect 6503 14504 7880 14532
rect 6503 14501 6515 14504
rect 6457 14495 6515 14501
rect 6748 14476 6776 14504
rect 1489 14467 1547 14473
rect 1489 14433 1501 14467
rect 1535 14464 1547 14467
rect 1765 14467 1823 14473
rect 1765 14464 1777 14467
rect 1535 14436 1777 14464
rect 1535 14433 1547 14436
rect 1489 14427 1547 14433
rect 1765 14433 1777 14436
rect 1811 14464 1823 14467
rect 2682 14464 2688 14476
rect 1811 14436 2688 14464
rect 1811 14433 1823 14436
rect 1765 14427 1823 14433
rect 2682 14424 2688 14436
rect 2740 14424 2746 14476
rect 3073 14467 3131 14473
rect 3073 14433 3085 14467
rect 3119 14464 3131 14467
rect 4706 14464 4712 14476
rect 3119 14436 4712 14464
rect 3119 14433 3131 14436
rect 3073 14427 3131 14433
rect 4706 14424 4712 14436
rect 4764 14424 4770 14476
rect 5534 14424 5540 14476
rect 5592 14464 5598 14476
rect 5721 14467 5779 14473
rect 5721 14464 5733 14467
rect 5592 14436 5733 14464
rect 5592 14424 5598 14436
rect 5721 14433 5733 14436
rect 5767 14433 5779 14467
rect 6181 14467 6239 14473
rect 5721 14427 5779 14433
rect 5828 14436 6040 14464
rect 3329 14399 3387 14405
rect 3329 14365 3341 14399
rect 3375 14396 3387 14399
rect 3786 14396 3792 14408
rect 3375 14368 3792 14396
rect 3375 14365 3387 14368
rect 3329 14359 3387 14365
rect 3786 14356 3792 14368
rect 3844 14396 3850 14408
rect 3881 14399 3939 14405
rect 3881 14396 3893 14399
rect 3844 14368 3893 14396
rect 3844 14356 3850 14368
rect 3881 14365 3893 14368
rect 3927 14365 3939 14399
rect 3881 14359 3939 14365
rect 4982 14356 4988 14408
rect 5040 14396 5046 14408
rect 5828 14396 5856 14436
rect 5040 14368 5856 14396
rect 5905 14399 5963 14405
rect 5040 14356 5046 14368
rect 5905 14365 5917 14399
rect 5951 14365 5963 14399
rect 6012 14396 6040 14436
rect 6181 14433 6193 14467
rect 6227 14464 6239 14467
rect 6362 14464 6368 14476
rect 6227 14436 6368 14464
rect 6227 14433 6239 14436
rect 6181 14427 6239 14433
rect 6362 14424 6368 14436
rect 6420 14424 6426 14476
rect 6730 14424 6736 14476
rect 6788 14424 6794 14476
rect 7190 14464 7196 14476
rect 7151 14436 7196 14464
rect 7190 14424 7196 14436
rect 7248 14424 7254 14476
rect 7852 14464 7880 14504
rect 8294 14492 8300 14544
rect 8352 14532 8358 14544
rect 9122 14532 9128 14544
rect 8352 14504 9128 14532
rect 8352 14492 8358 14504
rect 9122 14492 9128 14504
rect 9180 14492 9186 14544
rect 9508 14464 9536 14572
rect 9858 14560 9864 14572
rect 9916 14560 9922 14612
rect 9950 14560 9956 14612
rect 10008 14600 10014 14612
rect 10045 14603 10103 14609
rect 10045 14600 10057 14603
rect 10008 14572 10057 14600
rect 10008 14560 10014 14572
rect 10045 14569 10057 14572
rect 10091 14600 10103 14603
rect 10226 14600 10232 14612
rect 10091 14572 10232 14600
rect 10091 14569 10103 14572
rect 10045 14563 10103 14569
rect 10226 14560 10232 14572
rect 10284 14560 10290 14612
rect 10410 14600 10416 14612
rect 10371 14572 10416 14600
rect 10410 14560 10416 14572
rect 10468 14560 10474 14612
rect 14185 14603 14243 14609
rect 14185 14569 14197 14603
rect 14231 14569 14243 14603
rect 14550 14600 14556 14612
rect 14511 14572 14556 14600
rect 14185 14563 14243 14569
rect 9674 14492 9680 14544
rect 9732 14532 9738 14544
rect 11232 14535 11290 14541
rect 9732 14504 11008 14532
rect 9732 14492 9738 14504
rect 7852 14436 9536 14464
rect 9585 14467 9643 14473
rect 9585 14433 9597 14467
rect 9631 14464 9643 14467
rect 10594 14464 10600 14476
rect 9631 14436 10600 14464
rect 9631 14433 9643 14436
rect 9585 14427 9643 14433
rect 10594 14424 10600 14436
rect 10652 14424 10658 14476
rect 10689 14467 10747 14473
rect 10689 14433 10701 14467
rect 10735 14464 10747 14467
rect 10870 14464 10876 14476
rect 10735 14436 10876 14464
rect 10735 14433 10747 14436
rect 10689 14427 10747 14433
rect 10870 14424 10876 14436
rect 10928 14424 10934 14476
rect 10980 14473 11008 14504
rect 11232 14501 11244 14535
rect 11278 14532 11290 14535
rect 11698 14532 11704 14544
rect 11278 14504 11704 14532
rect 11278 14501 11290 14504
rect 11232 14495 11290 14501
rect 11698 14492 11704 14504
rect 11756 14492 11762 14544
rect 12526 14492 12532 14544
rect 12584 14532 12590 14544
rect 12621 14535 12679 14541
rect 12621 14532 12633 14535
rect 12584 14504 12633 14532
rect 12584 14492 12590 14504
rect 12621 14501 12633 14504
rect 12667 14532 12679 14535
rect 12986 14532 12992 14544
rect 12667 14504 12992 14532
rect 12667 14501 12679 14504
rect 12621 14495 12679 14501
rect 12986 14492 12992 14504
rect 13044 14492 13050 14544
rect 13722 14492 13728 14544
rect 13780 14532 13786 14544
rect 14200 14532 14228 14563
rect 14550 14560 14556 14572
rect 14608 14560 14614 14612
rect 13780 14504 14228 14532
rect 13780 14492 13786 14504
rect 14458 14492 14464 14544
rect 14516 14532 14522 14544
rect 14829 14535 14887 14541
rect 14829 14532 14841 14535
rect 14516 14504 14841 14532
rect 14516 14492 14522 14504
rect 14829 14501 14841 14504
rect 14875 14501 14887 14535
rect 14829 14495 14887 14501
rect 15105 14535 15163 14541
rect 15105 14501 15117 14535
rect 15151 14532 15163 14535
rect 15194 14532 15200 14544
rect 15151 14504 15200 14532
rect 15151 14501 15163 14504
rect 15105 14495 15163 14501
rect 15194 14492 15200 14504
rect 15252 14492 15258 14544
rect 15289 14535 15347 14541
rect 15289 14501 15301 14535
rect 15335 14532 15347 14535
rect 16117 14535 16175 14541
rect 16117 14532 16129 14535
rect 15335 14504 16129 14532
rect 15335 14501 15347 14504
rect 15289 14495 15347 14501
rect 16117 14501 16129 14504
rect 16163 14501 16175 14535
rect 16117 14495 16175 14501
rect 10965 14467 11023 14473
rect 10965 14433 10977 14467
rect 11011 14464 11023 14467
rect 11514 14464 11520 14476
rect 11011 14436 11520 14464
rect 11011 14433 11023 14436
rect 10965 14427 11023 14433
rect 6641 14399 6699 14405
rect 6641 14396 6653 14399
rect 6012 14368 6653 14396
rect 5905 14359 5963 14365
rect 6641 14365 6653 14368
rect 6687 14396 6699 14399
rect 7208 14396 7236 14424
rect 6687 14368 7236 14396
rect 6687 14365 6699 14368
rect 6641 14359 6699 14365
rect 5258 14328 5264 14340
rect 5219 14300 5264 14328
rect 5258 14288 5264 14300
rect 5316 14288 5322 14340
rect 5442 14288 5448 14340
rect 5500 14328 5506 14340
rect 5920 14328 5948 14359
rect 7282 14356 7288 14408
rect 7340 14396 7346 14408
rect 7377 14399 7435 14405
rect 7377 14396 7389 14399
rect 7340 14368 7389 14396
rect 7340 14356 7346 14368
rect 7377 14365 7389 14368
rect 7423 14365 7435 14399
rect 7377 14359 7435 14365
rect 8018 14356 8024 14408
rect 8076 14396 8082 14408
rect 8113 14399 8171 14405
rect 8113 14396 8125 14399
rect 8076 14368 8125 14396
rect 8076 14356 8082 14368
rect 8113 14365 8125 14368
rect 8159 14365 8171 14399
rect 8113 14359 8171 14365
rect 8297 14399 8355 14405
rect 8297 14365 8309 14399
rect 8343 14396 8355 14399
rect 8846 14396 8852 14408
rect 8343 14368 8852 14396
rect 8343 14365 8355 14368
rect 8297 14359 8355 14365
rect 5500 14300 5948 14328
rect 5500 14288 5506 14300
rect 8128 14260 8156 14359
rect 8846 14356 8852 14368
rect 8904 14356 8910 14408
rect 8941 14399 8999 14405
rect 8941 14365 8953 14399
rect 8987 14396 8999 14399
rect 9030 14396 9036 14408
rect 8987 14368 9036 14396
rect 8987 14365 8999 14368
rect 8941 14359 8999 14365
rect 9030 14356 9036 14368
rect 9088 14356 9094 14408
rect 9677 14399 9735 14405
rect 9677 14396 9689 14399
rect 9600 14368 9689 14396
rect 8481 14263 8539 14269
rect 8481 14260 8493 14263
rect 8128 14232 8493 14260
rect 8481 14229 8493 14232
rect 8527 14229 8539 14263
rect 9048 14260 9076 14356
rect 9600 14340 9628 14368
rect 9677 14365 9689 14368
rect 9723 14365 9735 14399
rect 9858 14396 9864 14408
rect 9819 14368 9864 14396
rect 9677 14359 9735 14365
rect 9858 14356 9864 14368
rect 9916 14356 9922 14408
rect 10321 14399 10379 14405
rect 10321 14365 10333 14399
rect 10367 14396 10379 14399
rect 10778 14396 10784 14408
rect 10367 14368 10784 14396
rect 10367 14365 10379 14368
rect 10321 14359 10379 14365
rect 10778 14356 10784 14368
rect 10836 14356 10842 14408
rect 9122 14288 9128 14340
rect 9180 14328 9186 14340
rect 9217 14331 9275 14337
rect 9217 14328 9229 14331
rect 9180 14300 9229 14328
rect 9180 14288 9186 14300
rect 9217 14297 9229 14300
rect 9263 14297 9275 14331
rect 9217 14291 9275 14297
rect 9582 14288 9588 14340
rect 9640 14288 9646 14340
rect 9968 14300 10548 14328
rect 9968 14260 9996 14300
rect 9048 14232 9996 14260
rect 10520 14260 10548 14300
rect 10778 14260 10784 14272
rect 10520 14232 10784 14260
rect 8481 14223 8539 14229
rect 10778 14220 10784 14232
rect 10836 14220 10842 14272
rect 10873 14263 10931 14269
rect 10873 14229 10885 14263
rect 10919 14260 10931 14263
rect 10980 14260 11008 14427
rect 11514 14424 11520 14436
rect 11572 14464 11578 14476
rect 11572 14436 12020 14464
rect 11572 14424 11578 14436
rect 11992 14396 12020 14436
rect 12158 14424 12164 14476
rect 12216 14464 12222 14476
rect 12434 14464 12440 14476
rect 12216 14436 12440 14464
rect 12216 14424 12222 14436
rect 12434 14424 12440 14436
rect 12492 14424 12498 14476
rect 12802 14464 12808 14476
rect 12763 14436 12808 14464
rect 12802 14424 12808 14436
rect 12860 14424 12866 14476
rect 13078 14473 13084 14476
rect 13072 14464 13084 14473
rect 13039 14436 13084 14464
rect 13072 14427 13084 14436
rect 13078 14424 13084 14427
rect 13136 14424 13142 14476
rect 15378 14424 15384 14476
rect 15436 14464 15442 14476
rect 15565 14467 15623 14473
rect 15565 14464 15577 14467
rect 15436 14436 15577 14464
rect 15436 14424 15442 14436
rect 15565 14433 15577 14436
rect 15611 14464 15623 14467
rect 16574 14464 16580 14476
rect 15611 14436 16580 14464
rect 15611 14433 15623 14436
rect 15565 14427 15623 14433
rect 16574 14424 16580 14436
rect 16632 14424 16638 14476
rect 12820 14396 12848 14424
rect 11992 14368 12848 14396
rect 14461 14399 14519 14405
rect 14461 14365 14473 14399
rect 14507 14396 14519 14399
rect 14918 14396 14924 14408
rect 14507 14368 14924 14396
rect 14507 14365 14519 14368
rect 14461 14359 14519 14365
rect 14918 14356 14924 14368
rect 14976 14356 14982 14408
rect 12345 14331 12403 14337
rect 12345 14297 12357 14331
rect 12391 14328 12403 14331
rect 12391 14300 12848 14328
rect 12391 14297 12403 14300
rect 12345 14291 12403 14297
rect 10919 14232 11008 14260
rect 12529 14263 12587 14269
rect 10919 14229 10931 14232
rect 10873 14223 10931 14229
rect 12529 14229 12541 14263
rect 12575 14260 12587 14263
rect 12618 14260 12624 14272
rect 12575 14232 12624 14260
rect 12575 14229 12587 14232
rect 12529 14223 12587 14229
rect 12618 14220 12624 14232
rect 12676 14220 12682 14272
rect 12820 14260 12848 14300
rect 15194 14288 15200 14340
rect 15252 14328 15258 14340
rect 15381 14331 15439 14337
rect 15381 14328 15393 14331
rect 15252 14300 15393 14328
rect 15252 14288 15258 14300
rect 15381 14297 15393 14300
rect 15427 14297 15439 14331
rect 15381 14291 15439 14297
rect 13078 14260 13084 14272
rect 12820 14232 13084 14260
rect 13078 14220 13084 14232
rect 13136 14220 13142 14272
rect 1104 14170 16008 14192
rect 1104 14118 3480 14170
rect 3532 14118 3544 14170
rect 3596 14118 3608 14170
rect 3660 14118 3672 14170
rect 3724 14118 8478 14170
rect 8530 14118 8542 14170
rect 8594 14118 8606 14170
rect 8658 14118 8670 14170
rect 8722 14118 13475 14170
rect 13527 14118 13539 14170
rect 13591 14118 13603 14170
rect 13655 14118 13667 14170
rect 13719 14118 16008 14170
rect 1104 14096 16008 14118
rect 1578 14016 1584 14068
rect 1636 14056 1642 14068
rect 1765 14059 1823 14065
rect 1765 14056 1777 14059
rect 1636 14028 1777 14056
rect 1636 14016 1642 14028
rect 1765 14025 1777 14028
rect 1811 14025 1823 14059
rect 1765 14019 1823 14025
rect 2133 14059 2191 14065
rect 2133 14025 2145 14059
rect 2179 14056 2191 14059
rect 2590 14056 2596 14068
rect 2179 14028 2596 14056
rect 2179 14025 2191 14028
rect 2133 14019 2191 14025
rect 2590 14016 2596 14028
rect 2648 14016 2654 14068
rect 4062 14056 4068 14068
rect 4023 14028 4068 14056
rect 4062 14016 4068 14028
rect 4120 14016 4126 14068
rect 4430 14016 4436 14068
rect 4488 14056 4494 14068
rect 4982 14056 4988 14068
rect 4488 14028 4988 14056
rect 4488 14016 4494 14028
rect 4982 14016 4988 14028
rect 5040 14056 5046 14068
rect 5261 14059 5319 14065
rect 5261 14056 5273 14059
rect 5040 14028 5273 14056
rect 5040 14016 5046 14028
rect 5261 14025 5273 14028
rect 5307 14056 5319 14059
rect 7009 14059 7067 14065
rect 5307 14028 6040 14056
rect 5307 14025 5319 14028
rect 5261 14019 5319 14025
rect 2038 13948 2044 14000
rect 2096 13988 2102 14000
rect 3142 13988 3148 14000
rect 2096 13960 3148 13988
rect 2096 13948 2102 13960
rect 3142 13948 3148 13960
rect 3200 13948 3206 14000
rect 4798 13948 4804 14000
rect 4856 13988 4862 14000
rect 5353 13991 5411 13997
rect 5353 13988 5365 13991
rect 4856 13960 5365 13988
rect 4856 13948 4862 13960
rect 5353 13957 5365 13960
rect 5399 13957 5411 13991
rect 6012 13988 6040 14028
rect 7009 14025 7021 14059
rect 7055 14056 7067 14059
rect 7282 14056 7288 14068
rect 7055 14028 7288 14056
rect 7055 14025 7067 14028
rect 7009 14019 7067 14025
rect 7282 14016 7288 14028
rect 7340 14016 7346 14068
rect 7466 14016 7472 14068
rect 7524 14016 7530 14068
rect 8846 14056 8852 14068
rect 8404 14028 8852 14056
rect 7484 13988 7512 14016
rect 6012 13960 7512 13988
rect 5353 13951 5411 13957
rect 2774 13880 2780 13932
rect 2832 13920 2838 13932
rect 3605 13923 3663 13929
rect 2832 13892 2877 13920
rect 2832 13880 2838 13892
rect 3605 13889 3617 13923
rect 3651 13920 3663 13923
rect 4706 13920 4712 13932
rect 3651 13892 4712 13920
rect 3651 13889 3663 13892
rect 3605 13883 3663 13889
rect 4706 13880 4712 13892
rect 4764 13920 4770 13932
rect 5442 13920 5448 13932
rect 4764 13892 5448 13920
rect 4764 13880 4770 13892
rect 5442 13880 5448 13892
rect 5500 13880 5506 13932
rect 5905 13923 5963 13929
rect 5905 13889 5917 13923
rect 5951 13920 5963 13923
rect 6822 13920 6828 13932
rect 5951 13892 6828 13920
rect 5951 13889 5963 13892
rect 5905 13883 5963 13889
rect 6822 13880 6828 13892
rect 6880 13880 6886 13932
rect 8404 13920 8432 14028
rect 8846 14016 8852 14028
rect 8904 14056 8910 14068
rect 9953 14059 10011 14065
rect 9953 14056 9965 14059
rect 8904 14028 9965 14056
rect 8904 14016 8910 14028
rect 9953 14025 9965 14028
rect 9999 14025 10011 14059
rect 9953 14019 10011 14025
rect 10594 14016 10600 14068
rect 10652 14056 10658 14068
rect 11701 14059 11759 14065
rect 11701 14056 11713 14059
rect 10652 14028 11713 14056
rect 10652 14016 10658 14028
rect 11701 14025 11713 14028
rect 11747 14025 11759 14059
rect 13354 14056 13360 14068
rect 13315 14028 13360 14056
rect 11701 14019 11759 14025
rect 13354 14016 13360 14028
rect 13412 14016 13418 14068
rect 13998 14016 14004 14068
rect 14056 14056 14062 14068
rect 14277 14059 14335 14065
rect 14277 14056 14289 14059
rect 14056 14028 14289 14056
rect 14056 14016 14062 14028
rect 14277 14025 14289 14028
rect 14323 14025 14335 14059
rect 14277 14019 14335 14025
rect 14826 14016 14832 14068
rect 14884 14056 14890 14068
rect 15102 14056 15108 14068
rect 14884 14028 15108 14056
rect 14884 14016 14890 14028
rect 15102 14016 15108 14028
rect 15160 14016 15166 14068
rect 9858 13988 9864 14000
rect 9771 13960 9864 13988
rect 9858 13948 9864 13960
rect 9916 13948 9922 14000
rect 11422 13988 11428 14000
rect 11383 13960 11428 13988
rect 11422 13948 11428 13960
rect 11480 13948 11486 14000
rect 13262 13948 13268 14000
rect 13320 13988 13326 14000
rect 13449 13991 13507 13997
rect 13449 13988 13461 13991
rect 13320 13960 13461 13988
rect 13320 13948 13326 13960
rect 13449 13957 13461 13960
rect 13495 13957 13507 13991
rect 13449 13951 13507 13957
rect 8312 13892 8432 13920
rect 1394 13852 1400 13864
rect 1355 13824 1400 13852
rect 1394 13812 1400 13824
rect 1452 13812 1458 13864
rect 1946 13852 1952 13864
rect 1907 13824 1952 13852
rect 1946 13812 1952 13824
rect 2004 13812 2010 13864
rect 5718 13852 5724 13864
rect 5679 13824 5724 13852
rect 5718 13812 5724 13824
rect 5776 13812 5782 13864
rect 6549 13855 6607 13861
rect 6549 13821 6561 13855
rect 6595 13852 6607 13855
rect 6638 13852 6644 13864
rect 6595 13824 6644 13852
rect 6595 13821 6607 13824
rect 6549 13815 6607 13821
rect 6638 13812 6644 13824
rect 6696 13812 6702 13864
rect 8133 13855 8191 13861
rect 6840 13824 8064 13852
rect 1581 13787 1639 13793
rect 1581 13753 1593 13787
rect 1627 13784 1639 13787
rect 1670 13784 1676 13796
rect 1627 13756 1676 13784
rect 1627 13753 1639 13756
rect 1581 13747 1639 13753
rect 1670 13744 1676 13756
rect 1728 13744 1734 13796
rect 2501 13787 2559 13793
rect 2501 13753 2513 13787
rect 2547 13784 2559 13787
rect 3329 13787 3387 13793
rect 2547 13756 2774 13784
rect 2547 13753 2559 13756
rect 2501 13747 2559 13753
rect 2590 13676 2596 13728
rect 2648 13716 2654 13728
rect 2746 13716 2774 13756
rect 3329 13753 3341 13787
rect 3375 13784 3387 13787
rect 4430 13784 4436 13796
rect 3375 13756 3924 13784
rect 4391 13756 4436 13784
rect 3375 13753 3387 13756
rect 3329 13747 3387 13753
rect 2961 13719 3019 13725
rect 2961 13716 2973 13719
rect 2648 13688 2693 13716
rect 2746 13688 2973 13716
rect 2648 13676 2654 13688
rect 2961 13685 2973 13688
rect 3007 13685 3019 13719
rect 3418 13716 3424 13728
rect 3379 13688 3424 13716
rect 2961 13679 3019 13685
rect 3418 13676 3424 13688
rect 3476 13676 3482 13728
rect 3896 13725 3924 13756
rect 4430 13744 4436 13756
rect 4488 13744 4494 13796
rect 5077 13787 5135 13793
rect 5077 13753 5089 13787
rect 5123 13784 5135 13787
rect 5534 13784 5540 13796
rect 5123 13756 5540 13784
rect 5123 13753 5135 13756
rect 5077 13747 5135 13753
rect 5534 13744 5540 13756
rect 5592 13744 5598 13796
rect 5902 13784 5908 13796
rect 5736 13756 5908 13784
rect 3881 13719 3939 13725
rect 3881 13685 3893 13719
rect 3927 13716 3939 13719
rect 4062 13716 4068 13728
rect 3927 13688 4068 13716
rect 3927 13685 3939 13688
rect 3881 13679 3939 13685
rect 4062 13676 4068 13688
rect 4120 13676 4126 13728
rect 4522 13716 4528 13728
rect 4483 13688 4528 13716
rect 4522 13676 4528 13688
rect 4580 13676 4586 13728
rect 5442 13676 5448 13728
rect 5500 13716 5506 13728
rect 5736 13716 5764 13756
rect 5902 13744 5908 13756
rect 5960 13784 5966 13796
rect 6840 13784 6868 13824
rect 5960 13756 6868 13784
rect 8036 13784 8064 13824
rect 8133 13821 8145 13855
rect 8179 13852 8191 13855
rect 8312 13852 8340 13892
rect 8179 13824 8340 13852
rect 8179 13821 8191 13824
rect 8133 13815 8191 13821
rect 8386 13812 8392 13864
rect 8444 13852 8450 13864
rect 8481 13855 8539 13861
rect 8481 13852 8493 13855
rect 8444 13824 8493 13852
rect 8444 13812 8450 13824
rect 8481 13821 8493 13824
rect 8527 13821 8539 13855
rect 8481 13815 8539 13821
rect 8748 13855 8806 13861
rect 8748 13821 8760 13855
rect 8794 13852 8806 13855
rect 9876 13852 9904 13948
rect 12253 13923 12311 13929
rect 12253 13920 12265 13923
rect 11256 13892 12265 13920
rect 11066 13855 11124 13861
rect 11066 13852 11078 13855
rect 8794 13824 9812 13852
rect 9876 13824 11078 13852
rect 8794 13821 8806 13824
rect 8748 13815 8806 13821
rect 9214 13784 9220 13796
rect 8036 13756 9220 13784
rect 5960 13744 5966 13756
rect 9214 13744 9220 13756
rect 9272 13744 9278 13796
rect 9784 13784 9812 13824
rect 11066 13821 11078 13824
rect 11112 13821 11124 13855
rect 11256 13852 11284 13892
rect 12253 13889 12265 13892
rect 12299 13889 12311 13923
rect 12253 13883 12311 13889
rect 12342 13880 12348 13932
rect 12400 13920 12406 13932
rect 12805 13923 12863 13929
rect 12400 13892 12756 13920
rect 12400 13880 12406 13892
rect 11066 13815 11124 13821
rect 11164 13824 11284 13852
rect 11333 13855 11391 13861
rect 10410 13784 10416 13796
rect 9784 13756 10416 13784
rect 10410 13744 10416 13756
rect 10468 13784 10474 13796
rect 11164 13784 11192 13824
rect 11333 13821 11345 13855
rect 11379 13852 11391 13855
rect 11514 13852 11520 13864
rect 11379 13824 11520 13852
rect 11379 13821 11391 13824
rect 11333 13815 11391 13821
rect 11514 13812 11520 13824
rect 11572 13812 11578 13864
rect 12161 13855 12219 13861
rect 12161 13821 12173 13855
rect 12207 13852 12219 13855
rect 12526 13852 12532 13864
rect 12207 13824 12532 13852
rect 12207 13821 12219 13824
rect 12161 13815 12219 13821
rect 12526 13812 12532 13824
rect 12584 13812 12590 13864
rect 12728 13852 12756 13892
rect 12805 13889 12817 13923
rect 12851 13920 12863 13923
rect 13078 13920 13084 13932
rect 12851 13892 13084 13920
rect 12851 13889 12863 13892
rect 12805 13883 12863 13889
rect 13078 13880 13084 13892
rect 13136 13920 13142 13932
rect 14001 13923 14059 13929
rect 14001 13920 14013 13923
rect 13136 13892 14013 13920
rect 13136 13880 13142 13892
rect 14001 13889 14013 13892
rect 14047 13889 14059 13923
rect 14550 13920 14556 13932
rect 14511 13892 14556 13920
rect 14001 13883 14059 13889
rect 14550 13880 14556 13892
rect 14608 13880 14614 13932
rect 13814 13852 13820 13864
rect 12728 13824 13820 13852
rect 13814 13812 13820 13824
rect 13872 13812 13878 13864
rect 10468 13756 11192 13784
rect 10468 13744 10474 13756
rect 12434 13744 12440 13796
rect 12492 13784 12498 13796
rect 12897 13787 12955 13793
rect 12897 13784 12909 13787
rect 12492 13756 12909 13784
rect 12492 13744 12498 13756
rect 12897 13753 12909 13756
rect 12943 13784 12955 13787
rect 13078 13784 13084 13796
rect 12943 13756 13084 13784
rect 12943 13753 12955 13756
rect 12897 13747 12955 13753
rect 13078 13744 13084 13756
rect 13136 13744 13142 13796
rect 13538 13744 13544 13796
rect 13596 13784 13602 13796
rect 13909 13787 13967 13793
rect 13909 13784 13921 13787
rect 13596 13756 13921 13784
rect 13596 13744 13602 13756
rect 13909 13753 13921 13756
rect 13955 13753 13967 13787
rect 13909 13747 13967 13753
rect 15102 13744 15108 13796
rect 15160 13784 15166 13796
rect 15473 13787 15531 13793
rect 15473 13784 15485 13787
rect 15160 13756 15485 13784
rect 15160 13744 15166 13756
rect 15473 13753 15485 13756
rect 15519 13753 15531 13787
rect 15473 13747 15531 13753
rect 15562 13744 15568 13796
rect 15620 13784 15626 13796
rect 15620 13756 15665 13784
rect 15620 13744 15626 13756
rect 5500 13688 5764 13716
rect 5500 13676 5506 13688
rect 5810 13676 5816 13728
rect 5868 13716 5874 13728
rect 6733 13719 6791 13725
rect 5868 13688 5913 13716
rect 5868 13676 5874 13688
rect 6733 13685 6745 13719
rect 6779 13716 6791 13719
rect 6914 13716 6920 13728
rect 6779 13688 6920 13716
rect 6779 13685 6791 13688
rect 6733 13679 6791 13685
rect 6914 13676 6920 13688
rect 6972 13716 6978 13728
rect 8202 13716 8208 13728
rect 6972 13688 8208 13716
rect 6972 13676 6978 13688
rect 8202 13676 8208 13688
rect 8260 13676 8266 13728
rect 9398 13676 9404 13728
rect 9456 13716 9462 13728
rect 11790 13716 11796 13728
rect 9456 13688 11796 13716
rect 9456 13676 9462 13688
rect 11790 13676 11796 13688
rect 11848 13676 11854 13728
rect 12069 13719 12127 13725
rect 12069 13685 12081 13719
rect 12115 13716 12127 13719
rect 12158 13716 12164 13728
rect 12115 13688 12164 13716
rect 12115 13685 12127 13688
rect 12069 13679 12127 13685
rect 12158 13676 12164 13688
rect 12216 13676 12222 13728
rect 12989 13719 13047 13725
rect 12989 13685 13001 13719
rect 13035 13716 13047 13719
rect 13630 13716 13636 13728
rect 13035 13688 13636 13716
rect 13035 13685 13047 13688
rect 12989 13679 13047 13685
rect 13630 13676 13636 13688
rect 13688 13676 13694 13728
rect 1104 13626 16008 13648
rect 1104 13574 5979 13626
rect 6031 13574 6043 13626
rect 6095 13574 6107 13626
rect 6159 13574 6171 13626
rect 6223 13574 10976 13626
rect 11028 13574 11040 13626
rect 11092 13574 11104 13626
rect 11156 13574 11168 13626
rect 11220 13574 16008 13626
rect 1104 13552 16008 13574
rect 2590 13472 2596 13524
rect 2648 13512 2654 13524
rect 2685 13515 2743 13521
rect 2685 13512 2697 13515
rect 2648 13484 2697 13512
rect 2648 13472 2654 13484
rect 2685 13481 2697 13484
rect 2731 13481 2743 13515
rect 2685 13475 2743 13481
rect 2866 13472 2872 13524
rect 2924 13512 2930 13524
rect 3053 13515 3111 13521
rect 3053 13512 3065 13515
rect 2924 13484 3065 13512
rect 2924 13472 2930 13484
rect 3053 13481 3065 13484
rect 3099 13481 3111 13515
rect 3053 13475 3111 13481
rect 3068 13444 3096 13475
rect 3418 13472 3424 13524
rect 3476 13512 3482 13524
rect 3878 13512 3884 13524
rect 3476 13484 3884 13512
rect 3476 13472 3482 13484
rect 3878 13472 3884 13484
rect 3936 13512 3942 13524
rect 3973 13515 4031 13521
rect 3973 13512 3985 13515
rect 3936 13484 3985 13512
rect 3936 13472 3942 13484
rect 3973 13481 3985 13484
rect 4019 13481 4031 13515
rect 3973 13475 4031 13481
rect 5445 13515 5503 13521
rect 5445 13481 5457 13515
rect 5491 13512 5503 13515
rect 5810 13512 5816 13524
rect 5491 13484 5816 13512
rect 5491 13481 5503 13484
rect 5445 13475 5503 13481
rect 5810 13472 5816 13484
rect 5868 13472 5874 13524
rect 6638 13512 6644 13524
rect 5920 13484 6644 13512
rect 5920 13453 5948 13484
rect 6638 13472 6644 13484
rect 6696 13472 6702 13524
rect 6822 13472 6828 13524
rect 6880 13512 6886 13524
rect 7653 13515 7711 13521
rect 7653 13512 7665 13515
rect 6880 13484 7665 13512
rect 6880 13472 6886 13484
rect 7653 13481 7665 13484
rect 7699 13481 7711 13515
rect 7653 13475 7711 13481
rect 8294 13472 8300 13524
rect 8352 13512 8358 13524
rect 8665 13515 8723 13521
rect 8665 13512 8677 13515
rect 8352 13484 8677 13512
rect 8352 13472 8358 13484
rect 8665 13481 8677 13484
rect 8711 13481 8723 13515
rect 8938 13512 8944 13524
rect 8851 13484 8944 13512
rect 8665 13475 8723 13481
rect 3513 13447 3571 13453
rect 3513 13444 3525 13447
rect 3068 13416 3525 13444
rect 3513 13413 3525 13416
rect 3559 13413 3571 13447
rect 5905 13447 5963 13453
rect 5905 13444 5917 13447
rect 3513 13407 3571 13413
rect 5644 13416 5917 13444
rect 1673 13379 1731 13385
rect 1673 13345 1685 13379
rect 1719 13376 1731 13379
rect 2130 13376 2136 13388
rect 1719 13348 2136 13376
rect 1719 13345 1731 13348
rect 1673 13339 1731 13345
rect 2130 13336 2136 13348
rect 2188 13336 2194 13388
rect 2682 13336 2688 13388
rect 2740 13376 2746 13388
rect 5258 13376 5264 13388
rect 2740 13348 5264 13376
rect 2740 13336 2746 13348
rect 5258 13336 5264 13348
rect 5316 13376 5322 13388
rect 5644 13376 5672 13416
rect 5905 13413 5917 13416
rect 5951 13413 5963 13447
rect 5905 13407 5963 13413
rect 6012 13416 7236 13444
rect 5810 13376 5816 13388
rect 5316 13348 5672 13376
rect 5771 13348 5816 13376
rect 5316 13336 5322 13348
rect 5810 13336 5816 13348
rect 5868 13336 5874 13388
rect 3142 13308 3148 13320
rect 3103 13280 3148 13308
rect 3142 13268 3148 13280
rect 3200 13268 3206 13320
rect 3329 13311 3387 13317
rect 3329 13277 3341 13311
rect 3375 13308 3387 13311
rect 4706 13308 4712 13320
rect 3375 13280 4712 13308
rect 3375 13277 3387 13280
rect 3329 13271 3387 13277
rect 4706 13268 4712 13280
rect 4764 13268 4770 13320
rect 4522 13200 4528 13252
rect 4580 13240 4586 13252
rect 5169 13243 5227 13249
rect 5169 13240 5181 13243
rect 4580 13212 5181 13240
rect 4580 13200 4586 13212
rect 5169 13209 5181 13212
rect 5215 13240 5227 13243
rect 6012 13240 6040 13416
rect 6529 13379 6587 13385
rect 6529 13376 6541 13379
rect 6196 13348 6541 13376
rect 6196 13320 6224 13348
rect 6529 13345 6541 13348
rect 6575 13345 6587 13379
rect 7208 13376 7236 13416
rect 7282 13404 7288 13456
rect 7340 13444 7346 13456
rect 7837 13447 7895 13453
rect 7837 13444 7849 13447
rect 7340 13416 7849 13444
rect 7340 13404 7346 13416
rect 7837 13413 7849 13416
rect 7883 13444 7895 13447
rect 8202 13444 8208 13456
rect 7883 13416 8208 13444
rect 7883 13413 7895 13416
rect 7837 13407 7895 13413
rect 8202 13404 8208 13416
rect 8260 13404 8266 13456
rect 8680 13444 8708 13475
rect 8938 13472 8944 13484
rect 8996 13512 9002 13524
rect 9398 13512 9404 13524
rect 8996 13484 9404 13512
rect 8996 13472 9002 13484
rect 9398 13472 9404 13484
rect 9456 13472 9462 13524
rect 9582 13512 9588 13524
rect 9543 13484 9588 13512
rect 9582 13472 9588 13484
rect 9640 13472 9646 13524
rect 10410 13512 10416 13524
rect 10371 13484 10416 13512
rect 10410 13472 10416 13484
rect 10468 13472 10474 13524
rect 10778 13472 10784 13524
rect 10836 13512 10842 13524
rect 11882 13512 11888 13524
rect 10836 13484 11888 13512
rect 10836 13472 10842 13484
rect 11882 13472 11888 13484
rect 11940 13472 11946 13524
rect 12158 13512 12164 13524
rect 12119 13484 12164 13512
rect 12158 13472 12164 13484
rect 12216 13472 12222 13524
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 13538 13512 13544 13524
rect 12492 13484 13544 13512
rect 12492 13472 12498 13484
rect 13538 13472 13544 13484
rect 13596 13472 13602 13524
rect 13630 13472 13636 13524
rect 13688 13512 13694 13524
rect 13909 13515 13967 13521
rect 13909 13512 13921 13515
rect 13688 13484 13921 13512
rect 13688 13472 13694 13484
rect 13909 13481 13921 13484
rect 13955 13481 13967 13515
rect 13909 13475 13967 13481
rect 13998 13472 14004 13524
rect 14056 13512 14062 13524
rect 14645 13515 14703 13521
rect 14645 13512 14657 13515
rect 14056 13484 14657 13512
rect 14056 13472 14062 13484
rect 14645 13481 14657 13484
rect 14691 13512 14703 13515
rect 14734 13512 14740 13524
rect 14691 13484 14740 13512
rect 14691 13481 14703 13484
rect 14645 13475 14703 13481
rect 14734 13472 14740 13484
rect 14792 13472 14798 13524
rect 15102 13521 15108 13524
rect 15059 13515 15108 13521
rect 15059 13481 15071 13515
rect 15105 13481 15108 13515
rect 15059 13475 15108 13481
rect 15102 13472 15108 13475
rect 15160 13472 15166 13524
rect 15378 13512 15384 13524
rect 15339 13484 15384 13512
rect 15378 13472 15384 13484
rect 15436 13472 15442 13524
rect 15473 13515 15531 13521
rect 15473 13481 15485 13515
rect 15519 13512 15531 13515
rect 15562 13512 15568 13524
rect 15519 13484 15568 13512
rect 15519 13481 15531 13484
rect 15473 13475 15531 13481
rect 15562 13472 15568 13484
rect 15620 13472 15626 13524
rect 9493 13447 9551 13453
rect 9493 13444 9505 13447
rect 8680 13416 9505 13444
rect 9493 13413 9505 13416
rect 9539 13413 9551 13447
rect 9493 13407 9551 13413
rect 9953 13447 10011 13453
rect 9953 13413 9965 13447
rect 9999 13444 10011 13447
rect 11422 13444 11428 13456
rect 9999 13416 11428 13444
rect 9999 13413 10011 13416
rect 9953 13407 10011 13413
rect 11422 13404 11428 13416
rect 11480 13404 11486 13456
rect 11514 13404 11520 13456
rect 11572 13453 11578 13456
rect 11572 13444 11584 13453
rect 11572 13416 12112 13444
rect 11572 13407 11584 13416
rect 11572 13404 11578 13407
rect 7374 13376 7380 13388
rect 7208 13348 7380 13376
rect 6529 13339 6587 13345
rect 7374 13336 7380 13348
rect 7432 13376 7438 13388
rect 10594 13376 10600 13388
rect 7432 13348 10600 13376
rect 7432 13336 7438 13348
rect 10594 13336 10600 13348
rect 10652 13336 10658 13388
rect 10704 13348 11928 13376
rect 6089 13311 6147 13317
rect 6089 13277 6101 13311
rect 6135 13308 6147 13311
rect 6178 13308 6184 13320
rect 6135 13280 6184 13308
rect 6135 13277 6147 13280
rect 6089 13271 6147 13277
rect 6178 13268 6184 13280
rect 6236 13268 6242 13320
rect 6273 13311 6331 13317
rect 6273 13277 6285 13311
rect 6319 13277 6331 13311
rect 6273 13271 6331 13277
rect 5215 13212 6040 13240
rect 5215 13209 5227 13212
rect 5169 13203 5227 13209
rect 1489 13175 1547 13181
rect 1489 13141 1501 13175
rect 1535 13172 1547 13175
rect 1578 13172 1584 13184
rect 1535 13144 1584 13172
rect 1535 13141 1547 13144
rect 1489 13135 1547 13141
rect 1578 13132 1584 13144
rect 1636 13132 1642 13184
rect 6288 13172 6316 13271
rect 9766 13268 9772 13320
rect 9824 13308 9830 13320
rect 10045 13311 10103 13317
rect 10045 13308 10057 13311
rect 9824 13280 10057 13308
rect 9824 13268 9830 13280
rect 10045 13277 10057 13280
rect 10091 13277 10103 13311
rect 10045 13271 10103 13277
rect 10229 13311 10287 13317
rect 10229 13277 10241 13311
rect 10275 13308 10287 13311
rect 10410 13308 10416 13320
rect 10275 13280 10416 13308
rect 10275 13277 10287 13280
rect 10229 13271 10287 13277
rect 10410 13268 10416 13280
rect 10468 13268 10474 13320
rect 9493 13243 9551 13249
rect 7208 13212 8064 13240
rect 6546 13172 6552 13184
rect 6288 13144 6552 13172
rect 6546 13132 6552 13144
rect 6604 13132 6610 13184
rect 6638 13132 6644 13184
rect 6696 13172 6702 13184
rect 7208 13172 7236 13212
rect 6696 13144 7236 13172
rect 6696 13132 6702 13144
rect 7558 13132 7564 13184
rect 7616 13172 7622 13184
rect 7929 13175 7987 13181
rect 7929 13172 7941 13175
rect 7616 13144 7941 13172
rect 7616 13132 7622 13144
rect 7929 13141 7941 13144
rect 7975 13141 7987 13175
rect 8036 13172 8064 13212
rect 9493 13209 9505 13243
rect 9539 13240 9551 13243
rect 10704 13240 10732 13348
rect 11790 13308 11796 13320
rect 11751 13280 11796 13308
rect 11790 13268 11796 13280
rect 11848 13268 11854 13320
rect 9539 13212 10732 13240
rect 11900 13240 11928 13348
rect 12084 13308 12112 13416
rect 12250 13404 12256 13456
rect 12308 13444 12314 13456
rect 12621 13447 12679 13453
rect 12621 13444 12633 13447
rect 12308 13416 12633 13444
rect 12308 13404 12314 13416
rect 12621 13413 12633 13416
rect 12667 13444 12679 13447
rect 14093 13447 14151 13453
rect 14093 13444 14105 13447
rect 12667 13416 14105 13444
rect 12667 13413 12679 13416
rect 12621 13407 12679 13413
rect 14093 13413 14105 13416
rect 14139 13413 14151 13447
rect 14366 13444 14372 13456
rect 14327 13416 14372 13444
rect 14093 13407 14151 13413
rect 14366 13404 14372 13416
rect 14424 13404 14430 13456
rect 12529 13379 12587 13385
rect 12529 13345 12541 13379
rect 12575 13376 12587 13379
rect 13354 13376 13360 13388
rect 12575 13348 13360 13376
rect 12575 13345 12587 13348
rect 12529 13339 12587 13345
rect 13354 13336 13360 13348
rect 13412 13336 13418 13388
rect 14988 13379 15046 13385
rect 14988 13345 15000 13379
rect 15034 13376 15046 13379
rect 15286 13376 15292 13388
rect 15034 13348 15292 13376
rect 15034 13345 15046 13348
rect 14988 13339 15046 13345
rect 15286 13336 15292 13348
rect 15344 13336 15350 13388
rect 15654 13376 15660 13388
rect 15615 13348 15660 13376
rect 15654 13336 15660 13348
rect 15712 13336 15718 13388
rect 12710 13308 12716 13320
rect 12084 13280 12716 13308
rect 12710 13268 12716 13280
rect 12768 13268 12774 13320
rect 12986 13308 12992 13320
rect 12947 13280 12992 13308
rect 12986 13268 12992 13280
rect 13044 13268 13050 13320
rect 13078 13268 13084 13320
rect 13136 13308 13142 13320
rect 13173 13311 13231 13317
rect 13173 13308 13185 13311
rect 13136 13280 13185 13308
rect 13136 13268 13142 13280
rect 13173 13277 13185 13280
rect 13219 13277 13231 13311
rect 13173 13271 13231 13277
rect 13262 13268 13268 13320
rect 13320 13308 13326 13320
rect 13449 13311 13507 13317
rect 13449 13308 13461 13311
rect 13320 13280 13461 13308
rect 13320 13268 13326 13280
rect 13449 13277 13461 13280
rect 13495 13277 13507 13311
rect 13449 13271 13507 13277
rect 13630 13240 13636 13252
rect 11900 13212 13636 13240
rect 9539 13209 9551 13212
rect 9493 13203 9551 13209
rect 13630 13200 13636 13212
rect 13688 13200 13694 13252
rect 10226 13172 10232 13184
rect 8036 13144 10232 13172
rect 7929 13135 7987 13141
rect 10226 13132 10232 13144
rect 10284 13132 10290 13184
rect 11882 13132 11888 13184
rect 11940 13172 11946 13184
rect 11977 13175 12035 13181
rect 11977 13172 11989 13175
rect 11940 13144 11989 13172
rect 11940 13132 11946 13144
rect 11977 13141 11989 13144
rect 12023 13172 12035 13175
rect 12066 13172 12072 13184
rect 12023 13144 12072 13172
rect 12023 13141 12035 13144
rect 11977 13135 12035 13141
rect 12066 13132 12072 13144
rect 12124 13132 12130 13184
rect 12894 13132 12900 13184
rect 12952 13172 12958 13184
rect 13078 13172 13084 13184
rect 12952 13144 13084 13172
rect 12952 13132 12958 13144
rect 13078 13132 13084 13144
rect 13136 13172 13142 13184
rect 13817 13175 13875 13181
rect 13817 13172 13829 13175
rect 13136 13144 13829 13172
rect 13136 13132 13142 13144
rect 13817 13141 13829 13144
rect 13863 13141 13875 13175
rect 14734 13172 14740 13184
rect 14695 13144 14740 13172
rect 13817 13135 13875 13141
rect 14734 13132 14740 13144
rect 14792 13132 14798 13184
rect 1104 13082 16008 13104
rect 1104 13030 3480 13082
rect 3532 13030 3544 13082
rect 3596 13030 3608 13082
rect 3660 13030 3672 13082
rect 3724 13030 8478 13082
rect 8530 13030 8542 13082
rect 8594 13030 8606 13082
rect 8658 13030 8670 13082
rect 8722 13030 13475 13082
rect 13527 13030 13539 13082
rect 13591 13030 13603 13082
rect 13655 13030 13667 13082
rect 13719 13030 16008 13082
rect 1104 13008 16008 13030
rect 1670 12928 1676 12980
rect 1728 12968 1734 12980
rect 1765 12971 1823 12977
rect 1765 12968 1777 12971
rect 1728 12940 1777 12968
rect 1728 12928 1734 12940
rect 1765 12937 1777 12940
rect 1811 12937 1823 12971
rect 1765 12931 1823 12937
rect 3142 12928 3148 12980
rect 3200 12968 3206 12980
rect 3237 12971 3295 12977
rect 3237 12968 3249 12971
rect 3200 12940 3249 12968
rect 3200 12928 3206 12940
rect 3237 12937 3249 12940
rect 3283 12937 3295 12971
rect 3970 12968 3976 12980
rect 3237 12931 3295 12937
rect 3344 12940 3976 12968
rect 1394 12900 1400 12912
rect 1355 12872 1400 12900
rect 1394 12860 1400 12872
rect 1452 12860 1458 12912
rect 2866 12860 2872 12912
rect 2924 12900 2930 12912
rect 3344 12900 3372 12940
rect 3970 12928 3976 12940
rect 4028 12968 4034 12980
rect 4706 12968 4712 12980
rect 4028 12940 4568 12968
rect 4667 12940 4712 12968
rect 4028 12928 4034 12940
rect 2924 12872 3372 12900
rect 4540 12900 4568 12940
rect 4706 12928 4712 12940
rect 4764 12928 4770 12980
rect 5718 12928 5724 12980
rect 5776 12968 5782 12980
rect 6457 12971 6515 12977
rect 6457 12968 6469 12971
rect 5776 12940 6469 12968
rect 5776 12928 5782 12940
rect 6457 12937 6469 12940
rect 6503 12937 6515 12971
rect 6457 12931 6515 12937
rect 7834 12928 7840 12980
rect 7892 12968 7898 12980
rect 8389 12971 8447 12977
rect 8389 12968 8401 12971
rect 7892 12940 8401 12968
rect 7892 12928 7898 12940
rect 8389 12937 8401 12940
rect 8435 12968 8447 12971
rect 9766 12968 9772 12980
rect 8435 12940 9674 12968
rect 9727 12940 9772 12968
rect 8435 12937 8447 12940
rect 8389 12931 8447 12937
rect 5534 12900 5540 12912
rect 4540 12872 5540 12900
rect 2924 12860 2930 12872
rect 5534 12860 5540 12872
rect 5592 12860 5598 12912
rect 6270 12860 6276 12912
rect 6328 12900 6334 12912
rect 6822 12900 6828 12912
rect 6328 12872 6828 12900
rect 6328 12860 6334 12872
rect 6822 12860 6828 12872
rect 6880 12900 6886 12912
rect 8113 12903 8171 12909
rect 6880 12872 7880 12900
rect 6880 12860 6886 12872
rect 2685 12835 2743 12841
rect 2685 12801 2697 12835
rect 2731 12832 2743 12835
rect 2731 12804 3464 12832
rect 2731 12801 2743 12804
rect 2685 12795 2743 12801
rect 1578 12764 1584 12776
rect 1539 12736 1584 12764
rect 1578 12724 1584 12736
rect 1636 12724 1642 12776
rect 1949 12767 2007 12773
rect 1949 12733 1961 12767
rect 1995 12733 2007 12767
rect 1949 12727 2007 12733
rect 1964 12696 1992 12727
rect 2774 12724 2780 12776
rect 2832 12764 2838 12776
rect 3329 12767 3387 12773
rect 3329 12764 3341 12767
rect 2832 12736 3341 12764
rect 2832 12724 2838 12736
rect 3329 12733 3341 12736
rect 3375 12733 3387 12767
rect 3329 12727 3387 12733
rect 3436 12708 3464 12804
rect 4338 12792 4344 12844
rect 4396 12832 4402 12844
rect 5445 12835 5503 12841
rect 5445 12832 5457 12835
rect 4396 12804 5457 12832
rect 4396 12792 4402 12804
rect 5445 12801 5457 12804
rect 5491 12832 5503 12835
rect 5994 12832 6000 12844
rect 5491 12804 6000 12832
rect 5491 12801 5503 12804
rect 5445 12795 5503 12801
rect 5994 12792 6000 12804
rect 6052 12792 6058 12844
rect 6178 12832 6184 12844
rect 6139 12804 6184 12832
rect 6178 12792 6184 12804
rect 6236 12832 6242 12844
rect 7852 12841 7880 12872
rect 8113 12869 8125 12903
rect 8159 12869 8171 12903
rect 9646 12900 9674 12940
rect 9766 12928 9772 12940
rect 9824 12928 9830 12980
rect 11698 12968 11704 12980
rect 11659 12940 11704 12968
rect 11698 12928 11704 12940
rect 11756 12928 11762 12980
rect 11882 12928 11888 12980
rect 11940 12968 11946 12980
rect 12894 12968 12900 12980
rect 11940 12940 12900 12968
rect 11940 12928 11946 12940
rect 12894 12928 12900 12940
rect 12952 12968 12958 12980
rect 12952 12940 13676 12968
rect 12952 12928 12958 12940
rect 10226 12900 10232 12912
rect 9646 12872 10232 12900
rect 8113 12863 8171 12869
rect 7009 12835 7067 12841
rect 7009 12832 7021 12835
rect 6236 12804 7021 12832
rect 6236 12792 6242 12804
rect 7009 12801 7021 12804
rect 7055 12801 7067 12835
rect 7009 12795 7067 12801
rect 7837 12835 7895 12841
rect 7837 12801 7849 12835
rect 7883 12801 7895 12835
rect 7837 12795 7895 12801
rect 5810 12724 5816 12776
rect 5868 12764 5874 12776
rect 5905 12767 5963 12773
rect 5905 12764 5917 12767
rect 5868 12736 5917 12764
rect 5868 12724 5874 12736
rect 5905 12733 5917 12736
rect 5951 12733 5963 12767
rect 5905 12727 5963 12733
rect 6362 12724 6368 12776
rect 6420 12764 6426 12776
rect 8128 12764 8156 12863
rect 10226 12860 10232 12872
rect 10284 12860 10290 12912
rect 11514 12900 11520 12912
rect 10428 12872 11520 12900
rect 10428 12841 10456 12872
rect 11514 12860 11520 12872
rect 11572 12900 11578 12912
rect 12529 12903 12587 12909
rect 11572 12872 12296 12900
rect 11572 12860 11578 12872
rect 12268 12841 12296 12872
rect 12529 12869 12541 12903
rect 12575 12900 12587 12903
rect 13648 12900 13676 12940
rect 13814 12928 13820 12980
rect 13872 12968 13878 12980
rect 14366 12968 14372 12980
rect 13872 12940 14372 12968
rect 13872 12928 13878 12940
rect 14366 12928 14372 12940
rect 14424 12928 14430 12980
rect 15654 12968 15660 12980
rect 15615 12940 15660 12968
rect 15654 12928 15660 12940
rect 15712 12928 15718 12980
rect 14185 12903 14243 12909
rect 14185 12900 14197 12903
rect 12575 12872 12664 12900
rect 13648 12872 14197 12900
rect 12575 12869 12587 12872
rect 12529 12863 12587 12869
rect 10413 12835 10471 12841
rect 10413 12801 10425 12835
rect 10459 12801 10471 12835
rect 10413 12795 10471 12801
rect 10873 12835 10931 12841
rect 10873 12801 10885 12835
rect 10919 12832 10931 12835
rect 12253 12835 12311 12841
rect 10919 12804 11551 12832
rect 10919 12801 10931 12804
rect 10873 12795 10931 12801
rect 11523 12776 11551 12804
rect 12253 12801 12265 12835
rect 12299 12801 12311 12835
rect 12253 12795 12311 12801
rect 6420 12736 8156 12764
rect 8297 12767 8355 12773
rect 6420 12724 6426 12736
rect 8297 12733 8309 12767
rect 8343 12764 8355 12767
rect 8938 12764 8944 12776
rect 8343 12736 8944 12764
rect 8343 12733 8355 12736
rect 8297 12727 8355 12733
rect 8938 12724 8944 12736
rect 8996 12764 9002 12776
rect 9493 12767 9551 12773
rect 9493 12764 9505 12767
rect 8996 12736 9505 12764
rect 8996 12724 9002 12736
rect 9493 12733 9505 12736
rect 9539 12733 9551 12767
rect 9493 12727 9551 12733
rect 10965 12767 11023 12773
rect 10965 12733 10977 12767
rect 11011 12764 11023 12767
rect 11422 12764 11428 12776
rect 11011 12736 11428 12764
rect 11011 12733 11023 12736
rect 10965 12727 11023 12733
rect 11422 12724 11428 12736
rect 11480 12724 11486 12776
rect 11514 12724 11520 12776
rect 11572 12724 11578 12776
rect 11606 12724 11612 12776
rect 11664 12764 11670 12776
rect 12069 12767 12127 12773
rect 12069 12764 12081 12767
rect 11664 12736 12081 12764
rect 11664 12724 11670 12736
rect 12069 12733 12081 12736
rect 12115 12733 12127 12767
rect 12069 12727 12127 12733
rect 1964 12668 3372 12696
rect 2406 12588 2412 12640
rect 2464 12628 2470 12640
rect 2682 12628 2688 12640
rect 2464 12600 2688 12628
rect 2464 12588 2470 12600
rect 2682 12588 2688 12600
rect 2740 12628 2746 12640
rect 2777 12631 2835 12637
rect 2777 12628 2789 12631
rect 2740 12600 2789 12628
rect 2740 12588 2746 12600
rect 2777 12597 2789 12600
rect 2823 12597 2835 12631
rect 2777 12591 2835 12597
rect 2866 12588 2872 12640
rect 2924 12628 2930 12640
rect 3344 12628 3372 12668
rect 3418 12656 3424 12708
rect 3476 12696 3482 12708
rect 3574 12699 3632 12705
rect 3574 12696 3586 12699
rect 3476 12668 3586 12696
rect 3476 12656 3482 12668
rect 3574 12665 3586 12668
rect 3620 12665 3632 12699
rect 3574 12659 3632 12665
rect 4154 12656 4160 12708
rect 4212 12696 4218 12708
rect 6822 12696 6828 12708
rect 4212 12668 6828 12696
rect 4212 12656 4218 12668
rect 6822 12656 6828 12668
rect 6880 12696 6886 12708
rect 7558 12696 7564 12708
rect 6880 12668 7564 12696
rect 6880 12656 6886 12668
rect 7558 12656 7564 12668
rect 7616 12656 7622 12708
rect 7742 12696 7748 12708
rect 7655 12668 7748 12696
rect 7742 12656 7748 12668
rect 7800 12696 7806 12708
rect 8573 12699 8631 12705
rect 8573 12696 8585 12699
rect 7800 12668 8585 12696
rect 7800 12656 7806 12668
rect 8573 12665 8585 12668
rect 8619 12665 8631 12699
rect 11330 12696 11336 12708
rect 8573 12659 8631 12665
rect 9692 12668 11336 12696
rect 4430 12628 4436 12640
rect 2924 12600 2969 12628
rect 3344 12600 4436 12628
rect 2924 12588 2930 12600
rect 4430 12588 4436 12600
rect 4488 12588 4494 12640
rect 5534 12628 5540 12640
rect 5495 12600 5540 12628
rect 5534 12588 5540 12600
rect 5592 12588 5598 12640
rect 6917 12631 6975 12637
rect 6917 12597 6929 12631
rect 6963 12628 6975 12631
rect 7098 12628 7104 12640
rect 6963 12600 7104 12628
rect 6963 12597 6975 12600
rect 6917 12591 6975 12597
rect 7098 12588 7104 12600
rect 7156 12588 7162 12640
rect 7282 12628 7288 12640
rect 7243 12600 7288 12628
rect 7282 12588 7288 12600
rect 7340 12588 7346 12640
rect 7653 12631 7711 12637
rect 7653 12597 7665 12631
rect 7699 12628 7711 12631
rect 7834 12628 7840 12640
rect 7699 12600 7840 12628
rect 7699 12597 7711 12600
rect 7653 12591 7711 12597
rect 7834 12588 7840 12600
rect 7892 12588 7898 12640
rect 9692 12637 9720 12668
rect 11330 12656 11336 12668
rect 11388 12656 11394 12708
rect 12084 12696 12112 12727
rect 12526 12724 12532 12776
rect 12584 12764 12590 12776
rect 12636 12764 12664 12872
rect 14185 12869 14197 12872
rect 14231 12900 14243 12903
rect 15194 12900 15200 12912
rect 14231 12872 15200 12900
rect 14231 12869 14243 12872
rect 14185 12863 14243 12869
rect 15194 12860 15200 12872
rect 15252 12860 15258 12912
rect 12710 12792 12716 12844
rect 12768 12832 12774 12844
rect 13081 12835 13139 12841
rect 13081 12832 13093 12835
rect 12768 12804 13093 12832
rect 12768 12792 12774 12804
rect 13081 12801 13093 12804
rect 13127 12801 13139 12835
rect 13354 12832 13360 12844
rect 13315 12804 13360 12832
rect 13081 12795 13139 12801
rect 13354 12792 13360 12804
rect 13412 12792 13418 12844
rect 15289 12835 15347 12841
rect 15289 12801 15301 12835
rect 15335 12832 15347 12835
rect 15470 12832 15476 12844
rect 15335 12804 15476 12832
rect 15335 12801 15347 12804
rect 15289 12795 15347 12801
rect 15470 12792 15476 12804
rect 15528 12792 15534 12844
rect 13633 12767 13691 12773
rect 13633 12764 13645 12767
rect 12584 12736 12664 12764
rect 12728 12736 13645 12764
rect 12584 12724 12590 12736
rect 12728 12696 12756 12736
rect 13633 12733 13645 12736
rect 13679 12764 13691 12767
rect 14826 12764 14832 12776
rect 13679 12736 14832 12764
rect 13679 12733 13691 12736
rect 13633 12727 13691 12733
rect 14826 12724 14832 12736
rect 14884 12724 14890 12776
rect 14921 12767 14979 12773
rect 14921 12733 14933 12767
rect 14967 12764 14979 12767
rect 15013 12767 15071 12773
rect 15013 12764 15025 12767
rect 14967 12736 15025 12764
rect 14967 12733 14979 12736
rect 14921 12727 14979 12733
rect 15013 12733 15025 12736
rect 15059 12764 15071 12767
rect 15102 12764 15108 12776
rect 15059 12736 15108 12764
rect 15059 12733 15071 12736
rect 15013 12727 15071 12733
rect 15102 12724 15108 12736
rect 15160 12724 15166 12776
rect 12894 12696 12900 12708
rect 11440 12668 11836 12696
rect 12084 12668 12756 12696
rect 12855 12668 12900 12696
rect 9677 12631 9735 12637
rect 9677 12597 9689 12631
rect 9723 12597 9735 12631
rect 10134 12628 10140 12640
rect 10095 12600 10140 12628
rect 9677 12591 9735 12597
rect 10134 12588 10140 12600
rect 10192 12588 10198 12640
rect 10226 12588 10232 12640
rect 10284 12628 10290 12640
rect 10284 12600 10329 12628
rect 10284 12588 10290 12600
rect 10594 12588 10600 12640
rect 10652 12628 10658 12640
rect 11440 12637 11468 12668
rect 11057 12631 11115 12637
rect 11057 12628 11069 12631
rect 10652 12600 11069 12628
rect 10652 12588 10658 12600
rect 11057 12597 11069 12600
rect 11103 12597 11115 12631
rect 11057 12591 11115 12597
rect 11425 12631 11483 12637
rect 11425 12597 11437 12631
rect 11471 12597 11483 12631
rect 11808 12628 11836 12668
rect 12894 12656 12900 12668
rect 12952 12696 12958 12708
rect 13817 12699 13875 12705
rect 13817 12696 13829 12699
rect 12952 12668 13829 12696
rect 12952 12656 12958 12668
rect 13817 12665 13829 12668
rect 13863 12665 13875 12699
rect 13817 12659 13875 12665
rect 14093 12699 14151 12705
rect 14093 12665 14105 12699
rect 14139 12696 14151 12699
rect 14182 12696 14188 12708
rect 14139 12668 14188 12696
rect 14139 12665 14151 12668
rect 14093 12659 14151 12665
rect 12161 12631 12219 12637
rect 12161 12628 12173 12631
rect 11808 12600 12173 12628
rect 11425 12591 11483 12597
rect 12161 12597 12173 12600
rect 12207 12597 12219 12631
rect 12986 12628 12992 12640
rect 12899 12600 12992 12628
rect 12161 12591 12219 12597
rect 12986 12588 12992 12600
rect 13044 12628 13050 12640
rect 14108 12628 14136 12659
rect 14182 12656 14188 12668
rect 14240 12656 14246 12708
rect 13044 12600 14136 12628
rect 13044 12588 13050 12600
rect 1104 12538 16008 12560
rect 1104 12486 5979 12538
rect 6031 12486 6043 12538
rect 6095 12486 6107 12538
rect 6159 12486 6171 12538
rect 6223 12486 10976 12538
rect 11028 12486 11040 12538
rect 11092 12486 11104 12538
rect 11156 12486 11168 12538
rect 11220 12486 16008 12538
rect 1104 12464 16008 12486
rect 1765 12427 1823 12433
rect 1765 12424 1777 12427
rect 1596 12396 1777 12424
rect 1596 12365 1624 12396
rect 1765 12393 1777 12396
rect 1811 12393 1823 12427
rect 3418 12424 3424 12436
rect 3379 12396 3424 12424
rect 1765 12387 1823 12393
rect 3418 12384 3424 12396
rect 3476 12384 3482 12436
rect 3970 12424 3976 12436
rect 3931 12396 3976 12424
rect 3970 12384 3976 12396
rect 4028 12384 4034 12436
rect 4798 12424 4804 12436
rect 4759 12396 4804 12424
rect 4798 12384 4804 12396
rect 4856 12384 4862 12436
rect 4893 12427 4951 12433
rect 4893 12393 4905 12427
rect 4939 12424 4951 12427
rect 5353 12427 5411 12433
rect 5353 12424 5365 12427
rect 4939 12396 5365 12424
rect 4939 12393 4951 12396
rect 4893 12387 4951 12393
rect 5353 12393 5365 12396
rect 5399 12393 5411 12427
rect 5353 12387 5411 12393
rect 5534 12384 5540 12436
rect 5592 12424 5598 12436
rect 5813 12427 5871 12433
rect 5813 12424 5825 12427
rect 5592 12396 5825 12424
rect 5592 12384 5598 12396
rect 5813 12393 5825 12396
rect 5859 12393 5871 12427
rect 5813 12387 5871 12393
rect 6733 12427 6791 12433
rect 6733 12393 6745 12427
rect 6779 12424 6791 12427
rect 7650 12424 7656 12436
rect 6779 12396 7656 12424
rect 6779 12393 6791 12396
rect 6733 12387 6791 12393
rect 7650 12384 7656 12396
rect 7708 12424 7714 12436
rect 8938 12424 8944 12436
rect 7708 12396 8064 12424
rect 8899 12396 8944 12424
rect 7708 12384 7714 12396
rect 1581 12359 1639 12365
rect 1581 12325 1593 12359
rect 1627 12325 1639 12359
rect 2774 12356 2780 12368
rect 1581 12319 1639 12325
rect 2056 12328 2780 12356
rect 1854 12248 1860 12300
rect 1912 12288 1918 12300
rect 2056 12297 2084 12328
rect 2774 12316 2780 12328
rect 2832 12316 2838 12368
rect 7530 12359 7588 12365
rect 7530 12356 7542 12359
rect 4724 12328 7542 12356
rect 2314 12297 2320 12300
rect 1949 12291 2007 12297
rect 1949 12288 1961 12291
rect 1912 12260 1961 12288
rect 1912 12248 1918 12260
rect 1949 12257 1961 12260
rect 1995 12257 2007 12291
rect 1949 12251 2007 12257
rect 2041 12291 2099 12297
rect 2041 12257 2053 12291
rect 2087 12257 2099 12291
rect 2308 12288 2320 12297
rect 2275 12260 2320 12288
rect 2041 12251 2099 12257
rect 2308 12251 2320 12260
rect 2314 12248 2320 12251
rect 2372 12248 2378 12300
rect 4724 12229 4752 12328
rect 7530 12325 7542 12328
rect 7576 12356 7588 12359
rect 7742 12356 7748 12368
rect 7576 12328 7748 12356
rect 7576 12325 7588 12328
rect 7530 12319 7588 12325
rect 7742 12316 7748 12328
rect 7800 12316 7806 12368
rect 8036 12356 8064 12396
rect 8938 12384 8944 12396
rect 8996 12384 9002 12436
rect 10410 12424 10416 12436
rect 9048 12396 10416 12424
rect 9048 12356 9076 12396
rect 10410 12384 10416 12396
rect 10468 12384 10474 12436
rect 10594 12424 10600 12436
rect 10555 12396 10600 12424
rect 10594 12384 10600 12396
rect 10652 12384 10658 12436
rect 11606 12424 11612 12436
rect 10704 12396 11612 12424
rect 8036 12328 9076 12356
rect 10042 12316 10048 12368
rect 10100 12356 10106 12368
rect 10704 12356 10732 12396
rect 11606 12384 11612 12396
rect 11664 12384 11670 12436
rect 12621 12427 12679 12433
rect 12621 12393 12633 12427
rect 12667 12424 12679 12427
rect 12710 12424 12716 12436
rect 12667 12396 12716 12424
rect 12667 12393 12679 12396
rect 12621 12387 12679 12393
rect 12710 12384 12716 12396
rect 12768 12384 12774 12436
rect 13998 12356 14004 12368
rect 10100 12328 10732 12356
rect 10796 12328 14004 12356
rect 10100 12316 10106 12328
rect 5534 12248 5540 12300
rect 5592 12288 5598 12300
rect 5721 12291 5779 12297
rect 5721 12288 5733 12291
rect 5592 12260 5733 12288
rect 5592 12248 5598 12260
rect 5721 12257 5733 12260
rect 5767 12288 5779 12291
rect 6178 12288 6184 12300
rect 5767 12260 6184 12288
rect 5767 12257 5779 12260
rect 5721 12251 5779 12257
rect 6178 12248 6184 12260
rect 6236 12248 6242 12300
rect 6454 12248 6460 12300
rect 6512 12288 6518 12300
rect 6825 12291 6883 12297
rect 6512 12260 6776 12288
rect 6512 12248 6518 12260
rect 4709 12223 4767 12229
rect 4709 12189 4721 12223
rect 4755 12189 4767 12223
rect 4709 12183 4767 12189
rect 5997 12223 6055 12229
rect 5997 12189 6009 12223
rect 6043 12220 6055 12223
rect 6270 12220 6276 12232
rect 6043 12192 6276 12220
rect 6043 12189 6055 12192
rect 5997 12183 6055 12189
rect 6270 12180 6276 12192
rect 6328 12220 6334 12232
rect 6638 12220 6644 12232
rect 6328 12192 6644 12220
rect 6328 12180 6334 12192
rect 6638 12180 6644 12192
rect 6696 12180 6702 12232
rect 6748 12220 6776 12260
rect 6825 12257 6837 12291
rect 6871 12288 6883 12291
rect 8294 12288 8300 12300
rect 6871 12260 8300 12288
rect 6871 12257 6883 12260
rect 6825 12251 6883 12257
rect 8294 12248 8300 12260
rect 8352 12248 8358 12300
rect 8757 12291 8815 12297
rect 8757 12257 8769 12291
rect 8803 12288 8815 12291
rect 8938 12288 8944 12300
rect 8803 12260 8944 12288
rect 8803 12257 8815 12260
rect 8757 12251 8815 12257
rect 8938 12248 8944 12260
rect 8996 12248 9002 12300
rect 9381 12291 9439 12297
rect 9381 12288 9393 12291
rect 9048 12260 9393 12288
rect 7285 12223 7343 12229
rect 7285 12220 7297 12223
rect 6748 12192 7297 12220
rect 7285 12189 7297 12192
rect 7331 12189 7343 12223
rect 9048 12220 9076 12260
rect 9381 12257 9393 12260
rect 9427 12257 9439 12291
rect 9381 12251 9439 12257
rect 7285 12183 7343 12189
rect 8680 12192 9076 12220
rect 5350 12112 5356 12164
rect 5408 12152 5414 12164
rect 5408 12124 7328 12152
rect 5408 12112 5414 12124
rect 1486 12084 1492 12096
rect 1447 12056 1492 12084
rect 1486 12044 1492 12056
rect 1544 12044 1550 12096
rect 2682 12044 2688 12096
rect 2740 12084 2746 12096
rect 3605 12087 3663 12093
rect 3605 12084 3617 12087
rect 2740 12056 3617 12084
rect 2740 12044 2746 12056
rect 3605 12053 3617 12056
rect 3651 12084 3663 12087
rect 4798 12084 4804 12096
rect 3651 12056 4804 12084
rect 3651 12053 3663 12056
rect 3605 12047 3663 12053
rect 4798 12044 4804 12056
rect 4856 12044 4862 12096
rect 5166 12044 5172 12096
rect 5224 12084 5230 12096
rect 5261 12087 5319 12093
rect 5261 12084 5273 12087
rect 5224 12056 5273 12084
rect 5224 12044 5230 12056
rect 5261 12053 5273 12056
rect 5307 12053 5319 12087
rect 6270 12084 6276 12096
rect 6231 12056 6276 12084
rect 5261 12047 5319 12053
rect 6270 12044 6276 12056
rect 6328 12044 6334 12096
rect 7098 12044 7104 12096
rect 7156 12084 7162 12096
rect 7193 12087 7251 12093
rect 7193 12084 7205 12087
rect 7156 12056 7205 12084
rect 7156 12044 7162 12056
rect 7193 12053 7205 12056
rect 7239 12053 7251 12087
rect 7300 12084 7328 12124
rect 8680 12093 8708 12192
rect 9122 12180 9128 12232
rect 9180 12220 9186 12232
rect 9180 12192 9225 12220
rect 9180 12180 9186 12192
rect 10410 12180 10416 12232
rect 10468 12220 10474 12232
rect 10796 12220 10824 12328
rect 13998 12316 14004 12328
rect 14056 12356 14062 12368
rect 14550 12356 14556 12368
rect 14056 12328 14556 12356
rect 14056 12316 14062 12328
rect 14550 12316 14556 12328
rect 14608 12316 14614 12368
rect 11514 12297 11520 12300
rect 11508 12288 11520 12297
rect 10468 12192 10824 12220
rect 11072 12260 11520 12288
rect 10468 12180 10474 12192
rect 10505 12155 10563 12161
rect 10505 12121 10517 12155
rect 10551 12152 10563 12155
rect 11072 12152 11100 12260
rect 11508 12251 11520 12260
rect 11514 12248 11520 12251
rect 11572 12248 11578 12300
rect 12897 12291 12955 12297
rect 12897 12257 12909 12291
rect 12943 12288 12955 12291
rect 13817 12291 13875 12297
rect 13817 12288 13829 12291
rect 12943 12260 13829 12288
rect 12943 12257 12955 12260
rect 12897 12251 12955 12257
rect 13817 12257 13829 12260
rect 13863 12288 13875 12291
rect 14918 12288 14924 12300
rect 13863 12260 14924 12288
rect 13863 12257 13875 12260
rect 13817 12251 13875 12257
rect 14918 12248 14924 12260
rect 14976 12288 14982 12300
rect 15102 12288 15108 12300
rect 14976 12260 15108 12288
rect 14976 12248 14982 12260
rect 15102 12248 15108 12260
rect 15160 12248 15166 12300
rect 11238 12220 11244 12232
rect 11199 12192 11244 12220
rect 11238 12180 11244 12192
rect 11296 12180 11302 12232
rect 12802 12180 12808 12232
rect 12860 12220 12866 12232
rect 13173 12223 13231 12229
rect 13173 12220 13185 12223
rect 12860 12192 13185 12220
rect 12860 12180 12866 12192
rect 13173 12189 13185 12192
rect 13219 12189 13231 12223
rect 13173 12183 13231 12189
rect 10551 12124 11100 12152
rect 10551 12121 10563 12124
rect 10505 12115 10563 12121
rect 8665 12087 8723 12093
rect 8665 12084 8677 12087
rect 7300 12056 8677 12084
rect 7193 12047 7251 12053
rect 8665 12053 8677 12056
rect 8711 12053 8723 12087
rect 8665 12047 8723 12053
rect 10778 12044 10784 12096
rect 10836 12084 10842 12096
rect 10873 12087 10931 12093
rect 10873 12084 10885 12087
rect 10836 12056 10885 12084
rect 10836 12044 10842 12056
rect 10873 12053 10885 12056
rect 10919 12053 10931 12087
rect 11054 12084 11060 12096
rect 11015 12056 11060 12084
rect 10873 12047 10931 12053
rect 11054 12044 11060 12056
rect 11112 12084 11118 12096
rect 11422 12084 11428 12096
rect 11112 12056 11428 12084
rect 11112 12044 11118 12056
rect 11422 12044 11428 12056
rect 11480 12044 11486 12096
rect 1104 11994 16008 12016
rect 1104 11942 3480 11994
rect 3532 11942 3544 11994
rect 3596 11942 3608 11994
rect 3660 11942 3672 11994
rect 3724 11942 8478 11994
rect 8530 11942 8542 11994
rect 8594 11942 8606 11994
rect 8658 11942 8670 11994
rect 8722 11942 13475 11994
rect 13527 11942 13539 11994
rect 13591 11942 13603 11994
rect 13655 11942 13667 11994
rect 13719 11942 16008 11994
rect 1104 11920 16008 11942
rect 3326 11840 3332 11892
rect 3384 11880 3390 11892
rect 3789 11883 3847 11889
rect 3789 11880 3801 11883
rect 3384 11852 3801 11880
rect 3384 11840 3390 11852
rect 3789 11849 3801 11852
rect 3835 11880 3847 11883
rect 4338 11880 4344 11892
rect 3835 11852 4344 11880
rect 3835 11849 3847 11852
rect 3789 11843 3847 11849
rect 4338 11840 4344 11852
rect 4396 11840 4402 11892
rect 4430 11840 4436 11892
rect 4488 11880 4494 11892
rect 4709 11883 4767 11889
rect 4709 11880 4721 11883
rect 4488 11852 4721 11880
rect 4488 11840 4494 11852
rect 4709 11849 4721 11852
rect 4755 11849 4767 11883
rect 4709 11843 4767 11849
rect 4798 11840 4804 11892
rect 4856 11880 4862 11892
rect 9674 11880 9680 11892
rect 4856 11852 9680 11880
rect 4856 11840 4862 11852
rect 9674 11840 9680 11852
rect 9732 11880 9738 11892
rect 9769 11883 9827 11889
rect 9769 11880 9781 11883
rect 9732 11852 9781 11880
rect 9732 11840 9738 11852
rect 9769 11849 9781 11852
rect 9815 11849 9827 11883
rect 9769 11843 9827 11849
rect 9953 11883 10011 11889
rect 9953 11849 9965 11883
rect 9999 11880 10011 11883
rect 10226 11880 10232 11892
rect 9999 11852 10232 11880
rect 9999 11849 10011 11852
rect 9953 11843 10011 11849
rect 10226 11840 10232 11852
rect 10284 11840 10290 11892
rect 2774 11772 2780 11824
rect 2832 11812 2838 11824
rect 5534 11812 5540 11824
rect 2832 11784 5540 11812
rect 2832 11772 2838 11784
rect 5534 11772 5540 11784
rect 5592 11772 5598 11824
rect 7484 11784 9674 11812
rect 3786 11744 3792 11756
rect 2700 11716 3792 11744
rect 2700 11688 2728 11716
rect 3786 11704 3792 11716
rect 3844 11744 3850 11756
rect 4433 11747 4491 11753
rect 4433 11744 4445 11747
rect 3844 11716 4445 11744
rect 3844 11704 3850 11716
rect 4433 11713 4445 11716
rect 4479 11713 4491 11747
rect 5166 11744 5172 11756
rect 5127 11716 5172 11744
rect 4433 11707 4491 11713
rect 5166 11704 5172 11716
rect 5224 11704 5230 11756
rect 5350 11744 5356 11756
rect 5311 11716 5356 11744
rect 5350 11704 5356 11716
rect 5408 11704 5414 11756
rect 5552 11744 5580 11772
rect 6454 11744 6460 11756
rect 5552 11716 6460 11744
rect 6454 11704 6460 11716
rect 6512 11704 6518 11756
rect 2521 11679 2579 11685
rect 2521 11645 2533 11679
rect 2567 11676 2579 11679
rect 2682 11676 2688 11688
rect 2567 11648 2688 11676
rect 2567 11645 2579 11648
rect 2521 11639 2579 11645
rect 2682 11636 2688 11648
rect 2740 11636 2746 11688
rect 2774 11636 2780 11688
rect 2832 11676 2838 11688
rect 5718 11676 5724 11688
rect 2832 11648 2877 11676
rect 5679 11648 5724 11676
rect 2832 11636 2838 11648
rect 5718 11636 5724 11648
rect 5776 11636 5782 11688
rect 6362 11636 6368 11688
rect 6420 11676 6426 11688
rect 7484 11676 7512 11784
rect 8202 11704 8208 11756
rect 8260 11744 8266 11756
rect 8481 11747 8539 11753
rect 8481 11744 8493 11747
rect 8260 11716 8493 11744
rect 8260 11704 8266 11716
rect 8481 11713 8493 11716
rect 8527 11713 8539 11747
rect 9646 11744 9674 11784
rect 10134 11772 10140 11824
rect 10192 11812 10198 11824
rect 10781 11815 10839 11821
rect 10781 11812 10793 11815
rect 10192 11784 10793 11812
rect 10192 11772 10198 11784
rect 10781 11781 10793 11784
rect 10827 11781 10839 11815
rect 10781 11775 10839 11781
rect 11238 11772 11244 11824
rect 11296 11812 11302 11824
rect 11790 11812 11796 11824
rect 11296 11784 11796 11812
rect 11296 11772 11302 11784
rect 11790 11772 11796 11784
rect 11848 11812 11854 11824
rect 11885 11815 11943 11821
rect 11885 11812 11897 11815
rect 11848 11784 11897 11812
rect 11848 11772 11854 11784
rect 11885 11781 11897 11784
rect 11931 11781 11943 11815
rect 11885 11775 11943 11781
rect 9646 11716 9996 11744
rect 8481 11707 8539 11713
rect 6420 11648 7512 11676
rect 6420 11636 6426 11648
rect 7926 11636 7932 11688
rect 7984 11676 7990 11688
rect 8110 11676 8116 11688
rect 7984 11648 8116 11676
rect 7984 11636 7990 11648
rect 8110 11636 8116 11648
rect 8168 11636 8174 11688
rect 8389 11679 8447 11685
rect 8389 11645 8401 11679
rect 8435 11676 8447 11679
rect 9766 11676 9772 11688
rect 8435 11648 9772 11676
rect 8435 11645 8447 11648
rect 8389 11639 8447 11645
rect 9766 11636 9772 11648
rect 9824 11636 9830 11688
rect 9968 11676 9996 11716
rect 10226 11704 10232 11756
rect 10284 11744 10290 11756
rect 10413 11747 10471 11753
rect 10413 11744 10425 11747
rect 10284 11716 10425 11744
rect 10284 11704 10290 11716
rect 10413 11713 10425 11716
rect 10459 11713 10471 11747
rect 10413 11707 10471 11713
rect 10597 11747 10655 11753
rect 10597 11713 10609 11747
rect 10643 11744 10655 11747
rect 11333 11747 11391 11753
rect 11333 11744 11345 11747
rect 10643 11716 11345 11744
rect 10643 11713 10655 11716
rect 10597 11707 10655 11713
rect 11333 11713 11345 11716
rect 11379 11744 11391 11747
rect 11514 11744 11520 11756
rect 11379 11716 11520 11744
rect 11379 11713 11391 11716
rect 11333 11707 11391 11713
rect 11514 11704 11520 11716
rect 11572 11704 11578 11756
rect 11054 11676 11060 11688
rect 9968 11648 11060 11676
rect 11054 11636 11060 11648
rect 11112 11636 11118 11688
rect 11422 11636 11428 11688
rect 11480 11676 11486 11688
rect 11701 11679 11759 11685
rect 11701 11676 11713 11679
rect 11480 11648 11713 11676
rect 11480 11636 11486 11648
rect 11701 11645 11713 11648
rect 11747 11645 11759 11679
rect 11701 11639 11759 11645
rect 4154 11608 4160 11620
rect 3528 11580 4160 11608
rect 1397 11543 1455 11549
rect 1397 11509 1409 11543
rect 1443 11540 1455 11543
rect 2314 11540 2320 11552
rect 1443 11512 2320 11540
rect 1443 11509 1455 11512
rect 1397 11503 1455 11509
rect 2314 11500 2320 11512
rect 2372 11500 2378 11552
rect 3142 11500 3148 11552
rect 3200 11540 3206 11552
rect 3528 11549 3556 11580
rect 4154 11568 4160 11580
rect 4212 11568 4218 11620
rect 5258 11568 5264 11620
rect 5316 11608 5322 11620
rect 6454 11608 6460 11620
rect 5316 11580 6460 11608
rect 5316 11568 5322 11580
rect 6454 11568 6460 11580
rect 6512 11568 6518 11620
rect 6638 11568 6644 11620
rect 6696 11617 6702 11620
rect 6696 11611 6760 11617
rect 6696 11577 6714 11611
rect 6748 11577 6760 11611
rect 6696 11571 6760 11577
rect 6696 11568 6702 11571
rect 6914 11568 6920 11620
rect 6972 11608 6978 11620
rect 10502 11608 10508 11620
rect 6972 11580 10508 11608
rect 6972 11568 6978 11580
rect 10502 11568 10508 11580
rect 10560 11568 10566 11620
rect 10686 11568 10692 11620
rect 10744 11608 10750 11620
rect 11241 11611 11299 11617
rect 11241 11608 11253 11611
rect 10744 11580 11253 11608
rect 10744 11568 10750 11580
rect 11241 11577 11253 11580
rect 11287 11608 11299 11611
rect 11977 11611 12035 11617
rect 11977 11608 11989 11611
rect 11287 11580 11989 11608
rect 11287 11577 11299 11580
rect 11241 11571 11299 11577
rect 11977 11577 11989 11580
rect 12023 11577 12035 11611
rect 11977 11571 12035 11577
rect 3513 11543 3571 11549
rect 3513 11540 3525 11543
rect 3200 11512 3525 11540
rect 3200 11500 3206 11512
rect 3513 11509 3525 11512
rect 3559 11509 3571 11543
rect 3878 11540 3884 11552
rect 3839 11512 3884 11540
rect 3513 11503 3571 11509
rect 3878 11500 3884 11512
rect 3936 11500 3942 11552
rect 4246 11540 4252 11552
rect 4207 11512 4252 11540
rect 4246 11500 4252 11512
rect 4304 11500 4310 11552
rect 4338 11500 4344 11552
rect 4396 11540 4402 11552
rect 5077 11543 5135 11549
rect 4396 11512 4441 11540
rect 4396 11500 4402 11512
rect 5077 11509 5089 11543
rect 5123 11540 5135 11543
rect 5442 11540 5448 11552
rect 5123 11512 5448 11540
rect 5123 11509 5135 11512
rect 5077 11503 5135 11509
rect 5442 11500 5448 11512
rect 5500 11500 5506 11552
rect 7742 11500 7748 11552
rect 7800 11540 7806 11552
rect 7837 11543 7895 11549
rect 7837 11540 7849 11543
rect 7800 11512 7849 11540
rect 7800 11500 7806 11512
rect 7837 11509 7849 11512
rect 7883 11509 7895 11543
rect 7837 11503 7895 11509
rect 7926 11500 7932 11552
rect 7984 11540 7990 11552
rect 8294 11540 8300 11552
rect 7984 11512 8029 11540
rect 8255 11512 8300 11540
rect 7984 11500 7990 11512
rect 8294 11500 8300 11512
rect 8352 11500 8358 11552
rect 8386 11500 8392 11552
rect 8444 11540 8450 11552
rect 8757 11543 8815 11549
rect 8757 11540 8769 11543
rect 8444 11512 8769 11540
rect 8444 11500 8450 11512
rect 8757 11509 8769 11512
rect 8803 11509 8815 11543
rect 8757 11503 8815 11509
rect 9214 11500 9220 11552
rect 9272 11540 9278 11552
rect 9582 11540 9588 11552
rect 9272 11512 9588 11540
rect 9272 11500 9278 11512
rect 9582 11500 9588 11512
rect 9640 11540 9646 11552
rect 10321 11543 10379 11549
rect 10321 11540 10333 11543
rect 9640 11512 10333 11540
rect 9640 11500 9646 11512
rect 10321 11509 10333 11512
rect 10367 11509 10379 11543
rect 10321 11503 10379 11509
rect 10778 11500 10784 11552
rect 10836 11540 10842 11552
rect 11149 11543 11207 11549
rect 11149 11540 11161 11543
rect 10836 11512 11161 11540
rect 10836 11500 10842 11512
rect 11149 11509 11161 11512
rect 11195 11540 11207 11543
rect 12161 11543 12219 11549
rect 12161 11540 12173 11543
rect 11195 11512 12173 11540
rect 11195 11509 11207 11512
rect 11149 11503 11207 11509
rect 12161 11509 12173 11512
rect 12207 11509 12219 11543
rect 12161 11503 12219 11509
rect 12437 11543 12495 11549
rect 12437 11509 12449 11543
rect 12483 11540 12495 11543
rect 12526 11540 12532 11552
rect 12483 11512 12532 11540
rect 12483 11509 12495 11512
rect 12437 11503 12495 11509
rect 12526 11500 12532 11512
rect 12584 11540 12590 11552
rect 12710 11540 12716 11552
rect 12584 11512 12716 11540
rect 12584 11500 12590 11512
rect 12710 11500 12716 11512
rect 12768 11500 12774 11552
rect 1104 11450 16008 11472
rect 1104 11398 5979 11450
rect 6031 11398 6043 11450
rect 6095 11398 6107 11450
rect 6159 11398 6171 11450
rect 6223 11398 10976 11450
rect 11028 11398 11040 11450
rect 11092 11398 11104 11450
rect 11156 11398 11168 11450
rect 11220 11398 16008 11450
rect 1104 11376 16008 11398
rect 1854 11336 1860 11348
rect 1815 11308 1860 11336
rect 1854 11296 1860 11308
rect 1912 11296 1918 11348
rect 2225 11339 2283 11345
rect 2225 11305 2237 11339
rect 2271 11336 2283 11339
rect 3878 11336 3884 11348
rect 2271 11308 3884 11336
rect 2271 11305 2283 11308
rect 2225 11299 2283 11305
rect 3878 11296 3884 11308
rect 3936 11296 3942 11348
rect 4246 11296 4252 11348
rect 4304 11336 4310 11348
rect 5353 11339 5411 11345
rect 5353 11336 5365 11339
rect 4304 11308 5365 11336
rect 4304 11296 4310 11308
rect 5353 11305 5365 11308
rect 5399 11305 5411 11339
rect 5353 11299 5411 11305
rect 5442 11296 5448 11348
rect 5500 11336 5506 11348
rect 6733 11339 6791 11345
rect 6733 11336 6745 11339
rect 5500 11308 6745 11336
rect 5500 11296 5506 11308
rect 6733 11305 6745 11308
rect 6779 11305 6791 11339
rect 7098 11336 7104 11348
rect 7059 11308 7104 11336
rect 6733 11299 6791 11305
rect 7098 11296 7104 11308
rect 7156 11296 7162 11348
rect 7193 11339 7251 11345
rect 7193 11305 7205 11339
rect 7239 11336 7251 11339
rect 7282 11336 7288 11348
rect 7239 11308 7288 11336
rect 7239 11305 7251 11308
rect 7193 11299 7251 11305
rect 7282 11296 7288 11308
rect 7340 11296 7346 11348
rect 7650 11336 7656 11348
rect 7611 11308 7656 11336
rect 7650 11296 7656 11308
rect 7708 11296 7714 11348
rect 9769 11339 9827 11345
rect 9769 11305 9781 11339
rect 9815 11336 9827 11339
rect 10042 11336 10048 11348
rect 9815 11308 10048 11336
rect 9815 11305 9827 11308
rect 9769 11299 9827 11305
rect 10042 11296 10048 11308
rect 10100 11336 10106 11348
rect 10229 11339 10287 11345
rect 10229 11336 10241 11339
rect 10100 11308 10241 11336
rect 10100 11296 10106 11308
rect 10229 11305 10241 11308
rect 10275 11305 10287 11339
rect 10229 11299 10287 11305
rect 10502 11296 10508 11348
rect 10560 11336 10566 11348
rect 14642 11336 14648 11348
rect 10560 11308 14648 11336
rect 10560 11296 10566 11308
rect 14642 11296 14648 11308
rect 14700 11296 14706 11348
rect 2314 11228 2320 11280
rect 2372 11268 2378 11280
rect 3237 11271 3295 11277
rect 2372 11240 2452 11268
rect 2372 11228 2378 11240
rect 1578 11200 1584 11212
rect 1539 11172 1584 11200
rect 1578 11160 1584 11172
rect 1636 11160 1642 11212
rect 2314 11132 2320 11144
rect 2275 11104 2320 11132
rect 2314 11092 2320 11104
rect 2372 11092 2378 11144
rect 2424 11141 2452 11240
rect 3237 11237 3249 11271
rect 3283 11268 3295 11271
rect 3326 11268 3332 11280
rect 3283 11240 3332 11268
rect 3283 11237 3295 11240
rect 3237 11231 3295 11237
rect 3326 11228 3332 11240
rect 3384 11228 3390 11280
rect 5016 11271 5074 11277
rect 5016 11268 5028 11271
rect 4264 11240 5028 11268
rect 3970 11160 3976 11212
rect 4028 11200 4034 11212
rect 4264 11200 4292 11240
rect 5016 11237 5028 11240
rect 5062 11268 5074 11271
rect 5062 11240 6040 11268
rect 5062 11237 5074 11240
rect 5016 11231 5074 11237
rect 4028 11172 4292 11200
rect 5261 11203 5319 11209
rect 4028 11160 4034 11172
rect 5261 11169 5273 11203
rect 5307 11200 5319 11203
rect 5534 11200 5540 11212
rect 5307 11172 5540 11200
rect 5307 11169 5319 11172
rect 5261 11163 5319 11169
rect 5534 11160 5540 11172
rect 5592 11160 5598 11212
rect 5718 11200 5724 11212
rect 5679 11172 5724 11200
rect 5718 11160 5724 11172
rect 5776 11160 5782 11212
rect 2409 11135 2467 11141
rect 2409 11101 2421 11135
rect 2455 11101 2467 11135
rect 2409 11095 2467 11101
rect 3142 11092 3148 11144
rect 3200 11132 3206 11144
rect 3329 11135 3387 11141
rect 3329 11132 3341 11135
rect 3200 11104 3341 11132
rect 3200 11092 3206 11104
rect 3329 11101 3341 11104
rect 3375 11101 3387 11135
rect 3329 11095 3387 11101
rect 3513 11135 3571 11141
rect 3513 11101 3525 11135
rect 3559 11132 3571 11135
rect 3988 11132 4016 11160
rect 6012 11144 6040 11240
rect 6270 11228 6276 11280
rect 6328 11268 6334 11280
rect 12894 11268 12900 11280
rect 6328 11240 12900 11268
rect 6328 11228 6334 11240
rect 12894 11228 12900 11240
rect 12952 11228 12958 11280
rect 6822 11160 6828 11212
rect 6880 11200 6886 11212
rect 8018 11200 8024 11212
rect 6880 11172 8024 11200
rect 6880 11160 6886 11172
rect 8018 11160 8024 11172
rect 8076 11160 8082 11212
rect 8297 11203 8355 11209
rect 8297 11169 8309 11203
rect 8343 11200 8355 11203
rect 8846 11200 8852 11212
rect 8343 11172 8852 11200
rect 8343 11169 8355 11172
rect 8297 11163 8355 11169
rect 8846 11160 8852 11172
rect 8904 11160 8910 11212
rect 9309 11203 9367 11209
rect 9309 11169 9321 11203
rect 9355 11200 9367 11203
rect 9582 11200 9588 11212
rect 9355 11172 9588 11200
rect 9355 11169 9367 11172
rect 9309 11163 9367 11169
rect 9582 11160 9588 11172
rect 9640 11200 9646 11212
rect 10042 11200 10048 11212
rect 9640 11172 10048 11200
rect 9640 11160 9646 11172
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 11514 11160 11520 11212
rect 11572 11200 11578 11212
rect 12158 11200 12164 11212
rect 11572 11172 12164 11200
rect 11572 11160 11578 11172
rect 12158 11160 12164 11172
rect 12216 11160 12222 11212
rect 12733 11203 12791 11209
rect 12733 11169 12745 11203
rect 12779 11200 12791 11203
rect 14182 11200 14188 11212
rect 12779 11172 14188 11200
rect 12779 11169 12791 11172
rect 12733 11163 12791 11169
rect 14182 11160 14188 11172
rect 14240 11160 14246 11212
rect 3559 11104 4016 11132
rect 5813 11135 5871 11141
rect 3559 11101 3571 11104
rect 3513 11095 3571 11101
rect 5813 11101 5825 11135
rect 5859 11101 5871 11135
rect 5994 11132 6000 11144
rect 5955 11104 6000 11132
rect 5813 11095 5871 11101
rect 1394 11064 1400 11076
rect 1355 11036 1400 11064
rect 1394 11024 1400 11036
rect 1452 11024 1458 11076
rect 3786 11024 3792 11076
rect 3844 11064 3850 11076
rect 3881 11067 3939 11073
rect 3881 11064 3893 11067
rect 3844 11036 3893 11064
rect 3844 11024 3850 11036
rect 3881 11033 3893 11036
rect 3927 11033 3939 11067
rect 5828 11064 5856 11095
rect 5994 11092 6000 11104
rect 6052 11092 6058 11144
rect 6273 11135 6331 11141
rect 6273 11101 6285 11135
rect 6319 11132 6331 11135
rect 6914 11132 6920 11144
rect 6319 11104 6920 11132
rect 6319 11101 6331 11104
rect 6273 11095 6331 11101
rect 6288 11064 6316 11095
rect 6914 11092 6920 11104
rect 6972 11092 6978 11144
rect 7377 11135 7435 11141
rect 7377 11101 7389 11135
rect 7423 11132 7435 11135
rect 7742 11132 7748 11144
rect 7423 11104 7748 11132
rect 7423 11101 7435 11104
rect 7377 11095 7435 11101
rect 7742 11092 7748 11104
rect 7800 11092 7806 11144
rect 8389 11135 8447 11141
rect 8389 11101 8401 11135
rect 8435 11101 8447 11135
rect 8389 11095 8447 11101
rect 8573 11135 8631 11141
rect 8573 11101 8585 11135
rect 8619 11132 8631 11135
rect 8938 11132 8944 11144
rect 8619 11104 8944 11132
rect 8619 11101 8631 11104
rect 8573 11095 8631 11101
rect 5828 11036 6316 11064
rect 3881 11027 3939 11033
rect 7282 11024 7288 11076
rect 7340 11064 7346 11076
rect 8202 11064 8208 11076
rect 7340 11036 8208 11064
rect 7340 11024 7346 11036
rect 8202 11024 8208 11036
rect 8260 11024 8266 11076
rect 8404 11064 8432 11095
rect 8938 11092 8944 11104
rect 8996 11132 9002 11144
rect 9493 11135 9551 11141
rect 9493 11132 9505 11135
rect 8996 11104 9505 11132
rect 8996 11092 9002 11104
rect 9493 11101 9505 11104
rect 9539 11101 9551 11135
rect 9674 11132 9680 11144
rect 9635 11104 9680 11132
rect 9493 11095 9551 11101
rect 9674 11092 9680 11104
rect 9732 11092 9738 11144
rect 11882 11132 11888 11144
rect 9968 11104 11888 11132
rect 8849 11067 8907 11073
rect 8849 11064 8861 11067
rect 8404 11036 8861 11064
rect 8849 11033 8861 11036
rect 8895 11064 8907 11067
rect 9968 11064 9996 11104
rect 11882 11092 11888 11104
rect 11940 11092 11946 11144
rect 12986 11132 12992 11144
rect 12947 11104 12992 11132
rect 12986 11092 12992 11104
rect 13044 11092 13050 11144
rect 10134 11064 10140 11076
rect 8895 11036 9996 11064
rect 10095 11036 10140 11064
rect 8895 11033 8907 11036
rect 8849 11027 8907 11033
rect 10134 11024 10140 11036
rect 10192 11024 10198 11076
rect 10318 11024 10324 11076
rect 10376 11064 10382 11076
rect 10778 11064 10784 11076
rect 10376 11036 10784 11064
rect 10376 11024 10382 11036
rect 10778 11024 10784 11036
rect 10836 11024 10842 11076
rect 11790 11064 11796 11076
rect 11348 11036 11796 11064
rect 2866 10996 2872 11008
rect 2827 10968 2872 10996
rect 2866 10956 2872 10968
rect 2924 10956 2930 11008
rect 6914 10956 6920 11008
rect 6972 10996 6978 11008
rect 7098 10996 7104 11008
rect 6972 10968 7104 10996
rect 6972 10956 6978 10968
rect 7098 10956 7104 10968
rect 7156 10956 7162 11008
rect 7926 10996 7932 11008
rect 7887 10968 7932 10996
rect 7926 10956 7932 10968
rect 7984 10956 7990 11008
rect 9122 10956 9128 11008
rect 9180 10996 9186 11008
rect 11348 10996 11376 11036
rect 11790 11024 11796 11036
rect 11848 11024 11854 11076
rect 11606 10996 11612 11008
rect 9180 10968 11376 10996
rect 11567 10968 11612 10996
rect 9180 10956 9186 10968
rect 11606 10956 11612 10968
rect 11664 10956 11670 11008
rect 1104 10906 16008 10928
rect 1104 10854 3480 10906
rect 3532 10854 3544 10906
rect 3596 10854 3608 10906
rect 3660 10854 3672 10906
rect 3724 10854 8478 10906
rect 8530 10854 8542 10906
rect 8594 10854 8606 10906
rect 8658 10854 8670 10906
rect 8722 10854 13475 10906
rect 13527 10854 13539 10906
rect 13591 10854 13603 10906
rect 13655 10854 13667 10906
rect 13719 10854 16008 10906
rect 1104 10832 16008 10854
rect 1489 10795 1547 10801
rect 1489 10761 1501 10795
rect 1535 10792 1547 10795
rect 1578 10792 1584 10804
rect 1535 10764 1584 10792
rect 1535 10761 1547 10764
rect 1489 10755 1547 10761
rect 1578 10752 1584 10764
rect 1636 10752 1642 10804
rect 2041 10795 2099 10801
rect 2041 10761 2053 10795
rect 2087 10792 2099 10795
rect 2314 10792 2320 10804
rect 2087 10764 2320 10792
rect 2087 10761 2099 10764
rect 2041 10755 2099 10761
rect 2314 10752 2320 10764
rect 2372 10752 2378 10804
rect 3970 10792 3976 10804
rect 3931 10764 3976 10792
rect 3970 10752 3976 10764
rect 4028 10752 4034 10804
rect 4338 10752 4344 10804
rect 4396 10792 4402 10804
rect 5445 10795 5503 10801
rect 5445 10792 5457 10795
rect 4396 10764 5457 10792
rect 4396 10752 4402 10764
rect 5445 10761 5457 10764
rect 5491 10761 5503 10795
rect 5445 10755 5503 10761
rect 7653 10795 7711 10801
rect 7653 10761 7665 10795
rect 7699 10792 7711 10795
rect 8202 10792 8208 10804
rect 7699 10764 8208 10792
rect 7699 10761 7711 10764
rect 7653 10755 7711 10761
rect 8202 10752 8208 10764
rect 8260 10752 8266 10804
rect 9674 10752 9680 10804
rect 9732 10792 9738 10804
rect 10689 10795 10747 10801
rect 10689 10792 10701 10795
rect 9732 10764 10701 10792
rect 9732 10752 9738 10764
rect 10689 10761 10701 10764
rect 10735 10761 10747 10795
rect 10689 10755 10747 10761
rect 10778 10752 10784 10804
rect 10836 10792 10842 10804
rect 12618 10792 12624 10804
rect 10836 10764 12624 10792
rect 10836 10752 10842 10764
rect 12618 10752 12624 10764
rect 12676 10752 12682 10804
rect 12986 10792 12992 10804
rect 12820 10764 12992 10792
rect 1688 10696 3464 10724
rect 1688 10597 1716 10696
rect 2682 10656 2688 10668
rect 2643 10628 2688 10656
rect 2682 10616 2688 10628
rect 2740 10616 2746 10668
rect 1673 10591 1731 10597
rect 1673 10557 1685 10591
rect 1719 10557 1731 10591
rect 1673 10551 1731 10557
rect 2409 10591 2467 10597
rect 2409 10557 2421 10591
rect 2455 10588 2467 10591
rect 2866 10588 2872 10600
rect 2455 10560 2872 10588
rect 2455 10557 2467 10560
rect 2409 10551 2467 10557
rect 2866 10548 2872 10560
rect 2924 10548 2930 10600
rect 3436 10588 3464 10696
rect 3513 10659 3571 10665
rect 3513 10625 3525 10659
rect 3559 10656 3571 10659
rect 3988 10656 4016 10752
rect 7834 10724 7840 10736
rect 5368 10696 7840 10724
rect 5368 10656 5396 10696
rect 7834 10684 7840 10696
rect 7892 10684 7898 10736
rect 12066 10724 12072 10736
rect 9232 10696 12072 10724
rect 3559 10628 4016 10656
rect 5276 10628 5396 10656
rect 3559 10625 3571 10628
rect 3513 10619 3571 10625
rect 5276 10588 5304 10628
rect 5534 10616 5540 10668
rect 5592 10616 5598 10668
rect 5994 10656 6000 10668
rect 5955 10628 6000 10656
rect 5994 10616 6000 10628
rect 6052 10616 6058 10668
rect 7101 10659 7159 10665
rect 7101 10625 7113 10659
rect 7147 10656 7159 10659
rect 7742 10656 7748 10668
rect 7147 10628 7748 10656
rect 7147 10625 7159 10628
rect 7101 10619 7159 10625
rect 7742 10616 7748 10628
rect 7800 10616 7806 10668
rect 9122 10656 9128 10668
rect 9083 10628 9128 10656
rect 9122 10616 9128 10628
rect 9180 10616 9186 10668
rect 3436 10560 5304 10588
rect 5353 10591 5411 10597
rect 5353 10557 5365 10591
rect 5399 10588 5411 10591
rect 5552 10588 5580 10616
rect 9232 10600 9260 10696
rect 12066 10684 12072 10696
rect 12124 10684 12130 10736
rect 12820 10724 12848 10764
rect 12986 10752 12992 10764
rect 13044 10752 13050 10804
rect 13906 10752 13912 10804
rect 13964 10792 13970 10804
rect 14182 10792 14188 10804
rect 13964 10764 14188 10792
rect 13964 10752 13970 10764
rect 14182 10752 14188 10764
rect 14240 10752 14246 10804
rect 12176 10696 12848 10724
rect 9769 10659 9827 10665
rect 9769 10625 9781 10659
rect 9815 10656 9827 10659
rect 10226 10656 10232 10668
rect 9815 10628 10232 10656
rect 9815 10625 9827 10628
rect 9769 10619 9827 10625
rect 10226 10616 10232 10628
rect 10284 10656 10290 10668
rect 10321 10659 10379 10665
rect 10321 10656 10333 10659
rect 10284 10628 10333 10656
rect 10284 10616 10290 10628
rect 10321 10625 10333 10628
rect 10367 10625 10379 10659
rect 10502 10656 10508 10668
rect 10463 10628 10508 10656
rect 10321 10619 10379 10625
rect 10502 10616 10508 10628
rect 10560 10656 10566 10668
rect 11241 10659 11299 10665
rect 11241 10656 11253 10659
rect 10560 10628 11253 10656
rect 10560 10616 10566 10628
rect 11241 10625 11253 10628
rect 11287 10625 11299 10659
rect 11241 10619 11299 10625
rect 11790 10616 11796 10668
rect 11848 10656 11854 10668
rect 12176 10656 12204 10696
rect 11848 10628 12204 10656
rect 11848 10616 11854 10628
rect 12250 10616 12256 10668
rect 12308 10656 12314 10668
rect 12820 10665 12848 10696
rect 12805 10659 12863 10665
rect 12308 10628 12353 10656
rect 12308 10616 12314 10628
rect 12805 10625 12817 10659
rect 12851 10625 12863 10659
rect 12805 10619 12863 10625
rect 7285 10591 7343 10597
rect 5399 10560 5580 10588
rect 5736 10560 7236 10588
rect 5399 10557 5411 10560
rect 5353 10551 5411 10557
rect 3237 10523 3295 10529
rect 3237 10489 3249 10523
rect 3283 10520 3295 10523
rect 3697 10523 3755 10529
rect 3697 10520 3709 10523
rect 3283 10492 3709 10520
rect 3283 10489 3295 10492
rect 3237 10483 3295 10489
rect 3697 10489 3709 10492
rect 3743 10520 3755 10523
rect 3878 10520 3884 10532
rect 3743 10492 3884 10520
rect 3743 10489 3755 10492
rect 3697 10483 3755 10489
rect 3878 10480 3884 10492
rect 3936 10480 3942 10532
rect 5108 10523 5166 10529
rect 5108 10489 5120 10523
rect 5154 10520 5166 10523
rect 5534 10520 5540 10532
rect 5154 10492 5540 10520
rect 5154 10489 5166 10492
rect 5108 10483 5166 10489
rect 5534 10480 5540 10492
rect 5592 10480 5598 10532
rect 2501 10455 2559 10461
rect 2501 10421 2513 10455
rect 2547 10452 2559 10455
rect 2869 10455 2927 10461
rect 2869 10452 2881 10455
rect 2547 10424 2881 10452
rect 2547 10421 2559 10424
rect 2501 10415 2559 10421
rect 2869 10421 2881 10424
rect 2915 10421 2927 10455
rect 3326 10452 3332 10464
rect 3287 10424 3332 10452
rect 2869 10415 2927 10421
rect 3326 10412 3332 10424
rect 3384 10412 3390 10464
rect 4890 10412 4896 10464
rect 4948 10452 4954 10464
rect 5736 10452 5764 10560
rect 5905 10523 5963 10529
rect 5905 10489 5917 10523
rect 5951 10520 5963 10523
rect 6638 10520 6644 10532
rect 5951 10492 6644 10520
rect 5951 10489 5963 10492
rect 5905 10483 5963 10489
rect 6638 10480 6644 10492
rect 6696 10480 6702 10532
rect 7208 10520 7236 10560
rect 7285 10557 7297 10591
rect 7331 10588 7343 10591
rect 7926 10588 7932 10600
rect 7331 10560 7932 10588
rect 7331 10557 7343 10560
rect 7285 10551 7343 10557
rect 7926 10548 7932 10560
rect 7984 10548 7990 10600
rect 8570 10548 8576 10600
rect 8628 10588 8634 10600
rect 8858 10591 8916 10597
rect 8858 10588 8870 10591
rect 8628 10560 8870 10588
rect 8628 10548 8634 10560
rect 8858 10557 8870 10560
rect 8904 10557 8916 10591
rect 9214 10588 9220 10600
rect 9175 10560 9220 10588
rect 8858 10551 8916 10557
rect 9214 10548 9220 10560
rect 9272 10548 9278 10600
rect 9493 10591 9551 10597
rect 9493 10557 9505 10591
rect 9539 10588 9551 10591
rect 9585 10591 9643 10597
rect 9585 10588 9597 10591
rect 9539 10560 9597 10588
rect 9539 10557 9551 10560
rect 9493 10551 9551 10557
rect 9585 10557 9597 10560
rect 9631 10588 9643 10591
rect 11054 10588 11060 10600
rect 9631 10560 11060 10588
rect 9631 10557 9643 10560
rect 9585 10551 9643 10557
rect 11054 10548 11060 10560
rect 11112 10548 11118 10600
rect 11149 10523 11207 10529
rect 11149 10520 11161 10523
rect 7208 10492 11161 10520
rect 11149 10489 11161 10492
rect 11195 10520 11207 10523
rect 11422 10520 11428 10532
rect 11195 10492 11428 10520
rect 11195 10489 11207 10492
rect 11149 10483 11207 10489
rect 11422 10480 11428 10492
rect 11480 10480 11486 10532
rect 12069 10523 12127 10529
rect 12069 10489 12081 10523
rect 12115 10520 12127 10523
rect 12894 10520 12900 10532
rect 12115 10492 12900 10520
rect 12115 10489 12127 10492
rect 12069 10483 12127 10489
rect 12894 10480 12900 10492
rect 12952 10480 12958 10532
rect 13072 10523 13130 10529
rect 13072 10489 13084 10523
rect 13118 10520 13130 10523
rect 13354 10520 13360 10532
rect 13118 10492 13360 10520
rect 13118 10489 13130 10492
rect 13072 10483 13130 10489
rect 13354 10480 13360 10492
rect 13412 10480 13418 10532
rect 4948 10424 5764 10452
rect 4948 10412 4954 10424
rect 5810 10412 5816 10464
rect 5868 10452 5874 10464
rect 6546 10452 6552 10464
rect 5868 10424 6552 10452
rect 5868 10412 5874 10424
rect 6546 10412 6552 10424
rect 6604 10412 6610 10464
rect 7190 10452 7196 10464
rect 7151 10424 7196 10452
rect 7190 10412 7196 10424
rect 7248 10412 7254 10464
rect 7742 10452 7748 10464
rect 7703 10424 7748 10452
rect 7742 10412 7748 10424
rect 7800 10412 7806 10464
rect 8386 10412 8392 10464
rect 8444 10452 8450 10464
rect 9122 10452 9128 10464
rect 8444 10424 9128 10452
rect 8444 10412 8450 10424
rect 9122 10412 9128 10424
rect 9180 10452 9186 10464
rect 9585 10455 9643 10461
rect 9585 10452 9597 10455
rect 9180 10424 9597 10452
rect 9180 10412 9186 10424
rect 9585 10421 9597 10424
rect 9631 10421 9643 10455
rect 9858 10452 9864 10464
rect 9819 10424 9864 10452
rect 9585 10415 9643 10421
rect 9858 10412 9864 10424
rect 9916 10412 9922 10464
rect 10042 10412 10048 10464
rect 10100 10452 10106 10464
rect 10229 10455 10287 10461
rect 10229 10452 10241 10455
rect 10100 10424 10241 10452
rect 10100 10412 10106 10424
rect 10229 10421 10241 10424
rect 10275 10421 10287 10455
rect 10229 10415 10287 10421
rect 10778 10412 10784 10464
rect 10836 10452 10842 10464
rect 11057 10455 11115 10461
rect 11057 10452 11069 10455
rect 10836 10424 11069 10452
rect 10836 10412 10842 10424
rect 11057 10421 11069 10424
rect 11103 10421 11115 10455
rect 11057 10415 11115 10421
rect 11330 10412 11336 10464
rect 11388 10452 11394 10464
rect 11701 10455 11759 10461
rect 11701 10452 11713 10455
rect 11388 10424 11713 10452
rect 11388 10412 11394 10424
rect 11701 10421 11713 10424
rect 11747 10421 11759 10455
rect 11701 10415 11759 10421
rect 12161 10455 12219 10461
rect 12161 10421 12173 10455
rect 12207 10452 12219 10455
rect 12434 10452 12440 10464
rect 12207 10424 12440 10452
rect 12207 10421 12219 10424
rect 12161 10415 12219 10421
rect 12434 10412 12440 10424
rect 12492 10412 12498 10464
rect 12621 10455 12679 10461
rect 12621 10421 12633 10455
rect 12667 10452 12679 10455
rect 13170 10452 13176 10464
rect 12667 10424 13176 10452
rect 12667 10421 12679 10424
rect 12621 10415 12679 10421
rect 13170 10412 13176 10424
rect 13228 10412 13234 10464
rect 14458 10452 14464 10464
rect 14419 10424 14464 10452
rect 14458 10412 14464 10424
rect 14516 10412 14522 10464
rect 14645 10455 14703 10461
rect 14645 10421 14657 10455
rect 14691 10452 14703 10455
rect 15102 10452 15108 10464
rect 14691 10424 15108 10452
rect 14691 10421 14703 10424
rect 14645 10415 14703 10421
rect 15102 10412 15108 10424
rect 15160 10412 15166 10464
rect 1104 10362 16008 10384
rect 1104 10310 5979 10362
rect 6031 10310 6043 10362
rect 6095 10310 6107 10362
rect 6159 10310 6171 10362
rect 6223 10310 10976 10362
rect 11028 10310 11040 10362
rect 11092 10310 11104 10362
rect 11156 10310 11168 10362
rect 11220 10310 16008 10362
rect 1104 10288 16008 10310
rect 1765 10251 1823 10257
rect 1765 10248 1777 10251
rect 1596 10220 1777 10248
rect 1596 10189 1624 10220
rect 1765 10217 1777 10220
rect 1811 10217 1823 10251
rect 1765 10211 1823 10217
rect 3326 10208 3332 10260
rect 3384 10248 3390 10260
rect 3881 10251 3939 10257
rect 3881 10248 3893 10251
rect 3384 10220 3893 10248
rect 3384 10208 3390 10220
rect 3881 10217 3893 10220
rect 3927 10217 3939 10251
rect 3881 10211 3939 10217
rect 5445 10251 5503 10257
rect 5445 10217 5457 10251
rect 5491 10248 5503 10251
rect 5718 10248 5724 10260
rect 5491 10220 5724 10248
rect 5491 10217 5503 10220
rect 5445 10211 5503 10217
rect 5718 10208 5724 10220
rect 5776 10208 5782 10260
rect 7190 10208 7196 10260
rect 7248 10248 7254 10260
rect 7929 10251 7987 10257
rect 7929 10248 7941 10251
rect 7248 10220 7941 10248
rect 7248 10208 7254 10220
rect 7929 10217 7941 10220
rect 7975 10217 7987 10251
rect 7929 10211 7987 10217
rect 8386 10208 8392 10260
rect 8444 10248 8450 10260
rect 8757 10251 8815 10257
rect 8444 10220 8489 10248
rect 8444 10208 8450 10220
rect 8757 10217 8769 10251
rect 8803 10248 8815 10251
rect 8846 10248 8852 10260
rect 8803 10220 8852 10248
rect 8803 10217 8815 10220
rect 8757 10211 8815 10217
rect 8846 10208 8852 10220
rect 8904 10208 8910 10260
rect 9493 10251 9551 10257
rect 9493 10217 9505 10251
rect 9539 10248 9551 10251
rect 9858 10248 9864 10260
rect 9539 10220 9864 10248
rect 9539 10217 9551 10220
rect 9493 10211 9551 10217
rect 9858 10208 9864 10220
rect 9916 10208 9922 10260
rect 11330 10248 11336 10260
rect 9968 10220 11336 10248
rect 1581 10183 1639 10189
rect 1581 10149 1593 10183
rect 1627 10149 1639 10183
rect 9968 10180 9996 10220
rect 11330 10208 11336 10220
rect 11388 10208 11394 10260
rect 11422 10208 11428 10260
rect 11480 10248 11486 10260
rect 13170 10248 13176 10260
rect 11480 10220 13176 10248
rect 11480 10208 11486 10220
rect 13170 10208 13176 10220
rect 13228 10208 13234 10260
rect 14458 10208 14464 10260
rect 14516 10248 14522 10260
rect 14737 10251 14795 10257
rect 14737 10248 14749 10251
rect 14516 10220 14749 10248
rect 14516 10208 14522 10220
rect 14737 10217 14749 10220
rect 14783 10217 14795 10251
rect 14737 10211 14795 10217
rect 15010 10208 15016 10260
rect 15068 10248 15074 10260
rect 15197 10251 15255 10257
rect 15197 10248 15209 10251
rect 15068 10220 15209 10248
rect 15068 10208 15074 10220
rect 15197 10217 15209 10220
rect 15243 10217 15255 10251
rect 15197 10211 15255 10217
rect 1581 10143 1639 10149
rect 2746 10152 9996 10180
rect 1949 10115 2007 10121
rect 1949 10081 1961 10115
rect 1995 10112 2007 10115
rect 2746 10112 2774 10152
rect 10502 10140 10508 10192
rect 10560 10180 10566 10192
rect 11158 10183 11216 10189
rect 11158 10180 11170 10183
rect 10560 10152 11170 10180
rect 10560 10140 10566 10152
rect 11158 10149 11170 10152
rect 11204 10180 11216 10183
rect 11204 10152 11376 10180
rect 11204 10149 11216 10152
rect 11158 10143 11216 10149
rect 1995 10084 2774 10112
rect 4249 10115 4307 10121
rect 1995 10081 2007 10084
rect 1949 10075 2007 10081
rect 4249 10081 4261 10115
rect 4295 10081 4307 10115
rect 4249 10075 4307 10081
rect 1394 9976 1400 9988
rect 1355 9948 1400 9976
rect 1394 9936 1400 9948
rect 1452 9936 1458 9988
rect 4264 9908 4292 10075
rect 5626 10072 5632 10124
rect 5684 10112 5690 10124
rect 5813 10115 5871 10121
rect 5813 10112 5825 10115
rect 5684 10084 5825 10112
rect 5684 10072 5690 10084
rect 5813 10081 5825 10084
rect 5859 10081 5871 10115
rect 5813 10075 5871 10081
rect 6080 10115 6138 10121
rect 6080 10081 6092 10115
rect 6126 10112 6138 10115
rect 7742 10112 7748 10124
rect 6126 10084 7748 10112
rect 6126 10081 6138 10084
rect 6080 10075 6138 10081
rect 7742 10072 7748 10084
rect 7800 10072 7806 10124
rect 8297 10115 8355 10121
rect 8297 10081 8309 10115
rect 8343 10112 8355 10115
rect 9214 10112 9220 10124
rect 8343 10084 9220 10112
rect 8343 10081 8355 10084
rect 8297 10075 8355 10081
rect 9214 10072 9220 10084
rect 9272 10072 9278 10124
rect 9585 10115 9643 10121
rect 9585 10081 9597 10115
rect 9631 10112 9643 10115
rect 9950 10112 9956 10124
rect 9631 10084 9956 10112
rect 9631 10081 9643 10084
rect 9585 10075 9643 10081
rect 9950 10072 9956 10084
rect 10008 10072 10014 10124
rect 4341 10047 4399 10053
rect 4341 10013 4353 10047
rect 4387 10013 4399 10047
rect 4341 10007 4399 10013
rect 4525 10047 4583 10053
rect 4525 10013 4537 10047
rect 4571 10044 4583 10047
rect 5534 10044 5540 10056
rect 4571 10016 5540 10044
rect 4571 10013 4583 10016
rect 4525 10007 4583 10013
rect 4356 9976 4384 10007
rect 5534 10004 5540 10016
rect 5592 10004 5598 10056
rect 8570 10044 8576 10056
rect 8483 10016 8576 10044
rect 8570 10004 8576 10016
rect 8628 10044 8634 10056
rect 8938 10044 8944 10056
rect 8628 10016 8944 10044
rect 8628 10004 8634 10016
rect 8938 10004 8944 10016
rect 8996 10044 9002 10056
rect 9401 10047 9459 10053
rect 9401 10044 9413 10047
rect 8996 10016 9413 10044
rect 8996 10004 9002 10016
rect 9401 10013 9413 10016
rect 9447 10044 9459 10047
rect 11348 10044 11376 10152
rect 11606 10140 11612 10192
rect 11664 10180 11670 10192
rect 12250 10180 12256 10192
rect 11664 10152 12256 10180
rect 11664 10140 11670 10152
rect 12250 10140 12256 10152
rect 12308 10180 12314 10192
rect 12630 10183 12688 10189
rect 12630 10180 12642 10183
rect 12308 10152 12642 10180
rect 12308 10140 12314 10152
rect 12630 10149 12642 10152
rect 12676 10149 12688 10183
rect 12630 10143 12688 10149
rect 13446 10140 13452 10192
rect 13504 10180 13510 10192
rect 13633 10183 13691 10189
rect 13633 10180 13645 10183
rect 13504 10152 13645 10180
rect 13504 10140 13510 10152
rect 13633 10149 13645 10152
rect 13679 10180 13691 10183
rect 15028 10180 15056 10208
rect 13679 10152 15056 10180
rect 13679 10149 13691 10152
rect 13633 10143 13691 10149
rect 15286 10140 15292 10192
rect 15344 10180 15350 10192
rect 15473 10183 15531 10189
rect 15473 10180 15485 10183
rect 15344 10152 15485 10180
rect 15344 10140 15350 10152
rect 15473 10149 15485 10152
rect 15519 10149 15531 10183
rect 15473 10143 15531 10149
rect 11425 10115 11483 10121
rect 11425 10081 11437 10115
rect 11471 10112 11483 10115
rect 11790 10112 11796 10124
rect 11471 10084 11796 10112
rect 11471 10081 11483 10084
rect 11425 10075 11483 10081
rect 11790 10072 11796 10084
rect 11848 10112 11854 10124
rect 12897 10115 12955 10121
rect 12897 10112 12909 10115
rect 11848 10084 12909 10112
rect 11848 10072 11854 10084
rect 12897 10081 12909 10084
rect 12943 10081 12955 10115
rect 12897 10075 12955 10081
rect 13725 10115 13783 10121
rect 13725 10081 13737 10115
rect 13771 10112 13783 10115
rect 15102 10112 15108 10124
rect 13771 10084 15108 10112
rect 13771 10081 13783 10084
rect 13725 10075 13783 10081
rect 15102 10072 15108 10084
rect 15160 10072 15166 10124
rect 9447 10016 9674 10044
rect 11348 10016 11560 10044
rect 9447 10013 9459 10016
rect 9401 10007 9459 10013
rect 4801 9979 4859 9985
rect 4801 9976 4813 9979
rect 4356 9948 4813 9976
rect 4801 9945 4813 9948
rect 4847 9976 4859 9979
rect 5810 9976 5816 9988
rect 4847 9948 5816 9976
rect 4847 9945 4859 9948
rect 4801 9939 4859 9945
rect 5810 9936 5816 9948
rect 5868 9936 5874 9988
rect 7193 9979 7251 9985
rect 7193 9945 7205 9979
rect 7239 9976 7251 9979
rect 7282 9976 7288 9988
rect 7239 9948 7288 9976
rect 7239 9945 7251 9948
rect 7193 9939 7251 9945
rect 7282 9936 7288 9948
rect 7340 9976 7346 9988
rect 7558 9976 7564 9988
rect 7340 9948 7564 9976
rect 7340 9936 7346 9948
rect 7558 9936 7564 9948
rect 7616 9936 7622 9988
rect 4985 9911 5043 9917
rect 4985 9908 4997 9911
rect 4264 9880 4997 9908
rect 4985 9877 4997 9880
rect 5031 9908 5043 9911
rect 6914 9908 6920 9920
rect 5031 9880 6920 9908
rect 5031 9877 5043 9880
rect 4985 9871 5043 9877
rect 6914 9868 6920 9880
rect 6972 9868 6978 9920
rect 9646 9908 9674 10016
rect 9953 9979 10011 9985
rect 9953 9945 9965 9979
rect 9999 9976 10011 9979
rect 10410 9976 10416 9988
rect 9999 9948 10416 9976
rect 9999 9945 10011 9948
rect 9953 9939 10011 9945
rect 10410 9936 10416 9948
rect 10468 9936 10474 9988
rect 11532 9985 11560 10016
rect 13354 10004 13360 10056
rect 13412 10044 13418 10056
rect 13449 10047 13507 10053
rect 13449 10044 13461 10047
rect 13412 10016 13461 10044
rect 13412 10004 13418 10016
rect 13449 10013 13461 10016
rect 13495 10013 13507 10047
rect 13449 10007 13507 10013
rect 11517 9979 11575 9985
rect 11517 9945 11529 9979
rect 11563 9945 11575 9979
rect 13262 9976 13268 9988
rect 11517 9939 11575 9945
rect 12912 9948 13268 9976
rect 10045 9911 10103 9917
rect 10045 9908 10057 9911
rect 9646 9880 10057 9908
rect 10045 9877 10057 9880
rect 10091 9877 10103 9911
rect 10045 9871 10103 9877
rect 12250 9868 12256 9920
rect 12308 9908 12314 9920
rect 12912 9908 12940 9948
rect 13262 9936 13268 9948
rect 13320 9936 13326 9988
rect 13464 9976 13492 10007
rect 13814 10004 13820 10056
rect 13872 10044 13878 10056
rect 14829 10047 14887 10053
rect 14829 10044 14841 10047
rect 13872 10016 14841 10044
rect 13872 10004 13878 10016
rect 14829 10013 14841 10016
rect 14875 10013 14887 10047
rect 14829 10007 14887 10013
rect 14921 10047 14979 10053
rect 14921 10013 14933 10047
rect 14967 10013 14979 10047
rect 14921 10007 14979 10013
rect 14936 9976 14964 10007
rect 15654 9976 15660 9988
rect 13464 9948 14964 9976
rect 15615 9948 15660 9976
rect 15654 9936 15660 9948
rect 15712 9936 15718 9988
rect 12308 9880 12940 9908
rect 12308 9868 12314 9880
rect 12986 9868 12992 9920
rect 13044 9908 13050 9920
rect 14090 9908 14096 9920
rect 13044 9880 13089 9908
rect 14051 9880 14096 9908
rect 13044 9868 13050 9880
rect 14090 9868 14096 9880
rect 14148 9868 14154 9920
rect 14182 9868 14188 9920
rect 14240 9908 14246 9920
rect 14369 9911 14427 9917
rect 14369 9908 14381 9911
rect 14240 9880 14381 9908
rect 14240 9868 14246 9880
rect 14369 9877 14381 9880
rect 14415 9877 14427 9911
rect 14369 9871 14427 9877
rect 1104 9818 16008 9840
rect 1104 9766 3480 9818
rect 3532 9766 3544 9818
rect 3596 9766 3608 9818
rect 3660 9766 3672 9818
rect 3724 9766 8478 9818
rect 8530 9766 8542 9818
rect 8594 9766 8606 9818
rect 8658 9766 8670 9818
rect 8722 9766 13475 9818
rect 13527 9766 13539 9818
rect 13591 9766 13603 9818
rect 13655 9766 13667 9818
rect 13719 9766 16008 9818
rect 1104 9744 16008 9766
rect 3878 9664 3884 9716
rect 3936 9704 3942 9716
rect 3936 9676 5488 9704
rect 3936 9664 3942 9676
rect 5460 9636 5488 9676
rect 5534 9664 5540 9716
rect 5592 9704 5598 9716
rect 6457 9707 6515 9713
rect 6457 9704 6469 9707
rect 5592 9676 6469 9704
rect 5592 9664 5598 9676
rect 6457 9673 6469 9676
rect 6503 9673 6515 9707
rect 7190 9704 7196 9716
rect 6457 9667 6515 9673
rect 6564 9676 7196 9704
rect 6564 9636 6592 9676
rect 7190 9664 7196 9676
rect 7248 9664 7254 9716
rect 9306 9664 9312 9716
rect 9364 9704 9370 9716
rect 13814 9704 13820 9716
rect 9364 9676 13820 9704
rect 9364 9664 9370 9676
rect 13814 9664 13820 9676
rect 13872 9664 13878 9716
rect 5460 9608 6592 9636
rect 8294 9596 8300 9648
rect 8352 9636 8358 9648
rect 8481 9639 8539 9645
rect 8481 9636 8493 9639
rect 8352 9608 8493 9636
rect 8352 9596 8358 9608
rect 8481 9605 8493 9608
rect 8527 9636 8539 9639
rect 9030 9636 9036 9648
rect 8527 9608 9036 9636
rect 8527 9605 8539 9608
rect 8481 9599 8539 9605
rect 9030 9596 9036 9608
rect 9088 9596 9094 9648
rect 9950 9636 9956 9648
rect 9911 9608 9956 9636
rect 9950 9596 9956 9608
rect 10008 9596 10014 9648
rect 10778 9636 10784 9648
rect 10336 9608 10784 9636
rect 4154 9528 4160 9580
rect 4212 9568 4218 9580
rect 4249 9571 4307 9577
rect 4249 9568 4261 9571
rect 4212 9540 4261 9568
rect 4212 9528 4218 9540
rect 4249 9537 4261 9540
rect 4295 9537 4307 9571
rect 5166 9568 5172 9580
rect 5127 9540 5172 9568
rect 4249 9531 4307 9537
rect 5166 9528 5172 9540
rect 5224 9568 5230 9580
rect 5905 9571 5963 9577
rect 5905 9568 5917 9571
rect 5224 9540 5917 9568
rect 5224 9528 5230 9540
rect 5905 9537 5917 9540
rect 5951 9537 5963 9571
rect 5905 9531 5963 9537
rect 5994 9528 6000 9580
rect 6052 9568 6058 9580
rect 6454 9568 6460 9580
rect 6052 9540 6460 9568
rect 6052 9528 6058 9540
rect 6454 9528 6460 9540
rect 6512 9528 6518 9580
rect 10336 9568 10364 9608
rect 10778 9596 10784 9608
rect 10836 9596 10842 9648
rect 12434 9596 12440 9648
rect 12492 9636 12498 9648
rect 12989 9639 13047 9645
rect 12989 9636 13001 9639
rect 12492 9608 13001 9636
rect 12492 9596 12498 9608
rect 12989 9605 13001 9608
rect 13035 9605 13047 9639
rect 12989 9599 13047 9605
rect 13924 9608 14412 9636
rect 13924 9580 13952 9608
rect 10502 9568 10508 9580
rect 7760 9540 10364 9568
rect 10463 9540 10508 9568
rect 4985 9503 5043 9509
rect 4985 9469 4997 9503
rect 5031 9500 5043 9503
rect 5350 9500 5356 9512
rect 5031 9472 5356 9500
rect 5031 9469 5043 9472
rect 4985 9463 5043 9469
rect 5350 9460 5356 9472
rect 5408 9500 5414 9512
rect 5813 9503 5871 9509
rect 5408 9472 5764 9500
rect 5408 9460 5414 9472
rect 4065 9435 4123 9441
rect 4065 9401 4077 9435
rect 4111 9432 4123 9435
rect 5736 9432 5764 9472
rect 5813 9469 5825 9503
rect 5859 9500 5871 9503
rect 6270 9500 6276 9512
rect 5859 9472 6276 9500
rect 5859 9469 5871 9472
rect 5813 9463 5871 9469
rect 6270 9460 6276 9472
rect 6328 9500 6334 9512
rect 6730 9500 6736 9512
rect 6328 9472 6736 9500
rect 6328 9460 6334 9472
rect 6730 9460 6736 9472
rect 6788 9460 6794 9512
rect 7760 9500 7788 9540
rect 10502 9528 10508 9540
rect 10560 9528 10566 9580
rect 12345 9571 12403 9577
rect 12345 9537 12357 9571
rect 12391 9568 12403 9571
rect 13262 9568 13268 9580
rect 12391 9540 13268 9568
rect 12391 9537 12403 9540
rect 12345 9531 12403 9537
rect 13262 9528 13268 9540
rect 13320 9528 13326 9580
rect 13633 9571 13691 9577
rect 13633 9537 13645 9571
rect 13679 9568 13691 9571
rect 13906 9568 13912 9580
rect 13679 9540 13912 9568
rect 13679 9537 13691 9540
rect 13633 9531 13691 9537
rect 13906 9528 13912 9540
rect 13964 9528 13970 9580
rect 14090 9528 14096 9580
rect 14148 9568 14154 9580
rect 14384 9577 14412 9608
rect 14277 9571 14335 9577
rect 14277 9568 14289 9571
rect 14148 9540 14289 9568
rect 14148 9528 14154 9540
rect 14277 9537 14289 9540
rect 14323 9537 14335 9571
rect 14277 9531 14335 9537
rect 14369 9571 14427 9577
rect 14369 9537 14381 9571
rect 14415 9537 14427 9571
rect 14369 9531 14427 9537
rect 7484 9472 7788 9500
rect 7837 9503 7895 9509
rect 7484 9432 7512 9472
rect 7837 9469 7849 9503
rect 7883 9500 7895 9503
rect 9674 9500 9680 9512
rect 7883 9472 9680 9500
rect 7883 9469 7895 9472
rect 7837 9463 7895 9469
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 9769 9503 9827 9509
rect 9769 9469 9781 9503
rect 9815 9500 9827 9503
rect 12802 9500 12808 9512
rect 9815 9472 12808 9500
rect 9815 9469 9827 9472
rect 9769 9463 9827 9469
rect 12802 9460 12808 9472
rect 12860 9460 12866 9512
rect 12894 9460 12900 9512
rect 12952 9500 12958 9512
rect 14182 9500 14188 9512
rect 12952 9472 13492 9500
rect 14143 9472 14188 9500
rect 12952 9460 12958 9472
rect 4111 9404 5396 9432
rect 5736 9404 7512 9432
rect 4111 9401 4123 9404
rect 4065 9395 4123 9401
rect 3326 9324 3332 9376
rect 3384 9364 3390 9376
rect 3697 9367 3755 9373
rect 3697 9364 3709 9367
rect 3384 9336 3709 9364
rect 3384 9324 3390 9336
rect 3697 9333 3709 9336
rect 3743 9333 3755 9367
rect 3697 9327 3755 9333
rect 4157 9367 4215 9373
rect 4157 9333 4169 9367
rect 4203 9364 4215 9367
rect 4525 9367 4583 9373
rect 4525 9364 4537 9367
rect 4203 9336 4537 9364
rect 4203 9333 4215 9336
rect 4157 9327 4215 9333
rect 4525 9333 4537 9336
rect 4571 9333 4583 9367
rect 4525 9327 4583 9333
rect 4893 9367 4951 9373
rect 4893 9333 4905 9367
rect 4939 9364 4951 9367
rect 4982 9364 4988 9376
rect 4939 9336 4988 9364
rect 4939 9333 4951 9336
rect 4893 9327 4951 9333
rect 4982 9324 4988 9336
rect 5040 9324 5046 9376
rect 5368 9373 5396 9404
rect 7558 9392 7564 9444
rect 7616 9441 7622 9444
rect 7616 9432 7628 9441
rect 7616 9404 7661 9432
rect 7616 9395 7628 9404
rect 7616 9392 7622 9395
rect 9490 9392 9496 9444
rect 9548 9432 9554 9444
rect 10778 9432 10784 9444
rect 9548 9404 10784 9432
rect 9548 9392 9554 9404
rect 10778 9392 10784 9404
rect 10836 9392 10842 9444
rect 12529 9435 12587 9441
rect 12529 9401 12541 9435
rect 12575 9432 12587 9435
rect 13357 9435 13415 9441
rect 13357 9432 13369 9435
rect 12575 9404 12848 9432
rect 12575 9401 12587 9404
rect 12529 9395 12587 9401
rect 12820 9376 12848 9404
rect 12912 9404 13369 9432
rect 5353 9367 5411 9373
rect 5353 9333 5365 9367
rect 5399 9333 5411 9367
rect 5718 9364 5724 9376
rect 5679 9336 5724 9364
rect 5353 9327 5411 9333
rect 5718 9324 5724 9336
rect 5776 9324 5782 9376
rect 5810 9324 5816 9376
rect 5868 9364 5874 9376
rect 6181 9367 6239 9373
rect 6181 9364 6193 9367
rect 5868 9336 6193 9364
rect 5868 9324 5874 9336
rect 6181 9333 6193 9336
rect 6227 9333 6239 9367
rect 6181 9327 6239 9333
rect 7190 9324 7196 9376
rect 7248 9364 7254 9376
rect 7466 9364 7472 9376
rect 7248 9336 7472 9364
rect 7248 9324 7254 9336
rect 7466 9324 7472 9336
rect 7524 9364 7530 9376
rect 9950 9364 9956 9376
rect 7524 9336 9956 9364
rect 7524 9324 7530 9336
rect 9950 9324 9956 9336
rect 10008 9324 10014 9376
rect 10318 9364 10324 9376
rect 10279 9336 10324 9364
rect 10318 9324 10324 9336
rect 10376 9324 10382 9376
rect 10413 9367 10471 9373
rect 10413 9333 10425 9367
rect 10459 9364 10471 9367
rect 10686 9364 10692 9376
rect 10459 9336 10692 9364
rect 10459 9333 10471 9336
rect 10413 9327 10471 9333
rect 10686 9324 10692 9336
rect 10744 9364 10750 9376
rect 10965 9367 11023 9373
rect 10965 9364 10977 9367
rect 10744 9336 10977 9364
rect 10744 9324 10750 9336
rect 10965 9333 10977 9336
rect 11011 9333 11023 9367
rect 10965 9327 11023 9333
rect 11241 9367 11299 9373
rect 11241 9333 11253 9367
rect 11287 9364 11299 9367
rect 11606 9364 11612 9376
rect 11287 9336 11612 9364
rect 11287 9333 11299 9336
rect 11241 9327 11299 9333
rect 11606 9324 11612 9336
rect 11664 9324 11670 9376
rect 12434 9324 12440 9376
rect 12492 9364 12498 9376
rect 12492 9336 12537 9364
rect 12492 9324 12498 9336
rect 12802 9324 12808 9376
rect 12860 9324 12866 9376
rect 12912 9373 12940 9404
rect 13357 9401 13369 9404
rect 13403 9401 13415 9435
rect 13464 9432 13492 9472
rect 14182 9460 14188 9472
rect 14240 9460 14246 9512
rect 13464 9404 13860 9432
rect 13357 9395 13415 9401
rect 12897 9367 12955 9373
rect 12897 9333 12909 9367
rect 12943 9333 12955 9367
rect 13446 9364 13452 9376
rect 13407 9336 13452 9364
rect 12897 9327 12955 9333
rect 13446 9324 13452 9336
rect 13504 9324 13510 9376
rect 13832 9373 13860 9404
rect 13817 9367 13875 9373
rect 13817 9333 13829 9367
rect 13863 9333 13875 9367
rect 13817 9327 13875 9333
rect 1104 9274 16008 9296
rect 1104 9222 5979 9274
rect 6031 9222 6043 9274
rect 6095 9222 6107 9274
rect 6159 9222 6171 9274
rect 6223 9222 10976 9274
rect 11028 9222 11040 9274
rect 11092 9222 11104 9274
rect 11156 9222 11168 9274
rect 11220 9222 16008 9274
rect 1104 9200 16008 9222
rect 3326 9160 3332 9172
rect 3287 9132 3332 9160
rect 3326 9120 3332 9132
rect 3384 9120 3390 9172
rect 5261 9163 5319 9169
rect 5261 9160 5273 9163
rect 3620 9132 5273 9160
rect 1394 9092 1400 9104
rect 1355 9064 1400 9092
rect 1394 9052 1400 9064
rect 1452 9052 1458 9104
rect 1578 9024 1584 9036
rect 1539 8996 1584 9024
rect 1578 8984 1584 8996
rect 1636 8984 1642 9036
rect 3620 8965 3648 9132
rect 5261 9129 5273 9132
rect 5307 9129 5319 9163
rect 5261 9123 5319 9129
rect 5276 9092 5304 9123
rect 6914 9120 6920 9172
rect 6972 9160 6978 9172
rect 7193 9163 7251 9169
rect 7193 9160 7205 9163
rect 6972 9132 7205 9160
rect 6972 9120 6978 9132
rect 7193 9129 7205 9132
rect 7239 9160 7251 9163
rect 8754 9160 8760 9172
rect 7239 9132 8760 9160
rect 7239 9129 7251 9132
rect 7193 9123 7251 9129
rect 8754 9120 8760 9132
rect 8812 9120 8818 9172
rect 9490 9160 9496 9172
rect 9451 9132 9496 9160
rect 9490 9120 9496 9132
rect 9548 9120 9554 9172
rect 9766 9120 9772 9172
rect 9824 9160 9830 9172
rect 9953 9163 10011 9169
rect 9953 9160 9965 9163
rect 9824 9132 9965 9160
rect 9824 9120 9830 9132
rect 9953 9129 9965 9132
rect 9999 9129 10011 9163
rect 9953 9123 10011 9129
rect 10134 9120 10140 9172
rect 10192 9160 10198 9172
rect 10321 9163 10379 9169
rect 10321 9160 10333 9163
rect 10192 9132 10333 9160
rect 10192 9120 10198 9132
rect 10321 9129 10333 9132
rect 10367 9129 10379 9163
rect 10321 9123 10379 9129
rect 10410 9120 10416 9172
rect 10468 9160 10474 9172
rect 12802 9160 12808 9172
rect 10468 9132 10513 9160
rect 10704 9132 12808 9160
rect 10468 9120 10474 9132
rect 5598 9095 5656 9101
rect 5598 9092 5610 9095
rect 5276 9064 5610 9092
rect 5598 9061 5610 9064
rect 5644 9061 5656 9095
rect 5598 9055 5656 9061
rect 7742 9052 7748 9104
rect 7800 9092 7806 9104
rect 7800 9064 10548 9092
rect 7800 9052 7806 9064
rect 4154 9033 4160 9036
rect 4148 9024 4160 9033
rect 4115 8996 4160 9024
rect 4148 8987 4160 8996
rect 4154 8984 4160 8987
rect 4212 8984 4218 9036
rect 6454 8984 6460 9036
rect 6512 9024 6518 9036
rect 8202 9024 8208 9036
rect 6512 8996 7144 9024
rect 8163 8996 8208 9024
rect 6512 8984 6518 8996
rect 7116 8965 7144 8996
rect 8202 8984 8208 8996
rect 8260 8984 8266 9036
rect 8941 9027 8999 9033
rect 8941 8993 8953 9027
rect 8987 9024 8999 9027
rect 9398 9024 9404 9036
rect 8987 8996 9404 9024
rect 8987 8993 8999 8996
rect 8941 8987 8999 8993
rect 9398 8984 9404 8996
rect 9456 9024 9462 9036
rect 9585 9027 9643 9033
rect 9585 9024 9597 9027
rect 9456 8996 9597 9024
rect 9456 8984 9462 8996
rect 9585 8993 9597 8996
rect 9631 8993 9643 9027
rect 9585 8987 9643 8993
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8925 3479 8959
rect 3421 8919 3479 8925
rect 3605 8959 3663 8965
rect 3605 8925 3617 8959
rect 3651 8925 3663 8959
rect 3605 8919 3663 8925
rect 3881 8959 3939 8965
rect 3881 8925 3893 8959
rect 3927 8925 3939 8959
rect 3881 8919 3939 8925
rect 5353 8959 5411 8965
rect 5353 8925 5365 8959
rect 5399 8925 5411 8959
rect 5353 8919 5411 8925
rect 6917 8959 6975 8965
rect 6917 8925 6929 8959
rect 6963 8925 6975 8959
rect 6917 8919 6975 8925
rect 7101 8959 7159 8965
rect 7101 8925 7113 8959
rect 7147 8956 7159 8959
rect 7926 8956 7932 8968
rect 7147 8928 7696 8956
rect 7887 8928 7932 8956
rect 7147 8925 7159 8928
rect 7101 8919 7159 8925
rect 3436 8888 3464 8919
rect 3786 8888 3792 8900
rect 3436 8860 3792 8888
rect 3786 8848 3792 8860
rect 3844 8848 3850 8900
rect 2866 8780 2872 8832
rect 2924 8820 2930 8832
rect 2961 8823 3019 8829
rect 2961 8820 2973 8823
rect 2924 8792 2973 8820
rect 2924 8780 2930 8792
rect 2961 8789 2973 8792
rect 3007 8789 3019 8823
rect 2961 8783 3019 8789
rect 3050 8780 3056 8832
rect 3108 8820 3114 8832
rect 3896 8820 3924 8919
rect 5368 8820 5396 8919
rect 6730 8888 6736 8900
rect 6643 8860 6736 8888
rect 6730 8848 6736 8860
rect 6788 8888 6794 8900
rect 6932 8888 6960 8919
rect 6788 8860 6960 8888
rect 6788 8848 6794 8860
rect 6454 8820 6460 8832
rect 3108 8792 6460 8820
rect 3108 8780 3114 8792
rect 6454 8780 6460 8792
rect 6512 8780 6518 8832
rect 7558 8820 7564 8832
rect 7519 8792 7564 8820
rect 7558 8780 7564 8792
rect 7616 8780 7622 8832
rect 7668 8820 7696 8928
rect 7926 8916 7932 8928
rect 7984 8916 7990 8968
rect 8110 8956 8116 8968
rect 8071 8928 8116 8956
rect 8110 8916 8116 8928
rect 8168 8916 8174 8968
rect 8754 8956 8760 8968
rect 8715 8928 8760 8956
rect 8754 8916 8760 8928
rect 8812 8916 8818 8968
rect 10520 8965 10548 9064
rect 9677 8959 9735 8965
rect 9677 8956 9689 8959
rect 9600 8928 9689 8956
rect 8573 8891 8631 8897
rect 8573 8857 8585 8891
rect 8619 8888 8631 8891
rect 8938 8888 8944 8900
rect 8619 8860 8944 8888
rect 8619 8857 8631 8860
rect 8573 8851 8631 8857
rect 8938 8848 8944 8860
rect 8996 8848 9002 8900
rect 9214 8848 9220 8900
rect 9272 8888 9278 8900
rect 9600 8888 9628 8928
rect 9677 8925 9689 8928
rect 9723 8925 9735 8959
rect 9677 8919 9735 8925
rect 10505 8959 10563 8965
rect 10505 8925 10517 8959
rect 10551 8925 10563 8959
rect 10505 8919 10563 8925
rect 10594 8916 10600 8968
rect 10652 8956 10658 8968
rect 10704 8956 10732 9132
rect 12802 9120 12808 9132
rect 12860 9120 12866 9172
rect 12986 9120 12992 9172
rect 13044 9160 13050 9172
rect 14458 9160 14464 9172
rect 13044 9132 14464 9160
rect 13044 9120 13050 9132
rect 14458 9120 14464 9132
rect 14516 9120 14522 9172
rect 10778 9052 10784 9104
rect 10836 9092 10842 9104
rect 15102 9092 15108 9104
rect 10836 9064 15108 9092
rect 10836 9052 10842 9064
rect 15102 9052 15108 9064
rect 15160 9052 15166 9104
rect 11048 9027 11106 9033
rect 11048 8993 11060 9027
rect 11094 9024 11106 9027
rect 11330 9024 11336 9036
rect 11094 8996 11336 9024
rect 11094 8993 11106 8996
rect 11048 8987 11106 8993
rect 11330 8984 11336 8996
rect 11388 8984 11394 9036
rect 12710 8984 12716 9036
rect 12768 9024 12774 9036
rect 12897 9027 12955 9033
rect 12897 9024 12909 9027
rect 12768 8996 12909 9024
rect 12768 8984 12774 8996
rect 12897 8993 12909 8996
rect 12943 9024 12955 9027
rect 13357 9027 13415 9033
rect 13357 9024 13369 9027
rect 12943 8996 13369 9024
rect 12943 8993 12955 8996
rect 12897 8987 12955 8993
rect 13357 8993 13369 8996
rect 13403 8993 13415 9027
rect 13357 8987 13415 8993
rect 10781 8959 10839 8965
rect 10781 8956 10793 8959
rect 10652 8928 10793 8956
rect 10652 8916 10658 8928
rect 10781 8925 10793 8928
rect 10827 8925 10839 8959
rect 12621 8959 12679 8965
rect 12621 8956 12633 8959
rect 10781 8919 10839 8925
rect 12176 8928 12633 8956
rect 9272 8860 9628 8888
rect 9272 8848 9278 8860
rect 7745 8823 7803 8829
rect 7745 8820 7757 8823
rect 7668 8792 7757 8820
rect 7745 8789 7757 8792
rect 7791 8820 7803 8823
rect 8846 8820 8852 8832
rect 7791 8792 8852 8820
rect 7791 8789 7803 8792
rect 7745 8783 7803 8789
rect 8846 8780 8852 8792
rect 8904 8780 8910 8832
rect 9030 8780 9036 8832
rect 9088 8820 9094 8832
rect 9125 8823 9183 8829
rect 9125 8820 9137 8823
rect 9088 8792 9137 8820
rect 9088 8780 9094 8792
rect 9125 8789 9137 8792
rect 9171 8789 9183 8823
rect 9125 8783 9183 8789
rect 9950 8780 9956 8832
rect 10008 8820 10014 8832
rect 11422 8820 11428 8832
rect 10008 8792 11428 8820
rect 10008 8780 10014 8792
rect 11422 8780 11428 8792
rect 11480 8820 11486 8832
rect 11790 8820 11796 8832
rect 11480 8792 11796 8820
rect 11480 8780 11486 8792
rect 11790 8780 11796 8792
rect 11848 8780 11854 8832
rect 11974 8780 11980 8832
rect 12032 8820 12038 8832
rect 12176 8829 12204 8928
rect 12621 8925 12633 8928
rect 12667 8925 12679 8959
rect 12621 8919 12679 8925
rect 12805 8959 12863 8965
rect 12805 8925 12817 8959
rect 12851 8925 12863 8959
rect 12805 8919 12863 8925
rect 12820 8888 12848 8919
rect 12544 8860 12848 8888
rect 12544 8832 12572 8860
rect 12161 8823 12219 8829
rect 12161 8820 12173 8823
rect 12032 8792 12173 8820
rect 12032 8780 12038 8792
rect 12161 8789 12173 8792
rect 12207 8789 12219 8823
rect 12161 8783 12219 8789
rect 12437 8823 12495 8829
rect 12437 8789 12449 8823
rect 12483 8820 12495 8823
rect 12526 8820 12532 8832
rect 12483 8792 12532 8820
rect 12483 8789 12495 8792
rect 12437 8783 12495 8789
rect 12526 8780 12532 8792
rect 12584 8780 12590 8832
rect 12894 8780 12900 8832
rect 12952 8820 12958 8832
rect 13265 8823 13323 8829
rect 13265 8820 13277 8823
rect 12952 8792 13277 8820
rect 12952 8780 12958 8792
rect 13265 8789 13277 8792
rect 13311 8789 13323 8823
rect 13265 8783 13323 8789
rect 1104 8730 16008 8752
rect 1104 8678 3480 8730
rect 3532 8678 3544 8730
rect 3596 8678 3608 8730
rect 3660 8678 3672 8730
rect 3724 8678 8478 8730
rect 8530 8678 8542 8730
rect 8594 8678 8606 8730
rect 8658 8678 8670 8730
rect 8722 8678 13475 8730
rect 13527 8678 13539 8730
rect 13591 8678 13603 8730
rect 13655 8678 13667 8730
rect 13719 8678 16008 8730
rect 1104 8656 16008 8678
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 1780 8588 3740 8616
rect 1780 8421 1808 8588
rect 3712 8548 3740 8588
rect 3786 8576 3792 8628
rect 3844 8616 3850 8628
rect 3973 8619 4031 8625
rect 3973 8616 3985 8619
rect 3844 8588 3985 8616
rect 3844 8576 3850 8588
rect 3973 8585 3985 8588
rect 4019 8585 4031 8619
rect 3973 8579 4031 8585
rect 4356 8588 8156 8616
rect 4356 8548 4384 8588
rect 5077 8551 5135 8557
rect 5077 8548 5089 8551
rect 3712 8520 4384 8548
rect 4448 8520 5089 8548
rect 4246 8480 4252 8492
rect 3804 8452 4252 8480
rect 1765 8415 1823 8421
rect 1765 8381 1777 8415
rect 1811 8381 1823 8415
rect 1765 8375 1823 8381
rect 2501 8415 2559 8421
rect 2501 8381 2513 8415
rect 2547 8381 2559 8415
rect 2501 8375 2559 8381
rect 2768 8415 2826 8421
rect 2768 8381 2780 8415
rect 2814 8412 2826 8415
rect 3804 8412 3832 8452
rect 4246 8440 4252 8452
rect 4304 8440 4310 8492
rect 4448 8489 4476 8520
rect 5077 8517 5089 8520
rect 5123 8517 5135 8551
rect 6270 8548 6276 8560
rect 6231 8520 6276 8548
rect 5077 8511 5135 8517
rect 6270 8508 6276 8520
rect 6328 8508 6334 8560
rect 8128 8548 8156 8588
rect 8202 8576 8208 8628
rect 8260 8616 8266 8628
rect 8481 8619 8539 8625
rect 8481 8616 8493 8619
rect 8260 8588 8493 8616
rect 8260 8576 8266 8588
rect 8481 8585 8493 8588
rect 8527 8585 8539 8619
rect 8481 8579 8539 8585
rect 9585 8619 9643 8625
rect 9585 8585 9597 8619
rect 9631 8616 9643 8619
rect 11330 8616 11336 8628
rect 9631 8588 11192 8616
rect 11291 8588 11336 8616
rect 9631 8585 9643 8588
rect 9585 8579 9643 8585
rect 9858 8548 9864 8560
rect 8128 8520 9864 8548
rect 9858 8508 9864 8520
rect 9916 8508 9922 8560
rect 9950 8508 9956 8560
rect 10008 8508 10014 8560
rect 11164 8548 11192 8588
rect 11330 8576 11336 8588
rect 11388 8576 11394 8628
rect 11790 8576 11796 8628
rect 11848 8616 11854 8628
rect 11885 8619 11943 8625
rect 11885 8616 11897 8619
rect 11848 8588 11897 8616
rect 11848 8576 11854 8588
rect 11885 8585 11897 8588
rect 11931 8585 11943 8619
rect 11885 8579 11943 8585
rect 11164 8520 11376 8548
rect 4433 8483 4491 8489
rect 4433 8449 4445 8483
rect 4479 8449 4491 8483
rect 4433 8443 4491 8449
rect 4525 8483 4583 8489
rect 4525 8449 4537 8483
rect 4571 8449 4583 8483
rect 5166 8480 5172 8492
rect 4525 8443 4583 8449
rect 4632 8452 5172 8480
rect 4154 8412 4160 8424
rect 2814 8384 3832 8412
rect 3896 8384 4160 8412
rect 2814 8381 2826 8384
rect 2768 8375 2826 8381
rect 2516 8344 2544 8375
rect 2958 8344 2964 8356
rect 2516 8316 2964 8344
rect 2958 8304 2964 8316
rect 3016 8304 3022 8356
rect 3896 8285 3924 8384
rect 4154 8372 4160 8384
rect 4212 8412 4218 8424
rect 4540 8412 4568 8443
rect 4212 8384 4568 8412
rect 4212 8372 4218 8384
rect 4632 8356 4660 8452
rect 5166 8440 5172 8452
rect 5224 8480 5230 8492
rect 5629 8483 5687 8489
rect 5629 8480 5641 8483
rect 5224 8452 5641 8480
rect 5224 8440 5230 8452
rect 5629 8449 5641 8452
rect 5675 8449 5687 8483
rect 5629 8443 5687 8449
rect 5718 8440 5724 8492
rect 5776 8480 5782 8492
rect 5905 8483 5963 8489
rect 5905 8480 5917 8483
rect 5776 8452 5917 8480
rect 5776 8440 5782 8452
rect 5905 8449 5917 8452
rect 5951 8449 5963 8483
rect 6454 8480 6460 8492
rect 6415 8452 6460 8480
rect 5905 8443 5963 8449
rect 6454 8440 6460 8452
rect 6512 8440 6518 8492
rect 9125 8483 9183 8489
rect 9125 8449 9137 8483
rect 9171 8480 9183 8483
rect 9214 8480 9220 8492
rect 9171 8452 9220 8480
rect 9171 8449 9183 8452
rect 9125 8443 9183 8449
rect 9214 8440 9220 8452
rect 9272 8440 9278 8492
rect 9968 8480 9996 8508
rect 9600 8452 9996 8480
rect 4246 8304 4252 8356
rect 4304 8344 4310 8356
rect 4614 8344 4620 8356
rect 4304 8316 4620 8344
rect 4304 8304 4310 8316
rect 4614 8304 4620 8316
rect 4672 8304 4678 8356
rect 5445 8347 5503 8353
rect 5445 8313 5457 8347
rect 5491 8344 5503 8347
rect 5626 8344 5632 8356
rect 5491 8316 5632 8344
rect 5491 8313 5503 8316
rect 5445 8307 5503 8313
rect 5626 8304 5632 8316
rect 5684 8304 5690 8356
rect 6472 8344 6500 8440
rect 6730 8421 6736 8424
rect 6724 8412 6736 8421
rect 6691 8384 6736 8412
rect 6724 8375 6736 8384
rect 6730 8372 6736 8375
rect 6788 8372 6794 8424
rect 7190 8372 7196 8424
rect 7248 8412 7254 8424
rect 7466 8412 7472 8424
rect 7248 8384 7472 8412
rect 7248 8372 7254 8384
rect 7466 8372 7472 8384
rect 7524 8412 7530 8424
rect 7929 8415 7987 8421
rect 7929 8412 7941 8415
rect 7524 8384 7941 8412
rect 7524 8372 7530 8384
rect 7929 8381 7941 8384
rect 7975 8381 7987 8415
rect 7929 8375 7987 8381
rect 8018 8372 8024 8424
rect 8076 8412 8082 8424
rect 8113 8415 8171 8421
rect 8113 8412 8125 8415
rect 8076 8384 8125 8412
rect 8076 8372 8082 8384
rect 8113 8381 8125 8384
rect 8159 8412 8171 8415
rect 8297 8415 8355 8421
rect 8297 8412 8309 8415
rect 8159 8384 8309 8412
rect 8159 8381 8171 8384
rect 8113 8375 8171 8381
rect 8297 8381 8309 8384
rect 8343 8381 8355 8415
rect 8297 8375 8355 8381
rect 8849 8415 8907 8421
rect 8849 8381 8861 8415
rect 8895 8412 8907 8415
rect 9600 8412 9628 8452
rect 8895 8384 9628 8412
rect 9677 8415 9735 8421
rect 8895 8381 8907 8384
rect 8849 8375 8907 8381
rect 9677 8381 9689 8415
rect 9723 8412 9735 8415
rect 9766 8412 9772 8424
rect 9723 8384 9772 8412
rect 9723 8381 9735 8384
rect 9677 8375 9735 8381
rect 6914 8344 6920 8356
rect 6472 8316 6920 8344
rect 6914 8304 6920 8316
rect 6972 8304 6978 8356
rect 7282 8304 7288 8356
rect 7340 8344 7346 8356
rect 8312 8344 8340 8375
rect 9766 8372 9772 8384
rect 9824 8372 9830 8424
rect 9953 8415 10011 8421
rect 9953 8381 9965 8415
rect 9999 8412 10011 8415
rect 10594 8412 10600 8424
rect 9999 8384 10600 8412
rect 9999 8381 10011 8384
rect 9953 8375 10011 8381
rect 8941 8347 8999 8353
rect 8941 8344 8953 8347
rect 7340 8316 7880 8344
rect 8312 8316 8953 8344
rect 7340 8304 7346 8316
rect 3881 8279 3939 8285
rect 3881 8245 3893 8279
rect 3927 8245 3939 8279
rect 4338 8276 4344 8288
rect 4299 8248 4344 8276
rect 3881 8239 3939 8245
rect 4338 8236 4344 8248
rect 4396 8236 4402 8288
rect 4985 8279 5043 8285
rect 4985 8245 4997 8279
rect 5031 8276 5043 8279
rect 5074 8276 5080 8288
rect 5031 8248 5080 8276
rect 5031 8245 5043 8248
rect 4985 8239 5043 8245
rect 5074 8236 5080 8248
rect 5132 8236 5138 8288
rect 5534 8236 5540 8288
rect 5592 8276 5598 8288
rect 7852 8285 7880 8316
rect 8941 8313 8953 8316
rect 8987 8344 8999 8347
rect 9585 8347 9643 8353
rect 9585 8344 9597 8347
rect 8987 8316 9597 8344
rect 8987 8313 8999 8316
rect 8941 8307 8999 8313
rect 9585 8313 9597 8316
rect 9631 8313 9643 8347
rect 9585 8307 9643 8313
rect 7837 8279 7895 8285
rect 5592 8248 5637 8276
rect 5592 8236 5598 8248
rect 7837 8245 7849 8279
rect 7883 8245 7895 8279
rect 9490 8276 9496 8288
rect 9451 8248 9496 8276
rect 7837 8239 7895 8245
rect 9490 8236 9496 8248
rect 9548 8236 9554 8288
rect 9674 8236 9680 8288
rect 9732 8276 9738 8288
rect 9861 8279 9919 8285
rect 9861 8276 9873 8279
rect 9732 8248 9873 8276
rect 9732 8236 9738 8248
rect 9861 8245 9873 8248
rect 9907 8276 9919 8279
rect 9968 8276 9996 8375
rect 10594 8372 10600 8384
rect 10652 8372 10658 8424
rect 10226 8353 10232 8356
rect 10220 8344 10232 8353
rect 10187 8316 10232 8344
rect 10220 8307 10232 8316
rect 10226 8304 10232 8307
rect 10284 8304 10290 8356
rect 9907 8248 9996 8276
rect 11348 8276 11376 8520
rect 11900 8412 11928 8579
rect 13262 8576 13268 8628
rect 13320 8616 13326 8628
rect 14277 8619 14335 8625
rect 14277 8616 14289 8619
rect 13320 8588 14289 8616
rect 13320 8576 13326 8588
rect 14277 8585 14289 8588
rect 14323 8585 14335 8619
rect 14277 8579 14335 8585
rect 11974 8440 11980 8492
rect 12032 8480 12038 8492
rect 12161 8483 12219 8489
rect 12161 8480 12173 8483
rect 12032 8452 12173 8480
rect 12032 8440 12038 8452
rect 12161 8449 12173 8452
rect 12207 8480 12219 8483
rect 12207 8452 13032 8480
rect 12207 8449 12219 8452
rect 12161 8443 12219 8449
rect 12345 8415 12403 8421
rect 12345 8412 12357 8415
rect 11900 8384 12357 8412
rect 12345 8381 12357 8384
rect 12391 8381 12403 8415
rect 12345 8375 12403 8381
rect 12802 8372 12808 8424
rect 12860 8412 12866 8424
rect 12897 8415 12955 8421
rect 12897 8412 12909 8415
rect 12860 8384 12909 8412
rect 12860 8372 12866 8384
rect 12897 8381 12909 8384
rect 12943 8381 12955 8415
rect 13004 8412 13032 8452
rect 13153 8415 13211 8421
rect 13153 8412 13165 8415
rect 13004 8384 13165 8412
rect 12897 8375 12955 8381
rect 13153 8381 13165 8384
rect 13199 8381 13211 8415
rect 13153 8375 13211 8381
rect 12437 8347 12495 8353
rect 12437 8313 12449 8347
rect 12483 8344 12495 8347
rect 13446 8344 13452 8356
rect 12483 8316 13452 8344
rect 12483 8313 12495 8316
rect 12437 8307 12495 8313
rect 11793 8279 11851 8285
rect 11793 8276 11805 8279
rect 11348 8248 11805 8276
rect 9907 8245 9919 8248
rect 9861 8239 9919 8245
rect 11793 8245 11805 8248
rect 11839 8276 11851 8279
rect 12452 8276 12480 8307
rect 13446 8304 13452 8316
rect 13504 8344 13510 8356
rect 14366 8344 14372 8356
rect 13504 8316 14372 8344
rect 13504 8304 13510 8316
rect 14366 8304 14372 8316
rect 14424 8304 14430 8356
rect 12802 8276 12808 8288
rect 11839 8248 12480 8276
rect 12763 8248 12808 8276
rect 11839 8245 11851 8248
rect 11793 8239 11851 8245
rect 12802 8236 12808 8248
rect 12860 8236 12866 8288
rect 1104 8186 16008 8208
rect 1104 8134 5979 8186
rect 6031 8134 6043 8186
rect 6095 8134 6107 8186
rect 6159 8134 6171 8186
rect 6223 8134 10976 8186
rect 11028 8134 11040 8186
rect 11092 8134 11104 8186
rect 11156 8134 11168 8186
rect 11220 8134 16008 8186
rect 1104 8112 16008 8134
rect 1486 8072 1492 8084
rect 1447 8044 1492 8072
rect 1486 8032 1492 8044
rect 1544 8032 1550 8084
rect 1765 8075 1823 8081
rect 1765 8072 1777 8075
rect 1596 8044 1777 8072
rect 1596 8013 1624 8044
rect 1765 8041 1777 8044
rect 1811 8041 1823 8075
rect 1765 8035 1823 8041
rect 4065 8075 4123 8081
rect 4065 8041 4077 8075
rect 4111 8072 4123 8075
rect 4338 8072 4344 8084
rect 4111 8044 4344 8072
rect 4111 8041 4123 8044
rect 4065 8035 4123 8041
rect 4338 8032 4344 8044
rect 4396 8032 4402 8084
rect 4433 8075 4491 8081
rect 4433 8041 4445 8075
rect 4479 8072 4491 8075
rect 4890 8072 4896 8084
rect 4479 8044 4896 8072
rect 4479 8041 4491 8044
rect 4433 8035 4491 8041
rect 4890 8032 4896 8044
rect 4948 8072 4954 8084
rect 5169 8075 5227 8081
rect 5169 8072 5181 8075
rect 4948 8044 5181 8072
rect 4948 8032 4954 8044
rect 5169 8041 5181 8044
rect 5215 8041 5227 8075
rect 5169 8035 5227 8041
rect 5442 8032 5448 8084
rect 5500 8072 5506 8084
rect 7098 8072 7104 8084
rect 5500 8044 7104 8072
rect 5500 8032 5506 8044
rect 7098 8032 7104 8044
rect 7156 8032 7162 8084
rect 7285 8075 7343 8081
rect 7285 8041 7297 8075
rect 7331 8072 7343 8075
rect 7558 8072 7564 8084
rect 7331 8044 7564 8072
rect 7331 8041 7343 8044
rect 7285 8035 7343 8041
rect 7558 8032 7564 8044
rect 7616 8032 7622 8084
rect 7745 8075 7803 8081
rect 7745 8041 7757 8075
rect 7791 8072 7803 8075
rect 8110 8072 8116 8084
rect 7791 8044 8116 8072
rect 7791 8041 7803 8044
rect 7745 8035 7803 8041
rect 8110 8032 8116 8044
rect 8168 8032 8174 8084
rect 8573 8075 8631 8081
rect 8220 8044 8432 8072
rect 1581 8007 1639 8013
rect 1581 7973 1593 8007
rect 1627 7973 1639 8007
rect 1581 7967 1639 7973
rect 2746 7976 7144 8004
rect 1949 7939 2007 7945
rect 1949 7905 1961 7939
rect 1995 7936 2007 7939
rect 2746 7936 2774 7976
rect 1995 7908 2774 7936
rect 3697 7939 3755 7945
rect 1995 7905 2007 7908
rect 1949 7899 2007 7905
rect 3697 7905 3709 7939
rect 3743 7936 3755 7939
rect 3973 7939 4031 7945
rect 3973 7936 3985 7939
rect 3743 7908 3985 7936
rect 3743 7905 3755 7908
rect 3697 7899 3755 7905
rect 3973 7905 3985 7908
rect 4019 7936 4031 7939
rect 4338 7936 4344 7948
rect 4019 7908 4344 7936
rect 4019 7905 4031 7908
rect 3973 7899 4031 7905
rect 4338 7896 4344 7908
rect 4396 7896 4402 7948
rect 4890 7936 4896 7948
rect 4851 7908 4896 7936
rect 4890 7896 4896 7908
rect 4948 7896 4954 7948
rect 6178 7896 6184 7948
rect 6236 7936 6242 7948
rect 6466 7939 6524 7945
rect 6466 7936 6478 7939
rect 6236 7908 6478 7936
rect 6236 7896 6242 7908
rect 6466 7905 6478 7908
rect 6512 7905 6524 7939
rect 6466 7899 6524 7905
rect 6733 7939 6791 7945
rect 6733 7905 6745 7939
rect 6779 7936 6791 7939
rect 6914 7936 6920 7948
rect 6779 7908 6920 7936
rect 6779 7905 6791 7908
rect 6733 7899 6791 7905
rect 6914 7896 6920 7908
rect 6972 7896 6978 7948
rect 2774 7828 2780 7880
rect 2832 7868 2838 7880
rect 4062 7868 4068 7880
rect 2832 7840 4068 7868
rect 2832 7828 2838 7840
rect 4062 7828 4068 7840
rect 4120 7828 4126 7880
rect 4522 7868 4528 7880
rect 4483 7840 4528 7868
rect 4522 7828 4528 7840
rect 4580 7828 4586 7880
rect 4614 7828 4620 7880
rect 4672 7868 4678 7880
rect 4672 7840 5396 7868
rect 4672 7828 4678 7840
rect 2958 7760 2964 7812
rect 3016 7800 3022 7812
rect 5368 7809 5396 7840
rect 5077 7803 5135 7809
rect 5077 7800 5089 7803
rect 3016 7772 5089 7800
rect 3016 7760 3022 7772
rect 5077 7769 5089 7772
rect 5123 7769 5135 7803
rect 5077 7763 5135 7769
rect 5353 7803 5411 7809
rect 5353 7769 5365 7803
rect 5399 7769 5411 7803
rect 7116 7800 7144 7976
rect 7190 7964 7196 8016
rect 7248 8004 7254 8016
rect 7377 8007 7435 8013
rect 7377 8004 7389 8007
rect 7248 7976 7389 8004
rect 7248 7964 7254 7976
rect 7377 7973 7389 7976
rect 7423 7973 7435 8007
rect 7377 7967 7435 7973
rect 7466 7964 7472 8016
rect 7524 8004 7530 8016
rect 8220 8004 8248 8044
rect 7524 7976 8248 8004
rect 7524 7964 7530 7976
rect 8294 7964 8300 8016
rect 8352 7964 8358 8016
rect 8021 7939 8079 7945
rect 8021 7905 8033 7939
rect 8067 7936 8079 7939
rect 8312 7936 8340 7964
rect 8067 7908 8340 7936
rect 8404 7936 8432 8044
rect 8573 8041 8585 8075
rect 8619 8072 8631 8075
rect 9125 8075 9183 8081
rect 9125 8072 9137 8075
rect 8619 8044 9137 8072
rect 8619 8041 8631 8044
rect 8573 8035 8631 8041
rect 9125 8041 9137 8044
rect 9171 8041 9183 8075
rect 9490 8072 9496 8084
rect 9451 8044 9496 8072
rect 9125 8035 9183 8041
rect 9490 8032 9496 8044
rect 9548 8032 9554 8084
rect 10873 8075 10931 8081
rect 10873 8041 10885 8075
rect 10919 8072 10931 8075
rect 11425 8075 11483 8081
rect 11425 8072 11437 8075
rect 10919 8044 11437 8072
rect 10919 8041 10931 8044
rect 10873 8035 10931 8041
rect 11425 8041 11437 8044
rect 11471 8041 11483 8075
rect 11425 8035 11483 8041
rect 12434 8032 12440 8084
rect 12492 8072 12498 8084
rect 12529 8075 12587 8081
rect 12529 8072 12541 8075
rect 12492 8044 12541 8072
rect 12492 8032 12498 8044
rect 12529 8041 12541 8044
rect 12575 8041 12587 8075
rect 12529 8035 12587 8041
rect 12802 8032 12808 8084
rect 12860 8072 12866 8084
rect 12989 8075 13047 8081
rect 12989 8072 13001 8075
rect 12860 8044 13001 8072
rect 12860 8032 12866 8044
rect 12989 8041 13001 8044
rect 13035 8041 13047 8075
rect 13354 8072 13360 8084
rect 13315 8044 13360 8072
rect 12989 8035 13047 8041
rect 13354 8032 13360 8044
rect 13412 8032 13418 8084
rect 13725 8075 13783 8081
rect 13725 8041 13737 8075
rect 13771 8072 13783 8075
rect 13998 8072 14004 8084
rect 13771 8044 14004 8072
rect 13771 8041 13783 8044
rect 13725 8035 13783 8041
rect 8481 8007 8539 8013
rect 8481 7973 8493 8007
rect 8527 8004 8539 8007
rect 9030 8004 9036 8016
rect 8527 7976 9036 8004
rect 8527 7973 8539 7976
rect 8481 7967 8539 7973
rect 9030 7964 9036 7976
rect 9088 7964 9094 8016
rect 11333 8007 11391 8013
rect 9140 7976 11284 8004
rect 9140 7936 9168 7976
rect 8404 7908 9168 7936
rect 8067 7905 8079 7908
rect 8021 7899 8079 7905
rect 9214 7896 9220 7948
rect 9272 7936 9278 7948
rect 10318 7936 10324 7948
rect 9272 7908 9720 7936
rect 9272 7896 9278 7908
rect 7193 7871 7251 7877
rect 7193 7837 7205 7871
rect 7239 7868 7251 7871
rect 7282 7868 7288 7880
rect 7239 7840 7288 7868
rect 7239 7837 7251 7840
rect 7193 7831 7251 7837
rect 7282 7828 7288 7840
rect 7340 7828 7346 7880
rect 7926 7828 7932 7880
rect 7984 7868 7990 7880
rect 8297 7871 8355 7877
rect 8297 7868 8309 7871
rect 7984 7840 8309 7868
rect 7984 7828 7990 7840
rect 8297 7837 8309 7840
rect 8343 7837 8355 7871
rect 8297 7831 8355 7837
rect 9306 7828 9312 7880
rect 9364 7868 9370 7880
rect 9582 7868 9588 7880
rect 9364 7840 9588 7868
rect 9364 7828 9370 7840
rect 9582 7828 9588 7840
rect 9640 7828 9646 7880
rect 9692 7877 9720 7908
rect 9784 7908 10324 7936
rect 9677 7871 9735 7877
rect 9677 7837 9689 7871
rect 9723 7837 9735 7871
rect 9677 7831 9735 7837
rect 8110 7800 8116 7812
rect 7116 7772 8116 7800
rect 5353 7763 5411 7769
rect 8110 7760 8116 7772
rect 8168 7760 8174 7812
rect 8386 7760 8392 7812
rect 8444 7800 8450 7812
rect 9784 7800 9812 7908
rect 10318 7896 10324 7908
rect 10376 7896 10382 7948
rect 10505 7939 10563 7945
rect 10505 7905 10517 7939
rect 10551 7936 10563 7939
rect 10594 7936 10600 7948
rect 10551 7908 10600 7936
rect 10551 7905 10563 7908
rect 10505 7899 10563 7905
rect 10594 7896 10600 7908
rect 10652 7896 10658 7948
rect 11256 7936 11284 7976
rect 11333 7973 11345 8007
rect 11379 8004 11391 8007
rect 12894 8004 12900 8016
rect 11379 7976 12756 8004
rect 12855 7976 12900 8004
rect 11379 7973 11391 7976
rect 11333 7967 11391 7973
rect 12161 7939 12219 7945
rect 11256 7908 12112 7936
rect 10226 7868 10232 7880
rect 10187 7840 10232 7868
rect 10226 7828 10232 7840
rect 10284 7828 10290 7880
rect 10410 7868 10416 7880
rect 10371 7840 10416 7868
rect 10410 7828 10416 7840
rect 10468 7828 10474 7880
rect 11330 7828 11336 7880
rect 11388 7868 11394 7880
rect 11517 7871 11575 7877
rect 11517 7868 11529 7871
rect 11388 7840 11529 7868
rect 11388 7828 11394 7840
rect 11517 7837 11529 7840
rect 11563 7837 11575 7871
rect 11974 7868 11980 7880
rect 11935 7840 11980 7868
rect 11517 7831 11575 7837
rect 11974 7828 11980 7840
rect 12032 7828 12038 7880
rect 12084 7877 12112 7908
rect 12161 7905 12173 7939
rect 12207 7936 12219 7939
rect 12728 7936 12756 7976
rect 12894 7964 12900 7976
rect 12952 7964 12958 8016
rect 13078 7936 13084 7948
rect 12207 7908 12664 7936
rect 12728 7908 13084 7936
rect 12207 7905 12219 7908
rect 12161 7899 12219 7905
rect 12069 7871 12127 7877
rect 12069 7837 12081 7871
rect 12115 7868 12127 7871
rect 12115 7840 12388 7868
rect 12115 7837 12127 7840
rect 12069 7831 12127 7837
rect 8444 7772 9812 7800
rect 8444 7760 8450 7772
rect 9858 7760 9864 7812
rect 9916 7800 9922 7812
rect 10965 7803 11023 7809
rect 10965 7800 10977 7803
rect 9916 7772 10977 7800
rect 9916 7760 9922 7772
rect 10965 7769 10977 7772
rect 11011 7769 11023 7803
rect 10965 7763 11023 7769
rect 3234 7692 3240 7744
rect 3292 7732 3298 7744
rect 3513 7735 3571 7741
rect 3513 7732 3525 7735
rect 3292 7704 3525 7732
rect 3292 7692 3298 7704
rect 3513 7701 3525 7704
rect 3559 7732 3571 7735
rect 5166 7732 5172 7744
rect 3559 7704 5172 7732
rect 3559 7701 3571 7704
rect 3513 7695 3571 7701
rect 5166 7692 5172 7704
rect 5224 7692 5230 7744
rect 5810 7692 5816 7744
rect 5868 7732 5874 7744
rect 6825 7735 6883 7741
rect 6825 7732 6837 7735
rect 5868 7704 6837 7732
rect 5868 7692 5874 7704
rect 6825 7701 6837 7704
rect 6871 7732 6883 7735
rect 7558 7732 7564 7744
rect 6871 7704 7564 7732
rect 6871 7701 6883 7704
rect 6825 7695 6883 7701
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 7837 7735 7895 7741
rect 7837 7701 7849 7735
rect 7883 7732 7895 7735
rect 8202 7732 8208 7744
rect 7883 7704 8208 7732
rect 7883 7701 7895 7704
rect 7837 7695 7895 7701
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 8846 7692 8852 7744
rect 8904 7732 8910 7744
rect 8941 7735 8999 7741
rect 8941 7732 8953 7735
rect 8904 7704 8953 7732
rect 8904 7692 8910 7704
rect 8941 7701 8953 7704
rect 8987 7701 8999 7735
rect 8941 7695 8999 7701
rect 9950 7692 9956 7744
rect 10008 7732 10014 7744
rect 10045 7735 10103 7741
rect 10045 7732 10057 7735
rect 10008 7704 10057 7732
rect 10008 7692 10014 7704
rect 10045 7701 10057 7704
rect 10091 7732 10103 7735
rect 12250 7732 12256 7744
rect 10091 7704 12256 7732
rect 10091 7701 10103 7704
rect 10045 7695 10103 7701
rect 12250 7692 12256 7704
rect 12308 7692 12314 7744
rect 12360 7732 12388 7840
rect 12636 7800 12664 7908
rect 13078 7896 13084 7908
rect 13136 7896 13142 7948
rect 12805 7871 12863 7877
rect 12805 7837 12817 7871
rect 12851 7868 12863 7871
rect 13262 7868 13268 7880
rect 12851 7840 13268 7868
rect 12851 7837 12863 7840
rect 12805 7831 12863 7837
rect 13262 7828 13268 7840
rect 13320 7828 13326 7880
rect 12710 7800 12716 7812
rect 12623 7772 12716 7800
rect 12710 7760 12716 7772
rect 12768 7800 12774 7812
rect 13740 7800 13768 8035
rect 13998 8032 14004 8044
rect 14056 8032 14062 8084
rect 12768 7772 13768 7800
rect 12768 7760 12774 7772
rect 12986 7732 12992 7744
rect 12360 7704 12992 7732
rect 12986 7692 12992 7704
rect 13044 7732 13050 7744
rect 13449 7735 13507 7741
rect 13449 7732 13461 7735
rect 13044 7704 13461 7732
rect 13044 7692 13050 7704
rect 13449 7701 13461 7704
rect 13495 7701 13507 7735
rect 13449 7695 13507 7701
rect 1104 7642 16008 7664
rect 1104 7590 3480 7642
rect 3532 7590 3544 7642
rect 3596 7590 3608 7642
rect 3660 7590 3672 7642
rect 3724 7590 8478 7642
rect 8530 7590 8542 7642
rect 8594 7590 8606 7642
rect 8658 7590 8670 7642
rect 8722 7590 13475 7642
rect 13527 7590 13539 7642
rect 13591 7590 13603 7642
rect 13655 7590 13667 7642
rect 13719 7590 16008 7642
rect 1104 7568 16008 7590
rect 2038 7488 2044 7540
rect 2096 7528 2102 7540
rect 2133 7531 2191 7537
rect 2133 7528 2145 7531
rect 2096 7500 2145 7528
rect 2096 7488 2102 7500
rect 2133 7497 2145 7500
rect 2179 7497 2191 7531
rect 2133 7491 2191 7497
rect 2314 7488 2320 7540
rect 2372 7528 2378 7540
rect 2774 7528 2780 7540
rect 2372 7500 2780 7528
rect 2372 7488 2378 7500
rect 2774 7488 2780 7500
rect 2832 7488 2838 7540
rect 2869 7531 2927 7537
rect 2869 7497 2881 7531
rect 2915 7528 2927 7531
rect 3234 7528 3240 7540
rect 2915 7500 3240 7528
rect 2915 7497 2927 7500
rect 2869 7491 2927 7497
rect 3234 7488 3240 7500
rect 3292 7488 3298 7540
rect 4433 7531 4491 7537
rect 4433 7497 4445 7531
rect 4479 7528 4491 7531
rect 4522 7528 4528 7540
rect 4479 7500 4528 7528
rect 4479 7497 4491 7500
rect 4433 7491 4491 7497
rect 4522 7488 4528 7500
rect 4580 7488 4586 7540
rect 5534 7528 5540 7540
rect 5495 7500 5540 7528
rect 5534 7488 5540 7500
rect 5592 7488 5598 7540
rect 5718 7488 5724 7540
rect 5776 7528 5782 7540
rect 6270 7528 6276 7540
rect 5776 7500 6276 7528
rect 5776 7488 5782 7500
rect 6270 7488 6276 7500
rect 6328 7528 6334 7540
rect 6641 7531 6699 7537
rect 6641 7528 6653 7531
rect 6328 7500 6653 7528
rect 6328 7488 6334 7500
rect 6641 7497 6653 7500
rect 6687 7497 6699 7531
rect 6641 7491 6699 7497
rect 6917 7531 6975 7537
rect 6917 7497 6929 7531
rect 6963 7528 6975 7531
rect 7190 7528 7196 7540
rect 6963 7500 7196 7528
rect 6963 7497 6975 7500
rect 6917 7491 6975 7497
rect 7190 7488 7196 7500
rect 7248 7528 7254 7540
rect 7650 7528 7656 7540
rect 7248 7500 7656 7528
rect 7248 7488 7254 7500
rect 7650 7488 7656 7500
rect 7708 7488 7714 7540
rect 7926 7488 7932 7540
rect 7984 7528 7990 7540
rect 8389 7531 8447 7537
rect 8389 7528 8401 7531
rect 7984 7500 8401 7528
rect 7984 7488 7990 7500
rect 8389 7497 8401 7500
rect 8435 7497 8447 7531
rect 9858 7528 9864 7540
rect 8389 7491 8447 7497
rect 9646 7500 9864 7528
rect 4341 7463 4399 7469
rect 4341 7429 4353 7463
rect 4387 7429 4399 7463
rect 4341 7423 4399 7429
rect 2866 7392 2872 7404
rect 2746 7364 2872 7392
rect 1949 7327 2007 7333
rect 1949 7293 1961 7327
rect 1995 7324 2007 7327
rect 2746 7324 2774 7364
rect 2866 7352 2872 7364
rect 2924 7352 2930 7404
rect 4356 7392 4384 7423
rect 8110 7420 8116 7472
rect 8168 7460 8174 7472
rect 8481 7463 8539 7469
rect 8481 7460 8493 7463
rect 8168 7432 8493 7460
rect 8168 7420 8174 7432
rect 8481 7429 8493 7432
rect 8527 7429 8539 7463
rect 9309 7463 9367 7469
rect 9309 7460 9321 7463
rect 8481 7423 8539 7429
rect 8588 7432 9321 7460
rect 5077 7395 5135 7401
rect 5077 7392 5089 7395
rect 4356 7364 5089 7392
rect 5077 7361 5089 7364
rect 5123 7392 5135 7395
rect 6178 7392 6184 7404
rect 5123 7364 6184 7392
rect 5123 7361 5135 7364
rect 5077 7355 5135 7361
rect 6178 7352 6184 7364
rect 6236 7352 6242 7404
rect 6914 7352 6920 7404
rect 6972 7392 6978 7404
rect 7009 7395 7067 7401
rect 7009 7392 7021 7395
rect 6972 7364 7021 7392
rect 6972 7352 6978 7364
rect 7009 7361 7021 7364
rect 7055 7361 7067 7395
rect 8588 7392 8616 7432
rect 9309 7429 9321 7432
rect 9355 7460 9367 7463
rect 9493 7463 9551 7469
rect 9493 7460 9505 7463
rect 9355 7432 9505 7460
rect 9355 7429 9367 7432
rect 9309 7423 9367 7429
rect 9493 7429 9505 7432
rect 9539 7460 9551 7463
rect 9646 7460 9674 7500
rect 9858 7488 9864 7500
rect 9916 7528 9922 7540
rect 10042 7528 10048 7540
rect 9916 7500 10048 7528
rect 9916 7488 9922 7500
rect 10042 7488 10048 7500
rect 10100 7488 10106 7540
rect 10318 7488 10324 7540
rect 10376 7528 10382 7540
rect 10778 7528 10784 7540
rect 10376 7500 10784 7528
rect 10376 7488 10382 7500
rect 10778 7488 10784 7500
rect 10836 7528 10842 7540
rect 11425 7531 11483 7537
rect 11425 7528 11437 7531
rect 10836 7500 11437 7528
rect 10836 7488 10842 7500
rect 11425 7497 11437 7500
rect 11471 7528 11483 7531
rect 11514 7528 11520 7540
rect 11471 7500 11520 7528
rect 11471 7497 11483 7500
rect 11425 7491 11483 7497
rect 11514 7488 11520 7500
rect 11572 7488 11578 7540
rect 9539 7432 9674 7460
rect 9539 7429 9551 7432
rect 9493 7423 9551 7429
rect 9030 7392 9036 7404
rect 7009 7355 7067 7361
rect 8036 7364 8616 7392
rect 8991 7364 9036 7392
rect 2958 7324 2964 7336
rect 1995 7296 2774 7324
rect 2919 7296 2964 7324
rect 1995 7293 2007 7296
rect 1949 7287 2007 7293
rect 2958 7284 2964 7296
rect 3016 7284 3022 7336
rect 4706 7284 4712 7336
rect 4764 7324 4770 7336
rect 4893 7327 4951 7333
rect 4893 7324 4905 7327
rect 4764 7296 4905 7324
rect 4764 7284 4770 7296
rect 4893 7293 4905 7296
rect 4939 7324 4951 7327
rect 5353 7327 5411 7333
rect 5353 7324 5365 7327
rect 4939 7296 5365 7324
rect 4939 7293 4951 7296
rect 4893 7287 4951 7293
rect 5353 7293 5365 7296
rect 5399 7324 5411 7327
rect 5534 7324 5540 7336
rect 5399 7296 5540 7324
rect 5399 7293 5411 7296
rect 5353 7287 5411 7293
rect 5534 7284 5540 7296
rect 5592 7284 5598 7336
rect 7558 7284 7564 7336
rect 7616 7324 7622 7336
rect 8036 7324 8064 7364
rect 9030 7352 9036 7364
rect 9088 7352 9094 7404
rect 9674 7352 9680 7404
rect 9732 7392 9738 7404
rect 9732 7364 9777 7392
rect 9732 7352 9738 7364
rect 11330 7352 11336 7404
rect 11388 7392 11394 7404
rect 11885 7395 11943 7401
rect 11885 7392 11897 7395
rect 11388 7364 11897 7392
rect 11388 7352 11394 7364
rect 11885 7361 11897 7364
rect 11931 7361 11943 7395
rect 12066 7392 12072 7404
rect 12027 7364 12072 7392
rect 11885 7355 11943 7361
rect 12066 7352 12072 7364
rect 12124 7352 12130 7404
rect 12618 7352 12624 7404
rect 12676 7392 12682 7404
rect 13262 7392 13268 7404
rect 12676 7364 13268 7392
rect 12676 7352 12682 7364
rect 13262 7352 13268 7364
rect 13320 7352 13326 7404
rect 8846 7324 8852 7336
rect 7616 7296 8064 7324
rect 8807 7296 8852 7324
rect 7616 7284 7622 7296
rect 8846 7284 8852 7296
rect 8904 7284 8910 7336
rect 8938 7284 8944 7336
rect 8996 7324 9002 7336
rect 11241 7327 11299 7333
rect 8996 7296 9041 7324
rect 9646 7296 10640 7324
rect 8996 7284 9002 7296
rect 3234 7265 3240 7268
rect 1581 7259 1639 7265
rect 1581 7225 1593 7259
rect 1627 7225 1639 7259
rect 3228 7256 3240 7265
rect 3195 7228 3240 7256
rect 1581 7219 1639 7225
rect 3228 7219 3240 7228
rect 1486 7188 1492 7200
rect 1447 7160 1492 7188
rect 1486 7148 1492 7160
rect 1544 7148 1550 7200
rect 1596 7188 1624 7219
rect 3234 7216 3240 7219
rect 3292 7216 3298 7268
rect 3418 7216 3424 7268
rect 3476 7256 3482 7268
rect 4801 7259 4859 7265
rect 4801 7256 4813 7259
rect 3476 7228 4813 7256
rect 3476 7216 3482 7228
rect 4801 7225 4813 7228
rect 4847 7256 4859 7259
rect 5074 7256 5080 7268
rect 4847 7228 5080 7256
rect 4847 7225 4859 7228
rect 4801 7219 4859 7225
rect 5074 7216 5080 7228
rect 5132 7216 5138 7268
rect 5166 7216 5172 7268
rect 5224 7256 5230 7268
rect 5224 7228 6592 7256
rect 5224 7216 5230 7228
rect 1765 7191 1823 7197
rect 1765 7188 1777 7191
rect 1596 7160 1777 7188
rect 1765 7157 1777 7160
rect 1811 7157 1823 7191
rect 2314 7188 2320 7200
rect 2275 7160 2320 7188
rect 1765 7151 1823 7157
rect 2314 7148 2320 7160
rect 2372 7148 2378 7200
rect 5258 7148 5264 7200
rect 5316 7188 5322 7200
rect 5810 7188 5816 7200
rect 5316 7160 5816 7188
rect 5316 7148 5322 7160
rect 5810 7148 5816 7160
rect 5868 7188 5874 7200
rect 5905 7191 5963 7197
rect 5905 7188 5917 7191
rect 5868 7160 5917 7188
rect 5868 7148 5874 7160
rect 5905 7157 5917 7160
rect 5951 7157 5963 7191
rect 5905 7151 5963 7157
rect 5997 7191 6055 7197
rect 5997 7157 6009 7191
rect 6043 7188 6055 7191
rect 6454 7188 6460 7200
rect 6043 7160 6460 7188
rect 6043 7157 6055 7160
rect 5997 7151 6055 7157
rect 6454 7148 6460 7160
rect 6512 7148 6518 7200
rect 6564 7188 6592 7228
rect 6822 7216 6828 7268
rect 6880 7256 6886 7268
rect 7254 7259 7312 7265
rect 7254 7256 7266 7259
rect 6880 7228 7266 7256
rect 6880 7216 6886 7228
rect 7254 7225 7266 7228
rect 7300 7225 7312 7259
rect 9646 7256 9674 7296
rect 7254 7219 7312 7225
rect 7392 7228 9674 7256
rect 9944 7259 10002 7265
rect 7392 7188 7420 7228
rect 9944 7225 9956 7259
rect 9990 7256 10002 7259
rect 10502 7256 10508 7268
rect 9990 7228 10508 7256
rect 9990 7225 10002 7228
rect 9944 7219 10002 7225
rect 10502 7216 10508 7228
rect 10560 7216 10566 7268
rect 10612 7256 10640 7296
rect 11241 7293 11253 7327
rect 11287 7324 11299 7327
rect 11606 7324 11612 7336
rect 11287 7296 11612 7324
rect 11287 7293 11299 7296
rect 11241 7287 11299 7293
rect 11606 7284 11612 7296
rect 11664 7284 11670 7336
rect 12158 7324 12164 7336
rect 12119 7296 12164 7324
rect 12158 7284 12164 7296
rect 12216 7324 12222 7336
rect 12216 7296 13032 7324
rect 12216 7284 12222 7296
rect 12710 7256 12716 7268
rect 10612 7228 12716 7256
rect 12710 7216 12716 7228
rect 12768 7216 12774 7268
rect 6564 7160 7420 7188
rect 7650 7148 7656 7200
rect 7708 7188 7714 7200
rect 10042 7188 10048 7200
rect 7708 7160 10048 7188
rect 7708 7148 7714 7160
rect 10042 7148 10048 7160
rect 10100 7148 10106 7200
rect 11057 7191 11115 7197
rect 11057 7157 11069 7191
rect 11103 7188 11115 7191
rect 11330 7188 11336 7200
rect 11103 7160 11336 7188
rect 11103 7157 11115 7160
rect 11057 7151 11115 7157
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 12526 7188 12532 7200
rect 12487 7160 12532 7188
rect 12526 7148 12532 7160
rect 12584 7148 12590 7200
rect 12618 7148 12624 7200
rect 12676 7188 12682 7200
rect 13004 7197 13032 7296
rect 12989 7191 13047 7197
rect 12676 7160 12721 7188
rect 12676 7148 12682 7160
rect 12989 7157 13001 7191
rect 13035 7188 13047 7191
rect 15838 7188 15844 7200
rect 13035 7160 15844 7188
rect 13035 7157 13047 7160
rect 12989 7151 13047 7157
rect 15838 7148 15844 7160
rect 15896 7148 15902 7200
rect 1104 7098 16008 7120
rect 1104 7046 5979 7098
rect 6031 7046 6043 7098
rect 6095 7046 6107 7098
rect 6159 7046 6171 7098
rect 6223 7046 10976 7098
rect 11028 7046 11040 7098
rect 11092 7046 11104 7098
rect 11156 7046 11168 7098
rect 11220 7046 16008 7098
rect 1104 7024 16008 7046
rect 3326 6944 3332 6996
rect 3384 6984 3390 6996
rect 7466 6984 7472 6996
rect 3384 6956 7472 6984
rect 3384 6944 3390 6956
rect 7466 6944 7472 6956
rect 7524 6944 7530 6996
rect 8202 6984 8208 6996
rect 7760 6956 8208 6984
rect 2498 6876 2504 6928
rect 2556 6916 2562 6928
rect 3418 6916 3424 6928
rect 2556 6888 3424 6916
rect 2556 6876 2562 6888
rect 3418 6876 3424 6888
rect 3476 6876 3482 6928
rect 4062 6876 4068 6928
rect 4120 6916 4126 6928
rect 4341 6919 4399 6925
rect 4341 6916 4353 6919
rect 4120 6888 4353 6916
rect 4120 6876 4126 6888
rect 4341 6885 4353 6888
rect 4387 6916 4399 6919
rect 4525 6919 4583 6925
rect 4525 6916 4537 6919
rect 4387 6888 4537 6916
rect 4387 6885 4399 6888
rect 4341 6879 4399 6885
rect 4525 6885 4537 6888
rect 4571 6916 4583 6919
rect 5534 6916 5540 6928
rect 4571 6888 5540 6916
rect 4571 6885 4583 6888
rect 4525 6879 4583 6885
rect 5534 6876 5540 6888
rect 5592 6916 5598 6928
rect 5905 6919 5963 6925
rect 5905 6916 5917 6919
rect 5592 6888 5917 6916
rect 5592 6876 5598 6888
rect 5905 6885 5917 6888
rect 5951 6885 5963 6919
rect 5905 6879 5963 6885
rect 1581 6851 1639 6857
rect 1581 6817 1593 6851
rect 1627 6848 1639 6851
rect 1762 6848 1768 6860
rect 1627 6820 1768 6848
rect 1627 6817 1639 6820
rect 1581 6811 1639 6817
rect 1762 6808 1768 6820
rect 1820 6808 1826 6860
rect 1946 6808 1952 6860
rect 2004 6848 2010 6860
rect 2113 6851 2171 6857
rect 2113 6848 2125 6851
rect 2004 6820 2125 6848
rect 2004 6808 2010 6820
rect 2113 6817 2125 6820
rect 2159 6817 2171 6851
rect 2113 6811 2171 6817
rect 2682 6808 2688 6860
rect 2740 6848 2746 6860
rect 4985 6851 5043 6857
rect 4985 6848 4997 6851
rect 2740 6820 4997 6848
rect 2740 6808 2746 6820
rect 4985 6817 4997 6820
rect 5031 6848 5043 6851
rect 5258 6848 5264 6860
rect 5031 6820 5264 6848
rect 5031 6817 5043 6820
rect 4985 6811 5043 6817
rect 5258 6808 5264 6820
rect 5316 6808 5322 6860
rect 5445 6851 5503 6857
rect 5445 6817 5457 6851
rect 5491 6848 5503 6851
rect 5718 6848 5724 6860
rect 5491 6820 5724 6848
rect 5491 6817 5503 6820
rect 5445 6811 5503 6817
rect 5718 6808 5724 6820
rect 5776 6808 5782 6860
rect 5997 6851 6055 6857
rect 5997 6817 6009 6851
rect 6043 6848 6055 6851
rect 6549 6851 6607 6857
rect 6043 6820 6408 6848
rect 6043 6817 6055 6820
rect 5997 6811 6055 6817
rect 1857 6783 1915 6789
rect 1857 6749 1869 6783
rect 1903 6749 1915 6783
rect 1857 6743 1915 6749
rect 1486 6644 1492 6656
rect 1447 6616 1492 6644
rect 1486 6604 1492 6616
rect 1544 6604 1550 6656
rect 1872 6644 1900 6743
rect 4890 6740 4896 6792
rect 4948 6780 4954 6792
rect 6181 6783 6239 6789
rect 4948 6752 5764 6780
rect 4948 6740 4954 6752
rect 3142 6672 3148 6724
rect 3200 6712 3206 6724
rect 3881 6715 3939 6721
rect 3881 6712 3893 6715
rect 3200 6684 3893 6712
rect 3200 6672 3206 6684
rect 3881 6681 3893 6684
rect 3927 6681 3939 6715
rect 3881 6675 3939 6681
rect 4522 6672 4528 6724
rect 4580 6712 4586 6724
rect 4801 6715 4859 6721
rect 4801 6712 4813 6715
rect 4580 6684 4813 6712
rect 4580 6672 4586 6684
rect 4801 6681 4813 6684
rect 4847 6712 4859 6715
rect 5537 6715 5595 6721
rect 4847 6684 5488 6712
rect 4847 6681 4859 6684
rect 4801 6675 4859 6681
rect 2958 6644 2964 6656
rect 1872 6616 2964 6644
rect 2958 6604 2964 6616
rect 3016 6604 3022 6656
rect 3234 6644 3240 6656
rect 3195 6616 3240 6644
rect 3234 6604 3240 6616
rect 3292 6604 3298 6656
rect 3697 6647 3755 6653
rect 3697 6613 3709 6647
rect 3743 6644 3755 6647
rect 4246 6644 4252 6656
rect 3743 6616 4252 6644
rect 3743 6613 3755 6616
rect 3697 6607 3755 6613
rect 4246 6604 4252 6616
rect 4304 6604 4310 6656
rect 5258 6644 5264 6656
rect 5219 6616 5264 6644
rect 5258 6604 5264 6616
rect 5316 6604 5322 6656
rect 5460 6644 5488 6684
rect 5537 6681 5549 6715
rect 5583 6712 5595 6715
rect 5626 6712 5632 6724
rect 5583 6684 5632 6712
rect 5583 6681 5595 6684
rect 5537 6675 5595 6681
rect 5626 6672 5632 6684
rect 5684 6672 5690 6724
rect 5736 6712 5764 6752
rect 6181 6749 6193 6783
rect 6227 6780 6239 6783
rect 6270 6780 6276 6792
rect 6227 6752 6276 6780
rect 6227 6749 6239 6752
rect 6181 6743 6239 6749
rect 6270 6740 6276 6752
rect 6328 6740 6334 6792
rect 6380 6780 6408 6820
rect 6549 6817 6561 6851
rect 6595 6848 6607 6851
rect 7760 6848 7788 6956
rect 8202 6944 8208 6956
rect 8260 6944 8266 6996
rect 8941 6987 8999 6993
rect 8941 6953 8953 6987
rect 8987 6984 8999 6987
rect 9030 6984 9036 6996
rect 8987 6956 9036 6984
rect 8987 6953 8999 6956
rect 8941 6947 8999 6953
rect 9030 6944 9036 6956
rect 9088 6944 9094 6996
rect 10410 6944 10416 6996
rect 10468 6984 10474 6996
rect 10597 6987 10655 6993
rect 10597 6984 10609 6987
rect 10468 6956 10609 6984
rect 10468 6944 10474 6956
rect 10597 6953 10609 6956
rect 10643 6953 10655 6987
rect 10597 6947 10655 6953
rect 11330 6944 11336 6996
rect 11388 6984 11394 6996
rect 11388 6956 11551 6984
rect 11388 6944 11394 6956
rect 7926 6876 7932 6928
rect 7984 6876 7990 6928
rect 9048 6916 9076 6944
rect 9370 6919 9428 6925
rect 9370 6916 9382 6919
rect 9048 6888 9382 6916
rect 9370 6885 9382 6888
rect 9416 6885 9428 6919
rect 9370 6879 9428 6885
rect 10686 6876 10692 6928
rect 10744 6916 10750 6928
rect 10965 6919 11023 6925
rect 10965 6916 10977 6919
rect 10744 6888 10977 6916
rect 10744 6876 10750 6888
rect 10965 6885 10977 6888
rect 11011 6885 11023 6919
rect 10965 6879 11023 6885
rect 6595 6820 7788 6848
rect 7828 6851 7886 6857
rect 6595 6817 6607 6820
rect 6549 6811 6607 6817
rect 7828 6817 7840 6851
rect 7874 6848 7886 6851
rect 7944 6848 7972 6876
rect 7874 6820 7972 6848
rect 9125 6851 9183 6857
rect 7874 6817 7886 6820
rect 7828 6811 7886 6817
rect 9125 6817 9137 6851
rect 9171 6848 9183 6851
rect 9674 6848 9680 6860
rect 9171 6820 9680 6848
rect 9171 6817 9183 6820
rect 9125 6811 9183 6817
rect 9674 6808 9680 6820
rect 9732 6848 9738 6860
rect 11523 6848 11551 6956
rect 12526 6944 12532 6996
rect 12584 6984 12590 6996
rect 13541 6987 13599 6993
rect 13541 6984 13553 6987
rect 12584 6956 13553 6984
rect 12584 6944 12590 6956
rect 13541 6953 13553 6956
rect 13587 6953 13599 6987
rect 13541 6947 13599 6953
rect 11865 6851 11923 6857
rect 11865 6848 11877 6851
rect 9732 6820 11468 6848
rect 11523 6820 11877 6848
rect 9732 6808 9738 6820
rect 6380 6752 6776 6780
rect 6748 6724 6776 6752
rect 6914 6740 6920 6792
rect 6972 6780 6978 6792
rect 7466 6780 7472 6792
rect 6972 6752 7328 6780
rect 7427 6752 7472 6780
rect 6972 6740 6978 6752
rect 6365 6715 6423 6721
rect 6365 6712 6377 6715
rect 5736 6684 6377 6712
rect 6365 6681 6377 6684
rect 6411 6681 6423 6715
rect 6730 6712 6736 6724
rect 6691 6684 6736 6712
rect 6365 6675 6423 6681
rect 6730 6672 6736 6684
rect 6788 6672 6794 6724
rect 7300 6712 7328 6752
rect 7466 6740 7472 6752
rect 7524 6740 7530 6792
rect 7561 6783 7619 6789
rect 7561 6749 7573 6783
rect 7607 6749 7619 6783
rect 7561 6743 7619 6749
rect 7576 6712 7604 6743
rect 10226 6740 10232 6792
rect 10284 6780 10290 6792
rect 10284 6752 10640 6780
rect 10284 6740 10290 6752
rect 10502 6712 10508 6724
rect 6840 6684 7144 6712
rect 7300 6684 7604 6712
rect 10463 6684 10508 6712
rect 6840 6644 6868 6684
rect 5460 6616 6868 6644
rect 6917 6647 6975 6653
rect 6917 6613 6929 6647
rect 6963 6644 6975 6647
rect 7006 6644 7012 6656
rect 6963 6616 7012 6644
rect 6963 6613 6975 6616
rect 6917 6607 6975 6613
rect 7006 6604 7012 6616
rect 7064 6604 7070 6656
rect 7116 6644 7144 6684
rect 10502 6672 10508 6684
rect 10560 6672 10566 6724
rect 10612 6712 10640 6752
rect 10686 6740 10692 6792
rect 10744 6780 10750 6792
rect 11057 6783 11115 6789
rect 11057 6780 11069 6783
rect 10744 6752 11069 6780
rect 10744 6740 10750 6752
rect 11057 6749 11069 6752
rect 11103 6749 11115 6783
rect 11057 6743 11115 6749
rect 11241 6783 11299 6789
rect 11241 6749 11253 6783
rect 11287 6780 11299 6783
rect 11330 6780 11336 6792
rect 11287 6752 11336 6780
rect 11287 6749 11299 6752
rect 11241 6743 11299 6749
rect 11330 6740 11336 6752
rect 11388 6740 11394 6792
rect 11440 6780 11468 6820
rect 11865 6817 11877 6820
rect 11911 6817 11923 6851
rect 11865 6811 11923 6817
rect 12710 6808 12716 6860
rect 12768 6848 12774 6860
rect 13449 6851 13507 6857
rect 13449 6848 13461 6851
rect 12768 6820 13461 6848
rect 12768 6808 12774 6820
rect 13449 6817 13461 6820
rect 13495 6817 13507 6851
rect 13449 6811 13507 6817
rect 11609 6783 11667 6789
rect 11609 6780 11621 6783
rect 11440 6752 11621 6780
rect 11609 6749 11621 6752
rect 11655 6749 11667 6783
rect 13633 6783 13691 6789
rect 13633 6780 13645 6783
rect 11609 6743 11667 6749
rect 13004 6752 13645 6780
rect 13004 6721 13032 6752
rect 13633 6749 13645 6752
rect 13679 6749 13691 6783
rect 13633 6743 13691 6749
rect 12989 6715 13047 6721
rect 10612 6684 11551 6712
rect 11238 6644 11244 6656
rect 7116 6616 11244 6644
rect 11238 6604 11244 6616
rect 11296 6604 11302 6656
rect 11422 6644 11428 6656
rect 11383 6616 11428 6644
rect 11422 6604 11428 6616
rect 11480 6604 11486 6656
rect 11523 6644 11551 6684
rect 12989 6681 13001 6715
rect 13035 6681 13047 6715
rect 12989 6675 13047 6681
rect 13004 6644 13032 6675
rect 13078 6672 13084 6724
rect 13136 6712 13142 6724
rect 13136 6684 13181 6712
rect 13136 6672 13142 6684
rect 11523 6616 13032 6644
rect 1104 6554 16008 6576
rect 1104 6502 3480 6554
rect 3532 6502 3544 6554
rect 3596 6502 3608 6554
rect 3660 6502 3672 6554
rect 3724 6502 8478 6554
rect 8530 6502 8542 6554
rect 8594 6502 8606 6554
rect 8658 6502 8670 6554
rect 8722 6502 13475 6554
rect 13527 6502 13539 6554
rect 13591 6502 13603 6554
rect 13655 6502 13667 6554
rect 13719 6502 16008 6554
rect 1104 6480 16008 6502
rect 1854 6400 1860 6452
rect 1912 6440 1918 6452
rect 2682 6440 2688 6452
rect 1912 6412 2688 6440
rect 1912 6400 1918 6412
rect 2682 6400 2688 6412
rect 2740 6440 2746 6452
rect 3237 6443 3295 6449
rect 3237 6440 3249 6443
rect 2740 6412 3249 6440
rect 2740 6400 2746 6412
rect 3237 6409 3249 6412
rect 3283 6409 3295 6443
rect 3237 6403 3295 6409
rect 3326 6400 3332 6452
rect 3384 6440 3390 6452
rect 3605 6443 3663 6449
rect 3605 6440 3617 6443
rect 3384 6412 3617 6440
rect 3384 6400 3390 6412
rect 3605 6409 3617 6412
rect 3651 6409 3663 6443
rect 3605 6403 3663 6409
rect 5258 6400 5264 6452
rect 5316 6440 5322 6452
rect 5534 6440 5540 6452
rect 5316 6412 5540 6440
rect 5316 6400 5322 6412
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 5810 6400 5816 6452
rect 5868 6440 5874 6452
rect 6270 6440 6276 6452
rect 5868 6412 6276 6440
rect 5868 6400 5874 6412
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 7006 6400 7012 6452
rect 7064 6440 7070 6452
rect 8110 6440 8116 6452
rect 7064 6412 8116 6440
rect 7064 6400 7070 6412
rect 8110 6400 8116 6412
rect 8168 6440 8174 6452
rect 8757 6443 8815 6449
rect 8757 6440 8769 6443
rect 8168 6412 8769 6440
rect 8168 6400 8174 6412
rect 8757 6409 8769 6412
rect 8803 6409 8815 6443
rect 9122 6440 9128 6452
rect 9083 6412 9128 6440
rect 8757 6403 8815 6409
rect 9122 6400 9128 6412
rect 9180 6400 9186 6452
rect 9309 6443 9367 6449
rect 9309 6409 9321 6443
rect 9355 6440 9367 6443
rect 10134 6440 10140 6452
rect 9355 6412 10140 6440
rect 9355 6409 9367 6412
rect 9309 6403 9367 6409
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 10594 6440 10600 6452
rect 10555 6412 10600 6440
rect 10594 6400 10600 6412
rect 10652 6400 10658 6452
rect 11606 6400 11612 6452
rect 11664 6440 11670 6452
rect 12529 6443 12587 6449
rect 11664 6412 12103 6440
rect 11664 6400 11670 6412
rect 2958 6332 2964 6384
rect 3016 6372 3022 6384
rect 3789 6375 3847 6381
rect 3789 6372 3801 6375
rect 3016 6344 3801 6372
rect 3016 6332 3022 6344
rect 3789 6341 3801 6344
rect 3835 6341 3847 6375
rect 3789 6335 3847 6341
rect 9398 6332 9404 6384
rect 9456 6372 9462 6384
rect 9582 6372 9588 6384
rect 9456 6344 9588 6372
rect 9456 6332 9462 6344
rect 9582 6332 9588 6344
rect 9640 6372 9646 6384
rect 11974 6372 11980 6384
rect 9640 6344 11980 6372
rect 9640 6332 9646 6344
rect 11974 6332 11980 6344
rect 12032 6332 12038 6384
rect 12075 6372 12103 6412
rect 12529 6409 12541 6443
rect 12575 6440 12587 6443
rect 12710 6440 12716 6452
rect 12575 6412 12716 6440
rect 12575 6409 12587 6412
rect 12529 6403 12587 6409
rect 12710 6400 12716 6412
rect 12768 6400 12774 6452
rect 13081 6443 13139 6449
rect 13081 6409 13093 6443
rect 13127 6440 13139 6443
rect 13354 6440 13360 6452
rect 13127 6412 13360 6440
rect 13127 6409 13139 6412
rect 13081 6403 13139 6409
rect 13354 6400 13360 6412
rect 13412 6440 13418 6452
rect 14090 6440 14096 6452
rect 13412 6412 14096 6440
rect 13412 6400 13418 6412
rect 14090 6400 14096 6412
rect 14148 6400 14154 6452
rect 14277 6443 14335 6449
rect 14277 6409 14289 6443
rect 14323 6440 14335 6443
rect 14550 6440 14556 6452
rect 14323 6412 14556 6440
rect 14323 6409 14335 6412
rect 14277 6403 14335 6409
rect 14550 6400 14556 6412
rect 14608 6400 14614 6452
rect 14734 6400 14740 6452
rect 14792 6440 14798 6452
rect 15197 6443 15255 6449
rect 15197 6440 15209 6443
rect 14792 6412 15209 6440
rect 14792 6400 14798 6412
rect 15197 6409 15209 6412
rect 15243 6409 15255 6443
rect 15197 6403 15255 6409
rect 13173 6375 13231 6381
rect 13173 6372 13185 6375
rect 12075 6344 13185 6372
rect 13173 6341 13185 6344
rect 13219 6341 13231 6375
rect 13173 6335 13231 6341
rect 4338 6304 4344 6316
rect 4299 6276 4344 6304
rect 4338 6264 4344 6276
rect 4396 6264 4402 6316
rect 5166 6304 5172 6316
rect 5127 6276 5172 6304
rect 5166 6264 5172 6276
rect 5224 6264 5230 6316
rect 5258 6264 5264 6316
rect 5316 6304 5322 6316
rect 5353 6307 5411 6313
rect 5353 6304 5365 6307
rect 5316 6276 5365 6304
rect 5316 6264 5322 6276
rect 5353 6273 5365 6276
rect 5399 6304 5411 6307
rect 6089 6307 6147 6313
rect 6089 6304 6101 6307
rect 5399 6276 6101 6304
rect 5399 6273 5411 6276
rect 5353 6267 5411 6273
rect 6089 6273 6101 6276
rect 6135 6273 6147 6307
rect 6546 6304 6552 6316
rect 6459 6276 6552 6304
rect 6089 6267 6147 6273
rect 6546 6264 6552 6276
rect 6604 6304 6610 6316
rect 6641 6307 6699 6313
rect 6641 6304 6653 6307
rect 6604 6276 6653 6304
rect 6604 6264 6610 6276
rect 6641 6273 6653 6276
rect 6687 6304 6699 6307
rect 6914 6304 6920 6316
rect 6687 6276 6920 6304
rect 6687 6273 6699 6276
rect 6641 6267 6699 6273
rect 6914 6264 6920 6276
rect 6972 6264 6978 6316
rect 8297 6307 8355 6313
rect 8297 6273 8309 6307
rect 8343 6304 8355 6307
rect 9674 6304 9680 6316
rect 8343 6276 9680 6304
rect 8343 6273 8355 6276
rect 8297 6267 8355 6273
rect 9674 6264 9680 6276
rect 9732 6264 9738 6316
rect 9953 6307 10011 6313
rect 9953 6273 9965 6307
rect 9999 6304 10011 6307
rect 10502 6304 10508 6316
rect 9999 6276 10508 6304
rect 9999 6273 10011 6276
rect 9953 6267 10011 6273
rect 10502 6264 10508 6276
rect 10560 6264 10566 6316
rect 11241 6307 11299 6313
rect 11241 6273 11253 6307
rect 11287 6304 11299 6307
rect 11330 6304 11336 6316
rect 11287 6276 11336 6304
rect 11287 6273 11299 6276
rect 11241 6267 11299 6273
rect 11330 6264 11336 6276
rect 11388 6304 11394 6316
rect 11885 6307 11943 6313
rect 11885 6304 11897 6307
rect 11388 6276 11897 6304
rect 11388 6264 11394 6276
rect 11885 6273 11897 6276
rect 11931 6273 11943 6307
rect 11885 6267 11943 6273
rect 13262 6264 13268 6316
rect 13320 6304 13326 6316
rect 13357 6307 13415 6313
rect 13357 6304 13369 6307
rect 13320 6276 13369 6304
rect 13320 6264 13326 6276
rect 13357 6273 13369 6276
rect 13403 6273 13415 6307
rect 13357 6267 13415 6273
rect 2961 6239 3019 6245
rect 2961 6205 2973 6239
rect 3007 6236 3019 6239
rect 3326 6236 3332 6248
rect 3007 6208 3332 6236
rect 3007 6205 3019 6208
rect 2961 6199 3019 6205
rect 3326 6196 3332 6208
rect 3384 6196 3390 6248
rect 5077 6239 5135 6245
rect 5077 6205 5089 6239
rect 5123 6236 5135 6239
rect 5123 6208 5764 6236
rect 5123 6205 5135 6208
rect 5077 6199 5135 6205
rect 1489 6171 1547 6177
rect 1489 6137 1501 6171
rect 1535 6168 1547 6171
rect 2222 6168 2228 6180
rect 1535 6140 2228 6168
rect 1535 6137 1547 6140
rect 1489 6131 1547 6137
rect 2222 6128 2228 6140
rect 2280 6128 2286 6180
rect 2682 6168 2688 6180
rect 2740 6177 2746 6180
rect 2652 6140 2688 6168
rect 2682 6128 2688 6140
rect 2740 6131 2752 6177
rect 4157 6171 4215 6177
rect 4157 6137 4169 6171
rect 4203 6168 4215 6171
rect 5736 6168 5764 6208
rect 5810 6196 5816 6248
rect 5868 6236 5874 6248
rect 5997 6239 6055 6245
rect 5997 6236 6009 6239
rect 5868 6208 6009 6236
rect 5868 6196 5874 6208
rect 5997 6205 6009 6208
rect 6043 6236 6055 6239
rect 7006 6236 7012 6248
rect 6043 6208 7012 6236
rect 6043 6205 6055 6208
rect 5997 6199 6055 6205
rect 7006 6196 7012 6208
rect 7064 6196 7070 6248
rect 9401 6239 9459 6245
rect 9401 6205 9413 6239
rect 9447 6205 9459 6239
rect 9401 6199 9459 6205
rect 6641 6171 6699 6177
rect 6641 6168 6653 6171
rect 4203 6140 5580 6168
rect 5736 6140 6653 6168
rect 4203 6137 4215 6140
rect 4157 6131 4215 6137
rect 2740 6128 2746 6131
rect 1578 6100 1584 6112
rect 1539 6072 1584 6100
rect 1578 6060 1584 6072
rect 1636 6100 1642 6112
rect 1946 6100 1952 6112
rect 1636 6072 1952 6100
rect 1636 6060 1642 6072
rect 1946 6060 1952 6072
rect 2004 6060 2010 6112
rect 2240 6100 2268 6128
rect 3053 6103 3111 6109
rect 3053 6100 3065 6103
rect 2240 6072 3065 6100
rect 3053 6069 3065 6072
rect 3099 6069 3111 6103
rect 3053 6063 3111 6069
rect 3142 6060 3148 6112
rect 3200 6100 3206 6112
rect 5552 6109 5580 6140
rect 6641 6137 6653 6140
rect 6687 6137 6699 6171
rect 6641 6131 6699 6137
rect 6733 6171 6791 6177
rect 6733 6137 6745 6171
rect 6779 6168 6791 6171
rect 7282 6168 7288 6180
rect 6779 6140 7288 6168
rect 6779 6137 6791 6140
rect 6733 6131 6791 6137
rect 7282 6128 7288 6140
rect 7340 6168 7346 6180
rect 7742 6168 7748 6180
rect 7340 6140 7748 6168
rect 7340 6128 7346 6140
rect 7742 6128 7748 6140
rect 7800 6128 7806 6180
rect 8018 6128 8024 6180
rect 8076 6177 8082 6180
rect 8076 6168 8088 6177
rect 8076 6140 8121 6168
rect 8076 6131 8088 6140
rect 8076 6128 8082 6131
rect 8202 6128 8208 6180
rect 8260 6168 8266 6180
rect 9416 6168 9444 6199
rect 9858 6196 9864 6248
rect 9916 6236 9922 6248
rect 10137 6239 10195 6245
rect 10137 6236 10149 6239
rect 9916 6208 10149 6236
rect 9916 6196 9922 6208
rect 10137 6205 10149 6208
rect 10183 6236 10195 6239
rect 10318 6236 10324 6248
rect 10183 6208 10324 6236
rect 10183 6205 10195 6208
rect 10137 6199 10195 6205
rect 10318 6196 10324 6208
rect 10376 6196 10382 6248
rect 10594 6196 10600 6248
rect 10652 6236 10658 6248
rect 11057 6239 11115 6245
rect 11057 6236 11069 6239
rect 10652 6208 11069 6236
rect 10652 6196 10658 6208
rect 11057 6205 11069 6208
rect 11103 6236 11115 6239
rect 11606 6236 11612 6248
rect 11103 6208 11612 6236
rect 11103 6205 11115 6208
rect 11057 6199 11115 6205
rect 11606 6196 11612 6208
rect 11664 6196 11670 6248
rect 12618 6236 12624 6248
rect 11992 6208 12624 6236
rect 11992 6168 12020 6208
rect 12618 6196 12624 6208
rect 12676 6236 12682 6248
rect 13280 6236 13308 6264
rect 12676 6208 13308 6236
rect 12676 6196 12682 6208
rect 8260 6140 9444 6168
rect 9508 6140 12020 6168
rect 12161 6171 12219 6177
rect 8260 6128 8266 6140
rect 3421 6103 3479 6109
rect 3421 6100 3433 6103
rect 3200 6072 3433 6100
rect 3200 6060 3206 6072
rect 3421 6069 3433 6072
rect 3467 6069 3479 6103
rect 3421 6063 3479 6069
rect 4249 6103 4307 6109
rect 4249 6069 4261 6103
rect 4295 6100 4307 6103
rect 4709 6103 4767 6109
rect 4709 6100 4721 6103
rect 4295 6072 4721 6100
rect 4295 6069 4307 6072
rect 4249 6063 4307 6069
rect 4709 6069 4721 6072
rect 4755 6069 4767 6103
rect 4709 6063 4767 6069
rect 5537 6103 5595 6109
rect 5537 6069 5549 6103
rect 5583 6069 5595 6103
rect 5537 6063 5595 6069
rect 5626 6060 5632 6112
rect 5684 6100 5690 6112
rect 5905 6103 5963 6109
rect 5905 6100 5917 6103
rect 5684 6072 5917 6100
rect 5684 6060 5690 6072
rect 5905 6069 5917 6072
rect 5951 6069 5963 6103
rect 5905 6063 5963 6069
rect 6822 6060 6828 6112
rect 6880 6100 6886 6112
rect 6917 6103 6975 6109
rect 6917 6100 6929 6103
rect 6880 6072 6929 6100
rect 6880 6060 6886 6072
rect 6917 6069 6929 6072
rect 6963 6069 6975 6103
rect 6917 6063 6975 6069
rect 7374 6060 7380 6112
rect 7432 6100 7438 6112
rect 7650 6100 7656 6112
rect 7432 6072 7656 6100
rect 7432 6060 7438 6072
rect 7650 6060 7656 6072
rect 7708 6100 7714 6112
rect 8389 6103 8447 6109
rect 8389 6100 8401 6103
rect 7708 6072 8401 6100
rect 7708 6060 7714 6072
rect 8389 6069 8401 6072
rect 8435 6069 8447 6103
rect 8389 6063 8447 6069
rect 8665 6103 8723 6109
rect 8665 6069 8677 6103
rect 8711 6100 8723 6103
rect 9030 6100 9036 6112
rect 8711 6072 9036 6100
rect 8711 6069 8723 6072
rect 8665 6063 8723 6069
rect 9030 6060 9036 6072
rect 9088 6060 9094 6112
rect 9306 6060 9312 6112
rect 9364 6100 9370 6112
rect 9508 6100 9536 6140
rect 12161 6137 12173 6171
rect 12207 6168 12219 6171
rect 12342 6168 12348 6180
rect 12207 6140 12348 6168
rect 12207 6137 12219 6140
rect 12161 6131 12219 6137
rect 12342 6128 12348 6140
rect 12400 6128 12406 6180
rect 9364 6072 9536 6100
rect 9585 6103 9643 6109
rect 9364 6060 9370 6072
rect 9585 6069 9597 6103
rect 9631 6100 9643 6103
rect 9766 6100 9772 6112
rect 9631 6072 9772 6100
rect 9631 6069 9643 6072
rect 9585 6063 9643 6069
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 10045 6103 10103 6109
rect 10045 6069 10057 6103
rect 10091 6100 10103 6103
rect 10134 6100 10140 6112
rect 10091 6072 10140 6100
rect 10091 6069 10103 6072
rect 10045 6063 10103 6069
rect 10134 6060 10140 6072
rect 10192 6060 10198 6112
rect 10505 6103 10563 6109
rect 10505 6069 10517 6103
rect 10551 6100 10563 6103
rect 10686 6100 10692 6112
rect 10551 6072 10692 6100
rect 10551 6069 10563 6072
rect 10505 6063 10563 6069
rect 10686 6060 10692 6072
rect 10744 6060 10750 6112
rect 10870 6060 10876 6112
rect 10928 6100 10934 6112
rect 10965 6103 11023 6109
rect 10965 6100 10977 6103
rect 10928 6072 10977 6100
rect 10928 6060 10934 6072
rect 10965 6069 10977 6072
rect 11011 6100 11023 6103
rect 11425 6103 11483 6109
rect 11425 6100 11437 6103
rect 11011 6072 11437 6100
rect 11011 6069 11023 6072
rect 10965 6063 11023 6069
rect 11425 6069 11437 6072
rect 11471 6069 11483 6103
rect 11425 6063 11483 6069
rect 11790 6060 11796 6112
rect 11848 6100 11854 6112
rect 12069 6103 12127 6109
rect 12069 6100 12081 6103
rect 11848 6072 12081 6100
rect 11848 6060 11854 6072
rect 12069 6069 12081 6072
rect 12115 6100 12127 6103
rect 12621 6103 12679 6109
rect 12621 6100 12633 6103
rect 12115 6072 12633 6100
rect 12115 6069 12127 6072
rect 12069 6063 12127 6069
rect 12621 6069 12633 6072
rect 12667 6100 12679 6103
rect 12805 6103 12863 6109
rect 12805 6100 12817 6103
rect 12667 6072 12817 6100
rect 12667 6069 12679 6072
rect 12621 6063 12679 6069
rect 12805 6069 12817 6072
rect 12851 6069 12863 6103
rect 15378 6100 15384 6112
rect 15339 6072 15384 6100
rect 12805 6063 12863 6069
rect 15378 6060 15384 6072
rect 15436 6060 15442 6112
rect 1104 6010 16008 6032
rect 1104 5958 5979 6010
rect 6031 5958 6043 6010
rect 6095 5958 6107 6010
rect 6159 5958 6171 6010
rect 6223 5958 10976 6010
rect 11028 5958 11040 6010
rect 11092 5958 11104 6010
rect 11156 5958 11168 6010
rect 11220 5958 16008 6010
rect 1104 5936 16008 5958
rect 1762 5896 1768 5908
rect 1723 5868 1768 5896
rect 1762 5856 1768 5868
rect 1820 5856 1826 5908
rect 2501 5899 2559 5905
rect 2501 5865 2513 5899
rect 2547 5896 2559 5899
rect 2961 5899 3019 5905
rect 2961 5896 2973 5899
rect 2547 5868 2973 5896
rect 2547 5865 2559 5868
rect 2501 5859 2559 5865
rect 2961 5865 2973 5868
rect 3007 5865 3019 5899
rect 2961 5859 3019 5865
rect 3421 5899 3479 5905
rect 3421 5865 3433 5899
rect 3467 5896 3479 5899
rect 3881 5899 3939 5905
rect 3881 5896 3893 5899
rect 3467 5868 3893 5896
rect 3467 5865 3479 5868
rect 3421 5859 3479 5865
rect 3881 5865 3893 5868
rect 3927 5865 3939 5899
rect 4246 5896 4252 5908
rect 4159 5868 4252 5896
rect 3881 5859 3939 5865
rect 4246 5856 4252 5868
rect 4304 5896 4310 5908
rect 5169 5899 5227 5905
rect 4304 5868 5120 5896
rect 4304 5856 4310 5868
rect 1578 5788 1584 5840
rect 1636 5828 1642 5840
rect 4338 5828 4344 5840
rect 1636 5800 4344 5828
rect 1636 5788 1642 5800
rect 1673 5763 1731 5769
rect 1673 5729 1685 5763
rect 1719 5729 1731 5763
rect 1673 5723 1731 5729
rect 1949 5763 2007 5769
rect 1949 5729 1961 5763
rect 1995 5760 2007 5763
rect 2130 5760 2136 5772
rect 1995 5732 2136 5760
rect 1995 5729 2007 5732
rect 1949 5723 2007 5729
rect 1688 5624 1716 5723
rect 2130 5720 2136 5732
rect 2188 5720 2194 5772
rect 2240 5701 2268 5800
rect 4338 5788 4344 5800
rect 4396 5788 4402 5840
rect 5092 5828 5120 5868
rect 5169 5865 5181 5899
rect 5215 5896 5227 5899
rect 5626 5896 5632 5908
rect 5215 5868 5632 5896
rect 5215 5865 5227 5868
rect 5169 5859 5227 5865
rect 5626 5856 5632 5868
rect 5684 5856 5690 5908
rect 5736 5868 6960 5896
rect 5736 5828 5764 5868
rect 5092 5800 5764 5828
rect 6396 5831 6454 5837
rect 6396 5797 6408 5831
rect 6442 5828 6454 5831
rect 6822 5828 6828 5840
rect 6442 5800 6828 5828
rect 6442 5797 6454 5800
rect 6396 5791 6454 5797
rect 6822 5788 6828 5800
rect 6880 5788 6886 5840
rect 6932 5828 6960 5868
rect 7466 5856 7472 5908
rect 7524 5896 7530 5908
rect 8113 5899 8171 5905
rect 8113 5896 8125 5899
rect 7524 5868 8125 5896
rect 7524 5856 7530 5868
rect 8113 5865 8125 5868
rect 8159 5865 8171 5899
rect 8113 5859 8171 5865
rect 9582 5856 9588 5908
rect 9640 5896 9646 5908
rect 9769 5899 9827 5905
rect 9640 5856 9674 5896
rect 9769 5865 9781 5899
rect 9815 5896 9827 5899
rect 9858 5896 9864 5908
rect 9815 5868 9864 5896
rect 9815 5865 9827 5868
rect 9769 5859 9827 5865
rect 9858 5856 9864 5868
rect 9916 5856 9922 5908
rect 11425 5899 11483 5905
rect 11425 5865 11437 5899
rect 11471 5896 11483 5899
rect 11698 5896 11704 5908
rect 11471 5868 11704 5896
rect 11471 5865 11483 5868
rect 11425 5859 11483 5865
rect 11698 5856 11704 5868
rect 11756 5856 11762 5908
rect 11793 5899 11851 5905
rect 11793 5865 11805 5899
rect 11839 5896 11851 5899
rect 12250 5896 12256 5908
rect 11839 5868 12256 5896
rect 11839 5865 11851 5868
rect 11793 5859 11851 5865
rect 12250 5856 12256 5868
rect 12308 5856 12314 5908
rect 12342 5856 12348 5908
rect 12400 5896 12406 5908
rect 12621 5899 12679 5905
rect 12621 5896 12633 5899
rect 12400 5868 12633 5896
rect 12400 5856 12406 5868
rect 12621 5865 12633 5868
rect 12667 5896 12679 5899
rect 12894 5896 12900 5908
rect 12667 5868 12900 5896
rect 12667 5865 12679 5868
rect 12621 5859 12679 5865
rect 12894 5856 12900 5868
rect 12952 5856 12958 5908
rect 14921 5899 14979 5905
rect 14921 5865 14933 5899
rect 14967 5896 14979 5899
rect 15746 5896 15752 5908
rect 14967 5868 15752 5896
rect 14967 5865 14979 5868
rect 14921 5859 14979 5865
rect 15746 5856 15752 5868
rect 15804 5856 15810 5908
rect 9306 5828 9312 5840
rect 6932 5800 9312 5828
rect 9306 5788 9312 5800
rect 9364 5788 9370 5840
rect 3329 5763 3387 5769
rect 3329 5729 3341 5763
rect 3375 5760 3387 5763
rect 3418 5760 3424 5772
rect 3375 5732 3424 5760
rect 3375 5729 3387 5732
rect 3329 5723 3387 5729
rect 3418 5720 3424 5732
rect 3476 5720 3482 5772
rect 4522 5760 4528 5772
rect 4356 5732 4528 5760
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5661 2283 5695
rect 2406 5692 2412 5704
rect 2367 5664 2412 5692
rect 2225 5655 2283 5661
rect 2406 5652 2412 5664
rect 2464 5652 2470 5704
rect 2682 5652 2688 5704
rect 2740 5692 2746 5704
rect 3605 5695 3663 5701
rect 3605 5692 3617 5695
rect 2740 5664 3617 5692
rect 2740 5652 2746 5664
rect 3605 5661 3617 5664
rect 3651 5692 3663 5695
rect 4154 5692 4160 5704
rect 3651 5664 4160 5692
rect 3651 5661 3663 5664
rect 3605 5655 3663 5661
rect 4154 5652 4160 5664
rect 4212 5652 4218 5704
rect 4356 5701 4384 5732
rect 4522 5720 4528 5732
rect 4580 5720 4586 5772
rect 4890 5760 4896 5772
rect 4851 5732 4896 5760
rect 4890 5720 4896 5732
rect 4948 5720 4954 5772
rect 6641 5763 6699 5769
rect 6641 5760 6653 5763
rect 5000 5732 6653 5760
rect 4341 5695 4399 5701
rect 4341 5661 4353 5695
rect 4387 5661 4399 5695
rect 4341 5655 4399 5661
rect 4433 5695 4491 5701
rect 4433 5661 4445 5695
rect 4479 5661 4491 5695
rect 5000 5692 5028 5732
rect 6641 5729 6653 5732
rect 6687 5729 6699 5763
rect 6641 5723 6699 5729
rect 6914 5720 6920 5772
rect 6972 5760 6978 5772
rect 7285 5763 7343 5769
rect 7285 5760 7297 5763
rect 6972 5732 7297 5760
rect 6972 5720 6978 5732
rect 7285 5729 7297 5732
rect 7331 5760 7343 5763
rect 7466 5760 7472 5772
rect 7331 5732 7472 5760
rect 7331 5729 7343 5732
rect 7285 5723 7343 5729
rect 7466 5720 7472 5732
rect 7524 5720 7530 5772
rect 8110 5720 8116 5772
rect 8168 5760 8174 5772
rect 8205 5763 8263 5769
rect 8205 5760 8217 5763
rect 8168 5732 8217 5760
rect 8168 5720 8174 5732
rect 8205 5729 8217 5732
rect 8251 5729 8263 5763
rect 8205 5723 8263 5729
rect 8757 5763 8815 5769
rect 8757 5729 8769 5763
rect 8803 5760 8815 5763
rect 8938 5760 8944 5772
rect 8803 5732 8944 5760
rect 8803 5729 8815 5732
rect 8757 5723 8815 5729
rect 8938 5720 8944 5732
rect 8996 5720 9002 5772
rect 9646 5760 9674 5856
rect 10229 5831 10287 5837
rect 10229 5797 10241 5831
rect 10275 5797 10287 5831
rect 10229 5791 10287 5797
rect 9766 5760 9772 5772
rect 9646 5732 9772 5760
rect 9766 5720 9772 5732
rect 9824 5720 9830 5772
rect 10137 5763 10195 5769
rect 10137 5729 10149 5763
rect 10183 5729 10195 5763
rect 10137 5723 10195 5729
rect 4433 5655 4491 5661
rect 4724 5664 5028 5692
rect 3878 5624 3884 5636
rect 1688 5596 3884 5624
rect 3878 5584 3884 5596
rect 3936 5584 3942 5636
rect 4448 5624 4476 5655
rect 4522 5624 4528 5636
rect 4448 5596 4528 5624
rect 4522 5584 4528 5596
rect 4580 5584 4586 5636
rect 1486 5556 1492 5568
rect 1447 5528 1492 5556
rect 1486 5516 1492 5528
rect 1544 5516 1550 5568
rect 2866 5556 2872 5568
rect 2827 5528 2872 5556
rect 2866 5516 2872 5528
rect 2924 5516 2930 5568
rect 3326 5516 3332 5568
rect 3384 5556 3390 5568
rect 4724 5565 4752 5664
rect 6730 5652 6736 5704
rect 6788 5692 6794 5704
rect 7377 5695 7435 5701
rect 7377 5692 7389 5695
rect 6788 5664 7389 5692
rect 6788 5652 6794 5664
rect 7377 5661 7389 5664
rect 7423 5661 7435 5695
rect 7377 5655 7435 5661
rect 7561 5695 7619 5701
rect 7561 5661 7573 5695
rect 7607 5692 7619 5695
rect 8018 5692 8024 5704
rect 7607 5664 8024 5692
rect 7607 5661 7619 5664
rect 7561 5655 7619 5661
rect 8018 5652 8024 5664
rect 8076 5692 8082 5704
rect 8297 5695 8355 5701
rect 8297 5692 8309 5695
rect 8076 5664 8309 5692
rect 8076 5652 8082 5664
rect 8297 5661 8309 5664
rect 8343 5661 8355 5695
rect 8297 5655 8355 5661
rect 9324 5664 9904 5692
rect 7006 5584 7012 5636
rect 7064 5624 7070 5636
rect 8573 5627 8631 5633
rect 8573 5624 8585 5627
rect 7064 5596 8585 5624
rect 7064 5584 7070 5596
rect 8573 5593 8585 5596
rect 8619 5593 8631 5627
rect 8573 5587 8631 5593
rect 8846 5584 8852 5636
rect 8904 5624 8910 5636
rect 9125 5627 9183 5633
rect 9125 5624 9137 5627
rect 8904 5596 9137 5624
rect 8904 5584 8910 5596
rect 9125 5593 9137 5596
rect 9171 5624 9183 5627
rect 9214 5624 9220 5636
rect 9171 5596 9220 5624
rect 9171 5593 9183 5596
rect 9125 5587 9183 5593
rect 9214 5584 9220 5596
rect 9272 5584 9278 5636
rect 9324 5568 9352 5664
rect 9398 5584 9404 5636
rect 9456 5624 9462 5636
rect 9456 5596 9812 5624
rect 9456 5584 9462 5596
rect 9784 5568 9812 5596
rect 4709 5559 4767 5565
rect 4709 5556 4721 5559
rect 3384 5528 4721 5556
rect 3384 5516 3390 5528
rect 4709 5525 4721 5528
rect 4755 5525 4767 5559
rect 4709 5519 4767 5525
rect 5261 5559 5319 5565
rect 5261 5525 5273 5559
rect 5307 5556 5319 5559
rect 5994 5556 6000 5568
rect 5307 5528 6000 5556
rect 5307 5525 5319 5528
rect 5261 5519 5319 5525
rect 5994 5516 6000 5528
rect 6052 5516 6058 5568
rect 6362 5516 6368 5568
rect 6420 5556 6426 5568
rect 6638 5556 6644 5568
rect 6420 5528 6644 5556
rect 6420 5516 6426 5528
rect 6638 5516 6644 5528
rect 6696 5556 6702 5568
rect 6733 5559 6791 5565
rect 6733 5556 6745 5559
rect 6696 5528 6745 5556
rect 6696 5516 6702 5528
rect 6733 5525 6745 5528
rect 6779 5525 6791 5559
rect 6914 5556 6920 5568
rect 6875 5528 6920 5556
rect 6733 5519 6791 5525
rect 6914 5516 6920 5528
rect 6972 5516 6978 5568
rect 7742 5556 7748 5568
rect 7703 5528 7748 5556
rect 7742 5516 7748 5528
rect 7800 5516 7806 5568
rect 8938 5556 8944 5568
rect 8899 5528 8944 5556
rect 8938 5516 8944 5528
rect 8996 5516 9002 5568
rect 9306 5556 9312 5568
rect 9267 5528 9312 5556
rect 9306 5516 9312 5528
rect 9364 5516 9370 5568
rect 9582 5556 9588 5568
rect 9543 5528 9588 5556
rect 9582 5516 9588 5528
rect 9640 5516 9646 5568
rect 9766 5516 9772 5568
rect 9824 5516 9830 5568
rect 9876 5556 9904 5664
rect 10152 5636 10180 5723
rect 10244 5692 10272 5791
rect 10318 5788 10324 5840
rect 10376 5828 10382 5840
rect 11149 5831 11207 5837
rect 11149 5828 11161 5831
rect 10376 5800 11161 5828
rect 10376 5788 10382 5800
rect 11149 5797 11161 5800
rect 11195 5797 11207 5831
rect 11149 5791 11207 5797
rect 11517 5831 11575 5837
rect 11517 5797 11529 5831
rect 11563 5828 11575 5831
rect 12802 5828 12808 5840
rect 11563 5800 12808 5828
rect 11563 5797 11575 5800
rect 11517 5791 11575 5797
rect 10235 5664 10272 5692
rect 10235 5636 10263 5664
rect 10318 5652 10324 5704
rect 10376 5692 10382 5704
rect 10376 5664 10421 5692
rect 10376 5652 10382 5664
rect 10134 5584 10140 5636
rect 10192 5584 10198 5636
rect 10226 5584 10232 5636
rect 10284 5584 10290 5636
rect 11532 5624 11560 5791
rect 12802 5788 12808 5800
rect 12860 5788 12866 5840
rect 14366 5828 14372 5840
rect 13004 5800 14372 5828
rect 11606 5720 11612 5772
rect 11664 5760 11670 5772
rect 12069 5763 12127 5769
rect 12069 5760 12081 5763
rect 11664 5732 12081 5760
rect 11664 5720 11670 5732
rect 12069 5729 12081 5732
rect 12115 5729 12127 5763
rect 13004 5760 13032 5800
rect 14366 5788 14372 5800
rect 14424 5788 14430 5840
rect 15654 5828 15660 5840
rect 15615 5800 15660 5828
rect 15654 5788 15660 5800
rect 15712 5788 15718 5840
rect 13354 5760 13360 5772
rect 12069 5723 12127 5729
rect 12360 5732 13032 5760
rect 13315 5732 13360 5760
rect 11974 5652 11980 5704
rect 12032 5692 12038 5704
rect 12360 5692 12388 5732
rect 13354 5720 13360 5732
rect 13412 5720 13418 5772
rect 14642 5720 14648 5772
rect 14700 5760 14706 5772
rect 14737 5763 14795 5769
rect 14737 5760 14749 5763
rect 14700 5732 14749 5760
rect 14700 5720 14706 5732
rect 14737 5729 14749 5732
rect 14783 5760 14795 5763
rect 14918 5760 14924 5772
rect 14783 5732 14924 5760
rect 14783 5729 14795 5732
rect 14737 5723 14795 5729
rect 14918 5720 14924 5732
rect 14976 5720 14982 5772
rect 15470 5760 15476 5772
rect 15431 5732 15476 5760
rect 15470 5720 15476 5732
rect 15528 5720 15534 5772
rect 12032 5664 12388 5692
rect 12032 5652 12038 5664
rect 12434 5652 12440 5704
rect 12492 5692 12498 5704
rect 12802 5692 12808 5704
rect 12492 5664 12808 5692
rect 12492 5652 12498 5664
rect 12802 5652 12808 5664
rect 12860 5652 12866 5704
rect 13081 5695 13139 5701
rect 13081 5661 13093 5695
rect 13127 5661 13139 5695
rect 13262 5692 13268 5704
rect 13223 5664 13268 5692
rect 13081 5655 13139 5661
rect 10336 5596 11560 5624
rect 13096 5624 13124 5655
rect 13262 5652 13268 5664
rect 13320 5652 13326 5704
rect 15105 5695 15163 5701
rect 15105 5661 15117 5695
rect 15151 5692 15163 5695
rect 15562 5692 15568 5704
rect 15151 5664 15568 5692
rect 15151 5661 15163 5664
rect 15105 5655 15163 5661
rect 15562 5652 15568 5664
rect 15620 5652 15626 5704
rect 13170 5624 13176 5636
rect 13096 5596 13176 5624
rect 10336 5556 10364 5596
rect 13170 5584 13176 5596
rect 13228 5584 13234 5636
rect 13725 5627 13783 5633
rect 13725 5593 13737 5627
rect 13771 5624 13783 5627
rect 15286 5624 15292 5636
rect 13771 5596 15292 5624
rect 13771 5593 13783 5596
rect 13725 5587 13783 5593
rect 15286 5584 15292 5596
rect 15344 5584 15350 5636
rect 10594 5556 10600 5568
rect 9876 5528 10364 5556
rect 10555 5528 10600 5556
rect 10594 5516 10600 5528
rect 10652 5516 10658 5568
rect 10873 5559 10931 5565
rect 10873 5525 10885 5559
rect 10919 5556 10931 5559
rect 10962 5556 10968 5568
rect 10919 5528 10968 5556
rect 10919 5525 10931 5528
rect 10873 5519 10931 5525
rect 10962 5516 10968 5528
rect 11020 5516 11026 5568
rect 11057 5559 11115 5565
rect 11057 5525 11069 5559
rect 11103 5556 11115 5559
rect 11330 5556 11336 5568
rect 11103 5528 11336 5556
rect 11103 5525 11115 5528
rect 11057 5519 11115 5525
rect 11330 5516 11336 5528
rect 11388 5556 11394 5568
rect 11514 5556 11520 5568
rect 11388 5528 11520 5556
rect 11388 5516 11394 5528
rect 11514 5516 11520 5528
rect 11572 5516 11578 5568
rect 11974 5556 11980 5568
rect 11935 5528 11980 5556
rect 11974 5516 11980 5528
rect 12032 5516 12038 5568
rect 12158 5516 12164 5568
rect 12216 5556 12222 5568
rect 12805 5559 12863 5565
rect 12805 5556 12817 5559
rect 12216 5528 12817 5556
rect 12216 5516 12222 5528
rect 12805 5525 12817 5528
rect 12851 5525 12863 5559
rect 13814 5556 13820 5568
rect 13775 5528 13820 5556
rect 12805 5519 12863 5525
rect 13814 5516 13820 5528
rect 13872 5516 13878 5568
rect 13906 5516 13912 5568
rect 13964 5556 13970 5568
rect 14001 5559 14059 5565
rect 14001 5556 14013 5559
rect 13964 5528 14013 5556
rect 13964 5516 13970 5528
rect 14001 5525 14013 5528
rect 14047 5525 14059 5559
rect 15194 5556 15200 5568
rect 15155 5528 15200 5556
rect 14001 5519 14059 5525
rect 15194 5516 15200 5528
rect 15252 5516 15258 5568
rect 1104 5466 16008 5488
rect 1104 5414 3480 5466
rect 3532 5414 3544 5466
rect 3596 5414 3608 5466
rect 3660 5414 3672 5466
rect 3724 5414 8478 5466
rect 8530 5414 8542 5466
rect 8594 5414 8606 5466
rect 8658 5414 8670 5466
rect 8722 5414 13475 5466
rect 13527 5414 13539 5466
rect 13591 5414 13603 5466
rect 13655 5414 13667 5466
rect 13719 5414 16008 5466
rect 1104 5392 16008 5414
rect 2406 5312 2412 5364
rect 2464 5352 2470 5364
rect 2501 5355 2559 5361
rect 2501 5352 2513 5355
rect 2464 5324 2513 5352
rect 2464 5312 2470 5324
rect 2501 5321 2513 5324
rect 2547 5321 2559 5355
rect 2501 5315 2559 5321
rect 4154 5312 4160 5364
rect 4212 5352 4218 5364
rect 5258 5352 5264 5364
rect 4212 5324 5264 5352
rect 4212 5312 4218 5324
rect 5258 5312 5264 5324
rect 5316 5312 5322 5364
rect 6457 5355 6515 5361
rect 6457 5321 6469 5355
rect 6503 5352 6515 5355
rect 6546 5352 6552 5364
rect 6503 5324 6552 5352
rect 6503 5321 6515 5324
rect 6457 5315 6515 5321
rect 6546 5312 6552 5324
rect 6604 5312 6610 5364
rect 6822 5312 6828 5364
rect 6880 5352 6886 5364
rect 6880 5324 7420 5352
rect 6880 5312 6886 5324
rect 1394 5284 1400 5296
rect 1355 5256 1400 5284
rect 1394 5244 1400 5256
rect 1452 5244 1458 5296
rect 2130 5244 2136 5296
rect 2188 5284 2194 5296
rect 2593 5287 2651 5293
rect 2593 5284 2605 5287
rect 2188 5256 2605 5284
rect 2188 5244 2194 5256
rect 2593 5253 2605 5256
rect 2639 5253 2651 5287
rect 7285 5287 7343 5293
rect 7285 5284 7297 5287
rect 2593 5247 2651 5253
rect 6012 5256 7297 5284
rect 1949 5219 2007 5225
rect 1949 5185 1961 5219
rect 1995 5216 2007 5219
rect 2682 5216 2688 5228
rect 1995 5188 2688 5216
rect 1995 5185 2007 5188
rect 1949 5179 2007 5185
rect 2682 5176 2688 5188
rect 2740 5176 2746 5228
rect 2866 5176 2872 5228
rect 2924 5216 2930 5228
rect 3053 5219 3111 5225
rect 3053 5216 3065 5219
rect 2924 5188 3065 5216
rect 2924 5176 2930 5188
rect 3053 5185 3065 5188
rect 3099 5185 3111 5219
rect 3234 5216 3240 5228
rect 3195 5188 3240 5216
rect 3053 5179 3111 5185
rect 3234 5176 3240 5188
rect 3292 5176 3298 5228
rect 3326 5176 3332 5228
rect 3384 5216 3390 5228
rect 6012 5225 6040 5256
rect 7285 5253 7297 5256
rect 7331 5253 7343 5287
rect 7285 5247 7343 5253
rect 5997 5219 6055 5225
rect 3384 5188 3832 5216
rect 3384 5176 3390 5188
rect 1486 5108 1492 5160
rect 1544 5148 1550 5160
rect 1581 5151 1639 5157
rect 1581 5148 1593 5151
rect 1544 5120 1593 5148
rect 1544 5108 1550 5120
rect 1581 5117 1593 5120
rect 1627 5117 1639 5151
rect 2958 5148 2964 5160
rect 2919 5120 2964 5148
rect 1581 5111 1639 5117
rect 2958 5108 2964 5120
rect 3016 5108 3022 5160
rect 3605 5151 3663 5157
rect 3605 5148 3617 5151
rect 3528 5120 3617 5148
rect 2038 5012 2044 5024
rect 1999 4984 2044 5012
rect 2038 4972 2044 4984
rect 2096 4972 2102 5024
rect 2130 4972 2136 5024
rect 2188 5012 2194 5024
rect 2188 4984 2233 5012
rect 2188 4972 2194 4984
rect 3326 4972 3332 5024
rect 3384 5012 3390 5024
rect 3421 5015 3479 5021
rect 3421 5012 3433 5015
rect 3384 4984 3433 5012
rect 3384 4972 3390 4984
rect 3421 4981 3433 4984
rect 3467 4981 3479 5015
rect 3528 5012 3556 5120
rect 3605 5117 3617 5120
rect 3651 5117 3663 5151
rect 3804 5148 3832 5188
rect 5997 5185 6009 5219
rect 6043 5185 6055 5219
rect 5997 5179 6055 5185
rect 6086 5176 6092 5228
rect 6144 5216 6150 5228
rect 6546 5216 6552 5228
rect 6144 5188 6552 5216
rect 6144 5176 6150 5188
rect 6546 5176 6552 5188
rect 6604 5176 6610 5228
rect 6914 5216 6920 5228
rect 6875 5188 6920 5216
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 7101 5219 7159 5225
rect 7101 5185 7113 5219
rect 7147 5216 7159 5219
rect 7392 5216 7420 5324
rect 7834 5312 7840 5364
rect 7892 5352 7898 5364
rect 8938 5352 8944 5364
rect 7892 5324 8944 5352
rect 7892 5312 7898 5324
rect 8938 5312 8944 5324
rect 8996 5312 9002 5364
rect 11054 5352 11060 5364
rect 11015 5324 11060 5352
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 13170 5312 13176 5364
rect 13228 5352 13234 5364
rect 13357 5355 13415 5361
rect 13357 5352 13369 5355
rect 13228 5324 13369 5352
rect 13228 5312 13234 5324
rect 13357 5321 13369 5324
rect 13403 5321 13415 5355
rect 13357 5315 13415 5321
rect 15381 5355 15439 5361
rect 15381 5321 15393 5355
rect 15427 5352 15439 5355
rect 15470 5352 15476 5364
rect 15427 5324 15476 5352
rect 15427 5321 15439 5324
rect 15381 5315 15439 5321
rect 8018 5244 8024 5296
rect 8076 5284 8082 5296
rect 8297 5287 8355 5293
rect 8297 5284 8309 5287
rect 8076 5256 8309 5284
rect 8076 5244 8082 5256
rect 8297 5253 8309 5256
rect 8343 5253 8355 5287
rect 8297 5247 8355 5253
rect 9950 5244 9956 5296
rect 10008 5244 10014 5296
rect 10045 5287 10103 5293
rect 10045 5253 10057 5287
rect 10091 5284 10103 5287
rect 10226 5284 10232 5296
rect 10091 5256 10232 5284
rect 10091 5253 10103 5256
rect 10045 5247 10103 5253
rect 10226 5244 10232 5256
rect 10284 5244 10290 5296
rect 11072 5284 11100 5312
rect 11072 5256 12020 5284
rect 7837 5219 7895 5225
rect 7837 5216 7849 5219
rect 7147 5188 7849 5216
rect 7147 5185 7159 5188
rect 7101 5179 7159 5185
rect 7837 5185 7849 5188
rect 7883 5185 7895 5219
rect 7837 5179 7895 5185
rect 9674 5176 9680 5228
rect 9732 5216 9738 5228
rect 9968 5216 9996 5244
rect 11992 5225 12020 5256
rect 10689 5219 10747 5225
rect 9732 5188 9777 5216
rect 9968 5188 10640 5216
rect 9732 5176 9738 5188
rect 4154 5157 4160 5160
rect 3881 5151 3939 5157
rect 3881 5148 3893 5151
rect 3804 5120 3893 5148
rect 3605 5111 3663 5117
rect 3881 5117 3893 5120
rect 3927 5117 3939 5151
rect 4148 5148 4160 5157
rect 4067 5120 4160 5148
rect 3881 5111 3939 5117
rect 4148 5111 4160 5120
rect 4212 5148 4218 5160
rect 4522 5148 4528 5160
rect 4212 5120 4528 5148
rect 3694 5080 3700 5092
rect 3655 5052 3700 5080
rect 3694 5040 3700 5052
rect 3752 5040 3758 5092
rect 3896 5080 3924 5111
rect 4154 5108 4160 5111
rect 4212 5108 4218 5120
rect 4522 5108 4528 5120
rect 4580 5108 4586 5160
rect 6730 5148 6736 5160
rect 5276 5120 6736 5148
rect 3970 5080 3976 5092
rect 3896 5052 3976 5080
rect 3970 5040 3976 5052
rect 4028 5040 4034 5092
rect 5276 5012 5304 5120
rect 6730 5108 6736 5120
rect 6788 5108 6794 5160
rect 6825 5151 6883 5157
rect 6825 5117 6837 5151
rect 6871 5148 6883 5151
rect 7742 5148 7748 5160
rect 6871 5120 7748 5148
rect 6871 5117 6883 5120
rect 6825 5111 6883 5117
rect 7742 5108 7748 5120
rect 7800 5108 7806 5160
rect 9766 5108 9772 5160
rect 9824 5148 9830 5160
rect 9953 5151 10011 5157
rect 9953 5148 9965 5151
rect 9824 5120 9965 5148
rect 9824 5108 9830 5120
rect 9953 5117 9965 5120
rect 9999 5117 10011 5151
rect 10502 5148 10508 5160
rect 10463 5120 10508 5148
rect 9953 5111 10011 5117
rect 10502 5108 10508 5120
rect 10560 5108 10566 5160
rect 10612 5148 10640 5188
rect 10689 5185 10701 5219
rect 10735 5216 10747 5219
rect 11977 5219 12035 5225
rect 10735 5188 11836 5216
rect 10735 5185 10747 5188
rect 10689 5179 10747 5185
rect 10873 5151 10931 5157
rect 10873 5148 10885 5151
rect 10612 5120 10885 5148
rect 10873 5117 10885 5120
rect 10919 5117 10931 5151
rect 10873 5111 10931 5117
rect 5905 5083 5963 5089
rect 5905 5049 5917 5083
rect 5951 5080 5963 5083
rect 6178 5080 6184 5092
rect 5951 5052 6184 5080
rect 5951 5049 5963 5052
rect 5905 5043 5963 5049
rect 6178 5040 6184 5052
rect 6236 5040 6242 5092
rect 6454 5040 6460 5092
rect 6512 5080 6518 5092
rect 6914 5080 6920 5092
rect 6512 5052 6920 5080
rect 6512 5040 6518 5052
rect 6914 5040 6920 5052
rect 6972 5080 6978 5092
rect 7190 5080 7196 5092
rect 6972 5052 7196 5080
rect 6972 5040 6978 5052
rect 7190 5040 7196 5052
rect 7248 5040 7254 5092
rect 7466 5040 7472 5092
rect 7524 5080 7530 5092
rect 7524 5052 8156 5080
rect 7524 5040 7530 5052
rect 8128 5024 8156 5052
rect 8846 5040 8852 5092
rect 8904 5080 8910 5092
rect 9410 5083 9468 5089
rect 9410 5080 9422 5083
rect 8904 5052 9422 5080
rect 8904 5040 8910 5052
rect 9410 5049 9422 5052
rect 9456 5049 9468 5083
rect 9410 5043 9468 5049
rect 11241 5083 11299 5089
rect 11241 5049 11253 5083
rect 11287 5080 11299 5083
rect 11606 5080 11612 5092
rect 11287 5052 11612 5080
rect 11287 5049 11299 5052
rect 11241 5043 11299 5049
rect 11606 5040 11612 5052
rect 11664 5040 11670 5092
rect 11808 5024 11836 5188
rect 11977 5185 11989 5219
rect 12023 5216 12035 5219
rect 13372 5216 13400 5315
rect 15470 5312 15476 5324
rect 15528 5312 15534 5364
rect 14829 5287 14887 5293
rect 14829 5253 14841 5287
rect 14875 5253 14887 5287
rect 14829 5247 14887 5253
rect 12023 5188 12112 5216
rect 13372 5188 13584 5216
rect 12023 5185 12035 5188
rect 11977 5179 12035 5185
rect 12084 5160 12112 5188
rect 12066 5108 12072 5160
rect 12124 5148 12130 5160
rect 13449 5151 13507 5157
rect 13449 5148 13461 5151
rect 12124 5120 13461 5148
rect 12124 5108 12130 5120
rect 13449 5117 13461 5120
rect 13495 5117 13507 5151
rect 13556 5148 13584 5188
rect 13705 5151 13763 5157
rect 13705 5148 13717 5151
rect 13556 5120 13717 5148
rect 13449 5111 13507 5117
rect 13705 5117 13717 5120
rect 13751 5117 13763 5151
rect 13705 5111 13763 5117
rect 12244 5083 12302 5089
rect 12244 5049 12256 5083
rect 12290 5080 12302 5083
rect 13170 5080 13176 5092
rect 12290 5052 13176 5080
rect 12290 5049 12302 5052
rect 12244 5043 12302 5049
rect 13170 5040 13176 5052
rect 13228 5040 13234 5092
rect 14844 5080 14872 5247
rect 15197 5151 15255 5157
rect 15197 5117 15209 5151
rect 15243 5148 15255 5151
rect 15286 5148 15292 5160
rect 15243 5120 15292 5148
rect 15243 5117 15255 5120
rect 15197 5111 15255 5117
rect 15286 5108 15292 5120
rect 15344 5108 15350 5160
rect 13648 5052 14872 5080
rect 3528 4984 5304 5012
rect 3421 4975 3479 4981
rect 5350 4972 5356 5024
rect 5408 5012 5414 5024
rect 5534 5012 5540 5024
rect 5408 4984 5453 5012
rect 5495 4984 5540 5012
rect 5408 4972 5414 4984
rect 5534 4972 5540 4984
rect 5592 4972 5598 5024
rect 6270 4972 6276 5024
rect 6328 5012 6334 5024
rect 7006 5012 7012 5024
rect 6328 4984 7012 5012
rect 6328 4972 6334 4984
rect 7006 4972 7012 4984
rect 7064 4972 7070 5024
rect 7374 4972 7380 5024
rect 7432 5012 7438 5024
rect 7653 5015 7711 5021
rect 7653 5012 7665 5015
rect 7432 4984 7665 5012
rect 7432 4972 7438 4984
rect 7653 4981 7665 4984
rect 7699 4981 7711 5015
rect 7653 4975 7711 4981
rect 7742 4972 7748 5024
rect 7800 5012 7806 5024
rect 8110 5012 8116 5024
rect 7800 4984 7845 5012
rect 8071 4984 8116 5012
rect 7800 4972 7806 4984
rect 8110 4972 8116 4984
rect 8168 4972 8174 5024
rect 8570 4972 8576 5024
rect 8628 5012 8634 5024
rect 9214 5012 9220 5024
rect 8628 4984 9220 5012
rect 8628 4972 8634 4984
rect 9214 4972 9220 4984
rect 9272 4972 9278 5024
rect 9306 4972 9312 5024
rect 9364 5012 9370 5024
rect 9769 5015 9827 5021
rect 9769 5012 9781 5015
rect 9364 4984 9781 5012
rect 9364 4972 9370 4984
rect 9769 4981 9781 4984
rect 9815 4981 9827 5015
rect 10410 5012 10416 5024
rect 10371 4984 10416 5012
rect 9769 4975 9827 4981
rect 10410 4972 10416 4984
rect 10468 4972 10474 5024
rect 11330 5012 11336 5024
rect 11291 4984 11336 5012
rect 11330 4972 11336 4984
rect 11388 4972 11394 5024
rect 11698 5012 11704 5024
rect 11659 4984 11704 5012
rect 11698 4972 11704 4984
rect 11756 4972 11762 5024
rect 11790 4972 11796 5024
rect 11848 5012 11854 5024
rect 13648 5012 13676 5052
rect 14918 5012 14924 5024
rect 11848 4984 13676 5012
rect 14879 4984 14924 5012
rect 11848 4972 11854 4984
rect 14918 4972 14924 4984
rect 14976 4972 14982 5024
rect 15010 4972 15016 5024
rect 15068 5012 15074 5024
rect 15473 5015 15531 5021
rect 15473 5012 15485 5015
rect 15068 4984 15485 5012
rect 15068 4972 15074 4984
rect 15473 4981 15485 4984
rect 15519 4981 15531 5015
rect 15473 4975 15531 4981
rect 1104 4922 16008 4944
rect 1104 4870 5979 4922
rect 6031 4870 6043 4922
rect 6095 4870 6107 4922
rect 6159 4870 6171 4922
rect 6223 4870 10976 4922
rect 11028 4870 11040 4922
rect 11092 4870 11104 4922
rect 11156 4870 11168 4922
rect 11220 4870 16008 4922
rect 1104 4848 16008 4870
rect 2038 4808 2044 4820
rect 1999 4780 2044 4808
rect 2038 4768 2044 4780
rect 2096 4768 2102 4820
rect 2130 4768 2136 4820
rect 2188 4808 2194 4820
rect 2869 4811 2927 4817
rect 2869 4808 2881 4811
rect 2188 4780 2881 4808
rect 2188 4768 2194 4780
rect 2869 4777 2881 4780
rect 2915 4777 2927 4811
rect 3694 4808 3700 4820
rect 2869 4771 2927 4777
rect 3252 4780 3700 4808
rect 2501 4743 2559 4749
rect 2501 4709 2513 4743
rect 2547 4740 2559 4743
rect 3252 4740 3280 4780
rect 3694 4768 3700 4780
rect 3752 4768 3758 4820
rect 3878 4808 3884 4820
rect 3839 4780 3884 4808
rect 3878 4768 3884 4780
rect 3936 4768 3942 4820
rect 5997 4811 6055 4817
rect 5997 4777 6009 4811
rect 6043 4777 6055 4811
rect 5997 4771 6055 4777
rect 6733 4811 6791 4817
rect 6733 4777 6745 4811
rect 6779 4808 6791 4811
rect 7190 4808 7196 4820
rect 6779 4780 7052 4808
rect 7151 4780 7196 4808
rect 6779 4777 6791 4780
rect 6733 4771 6791 4777
rect 2547 4712 3280 4740
rect 3329 4743 3387 4749
rect 2547 4709 2559 4712
rect 2501 4703 2559 4709
rect 3329 4709 3341 4743
rect 3375 4740 3387 4743
rect 3786 4740 3792 4752
rect 3375 4712 3792 4740
rect 3375 4709 3387 4712
rect 3329 4703 3387 4709
rect 3786 4700 3792 4712
rect 3844 4700 3850 4752
rect 4706 4740 4712 4752
rect 4141 4712 4712 4740
rect 1670 4672 1676 4684
rect 1631 4644 1676 4672
rect 1670 4632 1676 4644
rect 1728 4632 1734 4684
rect 1949 4675 2007 4681
rect 1949 4641 1961 4675
rect 1995 4641 2007 4675
rect 1949 4635 2007 4641
rect 1964 4536 1992 4635
rect 2130 4632 2136 4684
rect 2188 4672 2194 4684
rect 2409 4675 2467 4681
rect 2409 4672 2421 4675
rect 2188 4644 2421 4672
rect 2188 4632 2194 4644
rect 2409 4641 2421 4644
rect 2455 4641 2467 4675
rect 2409 4635 2467 4641
rect 3142 4632 3148 4684
rect 3200 4672 3206 4684
rect 3237 4675 3295 4681
rect 3237 4672 3249 4675
rect 3200 4644 3249 4672
rect 3200 4632 3206 4644
rect 3237 4641 3249 4644
rect 3283 4641 3295 4675
rect 3804 4672 3832 4700
rect 4141 4672 4169 4712
rect 4706 4700 4712 4712
rect 4764 4700 4770 4752
rect 5718 4700 5724 4752
rect 5776 4740 5782 4752
rect 6012 4740 6040 4771
rect 7024 4749 7052 4780
rect 7190 4768 7196 4780
rect 7248 4768 7254 4820
rect 7374 4808 7380 4820
rect 7335 4780 7380 4808
rect 7374 4768 7380 4780
rect 7432 4768 7438 4820
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 7745 4811 7803 4817
rect 7745 4808 7757 4811
rect 7708 4780 7757 4808
rect 7708 4768 7714 4780
rect 7745 4777 7757 4780
rect 7791 4777 7803 4811
rect 7745 4771 7803 4777
rect 7837 4811 7895 4817
rect 7837 4777 7849 4811
rect 7883 4808 7895 4811
rect 7926 4808 7932 4820
rect 7883 4780 7932 4808
rect 7883 4777 7895 4780
rect 7837 4771 7895 4777
rect 7009 4743 7067 4749
rect 5776 4712 5948 4740
rect 6012 4712 6960 4740
rect 5776 4700 5782 4712
rect 4246 4672 4252 4684
rect 3804 4644 4169 4672
rect 4207 4644 4252 4672
rect 3237 4635 3295 4641
rect 4246 4632 4252 4644
rect 4304 4632 4310 4684
rect 4341 4675 4399 4681
rect 4341 4641 4353 4675
rect 4387 4672 4399 4675
rect 4798 4672 4804 4684
rect 4387 4644 4804 4672
rect 4387 4641 4399 4644
rect 4341 4635 4399 4641
rect 4798 4632 4804 4644
rect 4856 4632 4862 4684
rect 4893 4675 4951 4681
rect 4893 4641 4905 4675
rect 4939 4672 4951 4675
rect 5074 4672 5080 4684
rect 4939 4644 5080 4672
rect 4939 4641 4951 4644
rect 4893 4635 4951 4641
rect 5074 4632 5080 4644
rect 5132 4632 5138 4684
rect 5169 4675 5227 4681
rect 5169 4641 5181 4675
rect 5215 4672 5227 4675
rect 5258 4672 5264 4684
rect 5215 4644 5264 4672
rect 5215 4641 5227 4644
rect 5169 4635 5227 4641
rect 5258 4632 5264 4644
rect 5316 4632 5322 4684
rect 5350 4632 5356 4684
rect 5408 4672 5414 4684
rect 5445 4675 5503 4681
rect 5445 4672 5457 4675
rect 5408 4644 5457 4672
rect 5408 4632 5414 4644
rect 5445 4641 5457 4644
rect 5491 4641 5503 4675
rect 5445 4635 5503 4641
rect 5537 4675 5595 4681
rect 5537 4641 5549 4675
rect 5583 4672 5595 4675
rect 5626 4672 5632 4684
rect 5583 4644 5632 4672
rect 5583 4641 5595 4644
rect 5537 4635 5595 4641
rect 5626 4632 5632 4644
rect 5684 4632 5690 4684
rect 5810 4672 5816 4684
rect 5771 4644 5816 4672
rect 5810 4632 5816 4644
rect 5868 4632 5874 4684
rect 5920 4672 5948 4712
rect 6365 4675 6423 4681
rect 6365 4672 6377 4675
rect 5920 4644 6377 4672
rect 6365 4641 6377 4644
rect 6411 4672 6423 4675
rect 6454 4672 6460 4684
rect 6411 4644 6460 4672
rect 6411 4641 6423 4644
rect 6365 4635 6423 4641
rect 6454 4632 6460 4644
rect 6512 4632 6518 4684
rect 6549 4675 6607 4681
rect 6549 4641 6561 4675
rect 6595 4641 6607 4675
rect 6932 4672 6960 4712
rect 7009 4709 7021 4743
rect 7055 4709 7067 4743
rect 7760 4740 7788 4771
rect 7926 4768 7932 4780
rect 7984 4768 7990 4820
rect 9953 4811 10011 4817
rect 9953 4777 9965 4811
rect 9999 4808 10011 4811
rect 10042 4808 10048 4820
rect 9999 4780 10048 4808
rect 9999 4777 10011 4780
rect 9953 4771 10011 4777
rect 10042 4768 10048 4780
rect 10100 4768 10106 4820
rect 12066 4768 12072 4820
rect 12124 4768 12130 4820
rect 13170 4808 13176 4820
rect 13131 4780 13176 4808
rect 13170 4768 13176 4780
rect 13228 4768 13234 4820
rect 13817 4811 13875 4817
rect 13817 4777 13829 4811
rect 13863 4808 13875 4811
rect 14918 4808 14924 4820
rect 13863 4780 14924 4808
rect 13863 4777 13875 4780
rect 13817 4771 13875 4777
rect 14918 4768 14924 4780
rect 14976 4768 14982 4820
rect 15473 4811 15531 4817
rect 15473 4777 15485 4811
rect 15519 4808 15531 4811
rect 15838 4808 15844 4820
rect 15519 4780 15844 4808
rect 15519 4777 15531 4780
rect 15473 4771 15531 4777
rect 15838 4768 15844 4780
rect 15896 4768 15902 4820
rect 9306 4740 9312 4752
rect 7760 4712 9168 4740
rect 9267 4712 9312 4740
rect 7009 4703 7067 4709
rect 7190 4672 7196 4684
rect 6932 4644 7196 4672
rect 6549 4635 6607 4641
rect 2685 4607 2743 4613
rect 2685 4573 2697 4607
rect 2731 4604 2743 4607
rect 3050 4604 3056 4616
rect 2731 4576 3056 4604
rect 2731 4573 2743 4576
rect 2685 4567 2743 4573
rect 3050 4564 3056 4576
rect 3108 4604 3114 4616
rect 3513 4607 3571 4613
rect 3513 4604 3525 4607
rect 3108 4576 3525 4604
rect 3108 4564 3114 4576
rect 3513 4573 3525 4576
rect 3559 4604 3571 4607
rect 4062 4604 4068 4616
rect 3559 4576 4068 4604
rect 3559 4573 3571 4576
rect 3513 4567 3571 4573
rect 4062 4564 4068 4576
rect 4120 4564 4126 4616
rect 4154 4564 4160 4616
rect 4212 4604 4218 4616
rect 4433 4607 4491 4613
rect 4433 4604 4445 4607
rect 4212 4576 4445 4604
rect 4212 4564 4218 4576
rect 4433 4573 4445 4576
rect 4479 4573 4491 4607
rect 6564 4604 6592 4635
rect 7190 4632 7196 4644
rect 7248 4632 7254 4684
rect 8570 4672 8576 4684
rect 8531 4644 8576 4672
rect 8570 4632 8576 4644
rect 8628 4632 8634 4684
rect 9140 4672 9168 4712
rect 9306 4700 9312 4712
rect 9364 4700 9370 4752
rect 10778 4740 10784 4752
rect 10244 4712 10784 4740
rect 9214 4672 9220 4684
rect 9140 4644 9220 4672
rect 9214 4632 9220 4644
rect 9272 4632 9278 4684
rect 9861 4675 9919 4681
rect 9861 4641 9873 4675
rect 9907 4672 9919 4675
rect 9907 4644 9996 4672
rect 9907 4641 9919 4644
rect 9861 4635 9919 4641
rect 7098 4604 7104 4616
rect 4433 4567 4491 4573
rect 4540 4576 5580 4604
rect 6564 4576 7104 4604
rect 4540 4536 4568 4576
rect 5552 4548 5580 4576
rect 7098 4564 7104 4576
rect 7156 4564 7162 4616
rect 8018 4604 8024 4616
rect 7979 4576 8024 4604
rect 8018 4564 8024 4576
rect 8076 4564 8082 4616
rect 8662 4604 8668 4616
rect 8623 4576 8668 4604
rect 8662 4564 8668 4576
rect 8720 4564 8726 4616
rect 8846 4604 8852 4616
rect 8807 4576 8852 4604
rect 8846 4564 8852 4576
rect 8904 4564 8910 4616
rect 1964 4508 4568 4536
rect 4614 4496 4620 4548
rect 4672 4536 4678 4548
rect 5261 4539 5319 4545
rect 5261 4536 5273 4539
rect 4672 4508 5273 4536
rect 4672 4496 4678 4508
rect 5261 4505 5273 4508
rect 5307 4505 5319 4539
rect 5261 4499 5319 4505
rect 5534 4496 5540 4548
rect 5592 4496 5598 4548
rect 5721 4539 5779 4545
rect 5721 4505 5733 4539
rect 5767 4536 5779 4539
rect 6822 4536 6828 4548
rect 5767 4508 6684 4536
rect 6783 4508 6828 4536
rect 5767 4505 5779 4508
rect 5721 4499 5779 4505
rect 1486 4468 1492 4480
rect 1447 4440 1492 4468
rect 1486 4428 1492 4440
rect 1544 4428 1550 4480
rect 1762 4468 1768 4480
rect 1723 4440 1768 4468
rect 1762 4428 1768 4440
rect 1820 4428 1826 4480
rect 4338 4428 4344 4480
rect 4396 4468 4402 4480
rect 4709 4471 4767 4477
rect 4709 4468 4721 4471
rect 4396 4440 4721 4468
rect 4396 4428 4402 4440
rect 4709 4437 4721 4440
rect 4755 4437 4767 4471
rect 4982 4468 4988 4480
rect 4943 4440 4988 4468
rect 4709 4431 4767 4437
rect 4982 4428 4988 4440
rect 5040 4428 5046 4480
rect 6181 4471 6239 4477
rect 6181 4437 6193 4471
rect 6227 4468 6239 4471
rect 6270 4468 6276 4480
rect 6227 4440 6276 4468
rect 6227 4437 6239 4440
rect 6181 4431 6239 4437
rect 6270 4428 6276 4440
rect 6328 4428 6334 4480
rect 6656 4468 6684 4508
rect 6822 4496 6828 4508
rect 6880 4496 6886 4548
rect 8294 4496 8300 4548
rect 8352 4536 8358 4548
rect 9125 4539 9183 4545
rect 9125 4536 9137 4539
rect 8352 4508 9137 4536
rect 8352 4496 8358 4508
rect 9125 4505 9137 4508
rect 9171 4505 9183 4539
rect 9968 4536 9996 4644
rect 10137 4607 10195 4613
rect 10137 4573 10149 4607
rect 10183 4604 10195 4607
rect 10244 4604 10272 4712
rect 10778 4700 10784 4712
rect 10836 4740 10842 4752
rect 11456 4743 11514 4749
rect 11456 4740 11468 4743
rect 10836 4712 11468 4740
rect 10836 4700 10842 4712
rect 11456 4709 11468 4712
rect 11502 4740 11514 4743
rect 11790 4740 11796 4752
rect 11502 4712 11796 4740
rect 11502 4709 11514 4712
rect 11456 4703 11514 4709
rect 11790 4700 11796 4712
rect 11848 4700 11854 4752
rect 12084 4740 12112 4768
rect 11900 4712 12112 4740
rect 13725 4743 13783 4749
rect 11701 4675 11759 4681
rect 11701 4641 11713 4675
rect 11747 4672 11759 4675
rect 11900 4672 11928 4712
rect 13725 4709 13737 4743
rect 13771 4740 13783 4743
rect 14550 4740 14556 4752
rect 13771 4712 14556 4740
rect 13771 4709 13783 4712
rect 13725 4703 13783 4709
rect 14550 4700 14556 4712
rect 14608 4700 14614 4752
rect 14734 4740 14740 4752
rect 14695 4712 14740 4740
rect 14734 4700 14740 4712
rect 14792 4740 14798 4752
rect 15286 4740 15292 4752
rect 14792 4712 15292 4740
rect 14792 4700 14798 4712
rect 15286 4700 15292 4712
rect 15344 4700 15350 4752
rect 12066 4681 12072 4684
rect 12060 4672 12072 4681
rect 11747 4644 11928 4672
rect 11979 4644 12072 4672
rect 11747 4641 11759 4644
rect 11701 4635 11759 4641
rect 11808 4613 11836 4644
rect 12060 4635 12072 4644
rect 12124 4672 12130 4684
rect 12124 4644 13952 4672
rect 12066 4632 12072 4635
rect 12124 4632 12130 4644
rect 13556 4613 13584 4644
rect 10183 4576 10272 4604
rect 11793 4607 11851 4613
rect 10183 4573 10195 4576
rect 10137 4567 10195 4573
rect 11793 4573 11805 4607
rect 11839 4604 11851 4607
rect 13541 4607 13599 4613
rect 11839 4576 11873 4604
rect 11839 4573 11851 4576
rect 11793 4567 11851 4573
rect 13541 4573 13553 4607
rect 13587 4573 13599 4607
rect 13924 4604 13952 4644
rect 14366 4632 14372 4684
rect 14424 4672 14430 4684
rect 14829 4675 14887 4681
rect 14829 4672 14841 4675
rect 14424 4644 14841 4672
rect 14424 4632 14430 4644
rect 14829 4641 14841 4644
rect 14875 4641 14887 4675
rect 14829 4635 14887 4641
rect 15565 4675 15623 4681
rect 15565 4641 15577 4675
rect 15611 4672 15623 4675
rect 15746 4672 15752 4684
rect 15611 4644 15752 4672
rect 15611 4641 15623 4644
rect 15565 4635 15623 4641
rect 15746 4632 15752 4644
rect 15804 4672 15810 4684
rect 16482 4672 16488 4684
rect 15804 4644 16488 4672
rect 15804 4632 15810 4644
rect 16482 4632 16488 4644
rect 16540 4632 16546 4684
rect 14182 4604 14188 4616
rect 13924 4576 14188 4604
rect 13541 4567 13599 4573
rect 14182 4564 14188 4576
rect 14240 4604 14246 4616
rect 14921 4607 14979 4613
rect 14921 4604 14933 4607
rect 14240 4576 14933 4604
rect 14240 4564 14246 4576
rect 14921 4573 14933 4576
rect 14967 4573 14979 4607
rect 14921 4567 14979 4573
rect 10686 4536 10692 4548
rect 9968 4508 10692 4536
rect 9125 4499 9183 4505
rect 10686 4496 10692 4508
rect 10744 4496 10750 4548
rect 13265 4539 13323 4545
rect 13265 4536 13277 4539
rect 12728 4508 13277 4536
rect 7098 4468 7104 4480
rect 6656 4440 7104 4468
rect 7098 4428 7104 4440
rect 7156 4428 7162 4480
rect 8202 4468 8208 4480
rect 8163 4440 8208 4468
rect 8202 4428 8208 4440
rect 8260 4428 8266 4480
rect 9493 4471 9551 4477
rect 9493 4437 9505 4471
rect 9539 4468 9551 4471
rect 9674 4468 9680 4480
rect 9539 4440 9680 4468
rect 9539 4437 9551 4440
rect 9493 4431 9551 4437
rect 9674 4428 9680 4440
rect 9732 4428 9738 4480
rect 10318 4468 10324 4480
rect 10279 4440 10324 4468
rect 10318 4428 10324 4440
rect 10376 4428 10382 4480
rect 12434 4428 12440 4480
rect 12492 4468 12498 4480
rect 12728 4468 12756 4508
rect 13265 4505 13277 4508
rect 13311 4505 13323 4539
rect 13265 4499 13323 4505
rect 12492 4440 12756 4468
rect 12492 4428 12498 4440
rect 13998 4428 14004 4480
rect 14056 4468 14062 4480
rect 14185 4471 14243 4477
rect 14185 4468 14197 4471
rect 14056 4440 14197 4468
rect 14056 4428 14062 4440
rect 14185 4437 14197 4440
rect 14231 4437 14243 4471
rect 14366 4468 14372 4480
rect 14327 4440 14372 4468
rect 14185 4431 14243 4437
rect 14366 4428 14372 4440
rect 14424 4428 14430 4480
rect 14642 4428 14648 4480
rect 14700 4468 14706 4480
rect 15197 4471 15255 4477
rect 15197 4468 15209 4471
rect 14700 4440 15209 4468
rect 14700 4428 14706 4440
rect 15197 4437 15209 4440
rect 15243 4437 15255 4471
rect 15197 4431 15255 4437
rect 1104 4378 16008 4400
rect 1104 4326 3480 4378
rect 3532 4326 3544 4378
rect 3596 4326 3608 4378
rect 3660 4326 3672 4378
rect 3724 4326 8478 4378
rect 8530 4326 8542 4378
rect 8594 4326 8606 4378
rect 8658 4326 8670 4378
rect 8722 4326 13475 4378
rect 13527 4326 13539 4378
rect 13591 4326 13603 4378
rect 13655 4326 13667 4378
rect 13719 4326 16008 4378
rect 1104 4304 16008 4326
rect 3050 4264 3056 4276
rect 3011 4236 3056 4264
rect 3050 4224 3056 4236
rect 3108 4224 3114 4276
rect 4062 4224 4068 4276
rect 4120 4264 4126 4276
rect 4120 4236 4476 4264
rect 4120 4224 4126 4236
rect 1394 4128 1400 4140
rect 1355 4100 1400 4128
rect 1394 4088 1400 4100
rect 1452 4088 1458 4140
rect 4448 4137 4476 4236
rect 4798 4224 4804 4276
rect 4856 4264 4862 4276
rect 5077 4267 5135 4273
rect 5077 4264 5089 4267
rect 4856 4236 5089 4264
rect 4856 4224 4862 4236
rect 5077 4233 5089 4236
rect 5123 4233 5135 4267
rect 5077 4227 5135 4233
rect 6481 4236 7696 4264
rect 4706 4156 4712 4208
rect 4764 4196 4770 4208
rect 4893 4199 4951 4205
rect 4893 4196 4905 4199
rect 4764 4168 4905 4196
rect 4764 4156 4770 4168
rect 4893 4165 4905 4168
rect 4939 4196 4951 4199
rect 6481 4196 6509 4236
rect 4939 4168 6509 4196
rect 7668 4196 7696 4236
rect 7742 4224 7748 4276
rect 7800 4264 7806 4276
rect 7929 4267 7987 4273
rect 7929 4264 7941 4267
rect 7800 4236 7941 4264
rect 7800 4224 7806 4236
rect 7929 4233 7941 4236
rect 7975 4233 7987 4267
rect 7929 4227 7987 4233
rect 8018 4224 8024 4276
rect 8076 4264 8082 4276
rect 8076 4236 8616 4264
rect 8076 4224 8082 4236
rect 7834 4196 7840 4208
rect 7668 4168 7840 4196
rect 4939 4165 4951 4168
rect 4893 4159 4951 4165
rect 7834 4156 7840 4168
rect 7892 4156 7898 4208
rect 4433 4131 4491 4137
rect 4433 4097 4445 4131
rect 4479 4097 4491 4131
rect 4433 4091 4491 4097
rect 1581 4063 1639 4069
rect 1581 4029 1593 4063
rect 1627 4060 1639 4063
rect 1762 4060 1768 4072
rect 1627 4032 1768 4060
rect 1627 4029 1639 4032
rect 1581 4023 1639 4029
rect 1762 4020 1768 4032
rect 1820 4020 1826 4072
rect 1854 4020 1860 4072
rect 1912 4060 1918 4072
rect 1949 4063 2007 4069
rect 1949 4060 1961 4063
rect 1912 4032 1961 4060
rect 1912 4020 1918 4032
rect 1949 4029 1961 4032
rect 1995 4029 2007 4063
rect 1949 4023 2007 4029
rect 2225 4063 2283 4069
rect 2225 4029 2237 4063
rect 2271 4060 2283 4063
rect 2314 4060 2320 4072
rect 2271 4032 2320 4060
rect 2271 4029 2283 4032
rect 2225 4023 2283 4029
rect 2314 4020 2320 4032
rect 2372 4020 2378 4072
rect 2409 4063 2467 4069
rect 2409 4029 2421 4063
rect 2455 4060 2467 4063
rect 2498 4060 2504 4072
rect 2455 4032 2504 4060
rect 2455 4029 2467 4032
rect 2409 4023 2467 4029
rect 2498 4020 2504 4032
rect 2556 4020 2562 4072
rect 2777 4063 2835 4069
rect 2777 4029 2789 4063
rect 2823 4060 2835 4063
rect 4338 4060 4344 4072
rect 2823 4032 4344 4060
rect 2823 4029 2835 4032
rect 2777 4023 2835 4029
rect 4338 4020 4344 4032
rect 4396 4020 4402 4072
rect 2961 3995 3019 4001
rect 2961 3961 2973 3995
rect 3007 3992 3019 3995
rect 3234 3992 3240 4004
rect 3007 3964 3240 3992
rect 3007 3961 3019 3964
rect 2961 3955 3019 3961
rect 3234 3952 3240 3964
rect 3292 3952 3298 4004
rect 4154 3952 4160 4004
rect 4212 4001 4218 4004
rect 4212 3992 4224 4001
rect 4448 3992 4476 4091
rect 4522 4088 4528 4140
rect 4580 4128 4586 4140
rect 5629 4131 5687 4137
rect 5629 4128 5641 4131
rect 4580 4100 5641 4128
rect 4580 4088 4586 4100
rect 5629 4097 5641 4100
rect 5675 4097 5687 4131
rect 6457 4131 6515 4137
rect 6457 4128 6469 4131
rect 5629 4091 5687 4097
rect 5736 4100 6469 4128
rect 4709 4063 4767 4069
rect 4709 4029 4721 4063
rect 4755 4060 4767 4063
rect 4982 4060 4988 4072
rect 4755 4032 4988 4060
rect 4755 4029 4767 4032
rect 4709 4023 4767 4029
rect 4982 4020 4988 4032
rect 5040 4020 5046 4072
rect 5736 4060 5764 4100
rect 6457 4097 6469 4100
rect 6503 4097 6515 4131
rect 6457 4091 6515 4097
rect 8202 4088 8208 4140
rect 8260 4128 8266 4140
rect 8588 4137 8616 4236
rect 10042 4224 10048 4276
rect 10100 4264 10106 4276
rect 11057 4267 11115 4273
rect 11057 4264 11069 4267
rect 10100 4236 11069 4264
rect 10100 4224 10106 4236
rect 11057 4233 11069 4236
rect 11103 4233 11115 4267
rect 11514 4264 11520 4276
rect 11057 4227 11115 4233
rect 11164 4236 11520 4264
rect 10318 4196 10324 4208
rect 9508 4168 10324 4196
rect 9508 4137 9536 4168
rect 10318 4156 10324 4168
rect 10376 4156 10382 4208
rect 10778 4196 10784 4208
rect 10704 4168 10784 4196
rect 8389 4131 8447 4137
rect 8389 4128 8401 4131
rect 8260 4100 8401 4128
rect 8260 4088 8266 4100
rect 8389 4097 8401 4100
rect 8435 4097 8447 4131
rect 8389 4091 8447 4097
rect 8573 4131 8631 4137
rect 8573 4097 8585 4131
rect 8619 4097 8631 4131
rect 8573 4091 8631 4097
rect 9493 4131 9551 4137
rect 9493 4097 9505 4131
rect 9539 4097 9551 4131
rect 9493 4091 9551 4097
rect 9585 4131 9643 4137
rect 9585 4097 9597 4131
rect 9631 4128 9643 4131
rect 9674 4128 9680 4140
rect 9631 4100 9680 4128
rect 9631 4097 9643 4100
rect 9585 4091 9643 4097
rect 9674 4088 9680 4100
rect 9732 4088 9738 4140
rect 10704 4137 10732 4168
rect 10778 4156 10784 4168
rect 10836 4156 10842 4208
rect 10689 4131 10747 4137
rect 10689 4097 10701 4131
rect 10735 4097 10747 4131
rect 11164 4128 11192 4236
rect 11514 4224 11520 4236
rect 11572 4224 11578 4276
rect 14918 4224 14924 4276
rect 14976 4224 14982 4276
rect 15102 4264 15108 4276
rect 15063 4236 15108 4264
rect 15102 4224 15108 4236
rect 15160 4224 15166 4276
rect 11238 4156 11244 4208
rect 11296 4196 11302 4208
rect 11296 4168 11468 4196
rect 11296 4156 11302 4168
rect 10689 4091 10747 4097
rect 10796 4100 11192 4128
rect 5092 4032 5764 4060
rect 6089 4063 6147 4069
rect 5092 3992 5120 4032
rect 6089 4029 6101 4063
rect 6135 4060 6147 4063
rect 6178 4060 6184 4072
rect 6135 4032 6184 4060
rect 6135 4029 6147 4032
rect 6089 4023 6147 4029
rect 6178 4020 6184 4032
rect 6236 4020 6242 4072
rect 6546 4020 6552 4072
rect 6604 4060 6610 4072
rect 6713 4063 6771 4069
rect 6713 4060 6725 4063
rect 6604 4032 6725 4060
rect 6604 4020 6610 4032
rect 6713 4029 6725 4032
rect 6759 4029 6771 4063
rect 6713 4023 6771 4029
rect 7558 4020 7564 4072
rect 7616 4060 7622 4072
rect 8757 4063 8815 4069
rect 8757 4060 8769 4063
rect 7616 4032 8769 4060
rect 7616 4020 7622 4032
rect 8757 4029 8769 4032
rect 8803 4029 8815 4063
rect 8757 4023 8815 4029
rect 8846 4020 8852 4072
rect 8904 4060 8910 4072
rect 9125 4063 9183 4069
rect 9125 4060 9137 4063
rect 8904 4032 9137 4060
rect 8904 4020 8910 4032
rect 9125 4029 9137 4032
rect 9171 4029 9183 4063
rect 9125 4023 9183 4029
rect 9398 4020 9404 4072
rect 9456 4060 9462 4072
rect 10410 4060 10416 4072
rect 9456 4032 10416 4060
rect 9456 4020 9462 4032
rect 10410 4020 10416 4032
rect 10468 4060 10474 4072
rect 10597 4063 10655 4069
rect 10597 4060 10609 4063
rect 10468 4032 10609 4060
rect 10468 4020 10474 4032
rect 10597 4029 10609 4032
rect 10643 4060 10655 4063
rect 10796 4060 10824 4100
rect 10643 4032 10824 4060
rect 10643 4029 10655 4032
rect 10597 4023 10655 4029
rect 10870 4020 10876 4072
rect 10928 4060 10934 4072
rect 11146 4060 11152 4072
rect 10928 4032 11152 4060
rect 10928 4020 10934 4032
rect 11146 4020 11152 4032
rect 11204 4020 11210 4072
rect 11333 4063 11391 4069
rect 11333 4029 11345 4063
rect 11379 4060 11391 4063
rect 11440 4060 11468 4168
rect 12066 4156 12072 4208
rect 12124 4196 12130 4208
rect 13170 4196 13176 4208
rect 12124 4168 12204 4196
rect 12124 4156 12130 4168
rect 12176 4137 12204 4168
rect 13004 4168 13176 4196
rect 12161 4131 12219 4137
rect 12161 4097 12173 4131
rect 12207 4097 12219 4131
rect 12161 4091 12219 4097
rect 12250 4088 12256 4140
rect 12308 4128 12314 4140
rect 13004 4137 13032 4168
rect 13170 4156 13176 4168
rect 13228 4196 13234 4208
rect 14936 4196 14964 4224
rect 13228 4168 14228 4196
rect 14936 4168 15056 4196
rect 13228 4156 13234 4168
rect 12989 4131 13047 4137
rect 12308 4100 12434 4128
rect 12308 4088 12314 4100
rect 11379 4032 11468 4060
rect 11379 4029 11391 4032
rect 11333 4023 11391 4029
rect 11514 4020 11520 4072
rect 11572 4060 11578 4072
rect 11882 4060 11888 4072
rect 11572 4032 11888 4060
rect 11572 4020 11578 4032
rect 11882 4020 11888 4032
rect 11940 4020 11946 4072
rect 12406 4060 12434 4100
rect 12989 4097 13001 4131
rect 13035 4097 13047 4131
rect 12989 4091 13047 4097
rect 13078 4088 13084 4140
rect 13136 4128 13142 4140
rect 13722 4128 13728 4140
rect 13136 4100 13728 4128
rect 13136 4088 13142 4100
rect 13722 4088 13728 4100
rect 13780 4088 13786 4140
rect 14200 4137 14228 4168
rect 14185 4131 14243 4137
rect 14185 4097 14197 4131
rect 14231 4097 14243 4131
rect 14185 4091 14243 4097
rect 14553 4131 14611 4137
rect 14553 4097 14565 4131
rect 14599 4128 14611 4131
rect 14918 4128 14924 4140
rect 14599 4100 14924 4128
rect 14599 4097 14611 4100
rect 14553 4091 14611 4097
rect 14918 4088 14924 4100
rect 14976 4088 14982 4140
rect 15028 4072 15056 4168
rect 15381 4131 15439 4137
rect 15381 4128 15393 4131
rect 15120 4100 15393 4128
rect 13998 4060 14004 4072
rect 12406 4032 13860 4060
rect 13959 4032 14004 4060
rect 4212 3964 4257 3992
rect 4448 3964 5120 3992
rect 5445 3995 5503 4001
rect 4212 3955 4224 3964
rect 5445 3961 5457 3995
rect 5491 3992 5503 3995
rect 5626 3992 5632 4004
rect 5491 3964 5632 3992
rect 5491 3961 5503 3964
rect 5445 3955 5503 3961
rect 4212 3952 4218 3955
rect 5626 3952 5632 3964
rect 5684 3952 5690 4004
rect 7098 3952 7104 4004
rect 7156 3992 7162 4004
rect 8941 3995 8999 4001
rect 8941 3992 8953 3995
rect 7156 3964 8953 3992
rect 7156 3952 7162 3964
rect 8941 3961 8953 3964
rect 8987 3961 8999 3995
rect 8941 3955 8999 3961
rect 9677 3995 9735 4001
rect 9677 3961 9689 3995
rect 9723 3992 9735 3995
rect 10962 3992 10968 4004
rect 9723 3964 10968 3992
rect 9723 3961 9735 3964
rect 9677 3955 9735 3961
rect 10962 3952 10968 3964
rect 11020 3992 11026 4004
rect 12066 3992 12072 4004
rect 11020 3964 12072 3992
rect 11020 3952 11026 3964
rect 12066 3952 12072 3964
rect 12124 3952 12130 4004
rect 12253 3995 12311 4001
rect 12253 3961 12265 3995
rect 12299 3992 12311 3995
rect 12526 3992 12532 4004
rect 12299 3964 12532 3992
rect 12299 3961 12311 3964
rect 12253 3955 12311 3961
rect 12526 3952 12532 3964
rect 12584 3952 12590 4004
rect 13173 3995 13231 4001
rect 13173 3992 13185 3995
rect 12728 3964 13185 3992
rect 1578 3884 1584 3936
rect 1636 3924 1642 3936
rect 1765 3927 1823 3933
rect 1765 3924 1777 3927
rect 1636 3896 1777 3924
rect 1636 3884 1642 3896
rect 1765 3893 1777 3896
rect 1811 3893 1823 3927
rect 1765 3887 1823 3893
rect 2041 3927 2099 3933
rect 2041 3893 2053 3927
rect 2087 3924 2099 3927
rect 2314 3924 2320 3936
rect 2087 3896 2320 3924
rect 2087 3893 2099 3896
rect 2041 3887 2099 3893
rect 2314 3884 2320 3896
rect 2372 3884 2378 3936
rect 2590 3924 2596 3936
rect 2551 3896 2596 3924
rect 2590 3884 2596 3896
rect 2648 3884 2654 3936
rect 3970 3884 3976 3936
rect 4028 3924 4034 3936
rect 4617 3927 4675 3933
rect 4617 3924 4629 3927
rect 4028 3896 4629 3924
rect 4028 3884 4034 3896
rect 4617 3893 4629 3896
rect 4663 3893 4675 3927
rect 4617 3887 4675 3893
rect 5534 3884 5540 3936
rect 5592 3924 5598 3936
rect 6181 3927 6239 3933
rect 5592 3896 5637 3924
rect 5592 3884 5598 3896
rect 6181 3893 6193 3927
rect 6227 3924 6239 3927
rect 7650 3924 7656 3936
rect 6227 3896 7656 3924
rect 6227 3893 6239 3896
rect 6181 3887 6239 3893
rect 7650 3884 7656 3896
rect 7708 3884 7714 3936
rect 7834 3924 7840 3936
rect 7795 3896 7840 3924
rect 7834 3884 7840 3896
rect 7892 3884 7898 3936
rect 7926 3884 7932 3936
rect 7984 3924 7990 3936
rect 8297 3927 8355 3933
rect 8297 3924 8309 3927
rect 7984 3896 8309 3924
rect 7984 3884 7990 3896
rect 8297 3893 8309 3896
rect 8343 3924 8355 3927
rect 9582 3924 9588 3936
rect 8343 3896 9588 3924
rect 8343 3893 8355 3896
rect 8297 3887 8355 3893
rect 9582 3884 9588 3896
rect 9640 3884 9646 3936
rect 9766 3884 9772 3936
rect 9824 3924 9830 3936
rect 10045 3927 10103 3933
rect 10045 3924 10057 3927
rect 9824 3896 10057 3924
rect 9824 3884 9830 3896
rect 10045 3893 10057 3896
rect 10091 3893 10103 3927
rect 10045 3887 10103 3893
rect 10134 3884 10140 3936
rect 10192 3924 10198 3936
rect 10502 3924 10508 3936
rect 10192 3896 10237 3924
rect 10463 3896 10508 3924
rect 10192 3884 10198 3896
rect 10502 3884 10508 3896
rect 10560 3884 10566 3936
rect 10870 3884 10876 3936
rect 10928 3924 10934 3936
rect 11514 3924 11520 3936
rect 10928 3896 11520 3924
rect 10928 3884 10934 3896
rect 11514 3884 11520 3896
rect 11572 3884 11578 3936
rect 11701 3927 11759 3933
rect 11701 3893 11713 3927
rect 11747 3924 11759 3927
rect 11790 3924 11796 3936
rect 11747 3896 11796 3924
rect 11747 3893 11759 3896
rect 11701 3887 11759 3893
rect 11790 3884 11796 3896
rect 11848 3884 11854 3936
rect 12158 3884 12164 3936
rect 12216 3924 12222 3936
rect 12728 3933 12756 3964
rect 13173 3961 13185 3964
rect 13219 3961 13231 3995
rect 13173 3955 13231 3961
rect 13354 3952 13360 4004
rect 13412 3992 13418 4004
rect 13412 3964 13676 3992
rect 13412 3952 13418 3964
rect 12345 3927 12403 3933
rect 12345 3924 12357 3927
rect 12216 3896 12357 3924
rect 12216 3884 12222 3896
rect 12345 3893 12357 3896
rect 12391 3893 12403 3927
rect 12345 3887 12403 3893
rect 12713 3927 12771 3933
rect 12713 3893 12725 3927
rect 12759 3893 12771 3927
rect 12713 3887 12771 3893
rect 12894 3884 12900 3936
rect 12952 3924 12958 3936
rect 13081 3927 13139 3933
rect 13081 3924 13093 3927
rect 12952 3896 13093 3924
rect 12952 3884 12958 3896
rect 13081 3893 13093 3896
rect 13127 3893 13139 3927
rect 13081 3887 13139 3893
rect 13262 3884 13268 3936
rect 13320 3924 13326 3936
rect 13648 3933 13676 3964
rect 13541 3927 13599 3933
rect 13541 3924 13553 3927
rect 13320 3896 13553 3924
rect 13320 3884 13326 3896
rect 13541 3893 13553 3896
rect 13587 3893 13599 3927
rect 13541 3887 13599 3893
rect 13633 3927 13691 3933
rect 13633 3893 13645 3927
rect 13679 3893 13691 3927
rect 13832 3924 13860 4032
rect 13998 4020 14004 4032
rect 14056 4020 14062 4072
rect 14093 4063 14151 4069
rect 14093 4029 14105 4063
rect 14139 4060 14151 4063
rect 14366 4060 14372 4072
rect 14139 4032 14372 4060
rect 14139 4029 14151 4032
rect 14093 4023 14151 4029
rect 14366 4020 14372 4032
rect 14424 4020 14430 4072
rect 15010 4020 15016 4072
rect 15068 4020 15074 4072
rect 14274 3952 14280 4004
rect 14332 3992 14338 4004
rect 14737 3995 14795 4001
rect 14737 3992 14749 3995
rect 14332 3964 14749 3992
rect 14332 3952 14338 3964
rect 14737 3961 14749 3964
rect 14783 3961 14795 3995
rect 14918 3992 14924 4004
rect 14879 3964 14924 3992
rect 14737 3955 14795 3961
rect 14918 3952 14924 3964
rect 14976 3952 14982 4004
rect 15120 3924 15148 4100
rect 15381 4097 15393 4100
rect 15427 4097 15439 4131
rect 15381 4091 15439 4097
rect 15562 4060 15568 4072
rect 15523 4032 15568 4060
rect 15562 4020 15568 4032
rect 15620 4020 15626 4072
rect 15197 3995 15255 4001
rect 15197 3961 15209 3995
rect 15243 3992 15255 3995
rect 15378 3992 15384 4004
rect 15243 3964 15384 3992
rect 15243 3961 15255 3964
rect 15197 3955 15255 3961
rect 15378 3952 15384 3964
rect 15436 3952 15442 4004
rect 13832 3896 15148 3924
rect 15396 3924 15424 3952
rect 16114 3924 16120 3936
rect 15396 3896 16120 3924
rect 13633 3887 13691 3893
rect 16114 3884 16120 3896
rect 16172 3884 16178 3936
rect 1104 3834 16008 3856
rect 1104 3782 5979 3834
rect 6031 3782 6043 3834
rect 6095 3782 6107 3834
rect 6159 3782 6171 3834
rect 6223 3782 10976 3834
rect 11028 3782 11040 3834
rect 11092 3782 11104 3834
rect 11156 3782 11168 3834
rect 11220 3782 16008 3834
rect 1104 3760 16008 3782
rect 3513 3723 3571 3729
rect 2148 3692 2774 3720
rect 1486 3612 1492 3664
rect 1544 3652 1550 3664
rect 1581 3655 1639 3661
rect 1581 3652 1593 3655
rect 1544 3624 1593 3652
rect 1544 3612 1550 3624
rect 1581 3621 1593 3624
rect 1627 3621 1639 3655
rect 1946 3652 1952 3664
rect 1907 3624 1952 3652
rect 1581 3615 1639 3621
rect 1946 3612 1952 3624
rect 2004 3612 2010 3664
rect 2038 3476 2044 3528
rect 2096 3516 2102 3528
rect 2148 3525 2176 3692
rect 2746 3652 2774 3692
rect 3513 3689 3525 3723
rect 3559 3720 3571 3723
rect 4154 3720 4160 3732
rect 3559 3692 4160 3720
rect 3559 3689 3571 3692
rect 3513 3683 3571 3689
rect 4154 3680 4160 3692
rect 4212 3680 4218 3732
rect 4341 3723 4399 3729
rect 4341 3689 4353 3723
rect 4387 3720 4399 3723
rect 4522 3720 4528 3732
rect 4387 3692 4528 3720
rect 4387 3689 4399 3692
rect 4341 3683 4399 3689
rect 4522 3680 4528 3692
rect 4580 3680 4586 3732
rect 5813 3723 5871 3729
rect 5813 3689 5825 3723
rect 5859 3689 5871 3723
rect 5813 3683 5871 3689
rect 3878 3652 3884 3664
rect 2746 3624 3884 3652
rect 3878 3612 3884 3624
rect 3936 3612 3942 3664
rect 4065 3655 4123 3661
rect 4065 3621 4077 3655
rect 4111 3652 4123 3655
rect 5828 3652 5856 3683
rect 6730 3680 6736 3732
rect 6788 3720 6794 3732
rect 8938 3720 8944 3732
rect 6788 3692 8800 3720
rect 8899 3692 8944 3720
rect 6788 3680 6794 3692
rect 4111 3624 5856 3652
rect 6181 3655 6239 3661
rect 4111 3621 4123 3624
rect 4065 3615 4123 3621
rect 6181 3621 6193 3655
rect 6227 3652 6239 3655
rect 6270 3652 6276 3664
rect 6227 3624 6276 3652
rect 6227 3621 6239 3624
rect 6181 3615 6239 3621
rect 6270 3612 6276 3624
rect 6328 3612 6334 3664
rect 8772 3652 8800 3692
rect 8938 3680 8944 3692
rect 8996 3680 9002 3732
rect 9766 3720 9772 3732
rect 9727 3692 9772 3720
rect 9766 3680 9772 3692
rect 9824 3680 9830 3732
rect 9858 3680 9864 3732
rect 9916 3720 9922 3732
rect 9916 3692 9961 3720
rect 9916 3680 9922 3692
rect 10870 3680 10876 3732
rect 10928 3720 10934 3732
rect 11333 3723 11391 3729
rect 11333 3720 11345 3723
rect 10928 3692 11345 3720
rect 10928 3680 10934 3692
rect 11333 3689 11345 3692
rect 11379 3689 11391 3723
rect 12161 3723 12219 3729
rect 12161 3720 12173 3723
rect 11333 3683 11391 3689
rect 11440 3692 12173 3720
rect 6748 3624 7604 3652
rect 8772 3624 9444 3652
rect 2400 3587 2458 3593
rect 2400 3553 2412 3587
rect 2446 3584 2458 3587
rect 4522 3584 4528 3596
rect 2446 3556 4528 3584
rect 2446 3553 2458 3556
rect 2400 3547 2458 3553
rect 4522 3544 4528 3556
rect 4580 3544 4586 3596
rect 5465 3587 5523 3593
rect 5465 3553 5477 3587
rect 5511 3584 5523 3587
rect 5810 3584 5816 3596
rect 5511 3556 5816 3584
rect 5511 3553 5523 3556
rect 5465 3547 5523 3553
rect 5810 3544 5816 3556
rect 5868 3544 5874 3596
rect 5902 3544 5908 3596
rect 5960 3584 5966 3596
rect 5997 3587 6055 3593
rect 5997 3584 6009 3587
rect 5960 3556 6009 3584
rect 5960 3544 5966 3556
rect 5997 3553 6009 3556
rect 6043 3553 6055 3587
rect 6748 3584 6776 3624
rect 5997 3547 6055 3553
rect 6104 3556 6776 3584
rect 6825 3587 6883 3593
rect 2133 3519 2191 3525
rect 2133 3516 2145 3519
rect 2096 3488 2145 3516
rect 2096 3476 2102 3488
rect 2133 3485 2145 3488
rect 2179 3485 2191 3519
rect 2133 3479 2191 3485
rect 3697 3519 3755 3525
rect 3697 3485 3709 3519
rect 3743 3516 3755 3519
rect 4706 3516 4712 3528
rect 3743 3488 4712 3516
rect 3743 3485 3755 3488
rect 3697 3479 3755 3485
rect 4706 3476 4712 3488
rect 4764 3476 4770 3528
rect 5721 3519 5779 3525
rect 5721 3485 5733 3519
rect 5767 3516 5779 3519
rect 6104 3516 6132 3556
rect 6825 3553 6837 3587
rect 6871 3553 6883 3587
rect 6825 3547 6883 3553
rect 5767 3488 6132 3516
rect 6365 3519 6423 3525
rect 5767 3485 5779 3488
rect 5721 3479 5779 3485
rect 6365 3485 6377 3519
rect 6411 3516 6423 3519
rect 6454 3516 6460 3528
rect 6411 3488 6460 3516
rect 6411 3485 6423 3488
rect 6365 3479 6423 3485
rect 3881 3451 3939 3457
rect 3881 3448 3893 3451
rect 3068 3420 3893 3448
rect 3068 3392 3096 3420
rect 3881 3417 3893 3420
rect 3927 3417 3939 3451
rect 3881 3411 3939 3417
rect 1486 3380 1492 3392
rect 1447 3352 1492 3380
rect 1486 3340 1492 3352
rect 1544 3340 1550 3392
rect 1857 3383 1915 3389
rect 1857 3349 1869 3383
rect 1903 3380 1915 3383
rect 2774 3380 2780 3392
rect 1903 3352 2780 3380
rect 1903 3349 1915 3352
rect 1857 3343 1915 3349
rect 2774 3340 2780 3352
rect 2832 3340 2838 3392
rect 3050 3340 3056 3392
rect 3108 3340 3114 3392
rect 4062 3340 4068 3392
rect 4120 3380 4126 3392
rect 5736 3380 5764 3479
rect 6454 3476 6460 3488
rect 6512 3476 6518 3528
rect 6840 3516 6868 3547
rect 6914 3544 6920 3596
rect 6972 3584 6978 3596
rect 6972 3556 7017 3584
rect 6972 3544 6978 3556
rect 7282 3544 7288 3596
rect 7340 3584 7346 3596
rect 7576 3593 7604 3624
rect 7469 3587 7527 3593
rect 7469 3584 7481 3587
rect 7340 3556 7481 3584
rect 7340 3544 7346 3556
rect 7469 3553 7481 3556
rect 7515 3553 7527 3587
rect 7469 3547 7527 3553
rect 7561 3587 7619 3593
rect 7561 3553 7573 3587
rect 7607 3553 7619 3587
rect 7561 3547 7619 3553
rect 7828 3587 7886 3593
rect 7828 3553 7840 3587
rect 7874 3584 7886 3587
rect 8294 3584 8300 3596
rect 7874 3556 8300 3584
rect 7874 3553 7886 3556
rect 7828 3547 7886 3553
rect 8294 3544 8300 3556
rect 8352 3544 8358 3596
rect 9122 3544 9128 3596
rect 9180 3584 9186 3596
rect 9309 3587 9367 3593
rect 9309 3584 9321 3587
rect 9180 3556 9321 3584
rect 9180 3544 9186 3556
rect 9309 3553 9321 3556
rect 9355 3553 9367 3587
rect 9416 3584 9444 3624
rect 9490 3612 9496 3664
rect 9548 3652 9554 3664
rect 10321 3655 10379 3661
rect 10321 3652 10333 3655
rect 9548 3624 10333 3652
rect 9548 3612 9554 3624
rect 10321 3621 10333 3624
rect 10367 3652 10379 3655
rect 10594 3652 10600 3664
rect 10367 3624 10600 3652
rect 10367 3621 10379 3624
rect 10321 3615 10379 3621
rect 10594 3612 10600 3624
rect 10652 3612 10658 3664
rect 11440 3652 11468 3692
rect 12161 3689 12173 3692
rect 12207 3689 12219 3723
rect 12161 3683 12219 3689
rect 12710 3680 12716 3732
rect 12768 3720 12774 3732
rect 12897 3723 12955 3729
rect 12897 3720 12909 3723
rect 12768 3692 12909 3720
rect 12768 3680 12774 3692
rect 12897 3689 12909 3692
rect 12943 3689 12955 3723
rect 12897 3683 12955 3689
rect 13078 3680 13084 3732
rect 13136 3720 13142 3732
rect 14921 3723 14979 3729
rect 14921 3720 14933 3723
rect 13136 3692 14933 3720
rect 13136 3680 13142 3692
rect 14921 3689 14933 3692
rect 14967 3689 14979 3723
rect 14921 3683 14979 3689
rect 15286 3680 15292 3732
rect 15344 3720 15350 3732
rect 15381 3723 15439 3729
rect 15381 3720 15393 3723
rect 15344 3692 15393 3720
rect 15344 3680 15350 3692
rect 15381 3689 15393 3692
rect 15427 3689 15439 3723
rect 15381 3683 15439 3689
rect 10897 3624 11468 3652
rect 11885 3655 11943 3661
rect 10897 3584 10925 3624
rect 11885 3621 11897 3655
rect 11931 3652 11943 3655
rect 12342 3652 12348 3664
rect 11931 3624 12348 3652
rect 11931 3621 11943 3624
rect 11885 3615 11943 3621
rect 12342 3612 12348 3624
rect 12400 3612 12406 3664
rect 12618 3612 12624 3664
rect 12676 3652 12682 3664
rect 14461 3655 14519 3661
rect 14461 3652 14473 3655
rect 12676 3624 14473 3652
rect 12676 3612 12682 3624
rect 14461 3621 14473 3624
rect 14507 3621 14519 3655
rect 14642 3652 14648 3664
rect 14603 3624 14648 3652
rect 14461 3615 14519 3621
rect 14642 3612 14648 3624
rect 14700 3612 14706 3664
rect 15010 3652 15016 3664
rect 14971 3624 15016 3652
rect 15010 3612 15016 3624
rect 15068 3612 15074 3664
rect 15194 3612 15200 3664
rect 15252 3652 15258 3664
rect 15473 3655 15531 3661
rect 15473 3652 15485 3655
rect 15252 3624 15485 3652
rect 15252 3612 15258 3624
rect 15473 3621 15485 3624
rect 15519 3621 15531 3655
rect 15473 3615 15531 3621
rect 11238 3584 11244 3596
rect 9416 3556 10925 3584
rect 11199 3556 11244 3584
rect 9309 3547 9367 3553
rect 11238 3544 11244 3556
rect 11296 3544 11302 3596
rect 11514 3544 11520 3596
rect 11572 3584 11578 3596
rect 11974 3584 11980 3596
rect 11572 3556 11980 3584
rect 11572 3544 11578 3556
rect 11974 3544 11980 3556
rect 12032 3584 12038 3596
rect 12253 3587 12311 3593
rect 12253 3584 12265 3587
rect 12032 3556 12265 3584
rect 12032 3544 12038 3556
rect 12253 3553 12265 3556
rect 12299 3553 12311 3587
rect 12802 3584 12808 3596
rect 12763 3556 12808 3584
rect 12253 3547 12311 3553
rect 12802 3544 12808 3556
rect 12860 3544 12866 3596
rect 12986 3544 12992 3596
rect 13044 3584 13050 3596
rect 13357 3587 13415 3593
rect 13357 3584 13369 3587
rect 13044 3556 13369 3584
rect 13044 3544 13050 3556
rect 13357 3553 13369 3556
rect 13403 3553 13415 3587
rect 13357 3547 13415 3553
rect 13541 3587 13599 3593
rect 13541 3553 13553 3587
rect 13587 3553 13599 3587
rect 13722 3584 13728 3596
rect 13683 3556 13728 3584
rect 13541 3547 13599 3553
rect 6748 3488 6868 3516
rect 7101 3519 7159 3525
rect 6270 3408 6276 3460
rect 6328 3448 6334 3460
rect 6748 3448 6776 3488
rect 7101 3485 7113 3519
rect 7147 3516 7159 3519
rect 7147 3488 7512 3516
rect 7147 3485 7159 3488
rect 7101 3479 7159 3485
rect 6328 3420 6776 3448
rect 6328 3408 6334 3420
rect 4120 3352 5764 3380
rect 4120 3340 4126 3352
rect 5994 3340 6000 3392
rect 6052 3380 6058 3392
rect 6457 3383 6515 3389
rect 6457 3380 6469 3383
rect 6052 3352 6469 3380
rect 6052 3340 6058 3352
rect 6457 3349 6469 3352
rect 6503 3349 6515 3383
rect 7282 3380 7288 3392
rect 7243 3352 7288 3380
rect 6457 3343 6515 3349
rect 7282 3340 7288 3352
rect 7340 3340 7346 3392
rect 7484 3380 7512 3488
rect 8938 3476 8944 3528
rect 8996 3516 9002 3528
rect 9766 3516 9772 3528
rect 8996 3488 9772 3516
rect 8996 3476 9002 3488
rect 9766 3476 9772 3488
rect 9824 3476 9830 3528
rect 9950 3516 9956 3528
rect 9911 3488 9956 3516
rect 9950 3476 9956 3488
rect 10008 3476 10014 3528
rect 10318 3476 10324 3528
rect 10376 3516 10382 3528
rect 10778 3516 10784 3528
rect 10376 3488 10784 3516
rect 10376 3476 10382 3488
rect 10778 3476 10784 3488
rect 10836 3516 10842 3528
rect 11425 3519 11483 3525
rect 11425 3516 11437 3519
rect 10836 3488 11437 3516
rect 10836 3476 10842 3488
rect 11425 3485 11437 3488
rect 11471 3485 11483 3519
rect 12618 3516 12624 3528
rect 12579 3488 12624 3516
rect 11425 3479 11483 3485
rect 12618 3476 12624 3488
rect 12676 3476 12682 3528
rect 13556 3516 13584 3547
rect 13722 3544 13728 3556
rect 13780 3544 13786 3596
rect 13906 3584 13912 3596
rect 13867 3556 13912 3584
rect 13906 3544 13912 3556
rect 13964 3544 13970 3596
rect 13814 3516 13820 3528
rect 13556 3488 13820 3516
rect 13814 3476 13820 3488
rect 13872 3476 13878 3528
rect 9214 3408 9220 3460
rect 9272 3448 9278 3460
rect 9272 3420 11008 3448
rect 9272 3408 9278 3420
rect 7834 3380 7840 3392
rect 7484 3352 7840 3380
rect 7834 3340 7840 3352
rect 7892 3340 7898 3392
rect 9122 3380 9128 3392
rect 9083 3352 9128 3380
rect 9122 3340 9128 3352
rect 9180 3340 9186 3392
rect 9398 3380 9404 3392
rect 9359 3352 9404 3380
rect 9398 3340 9404 3352
rect 9456 3340 9462 3392
rect 9582 3340 9588 3392
rect 9640 3380 9646 3392
rect 10594 3380 10600 3392
rect 9640 3352 10600 3380
rect 9640 3340 9646 3352
rect 10594 3340 10600 3352
rect 10652 3340 10658 3392
rect 10870 3380 10876 3392
rect 10831 3352 10876 3380
rect 10870 3340 10876 3352
rect 10928 3340 10934 3392
rect 10980 3380 11008 3420
rect 11238 3408 11244 3460
rect 11296 3448 11302 3460
rect 12250 3448 12256 3460
rect 11296 3420 12256 3448
rect 11296 3408 11302 3420
rect 12250 3408 12256 3420
rect 12308 3408 12314 3460
rect 12342 3408 12348 3460
rect 12400 3448 12406 3460
rect 13924 3448 13952 3544
rect 12400 3420 13952 3448
rect 12400 3408 12406 3420
rect 11793 3383 11851 3389
rect 11793 3380 11805 3383
rect 10980 3352 11805 3380
rect 11793 3349 11805 3352
rect 11839 3349 11851 3383
rect 11793 3343 11851 3349
rect 13265 3383 13323 3389
rect 13265 3349 13277 3383
rect 13311 3380 13323 3383
rect 13354 3380 13360 3392
rect 13311 3352 13360 3380
rect 13311 3349 13323 3352
rect 13265 3343 13323 3349
rect 13354 3340 13360 3352
rect 13412 3340 13418 3392
rect 14090 3380 14096 3392
rect 14051 3352 14096 3380
rect 14090 3340 14096 3352
rect 14148 3340 14154 3392
rect 1104 3290 16008 3312
rect 1104 3238 3480 3290
rect 3532 3238 3544 3290
rect 3596 3238 3608 3290
rect 3660 3238 3672 3290
rect 3724 3238 8478 3290
rect 8530 3238 8542 3290
rect 8594 3238 8606 3290
rect 8658 3238 8670 3290
rect 8722 3238 13475 3290
rect 13527 3238 13539 3290
rect 13591 3238 13603 3290
rect 13655 3238 13667 3290
rect 13719 3238 16008 3290
rect 1104 3216 16008 3238
rect 4246 3136 4252 3188
rect 4304 3176 4310 3188
rect 4341 3179 4399 3185
rect 4341 3176 4353 3179
rect 4304 3148 4353 3176
rect 4304 3136 4310 3148
rect 4341 3145 4353 3148
rect 4387 3145 4399 3179
rect 5534 3176 5540 3188
rect 5495 3148 5540 3176
rect 4341 3139 4399 3145
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 8294 3176 8300 3188
rect 8255 3148 8300 3176
rect 8294 3136 8300 3148
rect 8352 3136 8358 3188
rect 9674 3176 9680 3188
rect 8772 3148 9680 3176
rect 1394 3068 1400 3120
rect 1452 3108 1458 3120
rect 2133 3111 2191 3117
rect 2133 3108 2145 3111
rect 1452 3080 2145 3108
rect 1452 3068 1458 3080
rect 2133 3077 2145 3080
rect 2179 3077 2191 3111
rect 2133 3071 2191 3077
rect 2222 3068 2228 3120
rect 2280 3108 2286 3120
rect 2869 3111 2927 3117
rect 2869 3108 2881 3111
rect 2280 3080 2881 3108
rect 2280 3068 2286 3080
rect 2869 3077 2881 3080
rect 2915 3077 2927 3111
rect 2869 3071 2927 3077
rect 5810 3068 5816 3120
rect 5868 3108 5874 3120
rect 6362 3108 6368 3120
rect 5868 3080 6368 3108
rect 5868 3068 5874 3080
rect 1854 3000 1860 3052
rect 1912 3040 1918 3052
rect 2501 3043 2559 3049
rect 2501 3040 2513 3043
rect 1912 3012 2513 3040
rect 1912 3000 1918 3012
rect 2501 3009 2513 3012
rect 2547 3009 2559 3043
rect 2501 3003 2559 3009
rect 2682 3000 2688 3052
rect 2740 3040 2746 3052
rect 3237 3043 3295 3049
rect 3237 3040 3249 3043
rect 2740 3012 3249 3040
rect 2740 3000 2746 3012
rect 3237 3009 3249 3012
rect 3283 3009 3295 3043
rect 3237 3003 3295 3009
rect 3789 3043 3847 3049
rect 3789 3009 3801 3043
rect 3835 3040 3847 3043
rect 4522 3040 4528 3052
rect 3835 3012 4528 3040
rect 3835 3009 3847 3012
rect 3789 3003 3847 3009
rect 4522 3000 4528 3012
rect 4580 3000 4586 3052
rect 5077 3043 5135 3049
rect 5077 3009 5089 3043
rect 5123 3040 5135 3043
rect 5828 3040 5856 3068
rect 5994 3040 6000 3052
rect 5123 3012 5856 3040
rect 5955 3012 6000 3040
rect 5123 3009 5135 3012
rect 5077 3003 5135 3009
rect 5994 3000 6000 3012
rect 6052 3000 6058 3052
rect 6196 3049 6224 3080
rect 6362 3068 6368 3080
rect 6420 3108 6426 3120
rect 6549 3111 6607 3117
rect 6549 3108 6561 3111
rect 6420 3080 6561 3108
rect 6420 3068 6426 3080
rect 6549 3077 6561 3080
rect 6595 3077 6607 3111
rect 8772 3108 8800 3148
rect 9674 3136 9680 3148
rect 9732 3176 9738 3188
rect 9732 3148 12480 3176
rect 9732 3136 9738 3148
rect 6549 3071 6607 3077
rect 7944 3080 8800 3108
rect 7944 3049 7972 3080
rect 9692 3049 9720 3136
rect 11164 3049 11192 3148
rect 11425 3111 11483 3117
rect 11425 3077 11437 3111
rect 11471 3108 11483 3111
rect 11882 3108 11888 3120
rect 11471 3080 11888 3108
rect 11471 3077 11483 3080
rect 11425 3071 11483 3077
rect 11882 3068 11888 3080
rect 11940 3068 11946 3120
rect 11974 3068 11980 3120
rect 12032 3108 12038 3120
rect 12032 3080 12077 3108
rect 12032 3068 12038 3080
rect 6181 3043 6239 3049
rect 6181 3009 6193 3043
rect 6227 3009 6239 3043
rect 6181 3003 6239 3009
rect 7929 3043 7987 3049
rect 7929 3009 7941 3043
rect 7975 3009 7987 3043
rect 7929 3003 7987 3009
rect 9677 3043 9735 3049
rect 9677 3009 9689 3043
rect 9723 3009 9735 3043
rect 9677 3003 9735 3009
rect 11149 3043 11207 3049
rect 11149 3009 11161 3043
rect 11195 3009 11207 3043
rect 11149 3003 11207 3009
rect 12253 3043 12311 3049
rect 12253 3009 12265 3043
rect 12299 3040 12311 3043
rect 12452 3040 12480 3148
rect 14182 3136 14188 3188
rect 14240 3176 14246 3188
rect 14277 3179 14335 3185
rect 14277 3176 14289 3179
rect 14240 3148 14289 3176
rect 14240 3136 14246 3148
rect 14277 3145 14289 3148
rect 14323 3145 14335 3179
rect 14458 3176 14464 3188
rect 14419 3148 14464 3176
rect 14277 3139 14335 3145
rect 14458 3136 14464 3148
rect 14516 3136 14522 3188
rect 12897 3043 12955 3049
rect 12897 3040 12909 3043
rect 12299 3012 12388 3040
rect 12452 3012 12909 3040
rect 12299 3009 12311 3012
rect 12253 3003 12311 3009
rect 1578 2972 1584 2984
rect 1539 2944 1584 2972
rect 1578 2932 1584 2944
rect 1636 2932 1642 2984
rect 2314 2972 2320 2984
rect 2275 2944 2320 2972
rect 2314 2932 2320 2944
rect 2372 2932 2378 2984
rect 2590 2932 2596 2984
rect 2648 2972 2654 2984
rect 3053 2975 3111 2981
rect 3053 2972 3065 2975
rect 2648 2944 3065 2972
rect 2648 2932 2654 2944
rect 3053 2941 3065 2944
rect 3099 2941 3111 2975
rect 3053 2935 3111 2941
rect 3326 2932 3332 2984
rect 3384 2972 3390 2984
rect 3421 2975 3479 2981
rect 3421 2972 3433 2975
rect 3384 2944 3433 2972
rect 3384 2932 3390 2944
rect 3421 2941 3433 2944
rect 3467 2941 3479 2975
rect 3421 2935 3479 2941
rect 3973 2975 4031 2981
rect 3973 2941 3985 2975
rect 4019 2972 4031 2975
rect 4338 2972 4344 2984
rect 4019 2944 4344 2972
rect 4019 2941 4031 2944
rect 3973 2935 4031 2941
rect 4338 2932 4344 2944
rect 4396 2932 4402 2984
rect 4430 2932 4436 2984
rect 4488 2972 4494 2984
rect 4893 2975 4951 2981
rect 4893 2972 4905 2975
rect 4488 2944 4905 2972
rect 4488 2932 4494 2944
rect 4893 2941 4905 2944
rect 4939 2972 4951 2975
rect 5902 2972 5908 2984
rect 4939 2944 5908 2972
rect 4939 2941 4951 2944
rect 4893 2935 4951 2941
rect 5902 2932 5908 2944
rect 5960 2932 5966 2984
rect 7673 2975 7731 2981
rect 7673 2941 7685 2975
rect 7719 2972 7731 2975
rect 7834 2972 7840 2984
rect 7719 2944 7840 2972
rect 7719 2941 7731 2944
rect 7673 2935 7731 2941
rect 7834 2932 7840 2944
rect 7892 2932 7898 2984
rect 8205 2975 8263 2981
rect 8205 2941 8217 2975
rect 8251 2941 8263 2975
rect 8205 2935 8263 2941
rect 566 2864 572 2916
rect 624 2904 630 2916
rect 1397 2907 1455 2913
rect 1397 2904 1409 2907
rect 624 2876 1409 2904
rect 624 2864 630 2876
rect 1397 2873 1409 2876
rect 1443 2873 1455 2907
rect 1397 2867 1455 2873
rect 1949 2907 2007 2913
rect 1949 2873 1961 2907
rect 1995 2873 2007 2907
rect 1949 2867 2007 2873
rect 2685 2907 2743 2913
rect 2685 2873 2697 2907
rect 2731 2904 2743 2907
rect 3786 2904 3792 2916
rect 2731 2876 3792 2904
rect 2731 2873 2743 2876
rect 2685 2867 2743 2873
rect 1026 2796 1032 2848
rect 1084 2836 1090 2848
rect 1857 2839 1915 2845
rect 1857 2836 1869 2839
rect 1084 2808 1869 2836
rect 1084 2796 1090 2808
rect 1857 2805 1869 2808
rect 1903 2805 1915 2839
rect 1964 2836 1992 2867
rect 3786 2864 3792 2876
rect 3844 2864 3850 2916
rect 3881 2907 3939 2913
rect 3881 2873 3893 2907
rect 3927 2904 3939 2907
rect 3927 2876 4476 2904
rect 3927 2873 3939 2876
rect 3881 2867 3939 2873
rect 3510 2836 3516 2848
rect 1964 2808 3516 2836
rect 1857 2799 1915 2805
rect 3510 2796 3516 2808
rect 3568 2796 3574 2848
rect 4448 2845 4476 2876
rect 4706 2864 4712 2916
rect 4764 2904 4770 2916
rect 4764 2876 5396 2904
rect 4764 2864 4770 2876
rect 4433 2839 4491 2845
rect 4433 2805 4445 2839
rect 4479 2805 4491 2839
rect 4798 2836 4804 2848
rect 4759 2808 4804 2836
rect 4433 2799 4491 2805
rect 4798 2796 4804 2808
rect 4856 2796 4862 2848
rect 5258 2836 5264 2848
rect 5219 2808 5264 2836
rect 5258 2796 5264 2808
rect 5316 2796 5322 2848
rect 5368 2836 5396 2876
rect 5534 2864 5540 2916
rect 5592 2904 5598 2916
rect 8220 2904 8248 2935
rect 8478 2932 8484 2984
rect 8536 2972 8542 2984
rect 9122 2972 9128 2984
rect 8536 2944 9128 2972
rect 8536 2932 8542 2944
rect 9122 2932 9128 2944
rect 9180 2932 9186 2984
rect 9766 2932 9772 2984
rect 9824 2972 9830 2984
rect 11241 2975 11299 2981
rect 9824 2944 11008 2972
rect 9824 2932 9830 2944
rect 9030 2904 9036 2916
rect 5592 2876 8064 2904
rect 8220 2876 9036 2904
rect 5592 2864 5598 2876
rect 5905 2839 5963 2845
rect 5905 2836 5917 2839
rect 5368 2808 5917 2836
rect 5905 2805 5917 2808
rect 5951 2836 5963 2839
rect 6638 2836 6644 2848
rect 5951 2808 6644 2836
rect 5951 2805 5963 2808
rect 5905 2799 5963 2805
rect 6638 2796 6644 2808
rect 6696 2796 6702 2848
rect 8036 2845 8064 2876
rect 9030 2864 9036 2876
rect 9088 2864 9094 2916
rect 9432 2907 9490 2913
rect 9432 2873 9444 2907
rect 9478 2904 9490 2907
rect 9478 2876 9812 2904
rect 9478 2873 9490 2876
rect 9432 2867 9490 2873
rect 9784 2845 9812 2876
rect 10226 2864 10232 2916
rect 10284 2904 10290 2916
rect 10284 2876 10732 2904
rect 10284 2864 10290 2876
rect 8021 2839 8079 2845
rect 8021 2805 8033 2839
rect 8067 2805 8079 2839
rect 8021 2799 8079 2805
rect 9769 2839 9827 2845
rect 9769 2805 9781 2839
rect 9815 2836 9827 2839
rect 9950 2836 9956 2848
rect 9815 2808 9956 2836
rect 9815 2805 9827 2808
rect 9769 2799 9827 2805
rect 9950 2796 9956 2808
rect 10008 2836 10014 2848
rect 10594 2836 10600 2848
rect 10008 2808 10600 2836
rect 10008 2796 10014 2808
rect 10594 2796 10600 2808
rect 10652 2796 10658 2848
rect 10704 2836 10732 2876
rect 10778 2864 10784 2916
rect 10836 2904 10842 2916
rect 10882 2907 10940 2913
rect 10882 2904 10894 2907
rect 10836 2876 10894 2904
rect 10836 2864 10842 2876
rect 10882 2873 10894 2876
rect 10928 2873 10940 2907
rect 10980 2904 11008 2944
rect 11241 2941 11253 2975
rect 11287 2972 11299 2975
rect 11606 2972 11612 2984
rect 11287 2944 11612 2972
rect 11287 2941 11299 2944
rect 11241 2935 11299 2941
rect 11256 2904 11284 2935
rect 11606 2932 11612 2944
rect 11664 2932 11670 2984
rect 11698 2932 11704 2984
rect 11756 2972 11762 2984
rect 11793 2975 11851 2981
rect 11793 2972 11805 2975
rect 11756 2944 11805 2972
rect 11756 2932 11762 2944
rect 11793 2941 11805 2944
rect 11839 2941 11851 2975
rect 11793 2935 11851 2941
rect 11716 2904 11744 2932
rect 10980 2876 11284 2904
rect 11348 2876 11744 2904
rect 12360 2904 12388 3012
rect 12897 3009 12909 3012
rect 12943 3009 12955 3043
rect 15565 3043 15623 3049
rect 15565 3040 15577 3043
rect 12897 3003 12955 3009
rect 14568 3012 15577 3040
rect 12437 2975 12495 2981
rect 12437 2941 12449 2975
rect 12483 2972 12495 2975
rect 12483 2944 13308 2972
rect 12483 2941 12495 2944
rect 12437 2935 12495 2941
rect 12526 2904 12532 2916
rect 12360 2876 12532 2904
rect 10882 2867 10940 2873
rect 11348 2836 11376 2876
rect 12526 2864 12532 2876
rect 12584 2904 12590 2916
rect 13142 2907 13200 2913
rect 13142 2904 13154 2907
rect 12584 2876 13154 2904
rect 12584 2864 12590 2876
rect 13142 2873 13154 2876
rect 13188 2873 13200 2907
rect 13280 2904 13308 2944
rect 13446 2932 13452 2984
rect 13504 2972 13510 2984
rect 14568 2981 14596 3012
rect 15565 3009 15577 3012
rect 15611 3009 15623 3043
rect 15565 3003 15623 3009
rect 14553 2975 14611 2981
rect 14553 2972 14565 2975
rect 13504 2944 14565 2972
rect 13504 2932 13510 2944
rect 14553 2941 14565 2944
rect 14599 2941 14611 2975
rect 14553 2935 14611 2941
rect 14734 2932 14740 2984
rect 14792 2972 14798 2984
rect 15013 2975 15071 2981
rect 15013 2972 15025 2975
rect 14792 2944 15025 2972
rect 14792 2932 14798 2944
rect 15013 2941 15025 2944
rect 15059 2941 15071 2975
rect 15013 2935 15071 2941
rect 13998 2904 14004 2916
rect 13280 2876 14004 2904
rect 13142 2867 13200 2873
rect 13998 2864 14004 2876
rect 14056 2864 14062 2916
rect 15289 2907 15347 2913
rect 15289 2873 15301 2907
rect 15335 2904 15347 2907
rect 15470 2904 15476 2916
rect 15335 2876 15476 2904
rect 15335 2873 15347 2876
rect 15289 2867 15347 2873
rect 15470 2864 15476 2876
rect 15528 2864 15534 2916
rect 10704 2808 11376 2836
rect 11882 2796 11888 2848
rect 11940 2836 11946 2848
rect 12345 2839 12403 2845
rect 12345 2836 12357 2839
rect 11940 2808 12357 2836
rect 11940 2796 11946 2808
rect 12345 2805 12357 2808
rect 12391 2805 12403 2839
rect 12802 2836 12808 2848
rect 12763 2808 12808 2836
rect 12345 2799 12403 2805
rect 12802 2796 12808 2808
rect 12860 2796 12866 2848
rect 14734 2836 14740 2848
rect 14695 2808 14740 2836
rect 14734 2796 14740 2808
rect 14792 2796 14798 2848
rect 1104 2746 16008 2768
rect 1104 2694 5979 2746
rect 6031 2694 6043 2746
rect 6095 2694 6107 2746
rect 6159 2694 6171 2746
rect 6223 2694 10976 2746
rect 11028 2694 11040 2746
rect 11092 2694 11104 2746
rect 11156 2694 11168 2746
rect 11220 2694 16008 2746
rect 1104 2672 16008 2694
rect 1765 2635 1823 2641
rect 1765 2632 1777 2635
rect 1596 2604 1777 2632
rect 1596 2573 1624 2604
rect 1765 2601 1777 2604
rect 1811 2601 1823 2635
rect 3510 2632 3516 2644
rect 3471 2604 3516 2632
rect 1765 2595 1823 2601
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 3786 2592 3792 2644
rect 3844 2632 3850 2644
rect 3881 2635 3939 2641
rect 3881 2632 3893 2635
rect 3844 2604 3893 2632
rect 3844 2592 3850 2604
rect 3881 2601 3893 2604
rect 3927 2601 3939 2635
rect 3881 2595 3939 2601
rect 4338 2592 4344 2644
rect 4396 2632 4402 2644
rect 4525 2635 4583 2641
rect 4525 2632 4537 2635
rect 4396 2604 4537 2632
rect 4396 2592 4402 2604
rect 4525 2601 4537 2604
rect 4571 2601 4583 2635
rect 4525 2595 4583 2601
rect 4893 2635 4951 2641
rect 4893 2601 4905 2635
rect 4939 2632 4951 2635
rect 5258 2632 5264 2644
rect 4939 2604 5264 2632
rect 4939 2601 4951 2604
rect 4893 2595 4951 2601
rect 5258 2592 5264 2604
rect 5316 2592 5322 2644
rect 5537 2635 5595 2641
rect 5537 2601 5549 2635
rect 5583 2632 5595 2635
rect 5626 2632 5632 2644
rect 5583 2604 5632 2632
rect 5583 2601 5595 2604
rect 5537 2595 5595 2601
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 5810 2592 5816 2644
rect 5868 2632 5874 2644
rect 5997 2635 6055 2641
rect 5997 2632 6009 2635
rect 5868 2604 6009 2632
rect 5868 2592 5874 2604
rect 5997 2601 6009 2604
rect 6043 2601 6055 2635
rect 5997 2595 6055 2601
rect 6730 2592 6736 2644
rect 6788 2592 6794 2644
rect 7190 2592 7196 2644
rect 7248 2632 7254 2644
rect 9214 2632 9220 2644
rect 7248 2604 7880 2632
rect 9175 2604 9220 2632
rect 7248 2592 7254 2604
rect 1581 2567 1639 2573
rect 1581 2533 1593 2567
rect 1627 2533 1639 2567
rect 1581 2527 1639 2533
rect 2308 2567 2366 2573
rect 2308 2533 2320 2567
rect 2354 2564 2366 2567
rect 2354 2536 3832 2564
rect 2354 2533 2366 2536
rect 2308 2527 2366 2533
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2496 2007 2499
rect 2130 2496 2136 2508
rect 1995 2468 2136 2496
rect 1995 2465 2007 2468
rect 1949 2459 2007 2465
rect 2130 2456 2136 2468
rect 2188 2456 2194 2508
rect 3142 2456 3148 2508
rect 3200 2496 3206 2508
rect 3697 2499 3755 2505
rect 3697 2496 3709 2499
rect 3200 2468 3709 2496
rect 3200 2456 3206 2468
rect 3697 2465 3709 2468
rect 3743 2465 3755 2499
rect 3697 2459 3755 2465
rect 2038 2428 2044 2440
rect 1999 2400 2044 2428
rect 2038 2388 2044 2400
rect 2096 2388 2102 2440
rect 3804 2428 3832 2536
rect 4798 2524 4804 2576
rect 4856 2564 4862 2576
rect 5445 2567 5503 2573
rect 5445 2564 5457 2567
rect 4856 2536 5457 2564
rect 4856 2524 4862 2536
rect 5445 2533 5457 2536
rect 5491 2564 5503 2567
rect 5905 2567 5963 2573
rect 5491 2536 5856 2564
rect 5491 2533 5503 2536
rect 5445 2527 5503 2533
rect 4062 2496 4068 2508
rect 4023 2468 4068 2496
rect 4062 2456 4068 2468
rect 4120 2456 4126 2508
rect 4341 2499 4399 2505
rect 4341 2465 4353 2499
rect 4387 2496 4399 2499
rect 5534 2496 5540 2508
rect 4387 2468 5540 2496
rect 4387 2465 4399 2468
rect 4341 2459 4399 2465
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 5828 2496 5856 2536
rect 5905 2533 5917 2567
rect 5951 2564 5963 2567
rect 6748 2564 6776 2592
rect 5951 2536 6776 2564
rect 7101 2567 7159 2573
rect 5951 2533 5963 2536
rect 5905 2527 5963 2533
rect 7101 2533 7113 2567
rect 7147 2564 7159 2567
rect 7282 2564 7288 2576
rect 7147 2536 7288 2564
rect 7147 2533 7159 2536
rect 7101 2527 7159 2533
rect 7282 2524 7288 2536
rect 7340 2524 7346 2576
rect 7852 2573 7880 2604
rect 9214 2592 9220 2604
rect 9272 2592 9278 2644
rect 9585 2635 9643 2641
rect 9585 2601 9597 2635
rect 9631 2632 9643 2635
rect 10045 2635 10103 2641
rect 10045 2632 10057 2635
rect 9631 2604 10057 2632
rect 9631 2601 9643 2604
rect 9585 2595 9643 2601
rect 10045 2601 10057 2604
rect 10091 2601 10103 2635
rect 10045 2595 10103 2601
rect 10413 2635 10471 2641
rect 10413 2601 10425 2635
rect 10459 2632 10471 2635
rect 10873 2635 10931 2641
rect 10873 2632 10885 2635
rect 10459 2604 10885 2632
rect 10459 2601 10471 2604
rect 10413 2595 10471 2601
rect 10873 2601 10885 2604
rect 10919 2601 10931 2635
rect 10873 2595 10931 2601
rect 11241 2635 11299 2641
rect 11241 2601 11253 2635
rect 11287 2632 11299 2635
rect 11330 2632 11336 2644
rect 11287 2604 11336 2632
rect 11287 2601 11299 2604
rect 11241 2595 11299 2601
rect 11330 2592 11336 2604
rect 11388 2592 11394 2644
rect 12437 2635 12495 2641
rect 12437 2601 12449 2635
rect 12483 2632 12495 2635
rect 12618 2632 12624 2644
rect 12483 2604 12624 2632
rect 12483 2601 12495 2604
rect 12437 2595 12495 2601
rect 12618 2592 12624 2604
rect 12676 2592 12682 2644
rect 12802 2592 12808 2644
rect 12860 2632 12866 2644
rect 13265 2635 13323 2641
rect 13265 2632 13277 2635
rect 12860 2604 13277 2632
rect 12860 2592 12866 2604
rect 13265 2601 13277 2604
rect 13311 2601 13323 2635
rect 13265 2595 13323 2601
rect 13354 2592 13360 2644
rect 13412 2632 13418 2644
rect 14182 2632 14188 2644
rect 13412 2604 13457 2632
rect 14143 2604 14188 2632
rect 13412 2592 13418 2604
rect 14182 2592 14188 2604
rect 14240 2592 14246 2644
rect 7837 2567 7895 2573
rect 7837 2533 7849 2567
rect 7883 2533 7895 2567
rect 8478 2564 8484 2576
rect 7837 2527 7895 2533
rect 7944 2536 8484 2564
rect 6270 2496 6276 2508
rect 5828 2468 6276 2496
rect 6270 2456 6276 2468
rect 6328 2456 6334 2508
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2496 6791 2499
rect 7469 2499 7527 2505
rect 6779 2468 7420 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 4614 2428 4620 2440
rect 3804 2400 4620 2428
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 4982 2428 4988 2440
rect 4943 2400 4988 2428
rect 4982 2388 4988 2400
rect 5040 2388 5046 2440
rect 5169 2431 5227 2437
rect 5169 2397 5181 2431
rect 5215 2428 5227 2431
rect 6181 2431 6239 2437
rect 6181 2428 6193 2431
rect 5215 2400 6193 2428
rect 5215 2397 5227 2400
rect 5169 2391 5227 2397
rect 6181 2397 6193 2400
rect 6227 2428 6239 2431
rect 6362 2428 6368 2440
rect 6227 2400 6368 2428
rect 6227 2397 6239 2400
rect 6181 2391 6239 2397
rect 6362 2388 6368 2400
rect 6420 2388 6426 2440
rect 198 2320 204 2372
rect 256 2360 262 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 256 2332 1409 2360
rect 256 2320 262 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 1397 2323 1455 2329
rect 4798 2320 4804 2372
rect 4856 2360 4862 2372
rect 4856 2332 5580 2360
rect 4856 2320 4862 2332
rect 3421 2295 3479 2301
rect 3421 2261 3433 2295
rect 3467 2292 3479 2295
rect 4154 2292 4160 2304
rect 3467 2264 4160 2292
rect 3467 2261 3479 2264
rect 3421 2255 3479 2261
rect 4154 2252 4160 2264
rect 4212 2252 4218 2304
rect 4249 2295 4307 2301
rect 4249 2261 4261 2295
rect 4295 2292 4307 2295
rect 4338 2292 4344 2304
rect 4295 2264 4344 2292
rect 4295 2261 4307 2264
rect 4249 2255 4307 2261
rect 4338 2252 4344 2264
rect 4396 2252 4402 2304
rect 5552 2292 5580 2332
rect 5626 2320 5632 2372
rect 5684 2360 5690 2372
rect 7285 2363 7343 2369
rect 7285 2360 7297 2363
rect 5684 2332 7297 2360
rect 5684 2320 5690 2332
rect 7285 2329 7297 2332
rect 7331 2329 7343 2363
rect 7392 2360 7420 2468
rect 7469 2465 7481 2499
rect 7515 2496 7527 2499
rect 7944 2496 7972 2536
rect 8478 2524 8484 2536
rect 8536 2524 8542 2576
rect 8772 2536 9352 2564
rect 7515 2468 7972 2496
rect 8389 2499 8447 2505
rect 7515 2465 7527 2468
rect 7469 2459 7527 2465
rect 8389 2465 8401 2499
rect 8435 2496 8447 2499
rect 8772 2496 8800 2536
rect 9048 2508 9076 2536
rect 8435 2468 8800 2496
rect 8435 2465 8447 2468
rect 8389 2459 8447 2465
rect 8846 2456 8852 2508
rect 8904 2496 8910 2508
rect 8941 2499 8999 2505
rect 8941 2496 8953 2499
rect 8904 2468 8953 2496
rect 8904 2456 8910 2468
rect 8941 2465 8953 2468
rect 8987 2465 8999 2499
rect 8941 2459 8999 2465
rect 9030 2456 9036 2508
rect 9088 2456 9094 2508
rect 9324 2496 9352 2536
rect 9398 2524 9404 2576
rect 9456 2564 9462 2576
rect 9677 2567 9735 2573
rect 9677 2564 9689 2567
rect 9456 2536 9689 2564
rect 9456 2524 9462 2536
rect 9677 2533 9689 2536
rect 9723 2533 9735 2567
rect 11885 2567 11943 2573
rect 11885 2564 11897 2567
rect 9677 2527 9735 2533
rect 9784 2536 11897 2564
rect 9784 2496 9812 2536
rect 11885 2533 11897 2536
rect 11931 2533 11943 2567
rect 11885 2527 11943 2533
rect 13170 2524 13176 2576
rect 13228 2564 13234 2576
rect 14277 2567 14335 2573
rect 14277 2564 14289 2567
rect 13228 2536 14289 2564
rect 13228 2524 13234 2536
rect 14277 2533 14289 2536
rect 14323 2564 14335 2567
rect 14734 2564 14740 2576
rect 14323 2536 14740 2564
rect 14323 2533 14335 2536
rect 14277 2527 14335 2533
rect 14734 2524 14740 2536
rect 14792 2524 14798 2576
rect 9324 2468 9812 2496
rect 10505 2499 10563 2505
rect 10505 2465 10517 2499
rect 10551 2496 10563 2499
rect 10870 2496 10876 2508
rect 10551 2468 10876 2496
rect 10551 2465 10563 2468
rect 10505 2459 10563 2465
rect 10870 2456 10876 2468
rect 10928 2456 10934 2508
rect 10980 2468 11468 2496
rect 7650 2428 7656 2440
rect 7611 2400 7656 2428
rect 7650 2388 7656 2400
rect 7708 2388 7714 2440
rect 8294 2388 8300 2440
rect 8352 2428 8358 2440
rect 9769 2431 9827 2437
rect 9769 2428 9781 2431
rect 8352 2400 9781 2428
rect 8352 2388 8358 2400
rect 9769 2397 9781 2400
rect 9815 2397 9827 2431
rect 9769 2391 9827 2397
rect 10594 2388 10600 2440
rect 10652 2428 10658 2440
rect 10652 2400 10697 2428
rect 10652 2388 10658 2400
rect 10778 2388 10784 2440
rect 10836 2428 10842 2440
rect 10980 2428 11008 2468
rect 11330 2428 11336 2440
rect 10836 2400 11008 2428
rect 11291 2400 11336 2428
rect 10836 2388 10842 2400
rect 11330 2388 11336 2400
rect 11388 2388 11394 2440
rect 11440 2437 11468 2468
rect 11974 2456 11980 2508
rect 12032 2496 12038 2508
rect 12529 2499 12587 2505
rect 12529 2496 12541 2499
rect 12032 2468 12541 2496
rect 12032 2456 12038 2468
rect 12529 2465 12541 2468
rect 12575 2465 12587 2499
rect 12529 2459 12587 2465
rect 12710 2456 12716 2508
rect 12768 2496 12774 2508
rect 13909 2499 13967 2505
rect 13909 2496 13921 2499
rect 12768 2468 13921 2496
rect 12768 2456 12774 2468
rect 13909 2465 13921 2468
rect 13955 2496 13967 2499
rect 14090 2496 14096 2508
rect 13955 2468 14096 2496
rect 13955 2465 13967 2468
rect 13909 2459 13967 2465
rect 14090 2456 14096 2468
rect 14148 2456 14154 2508
rect 14826 2496 14832 2508
rect 14787 2468 14832 2496
rect 14826 2456 14832 2468
rect 14884 2456 14890 2508
rect 15470 2496 15476 2508
rect 15431 2468 15476 2496
rect 15470 2456 15476 2468
rect 15528 2456 15534 2508
rect 11425 2431 11483 2437
rect 11425 2397 11437 2431
rect 11471 2397 11483 2431
rect 12618 2428 12624 2440
rect 12579 2400 12624 2428
rect 11425 2391 11483 2397
rect 12618 2388 12624 2400
rect 12676 2388 12682 2440
rect 13541 2431 13599 2437
rect 13541 2397 13553 2431
rect 13587 2397 13599 2431
rect 13541 2391 13599 2397
rect 11790 2360 11796 2372
rect 7392 2332 11796 2360
rect 7285 2323 7343 2329
rect 11790 2320 11796 2332
rect 11848 2320 11854 2372
rect 12069 2363 12127 2369
rect 12069 2329 12081 2363
rect 12115 2360 12127 2363
rect 12434 2360 12440 2372
rect 12115 2332 12440 2360
rect 12115 2329 12127 2332
rect 12069 2323 12127 2329
rect 12434 2320 12440 2332
rect 12492 2320 12498 2372
rect 12894 2360 12900 2372
rect 12855 2332 12900 2360
rect 12894 2320 12900 2332
rect 12952 2320 12958 2372
rect 13556 2360 13584 2391
rect 13998 2388 14004 2440
rect 14056 2428 14062 2440
rect 14553 2431 14611 2437
rect 14553 2428 14565 2431
rect 14056 2400 14565 2428
rect 14056 2388 14062 2400
rect 14553 2397 14565 2400
rect 14599 2428 14611 2431
rect 15102 2428 15108 2440
rect 14599 2400 15108 2428
rect 14599 2397 14611 2400
rect 14553 2391 14611 2397
rect 15102 2388 15108 2400
rect 15160 2388 15166 2440
rect 14274 2360 14280 2372
rect 13556 2332 14280 2360
rect 14274 2320 14280 2332
rect 14332 2320 14338 2372
rect 6641 2295 6699 2301
rect 6641 2292 6653 2295
rect 5552 2264 6653 2292
rect 6641 2261 6653 2264
rect 6687 2261 6699 2295
rect 6641 2255 6699 2261
rect 6730 2252 6736 2304
rect 6788 2292 6794 2304
rect 7009 2295 7067 2301
rect 7009 2292 7021 2295
rect 6788 2264 7021 2292
rect 6788 2252 6794 2264
rect 7009 2261 7021 2264
rect 7055 2261 7067 2295
rect 7009 2255 7067 2261
rect 7098 2252 7104 2304
rect 7156 2292 7162 2304
rect 8113 2295 8171 2301
rect 8113 2292 8125 2295
rect 7156 2264 8125 2292
rect 7156 2252 7162 2264
rect 8113 2261 8125 2264
rect 8159 2261 8171 2295
rect 8113 2255 8171 2261
rect 8849 2295 8907 2301
rect 8849 2261 8861 2295
rect 8895 2292 8907 2295
rect 9306 2292 9312 2304
rect 8895 2264 9312 2292
rect 8895 2261 8907 2264
rect 8849 2255 8907 2261
rect 9306 2252 9312 2264
rect 9364 2252 9370 2304
rect 12250 2252 12256 2304
rect 12308 2292 12314 2304
rect 13817 2295 13875 2301
rect 13817 2292 13829 2295
rect 12308 2264 13829 2292
rect 12308 2252 12314 2264
rect 13817 2261 13829 2264
rect 13863 2261 13875 2295
rect 13817 2255 13875 2261
rect 15657 2295 15715 2301
rect 15657 2261 15669 2295
rect 15703 2292 15715 2295
rect 16942 2292 16948 2304
rect 15703 2264 16948 2292
rect 15703 2261 15715 2264
rect 15657 2255 15715 2261
rect 16942 2252 16948 2264
rect 17000 2252 17006 2304
rect 1104 2202 16008 2224
rect 1104 2150 3480 2202
rect 3532 2150 3544 2202
rect 3596 2150 3608 2202
rect 3660 2150 3672 2202
rect 3724 2150 8478 2202
rect 8530 2150 8542 2202
rect 8594 2150 8606 2202
rect 8658 2150 8670 2202
rect 8722 2150 13475 2202
rect 13527 2150 13539 2202
rect 13591 2150 13603 2202
rect 13655 2150 13667 2202
rect 13719 2150 16008 2202
rect 1104 2128 16008 2150
rect 4982 2048 4988 2100
rect 5040 2088 5046 2100
rect 6546 2088 6552 2100
rect 5040 2060 6552 2088
rect 5040 2048 5046 2060
rect 6546 2048 6552 2060
rect 6604 2048 6610 2100
rect 12618 2088 12624 2100
rect 7944 2060 12624 2088
rect 4154 1980 4160 2032
rect 4212 2020 4218 2032
rect 7944 2020 7972 2060
rect 12618 2048 12624 2060
rect 12676 2048 12682 2100
rect 14642 2020 14648 2032
rect 4212 1992 7972 2020
rect 12406 1992 14648 2020
rect 4212 1980 4218 1992
rect 4062 1912 4068 1964
rect 4120 1952 4126 1964
rect 12406 1952 12434 1992
rect 14642 1980 14648 1992
rect 14700 1980 14706 2032
rect 4120 1924 12434 1952
rect 4120 1912 4126 1924
rect 3602 1844 3608 1896
rect 3660 1884 3666 1896
rect 5350 1884 5356 1896
rect 3660 1856 5356 1884
rect 3660 1844 3666 1856
rect 5350 1844 5356 1856
rect 5408 1844 5414 1896
rect 11882 1844 11888 1896
rect 11940 1884 11946 1896
rect 13814 1884 13820 1896
rect 11940 1856 13820 1884
rect 11940 1844 11946 1856
rect 13814 1844 13820 1856
rect 13872 1844 13878 1896
rect 5994 1436 6000 1488
rect 6052 1476 6058 1488
rect 7650 1476 7656 1488
rect 6052 1448 7656 1476
rect 6052 1436 6058 1448
rect 7650 1436 7656 1448
rect 7708 1436 7714 1488
rect 5166 1368 5172 1420
rect 5224 1408 5230 1420
rect 6730 1408 6736 1420
rect 5224 1380 6736 1408
rect 5224 1368 5230 1380
rect 6730 1368 6736 1380
rect 6788 1368 6794 1420
<< via1 >>
rect 3976 17552 4028 17604
rect 7748 17552 7800 17604
rect 4344 17484 4396 17536
rect 7472 17484 7524 17536
rect 3480 17382 3532 17434
rect 3544 17382 3596 17434
rect 3608 17382 3660 17434
rect 3672 17382 3724 17434
rect 8478 17382 8530 17434
rect 8542 17382 8594 17434
rect 8606 17382 8658 17434
rect 8670 17382 8722 17434
rect 13475 17382 13527 17434
rect 13539 17382 13591 17434
rect 13603 17382 13655 17434
rect 13667 17382 13719 17434
rect 940 17280 992 17332
rect 7104 17280 7156 17332
rect 7380 17280 7432 17332
rect 12624 17280 12676 17332
rect 13912 17280 13964 17332
rect 14832 17280 14884 17332
rect 15016 17323 15068 17332
rect 15016 17289 15025 17323
rect 15025 17289 15059 17323
rect 15059 17289 15068 17323
rect 15016 17280 15068 17289
rect 572 17212 624 17264
rect 1492 17212 1544 17264
rect 2228 17212 2280 17264
rect 4620 17255 4672 17264
rect 4620 17221 4629 17255
rect 4629 17221 4663 17255
rect 4663 17221 4672 17255
rect 4620 17212 4672 17221
rect 5080 17255 5132 17264
rect 5080 17221 5089 17255
rect 5089 17221 5123 17255
rect 5123 17221 5132 17255
rect 5080 17212 5132 17221
rect 5448 17255 5500 17264
rect 5448 17221 5457 17255
rect 5457 17221 5491 17255
rect 5491 17221 5500 17255
rect 5448 17212 5500 17221
rect 5908 17255 5960 17264
rect 5908 17221 5917 17255
rect 5917 17221 5951 17255
rect 5951 17221 5960 17255
rect 5908 17212 5960 17221
rect 6276 17212 6328 17264
rect 6736 17212 6788 17264
rect 1768 17144 1820 17196
rect 7840 17212 7892 17264
rect 9220 17212 9272 17264
rect 12164 17212 12216 17264
rect 14280 17212 14332 17264
rect 3976 17119 4028 17128
rect 3976 17085 3985 17119
rect 3985 17085 4019 17119
rect 4019 17085 4028 17119
rect 3976 17076 4028 17085
rect 7564 17076 7616 17128
rect 9128 17144 9180 17196
rect 11060 17144 11112 17196
rect 8852 17076 8904 17128
rect 1676 17008 1728 17060
rect 2136 17008 2188 17060
rect 2228 17008 2280 17060
rect 2688 17051 2740 17060
rect 2688 17017 2697 17051
rect 2697 17017 2731 17051
rect 2731 17017 2740 17051
rect 2688 17008 2740 17017
rect 2872 17008 2924 17060
rect 4344 17051 4396 17060
rect 4344 17017 4353 17051
rect 4353 17017 4387 17051
rect 4387 17017 4396 17051
rect 4344 17008 4396 17017
rect 4804 17051 4856 17060
rect 4804 17017 4813 17051
rect 4813 17017 4847 17051
rect 4847 17017 4856 17051
rect 4804 17008 4856 17017
rect 5080 17008 5132 17060
rect 5632 17051 5684 17060
rect 5632 17017 5641 17051
rect 5641 17017 5675 17051
rect 5675 17017 5684 17051
rect 5632 17008 5684 17017
rect 5816 17008 5868 17060
rect 6736 17051 6788 17060
rect 6736 17017 6745 17051
rect 6745 17017 6779 17051
rect 6779 17017 6788 17051
rect 6736 17008 6788 17017
rect 7104 17051 7156 17060
rect 7104 17017 7113 17051
rect 7113 17017 7147 17051
rect 7147 17017 7156 17051
rect 7104 17008 7156 17017
rect 7656 17051 7708 17060
rect 5448 16940 5500 16992
rect 7656 17017 7665 17051
rect 7665 17017 7699 17051
rect 7699 17017 7708 17051
rect 7656 17008 7708 17017
rect 8024 17051 8076 17060
rect 8024 17017 8033 17051
rect 8033 17017 8067 17051
rect 8067 17017 8076 17051
rect 8024 17008 8076 17017
rect 8116 17008 8168 17060
rect 8208 16940 8260 16992
rect 9128 17008 9180 17060
rect 10508 17076 10560 17128
rect 12256 17076 12308 17128
rect 9772 17008 9824 17060
rect 11796 17008 11848 17060
rect 11980 17008 12032 17060
rect 9864 16940 9916 16992
rect 10784 16983 10836 16992
rect 10784 16949 10793 16983
rect 10793 16949 10827 16983
rect 10827 16949 10836 16983
rect 10784 16940 10836 16949
rect 11520 16983 11572 16992
rect 11520 16949 11529 16983
rect 11529 16949 11563 16983
rect 11563 16949 11572 16983
rect 11520 16940 11572 16949
rect 12256 16940 12308 16992
rect 13912 17144 13964 17196
rect 13268 17076 13320 17128
rect 12900 17008 12952 17060
rect 12716 16983 12768 16992
rect 12716 16949 12725 16983
rect 12725 16949 12759 16983
rect 12759 16949 12768 16983
rect 12716 16940 12768 16949
rect 12992 16940 13044 16992
rect 13820 16940 13872 16992
rect 14556 17076 14608 17128
rect 14188 16940 14240 16992
rect 15292 16940 15344 16992
rect 5979 16838 6031 16890
rect 6043 16838 6095 16890
rect 6107 16838 6159 16890
rect 6171 16838 6223 16890
rect 10976 16838 11028 16890
rect 11040 16838 11092 16890
rect 11104 16838 11156 16890
rect 11168 16838 11220 16890
rect 1860 16779 1912 16788
rect 1860 16745 1869 16779
rect 1869 16745 1903 16779
rect 1903 16745 1912 16779
rect 1860 16736 1912 16745
rect 2136 16779 2188 16788
rect 2136 16745 2145 16779
rect 2145 16745 2179 16779
rect 2179 16745 2188 16779
rect 2136 16736 2188 16745
rect 1400 16711 1452 16720
rect 1400 16677 1409 16711
rect 1409 16677 1443 16711
rect 1443 16677 1452 16711
rect 1400 16668 1452 16677
rect 2596 16711 2648 16720
rect 2596 16677 2605 16711
rect 2605 16677 2639 16711
rect 2639 16677 2648 16711
rect 3056 16711 3108 16720
rect 2596 16668 2648 16677
rect 3056 16677 3065 16711
rect 3065 16677 3099 16711
rect 3099 16677 3108 16711
rect 3056 16668 3108 16677
rect 3332 16668 3384 16720
rect 3884 16711 3936 16720
rect 3884 16677 3893 16711
rect 3893 16677 3927 16711
rect 3927 16677 3936 16711
rect 3884 16668 3936 16677
rect 4252 16711 4304 16720
rect 4252 16677 4261 16711
rect 4261 16677 4295 16711
rect 4295 16677 4304 16711
rect 4252 16668 4304 16677
rect 5080 16779 5132 16788
rect 5080 16745 5089 16779
rect 5089 16745 5123 16779
rect 5123 16745 5132 16779
rect 5080 16736 5132 16745
rect 1584 16643 1636 16652
rect 1584 16609 1593 16643
rect 1593 16609 1627 16643
rect 1627 16609 1636 16643
rect 1584 16600 1636 16609
rect 1952 16643 2004 16652
rect 1952 16609 1961 16643
rect 1961 16609 1995 16643
rect 1995 16609 2004 16643
rect 1952 16600 2004 16609
rect 2412 16600 2464 16652
rect 3240 16643 3292 16652
rect 3240 16609 3249 16643
rect 3249 16609 3283 16643
rect 3283 16609 3292 16643
rect 3240 16600 3292 16609
rect 3792 16600 3844 16652
rect 3976 16600 4028 16652
rect 4896 16600 4948 16652
rect 8116 16736 8168 16788
rect 8300 16736 8352 16788
rect 5540 16668 5592 16720
rect 6644 16668 6696 16720
rect 11888 16736 11940 16788
rect 13912 16736 13964 16788
rect 14648 16736 14700 16788
rect 16948 16736 17000 16788
rect 5448 16600 5500 16652
rect 12164 16668 12216 16720
rect 12532 16668 12584 16720
rect 8300 16600 8352 16652
rect 8944 16643 8996 16652
rect 8944 16609 8953 16643
rect 8953 16609 8987 16643
rect 8987 16609 8996 16643
rect 8944 16600 8996 16609
rect 2780 16464 2832 16516
rect 2412 16439 2464 16448
rect 2412 16405 2421 16439
rect 2421 16405 2455 16439
rect 2455 16405 2464 16439
rect 2412 16396 2464 16405
rect 6644 16464 6696 16516
rect 6368 16396 6420 16448
rect 8852 16464 8904 16516
rect 9956 16600 10008 16652
rect 10416 16600 10468 16652
rect 11704 16600 11756 16652
rect 13820 16643 13872 16652
rect 13820 16609 13838 16643
rect 13838 16609 13872 16643
rect 13820 16600 13872 16609
rect 14464 16600 14516 16652
rect 14740 16643 14792 16652
rect 14740 16609 14749 16643
rect 14749 16609 14783 16643
rect 14783 16609 14792 16643
rect 14740 16600 14792 16609
rect 15292 16600 15344 16652
rect 15476 16643 15528 16652
rect 15476 16609 15485 16643
rect 15485 16609 15519 16643
rect 15519 16609 15528 16643
rect 15476 16600 15528 16609
rect 9128 16575 9180 16584
rect 9128 16541 9137 16575
rect 9137 16541 9171 16575
rect 9171 16541 9180 16575
rect 9128 16532 9180 16541
rect 14188 16532 14240 16584
rect 7012 16396 7064 16448
rect 10048 16396 10100 16448
rect 10508 16439 10560 16448
rect 10508 16405 10517 16439
rect 10517 16405 10551 16439
rect 10551 16405 10560 16439
rect 10508 16396 10560 16405
rect 10692 16396 10744 16448
rect 11060 16439 11112 16448
rect 11060 16405 11069 16439
rect 11069 16405 11103 16439
rect 11103 16405 11112 16439
rect 11060 16396 11112 16405
rect 11152 16396 11204 16448
rect 12072 16396 12124 16448
rect 13176 16396 13228 16448
rect 13360 16396 13412 16448
rect 16028 16464 16080 16516
rect 15200 16439 15252 16448
rect 15200 16405 15209 16439
rect 15209 16405 15243 16439
rect 15243 16405 15252 16439
rect 15200 16396 15252 16405
rect 3480 16294 3532 16346
rect 3544 16294 3596 16346
rect 3608 16294 3660 16346
rect 3672 16294 3724 16346
rect 8478 16294 8530 16346
rect 8542 16294 8594 16346
rect 8606 16294 8658 16346
rect 8670 16294 8722 16346
rect 13475 16294 13527 16346
rect 13539 16294 13591 16346
rect 13603 16294 13655 16346
rect 13667 16294 13719 16346
rect 2688 16192 2740 16244
rect 2780 16192 2832 16244
rect 3240 16192 3292 16244
rect 3792 16192 3844 16244
rect 3976 16192 4028 16244
rect 4252 16192 4304 16244
rect 2964 16124 3016 16176
rect 2044 15988 2096 16040
rect 2964 15988 3016 16040
rect 4160 16124 4212 16176
rect 4804 16192 4856 16244
rect 5632 16235 5684 16244
rect 5632 16201 5641 16235
rect 5641 16201 5675 16235
rect 5675 16201 5684 16235
rect 5632 16192 5684 16201
rect 5816 16192 5868 16244
rect 6460 16192 6512 16244
rect 7012 16192 7064 16244
rect 7104 16192 7156 16244
rect 7472 16192 7524 16244
rect 7748 16192 7800 16244
rect 8300 16192 8352 16244
rect 9588 16235 9640 16244
rect 9588 16201 9597 16235
rect 9597 16201 9631 16235
rect 9631 16201 9640 16235
rect 9588 16192 9640 16201
rect 3240 16056 3292 16108
rect 3424 16031 3476 16040
rect 3424 15997 3433 16031
rect 3433 15997 3467 16031
rect 3467 15997 3476 16031
rect 3976 16056 4028 16108
rect 3424 15988 3476 15997
rect 2596 15852 2648 15904
rect 2872 15852 2924 15904
rect 3424 15852 3476 15904
rect 3976 15852 4028 15904
rect 5724 16031 5776 16040
rect 4344 15852 4396 15904
rect 5080 15895 5132 15904
rect 5080 15861 5089 15895
rect 5089 15861 5123 15895
rect 5123 15861 5132 15895
rect 5080 15852 5132 15861
rect 5724 15997 5733 16031
rect 5733 15997 5767 16031
rect 5767 15997 5776 16031
rect 5724 15988 5776 15997
rect 6736 16124 6788 16176
rect 8024 16124 8076 16176
rect 10324 16192 10376 16244
rect 10876 16192 10928 16244
rect 6644 16056 6696 16108
rect 7656 16056 7708 16108
rect 8852 16099 8904 16108
rect 7288 15920 7340 15972
rect 7472 16031 7524 16040
rect 7472 15997 7481 16031
rect 7481 15997 7515 16031
rect 7515 15997 7524 16031
rect 7472 15988 7524 15997
rect 7840 15988 7892 16040
rect 8300 16031 8352 16040
rect 7932 15920 7984 15972
rect 8300 15997 8309 16031
rect 8309 15997 8343 16031
rect 8343 15997 8352 16031
rect 8300 15988 8352 15997
rect 8852 16065 8861 16099
rect 8861 16065 8895 16099
rect 8895 16065 8904 16099
rect 8852 16056 8904 16065
rect 11704 16124 11756 16176
rect 10232 16056 10284 16108
rect 10784 16056 10836 16108
rect 11060 16099 11112 16108
rect 11060 16065 11069 16099
rect 11069 16065 11103 16099
rect 11103 16065 11112 16099
rect 11060 16056 11112 16065
rect 11152 16031 11204 16040
rect 8760 15920 8812 15972
rect 9772 15920 9824 15972
rect 9956 15920 10008 15972
rect 11152 15997 11161 16031
rect 11161 15997 11195 16031
rect 11195 15997 11204 16031
rect 11152 15988 11204 15997
rect 11704 15988 11756 16040
rect 11980 16192 12032 16244
rect 13268 16192 13320 16244
rect 15752 16192 15804 16244
rect 11612 15920 11664 15972
rect 5632 15852 5684 15904
rect 5816 15852 5868 15904
rect 7196 15852 7248 15904
rect 9220 15852 9272 15904
rect 9404 15895 9456 15904
rect 9404 15861 9413 15895
rect 9413 15861 9447 15895
rect 9447 15861 9456 15895
rect 9404 15852 9456 15861
rect 10324 15895 10376 15904
rect 10324 15861 10333 15895
rect 10333 15861 10367 15895
rect 10367 15861 10376 15895
rect 10324 15852 10376 15861
rect 11336 15852 11388 15904
rect 11704 15852 11756 15904
rect 12072 15852 12124 15904
rect 13360 15988 13412 16040
rect 12532 15920 12584 15972
rect 12808 15920 12860 15972
rect 13912 15988 13964 16040
rect 14924 15988 14976 16040
rect 14188 15920 14240 15972
rect 15292 15963 15344 15972
rect 15292 15929 15301 15963
rect 15301 15929 15335 15963
rect 15335 15929 15344 15963
rect 15292 15920 15344 15929
rect 13820 15852 13872 15904
rect 14372 15852 14424 15904
rect 15016 15852 15068 15904
rect 5979 15750 6031 15802
rect 6043 15750 6095 15802
rect 6107 15750 6159 15802
rect 6171 15750 6223 15802
rect 10976 15750 11028 15802
rect 11040 15750 11092 15802
rect 11104 15750 11156 15802
rect 11168 15750 11220 15802
rect 1492 15691 1544 15700
rect 1492 15657 1501 15691
rect 1501 15657 1535 15691
rect 1535 15657 1544 15691
rect 1492 15648 1544 15657
rect 1952 15648 2004 15700
rect 2136 15512 2188 15564
rect 3148 15580 3200 15632
rect 5080 15648 5132 15700
rect 7012 15648 7064 15700
rect 7196 15691 7248 15700
rect 7196 15657 7205 15691
rect 7205 15657 7239 15691
rect 7239 15657 7248 15691
rect 7196 15648 7248 15657
rect 7288 15691 7340 15700
rect 7288 15657 7297 15691
rect 7297 15657 7331 15691
rect 7331 15657 7340 15691
rect 7288 15648 7340 15657
rect 7472 15648 7524 15700
rect 8300 15648 8352 15700
rect 9036 15648 9088 15700
rect 9404 15648 9456 15700
rect 9956 15691 10008 15700
rect 9956 15657 9965 15691
rect 9965 15657 9999 15691
rect 9999 15657 10008 15691
rect 9956 15648 10008 15657
rect 10324 15691 10376 15700
rect 10324 15657 10333 15691
rect 10333 15657 10367 15691
rect 10367 15657 10376 15691
rect 10324 15648 10376 15657
rect 10692 15648 10744 15700
rect 11704 15648 11756 15700
rect 11336 15580 11388 15632
rect 12532 15648 12584 15700
rect 13728 15648 13780 15700
rect 14004 15648 14056 15700
rect 2504 15555 2556 15564
rect 2504 15521 2513 15555
rect 2513 15521 2547 15555
rect 2547 15521 2556 15555
rect 2504 15512 2556 15521
rect 6092 15512 6144 15564
rect 6276 15512 6328 15564
rect 6460 15512 6512 15564
rect 6828 15555 6880 15564
rect 6828 15521 6837 15555
rect 6837 15521 6871 15555
rect 6871 15521 6880 15555
rect 6828 15512 6880 15521
rect 8300 15512 8352 15564
rect 8760 15555 8812 15564
rect 8760 15521 8769 15555
rect 8769 15521 8803 15555
rect 8803 15521 8812 15555
rect 8760 15512 8812 15521
rect 9312 15512 9364 15564
rect 9864 15512 9916 15564
rect 10784 15512 10836 15564
rect 1584 15376 1636 15428
rect 204 15308 256 15360
rect 4896 15376 4948 15428
rect 2780 15351 2832 15360
rect 2780 15317 2789 15351
rect 2789 15317 2823 15351
rect 2823 15317 2832 15351
rect 2780 15308 2832 15317
rect 3332 15308 3384 15360
rect 4160 15308 4212 15360
rect 4620 15308 4672 15360
rect 5540 15308 5592 15360
rect 6736 15487 6788 15496
rect 6736 15453 6745 15487
rect 6745 15453 6779 15487
rect 6779 15453 6788 15487
rect 6736 15444 6788 15453
rect 7748 15487 7800 15496
rect 7748 15453 7757 15487
rect 7757 15453 7791 15487
rect 7791 15453 7800 15487
rect 7748 15444 7800 15453
rect 8944 15444 8996 15496
rect 10508 15444 10560 15496
rect 11704 15487 11756 15496
rect 11704 15453 11713 15487
rect 11713 15453 11747 15487
rect 11747 15453 11756 15487
rect 13268 15580 13320 15632
rect 12900 15512 12952 15564
rect 13176 15512 13228 15564
rect 14004 15555 14056 15564
rect 14004 15521 14013 15555
rect 14013 15521 14047 15555
rect 14047 15521 14056 15555
rect 14004 15512 14056 15521
rect 11704 15444 11756 15453
rect 12440 15487 12492 15496
rect 12440 15453 12449 15487
rect 12449 15453 12483 15487
rect 12483 15453 12492 15487
rect 12440 15444 12492 15453
rect 13084 15444 13136 15496
rect 13820 15444 13872 15496
rect 14280 15444 14332 15496
rect 15016 15512 15068 15564
rect 15108 15444 15160 15496
rect 7932 15376 7984 15428
rect 10600 15376 10652 15428
rect 12992 15419 13044 15428
rect 12992 15385 13001 15419
rect 13001 15385 13035 15419
rect 13035 15385 13044 15419
rect 12992 15376 13044 15385
rect 15660 15580 15712 15632
rect 7840 15308 7892 15360
rect 10140 15308 10192 15360
rect 11796 15308 11848 15360
rect 13912 15351 13964 15360
rect 13912 15317 13921 15351
rect 13921 15317 13955 15351
rect 13955 15317 13964 15351
rect 13912 15308 13964 15317
rect 15292 15308 15344 15360
rect 3480 15206 3532 15258
rect 3544 15206 3596 15258
rect 3608 15206 3660 15258
rect 3672 15206 3724 15258
rect 8478 15206 8530 15258
rect 8542 15206 8594 15258
rect 8606 15206 8658 15258
rect 8670 15206 8722 15258
rect 13475 15206 13527 15258
rect 13539 15206 13591 15258
rect 13603 15206 13655 15258
rect 13667 15206 13719 15258
rect 2228 15104 2280 15156
rect 2872 15104 2924 15156
rect 4068 15104 4120 15156
rect 2964 15036 3016 15088
rect 2780 15011 2832 15020
rect 2780 14977 2789 15011
rect 2789 14977 2823 15011
rect 2823 14977 2832 15011
rect 2780 14968 2832 14977
rect 3148 15011 3200 15020
rect 3148 14977 3157 15011
rect 3157 14977 3191 15011
rect 3191 14977 3200 15011
rect 3148 14968 3200 14977
rect 1584 14875 1636 14884
rect 1584 14841 1593 14875
rect 1593 14841 1627 14875
rect 1627 14841 1636 14875
rect 1584 14832 1636 14841
rect 3792 15036 3844 15088
rect 6368 15104 6420 15156
rect 6828 15104 6880 15156
rect 7748 15147 7800 15156
rect 7748 15113 7757 15147
rect 7757 15113 7791 15147
rect 7791 15113 7800 15147
rect 7748 15104 7800 15113
rect 8300 15104 8352 15156
rect 9128 15104 9180 15156
rect 10876 15104 10928 15156
rect 11704 15104 11756 15156
rect 12440 15104 12492 15156
rect 13084 15104 13136 15156
rect 14096 15104 14148 15156
rect 3884 15011 3936 15020
rect 3884 14977 3893 15011
rect 3893 14977 3927 15011
rect 3927 14977 3936 15011
rect 3884 14968 3936 14977
rect 6276 15036 6328 15088
rect 7104 15036 7156 15088
rect 9588 15036 9640 15088
rect 9680 15036 9732 15088
rect 6092 14968 6144 15020
rect 7288 15011 7340 15020
rect 7288 14977 7297 15011
rect 7297 14977 7331 15011
rect 7331 14977 7340 15011
rect 11980 15036 12032 15088
rect 12716 15036 12768 15088
rect 16120 15147 16172 15156
rect 16120 15113 16129 15147
rect 16129 15113 16163 15147
rect 16163 15113 16172 15147
rect 16120 15104 16172 15113
rect 14280 15036 14332 15088
rect 7288 14968 7340 14977
rect 13084 14968 13136 15020
rect 13268 14968 13320 15020
rect 13728 14968 13780 15020
rect 14740 14968 14792 15020
rect 15108 14968 15160 15020
rect 15292 14968 15344 15020
rect 6828 14900 6880 14952
rect 7104 14943 7156 14952
rect 7104 14909 7113 14943
rect 7113 14909 7147 14943
rect 7147 14909 7156 14943
rect 7104 14900 7156 14909
rect 8760 14900 8812 14952
rect 8944 14943 8996 14952
rect 8944 14909 8953 14943
rect 8953 14909 8987 14943
rect 8987 14909 8996 14943
rect 8944 14900 8996 14909
rect 9312 14900 9364 14952
rect 9588 14900 9640 14952
rect 9772 14900 9824 14952
rect 10232 14943 10284 14952
rect 10232 14909 10266 14943
rect 10266 14909 10284 14943
rect 10232 14900 10284 14909
rect 11428 14900 11480 14952
rect 12716 14900 12768 14952
rect 13360 14900 13412 14952
rect 1492 14807 1544 14816
rect 1492 14773 1501 14807
rect 1501 14773 1535 14807
rect 1535 14773 1544 14807
rect 1492 14764 1544 14773
rect 2136 14807 2188 14816
rect 2136 14773 2145 14807
rect 2145 14773 2179 14807
rect 2179 14773 2188 14807
rect 2136 14764 2188 14773
rect 2596 14807 2648 14816
rect 2596 14773 2605 14807
rect 2605 14773 2639 14807
rect 2639 14773 2648 14807
rect 2596 14764 2648 14773
rect 2964 14764 3016 14816
rect 3700 14807 3752 14816
rect 3700 14773 3709 14807
rect 3709 14773 3743 14807
rect 3743 14773 3752 14807
rect 3700 14764 3752 14773
rect 4068 14764 4120 14816
rect 4528 14832 4580 14884
rect 5264 14832 5316 14884
rect 5724 14832 5776 14884
rect 6460 14832 6512 14884
rect 6644 14832 6696 14884
rect 10140 14832 10192 14884
rect 4988 14764 5040 14816
rect 5816 14764 5868 14816
rect 6828 14764 6880 14816
rect 7564 14764 7616 14816
rect 8944 14764 8996 14816
rect 9496 14807 9548 14816
rect 9496 14773 9505 14807
rect 9505 14773 9539 14807
rect 9539 14773 9548 14807
rect 9496 14764 9548 14773
rect 9588 14764 9640 14816
rect 11612 14764 11664 14816
rect 11796 14807 11848 14816
rect 11796 14773 11805 14807
rect 11805 14773 11839 14807
rect 11839 14773 11848 14807
rect 11796 14764 11848 14773
rect 11980 14764 12032 14816
rect 12164 14764 12216 14816
rect 12440 14807 12492 14816
rect 12440 14773 12449 14807
rect 12449 14773 12483 14807
rect 12483 14773 12492 14807
rect 12440 14764 12492 14773
rect 13268 14764 13320 14816
rect 14556 14764 14608 14816
rect 5979 14662 6031 14714
rect 6043 14662 6095 14714
rect 6107 14662 6159 14714
rect 6171 14662 6223 14714
rect 10976 14662 11028 14714
rect 11040 14662 11092 14714
rect 11104 14662 11156 14714
rect 11168 14662 11220 14714
rect 1676 14560 1728 14612
rect 2780 14560 2832 14612
rect 3700 14560 3752 14612
rect 6368 14603 6420 14612
rect 6368 14569 6377 14603
rect 6377 14569 6411 14603
rect 6411 14569 6420 14603
rect 6368 14560 6420 14569
rect 6552 14560 6604 14612
rect 6736 14560 6788 14612
rect 8208 14560 8260 14612
rect 8760 14603 8812 14612
rect 8760 14569 8769 14603
rect 8769 14569 8803 14603
rect 8803 14569 8812 14603
rect 8760 14560 8812 14569
rect 9404 14560 9456 14612
rect 3884 14492 3936 14544
rect 2688 14424 2740 14476
rect 4712 14424 4764 14476
rect 5540 14424 5592 14476
rect 3792 14356 3844 14408
rect 4988 14356 5040 14408
rect 6368 14424 6420 14476
rect 6736 14424 6788 14476
rect 7196 14467 7248 14476
rect 7196 14433 7205 14467
rect 7205 14433 7239 14467
rect 7239 14433 7248 14467
rect 7196 14424 7248 14433
rect 8300 14492 8352 14544
rect 9128 14492 9180 14544
rect 9864 14560 9916 14612
rect 9956 14560 10008 14612
rect 10232 14560 10284 14612
rect 10416 14603 10468 14612
rect 10416 14569 10425 14603
rect 10425 14569 10459 14603
rect 10459 14569 10468 14603
rect 10416 14560 10468 14569
rect 14556 14603 14608 14612
rect 9680 14492 9732 14544
rect 10600 14424 10652 14476
rect 10876 14424 10928 14476
rect 11704 14492 11756 14544
rect 12532 14492 12584 14544
rect 12992 14492 13044 14544
rect 13728 14492 13780 14544
rect 14556 14569 14565 14603
rect 14565 14569 14599 14603
rect 14599 14569 14608 14603
rect 14556 14560 14608 14569
rect 14464 14492 14516 14544
rect 15200 14492 15252 14544
rect 5264 14331 5316 14340
rect 5264 14297 5273 14331
rect 5273 14297 5307 14331
rect 5307 14297 5316 14331
rect 5264 14288 5316 14297
rect 5448 14288 5500 14340
rect 7288 14356 7340 14408
rect 8024 14356 8076 14408
rect 8852 14356 8904 14408
rect 9036 14356 9088 14408
rect 9864 14399 9916 14408
rect 9864 14365 9873 14399
rect 9873 14365 9907 14399
rect 9907 14365 9916 14399
rect 9864 14356 9916 14365
rect 10784 14356 10836 14408
rect 9128 14288 9180 14340
rect 9588 14288 9640 14340
rect 10784 14220 10836 14272
rect 11520 14424 11572 14476
rect 12164 14424 12216 14476
rect 12440 14424 12492 14476
rect 12808 14467 12860 14476
rect 12808 14433 12817 14467
rect 12817 14433 12851 14467
rect 12851 14433 12860 14467
rect 12808 14424 12860 14433
rect 13084 14467 13136 14476
rect 13084 14433 13118 14467
rect 13118 14433 13136 14467
rect 13084 14424 13136 14433
rect 15384 14424 15436 14476
rect 16580 14424 16632 14476
rect 14924 14356 14976 14408
rect 12624 14220 12676 14272
rect 15200 14288 15252 14340
rect 13084 14220 13136 14272
rect 3480 14118 3532 14170
rect 3544 14118 3596 14170
rect 3608 14118 3660 14170
rect 3672 14118 3724 14170
rect 8478 14118 8530 14170
rect 8542 14118 8594 14170
rect 8606 14118 8658 14170
rect 8670 14118 8722 14170
rect 13475 14118 13527 14170
rect 13539 14118 13591 14170
rect 13603 14118 13655 14170
rect 13667 14118 13719 14170
rect 1584 14016 1636 14068
rect 2596 14016 2648 14068
rect 4068 14059 4120 14068
rect 4068 14025 4077 14059
rect 4077 14025 4111 14059
rect 4111 14025 4120 14059
rect 4068 14016 4120 14025
rect 4436 14016 4488 14068
rect 4988 14016 5040 14068
rect 2044 13948 2096 14000
rect 3148 13948 3200 14000
rect 4804 13948 4856 14000
rect 7288 14016 7340 14068
rect 7472 14016 7524 14068
rect 2780 13923 2832 13932
rect 2780 13889 2789 13923
rect 2789 13889 2823 13923
rect 2823 13889 2832 13923
rect 2780 13880 2832 13889
rect 4712 13923 4764 13932
rect 4712 13889 4721 13923
rect 4721 13889 4755 13923
rect 4755 13889 4764 13923
rect 4712 13880 4764 13889
rect 5448 13880 5500 13932
rect 6828 13880 6880 13932
rect 8852 14016 8904 14068
rect 10600 14016 10652 14068
rect 13360 14059 13412 14068
rect 13360 14025 13369 14059
rect 13369 14025 13403 14059
rect 13403 14025 13412 14059
rect 13360 14016 13412 14025
rect 14004 14016 14056 14068
rect 14832 14016 14884 14068
rect 15108 14016 15160 14068
rect 9864 13991 9916 14000
rect 9864 13957 9873 13991
rect 9873 13957 9907 13991
rect 9907 13957 9916 13991
rect 9864 13948 9916 13957
rect 11428 13991 11480 14000
rect 11428 13957 11437 13991
rect 11437 13957 11471 13991
rect 11471 13957 11480 13991
rect 11428 13948 11480 13957
rect 13268 13948 13320 14000
rect 1400 13855 1452 13864
rect 1400 13821 1409 13855
rect 1409 13821 1443 13855
rect 1443 13821 1452 13855
rect 1400 13812 1452 13821
rect 1952 13855 2004 13864
rect 1952 13821 1961 13855
rect 1961 13821 1995 13855
rect 1995 13821 2004 13855
rect 1952 13812 2004 13821
rect 5724 13855 5776 13864
rect 5724 13821 5733 13855
rect 5733 13821 5767 13855
rect 5767 13821 5776 13855
rect 5724 13812 5776 13821
rect 6644 13812 6696 13864
rect 1676 13744 1728 13796
rect 2596 13719 2648 13728
rect 2596 13685 2605 13719
rect 2605 13685 2639 13719
rect 2639 13685 2648 13719
rect 4436 13787 4488 13796
rect 2596 13676 2648 13685
rect 3424 13719 3476 13728
rect 3424 13685 3433 13719
rect 3433 13685 3467 13719
rect 3467 13685 3476 13719
rect 3424 13676 3476 13685
rect 4436 13753 4445 13787
rect 4445 13753 4479 13787
rect 4479 13753 4488 13787
rect 4436 13744 4488 13753
rect 5540 13744 5592 13796
rect 4068 13676 4120 13728
rect 4528 13719 4580 13728
rect 4528 13685 4537 13719
rect 4537 13685 4571 13719
rect 4571 13685 4580 13719
rect 4528 13676 4580 13685
rect 5448 13676 5500 13728
rect 5908 13744 5960 13796
rect 8392 13855 8444 13864
rect 8392 13821 8401 13855
rect 8401 13821 8435 13855
rect 8435 13821 8444 13855
rect 8392 13812 8444 13821
rect 9220 13744 9272 13796
rect 12348 13880 12400 13932
rect 10416 13744 10468 13796
rect 11520 13812 11572 13864
rect 12532 13812 12584 13864
rect 13084 13880 13136 13932
rect 14556 13923 14608 13932
rect 14556 13889 14565 13923
rect 14565 13889 14599 13923
rect 14599 13889 14608 13923
rect 14556 13880 14608 13889
rect 13820 13855 13872 13864
rect 13820 13821 13829 13855
rect 13829 13821 13863 13855
rect 13863 13821 13872 13855
rect 13820 13812 13872 13821
rect 12440 13744 12492 13796
rect 13084 13744 13136 13796
rect 13544 13744 13596 13796
rect 15108 13744 15160 13796
rect 15568 13787 15620 13796
rect 15568 13753 15577 13787
rect 15577 13753 15611 13787
rect 15611 13753 15620 13787
rect 15568 13744 15620 13753
rect 5816 13719 5868 13728
rect 5816 13685 5825 13719
rect 5825 13685 5859 13719
rect 5859 13685 5868 13719
rect 5816 13676 5868 13685
rect 6920 13676 6972 13728
rect 8208 13676 8260 13728
rect 9404 13676 9456 13728
rect 11796 13676 11848 13728
rect 12164 13676 12216 13728
rect 13636 13676 13688 13728
rect 5979 13574 6031 13626
rect 6043 13574 6095 13626
rect 6107 13574 6159 13626
rect 6171 13574 6223 13626
rect 10976 13574 11028 13626
rect 11040 13574 11092 13626
rect 11104 13574 11156 13626
rect 11168 13574 11220 13626
rect 2596 13472 2648 13524
rect 2872 13472 2924 13524
rect 3424 13472 3476 13524
rect 3884 13472 3936 13524
rect 5816 13472 5868 13524
rect 6644 13472 6696 13524
rect 6828 13472 6880 13524
rect 8300 13472 8352 13524
rect 8944 13515 8996 13524
rect 2136 13336 2188 13388
rect 2688 13336 2740 13388
rect 5264 13336 5316 13388
rect 5816 13379 5868 13388
rect 5816 13345 5825 13379
rect 5825 13345 5859 13379
rect 5859 13345 5868 13379
rect 5816 13336 5868 13345
rect 3148 13311 3200 13320
rect 3148 13277 3157 13311
rect 3157 13277 3191 13311
rect 3191 13277 3200 13311
rect 3148 13268 3200 13277
rect 4712 13268 4764 13320
rect 4528 13200 4580 13252
rect 7288 13404 7340 13456
rect 8208 13404 8260 13456
rect 8944 13481 8953 13515
rect 8953 13481 8987 13515
rect 8987 13481 8996 13515
rect 8944 13472 8996 13481
rect 9404 13472 9456 13524
rect 9588 13515 9640 13524
rect 9588 13481 9597 13515
rect 9597 13481 9631 13515
rect 9631 13481 9640 13515
rect 9588 13472 9640 13481
rect 10416 13515 10468 13524
rect 10416 13481 10425 13515
rect 10425 13481 10459 13515
rect 10459 13481 10468 13515
rect 10416 13472 10468 13481
rect 10784 13472 10836 13524
rect 11888 13472 11940 13524
rect 12164 13515 12216 13524
rect 12164 13481 12173 13515
rect 12173 13481 12207 13515
rect 12207 13481 12216 13515
rect 12164 13472 12216 13481
rect 12440 13472 12492 13524
rect 13544 13515 13596 13524
rect 13544 13481 13553 13515
rect 13553 13481 13587 13515
rect 13587 13481 13596 13515
rect 13544 13472 13596 13481
rect 13636 13472 13688 13524
rect 14004 13472 14056 13524
rect 14740 13472 14792 13524
rect 15108 13472 15160 13524
rect 15384 13515 15436 13524
rect 15384 13481 15393 13515
rect 15393 13481 15427 13515
rect 15427 13481 15436 13515
rect 15384 13472 15436 13481
rect 15568 13472 15620 13524
rect 11428 13404 11480 13456
rect 11520 13447 11572 13456
rect 11520 13413 11538 13447
rect 11538 13413 11572 13447
rect 11520 13404 11572 13413
rect 7380 13336 7432 13388
rect 10600 13336 10652 13388
rect 6184 13268 6236 13320
rect 1584 13132 1636 13184
rect 9772 13268 9824 13320
rect 10416 13268 10468 13320
rect 6552 13132 6604 13184
rect 6644 13132 6696 13184
rect 7564 13132 7616 13184
rect 11796 13311 11848 13320
rect 11796 13277 11805 13311
rect 11805 13277 11839 13311
rect 11839 13277 11848 13311
rect 11796 13268 11848 13277
rect 12256 13404 12308 13456
rect 14372 13447 14424 13456
rect 14372 13413 14381 13447
rect 14381 13413 14415 13447
rect 14415 13413 14424 13447
rect 14372 13404 14424 13413
rect 13360 13336 13412 13388
rect 15292 13336 15344 13388
rect 15660 13379 15712 13388
rect 15660 13345 15669 13379
rect 15669 13345 15703 13379
rect 15703 13345 15712 13379
rect 15660 13336 15712 13345
rect 12716 13311 12768 13320
rect 12716 13277 12725 13311
rect 12725 13277 12759 13311
rect 12759 13277 12768 13311
rect 12716 13268 12768 13277
rect 12992 13311 13044 13320
rect 12992 13277 13001 13311
rect 13001 13277 13035 13311
rect 13035 13277 13044 13311
rect 12992 13268 13044 13277
rect 13084 13268 13136 13320
rect 13268 13268 13320 13320
rect 13636 13200 13688 13252
rect 10232 13132 10284 13184
rect 11888 13132 11940 13184
rect 12072 13132 12124 13184
rect 12900 13132 12952 13184
rect 13084 13132 13136 13184
rect 14740 13175 14792 13184
rect 14740 13141 14749 13175
rect 14749 13141 14783 13175
rect 14783 13141 14792 13175
rect 14740 13132 14792 13141
rect 3480 13030 3532 13082
rect 3544 13030 3596 13082
rect 3608 13030 3660 13082
rect 3672 13030 3724 13082
rect 8478 13030 8530 13082
rect 8542 13030 8594 13082
rect 8606 13030 8658 13082
rect 8670 13030 8722 13082
rect 13475 13030 13527 13082
rect 13539 13030 13591 13082
rect 13603 13030 13655 13082
rect 13667 13030 13719 13082
rect 1676 12928 1728 12980
rect 3148 12928 3200 12980
rect 1400 12903 1452 12912
rect 1400 12869 1409 12903
rect 1409 12869 1443 12903
rect 1443 12869 1452 12903
rect 1400 12860 1452 12869
rect 2872 12860 2924 12912
rect 3976 12928 4028 12980
rect 4712 12971 4764 12980
rect 4712 12937 4721 12971
rect 4721 12937 4755 12971
rect 4755 12937 4764 12971
rect 4712 12928 4764 12937
rect 5724 12928 5776 12980
rect 7840 12928 7892 12980
rect 9772 12971 9824 12980
rect 5540 12860 5592 12912
rect 6276 12860 6328 12912
rect 6828 12860 6880 12912
rect 1584 12767 1636 12776
rect 1584 12733 1593 12767
rect 1593 12733 1627 12767
rect 1627 12733 1636 12767
rect 1584 12724 1636 12733
rect 2780 12724 2832 12776
rect 4344 12792 4396 12844
rect 6000 12835 6052 12844
rect 6000 12801 6009 12835
rect 6009 12801 6043 12835
rect 6043 12801 6052 12835
rect 6000 12792 6052 12801
rect 6184 12835 6236 12844
rect 6184 12801 6193 12835
rect 6193 12801 6227 12835
rect 6227 12801 6236 12835
rect 9772 12937 9781 12971
rect 9781 12937 9815 12971
rect 9815 12937 9824 12971
rect 9772 12928 9824 12937
rect 11704 12971 11756 12980
rect 11704 12937 11713 12971
rect 11713 12937 11747 12971
rect 11747 12937 11756 12971
rect 11704 12928 11756 12937
rect 11888 12928 11940 12980
rect 12900 12928 12952 12980
rect 6184 12792 6236 12801
rect 5816 12724 5868 12776
rect 6368 12724 6420 12776
rect 10232 12860 10284 12912
rect 11520 12860 11572 12912
rect 13820 12928 13872 12980
rect 14372 12971 14424 12980
rect 14372 12937 14381 12971
rect 14381 12937 14415 12971
rect 14415 12937 14424 12971
rect 14372 12928 14424 12937
rect 15660 12971 15712 12980
rect 15660 12937 15669 12971
rect 15669 12937 15703 12971
rect 15703 12937 15712 12971
rect 15660 12928 15712 12937
rect 8944 12724 8996 12776
rect 11428 12724 11480 12776
rect 11520 12724 11572 12776
rect 11612 12724 11664 12776
rect 2412 12588 2464 12640
rect 2688 12588 2740 12640
rect 2872 12631 2924 12640
rect 2872 12597 2881 12631
rect 2881 12597 2915 12631
rect 2915 12597 2924 12631
rect 3424 12656 3476 12708
rect 4160 12656 4212 12708
rect 6828 12699 6880 12708
rect 6828 12665 6837 12699
rect 6837 12665 6871 12699
rect 6871 12665 6880 12699
rect 6828 12656 6880 12665
rect 7564 12656 7616 12708
rect 7748 12699 7800 12708
rect 7748 12665 7757 12699
rect 7757 12665 7791 12699
rect 7791 12665 7800 12699
rect 7748 12656 7800 12665
rect 2872 12588 2924 12597
rect 4436 12588 4488 12640
rect 5540 12631 5592 12640
rect 5540 12597 5549 12631
rect 5549 12597 5583 12631
rect 5583 12597 5592 12631
rect 5540 12588 5592 12597
rect 7104 12588 7156 12640
rect 7288 12631 7340 12640
rect 7288 12597 7297 12631
rect 7297 12597 7331 12631
rect 7331 12597 7340 12631
rect 7288 12588 7340 12597
rect 7840 12588 7892 12640
rect 11336 12656 11388 12708
rect 12532 12724 12584 12776
rect 15200 12860 15252 12912
rect 12716 12792 12768 12844
rect 13360 12835 13412 12844
rect 13360 12801 13369 12835
rect 13369 12801 13403 12835
rect 13403 12801 13412 12835
rect 13360 12792 13412 12801
rect 15476 12792 15528 12844
rect 14832 12724 14884 12776
rect 15108 12724 15160 12776
rect 12900 12699 12952 12708
rect 10140 12631 10192 12640
rect 10140 12597 10149 12631
rect 10149 12597 10183 12631
rect 10183 12597 10192 12631
rect 10140 12588 10192 12597
rect 10232 12631 10284 12640
rect 10232 12597 10241 12631
rect 10241 12597 10275 12631
rect 10275 12597 10284 12631
rect 10232 12588 10284 12597
rect 10600 12588 10652 12640
rect 12900 12665 12909 12699
rect 12909 12665 12943 12699
rect 12943 12665 12952 12699
rect 12900 12656 12952 12665
rect 12992 12631 13044 12640
rect 12992 12597 13001 12631
rect 13001 12597 13035 12631
rect 13035 12597 13044 12631
rect 14188 12656 14240 12708
rect 12992 12588 13044 12597
rect 5979 12486 6031 12538
rect 6043 12486 6095 12538
rect 6107 12486 6159 12538
rect 6171 12486 6223 12538
rect 10976 12486 11028 12538
rect 11040 12486 11092 12538
rect 11104 12486 11156 12538
rect 11168 12486 11220 12538
rect 3424 12427 3476 12436
rect 3424 12393 3433 12427
rect 3433 12393 3467 12427
rect 3467 12393 3476 12427
rect 3424 12384 3476 12393
rect 3976 12427 4028 12436
rect 3976 12393 3985 12427
rect 3985 12393 4019 12427
rect 4019 12393 4028 12427
rect 3976 12384 4028 12393
rect 4804 12427 4856 12436
rect 4804 12393 4813 12427
rect 4813 12393 4847 12427
rect 4847 12393 4856 12427
rect 4804 12384 4856 12393
rect 5540 12384 5592 12436
rect 7656 12384 7708 12436
rect 8944 12427 8996 12436
rect 1860 12248 1912 12300
rect 2780 12316 2832 12368
rect 2320 12291 2372 12300
rect 2320 12257 2354 12291
rect 2354 12257 2372 12291
rect 2320 12248 2372 12257
rect 7748 12316 7800 12368
rect 8944 12393 8953 12427
rect 8953 12393 8987 12427
rect 8987 12393 8996 12427
rect 8944 12384 8996 12393
rect 10416 12384 10468 12436
rect 10600 12427 10652 12436
rect 10600 12393 10609 12427
rect 10609 12393 10643 12427
rect 10643 12393 10652 12427
rect 10600 12384 10652 12393
rect 10048 12316 10100 12368
rect 11612 12384 11664 12436
rect 12716 12384 12768 12436
rect 5540 12248 5592 12300
rect 6184 12248 6236 12300
rect 6460 12248 6512 12300
rect 6276 12180 6328 12232
rect 6644 12223 6696 12232
rect 6644 12189 6653 12223
rect 6653 12189 6687 12223
rect 6687 12189 6696 12223
rect 6644 12180 6696 12189
rect 8300 12248 8352 12300
rect 8944 12248 8996 12300
rect 5356 12112 5408 12164
rect 1492 12087 1544 12096
rect 1492 12053 1501 12087
rect 1501 12053 1535 12087
rect 1535 12053 1544 12087
rect 1492 12044 1544 12053
rect 2688 12044 2740 12096
rect 4804 12044 4856 12096
rect 5172 12044 5224 12096
rect 6276 12087 6328 12096
rect 6276 12053 6285 12087
rect 6285 12053 6319 12087
rect 6319 12053 6328 12087
rect 6276 12044 6328 12053
rect 7104 12044 7156 12096
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 10416 12180 10468 12232
rect 14004 12316 14056 12368
rect 14556 12316 14608 12368
rect 11520 12291 11572 12300
rect 11520 12257 11554 12291
rect 11554 12257 11572 12291
rect 11520 12248 11572 12257
rect 14924 12248 14976 12300
rect 15108 12248 15160 12300
rect 11244 12223 11296 12232
rect 11244 12189 11253 12223
rect 11253 12189 11287 12223
rect 11287 12189 11296 12223
rect 11244 12180 11296 12189
rect 12808 12180 12860 12232
rect 10784 12044 10836 12096
rect 11060 12087 11112 12096
rect 11060 12053 11069 12087
rect 11069 12053 11103 12087
rect 11103 12053 11112 12087
rect 11060 12044 11112 12053
rect 11428 12044 11480 12096
rect 3480 11942 3532 11994
rect 3544 11942 3596 11994
rect 3608 11942 3660 11994
rect 3672 11942 3724 11994
rect 8478 11942 8530 11994
rect 8542 11942 8594 11994
rect 8606 11942 8658 11994
rect 8670 11942 8722 11994
rect 13475 11942 13527 11994
rect 13539 11942 13591 11994
rect 13603 11942 13655 11994
rect 13667 11942 13719 11994
rect 3332 11840 3384 11892
rect 4344 11840 4396 11892
rect 4436 11840 4488 11892
rect 4804 11840 4856 11892
rect 9680 11840 9732 11892
rect 10232 11840 10284 11892
rect 2780 11772 2832 11824
rect 5540 11815 5592 11824
rect 5540 11781 5549 11815
rect 5549 11781 5583 11815
rect 5583 11781 5592 11815
rect 5540 11772 5592 11781
rect 3792 11704 3844 11756
rect 5172 11747 5224 11756
rect 5172 11713 5181 11747
rect 5181 11713 5215 11747
rect 5215 11713 5224 11747
rect 5172 11704 5224 11713
rect 5356 11747 5408 11756
rect 5356 11713 5365 11747
rect 5365 11713 5399 11747
rect 5399 11713 5408 11747
rect 5356 11704 5408 11713
rect 6460 11747 6512 11756
rect 6460 11713 6469 11747
rect 6469 11713 6503 11747
rect 6503 11713 6512 11747
rect 6460 11704 6512 11713
rect 2688 11636 2740 11688
rect 2780 11679 2832 11688
rect 2780 11645 2789 11679
rect 2789 11645 2823 11679
rect 2823 11645 2832 11679
rect 5724 11679 5776 11688
rect 2780 11636 2832 11645
rect 5724 11645 5733 11679
rect 5733 11645 5767 11679
rect 5767 11645 5776 11679
rect 5724 11636 5776 11645
rect 6368 11636 6420 11688
rect 8208 11704 8260 11756
rect 10140 11772 10192 11824
rect 11244 11772 11296 11824
rect 11796 11772 11848 11824
rect 7932 11636 7984 11688
rect 8116 11636 8168 11688
rect 9772 11636 9824 11688
rect 10232 11704 10284 11756
rect 11520 11704 11572 11756
rect 11060 11636 11112 11688
rect 11428 11636 11480 11688
rect 2320 11500 2372 11552
rect 3148 11500 3200 11552
rect 4160 11568 4212 11620
rect 5264 11568 5316 11620
rect 6460 11568 6512 11620
rect 6644 11568 6696 11620
rect 6920 11568 6972 11620
rect 10508 11568 10560 11620
rect 10692 11568 10744 11620
rect 3884 11543 3936 11552
rect 3884 11509 3893 11543
rect 3893 11509 3927 11543
rect 3927 11509 3936 11543
rect 3884 11500 3936 11509
rect 4252 11543 4304 11552
rect 4252 11509 4261 11543
rect 4261 11509 4295 11543
rect 4295 11509 4304 11543
rect 4252 11500 4304 11509
rect 4344 11543 4396 11552
rect 4344 11509 4353 11543
rect 4353 11509 4387 11543
rect 4387 11509 4396 11543
rect 4344 11500 4396 11509
rect 5448 11500 5500 11552
rect 7748 11500 7800 11552
rect 7932 11543 7984 11552
rect 7932 11509 7941 11543
rect 7941 11509 7975 11543
rect 7975 11509 7984 11543
rect 8300 11543 8352 11552
rect 7932 11500 7984 11509
rect 8300 11509 8309 11543
rect 8309 11509 8343 11543
rect 8343 11509 8352 11543
rect 8300 11500 8352 11509
rect 8392 11500 8444 11552
rect 9220 11500 9272 11552
rect 9588 11543 9640 11552
rect 9588 11509 9597 11543
rect 9597 11509 9631 11543
rect 9631 11509 9640 11543
rect 9588 11500 9640 11509
rect 10784 11500 10836 11552
rect 12532 11500 12584 11552
rect 12716 11500 12768 11552
rect 5979 11398 6031 11450
rect 6043 11398 6095 11450
rect 6107 11398 6159 11450
rect 6171 11398 6223 11450
rect 10976 11398 11028 11450
rect 11040 11398 11092 11450
rect 11104 11398 11156 11450
rect 11168 11398 11220 11450
rect 1860 11339 1912 11348
rect 1860 11305 1869 11339
rect 1869 11305 1903 11339
rect 1903 11305 1912 11339
rect 1860 11296 1912 11305
rect 3884 11296 3936 11348
rect 4252 11296 4304 11348
rect 5448 11296 5500 11348
rect 7104 11339 7156 11348
rect 7104 11305 7113 11339
rect 7113 11305 7147 11339
rect 7147 11305 7156 11339
rect 7104 11296 7156 11305
rect 7288 11296 7340 11348
rect 7656 11339 7708 11348
rect 7656 11305 7665 11339
rect 7665 11305 7699 11339
rect 7699 11305 7708 11339
rect 7656 11296 7708 11305
rect 10048 11296 10100 11348
rect 10508 11296 10560 11348
rect 14648 11296 14700 11348
rect 2320 11228 2372 11280
rect 1584 11203 1636 11212
rect 1584 11169 1593 11203
rect 1593 11169 1627 11203
rect 1627 11169 1636 11203
rect 1584 11160 1636 11169
rect 2320 11135 2372 11144
rect 2320 11101 2329 11135
rect 2329 11101 2363 11135
rect 2363 11101 2372 11135
rect 2320 11092 2372 11101
rect 3332 11228 3384 11280
rect 3976 11160 4028 11212
rect 5540 11160 5592 11212
rect 5724 11203 5776 11212
rect 5724 11169 5733 11203
rect 5733 11169 5767 11203
rect 5767 11169 5776 11203
rect 5724 11160 5776 11169
rect 3148 11092 3200 11144
rect 6276 11228 6328 11280
rect 12900 11228 12952 11280
rect 6828 11160 6880 11212
rect 8024 11160 8076 11212
rect 8852 11160 8904 11212
rect 9588 11160 9640 11212
rect 10048 11160 10100 11212
rect 11520 11160 11572 11212
rect 12164 11160 12216 11212
rect 14188 11160 14240 11212
rect 6000 11135 6052 11144
rect 1400 11067 1452 11076
rect 1400 11033 1409 11067
rect 1409 11033 1443 11067
rect 1443 11033 1452 11067
rect 1400 11024 1452 11033
rect 3792 11024 3844 11076
rect 6000 11101 6009 11135
rect 6009 11101 6043 11135
rect 6043 11101 6052 11135
rect 6000 11092 6052 11101
rect 6920 11092 6972 11144
rect 7748 11092 7800 11144
rect 7288 11024 7340 11076
rect 8208 11024 8260 11076
rect 8944 11092 8996 11144
rect 9680 11135 9732 11144
rect 9680 11101 9689 11135
rect 9689 11101 9723 11135
rect 9723 11101 9732 11135
rect 9680 11092 9732 11101
rect 11888 11092 11940 11144
rect 12992 11135 13044 11144
rect 12992 11101 13001 11135
rect 13001 11101 13035 11135
rect 13035 11101 13044 11135
rect 12992 11092 13044 11101
rect 10140 11067 10192 11076
rect 10140 11033 10149 11067
rect 10149 11033 10183 11067
rect 10183 11033 10192 11067
rect 10140 11024 10192 11033
rect 10324 11024 10376 11076
rect 10784 11024 10836 11076
rect 2872 10999 2924 11008
rect 2872 10965 2881 10999
rect 2881 10965 2915 10999
rect 2915 10965 2924 10999
rect 2872 10956 2924 10965
rect 6920 10956 6972 11008
rect 7104 10956 7156 11008
rect 7932 10999 7984 11008
rect 7932 10965 7941 10999
rect 7941 10965 7975 10999
rect 7975 10965 7984 10999
rect 7932 10956 7984 10965
rect 9128 10956 9180 11008
rect 11796 11024 11848 11076
rect 11612 10999 11664 11008
rect 11612 10965 11621 10999
rect 11621 10965 11655 10999
rect 11655 10965 11664 10999
rect 11612 10956 11664 10965
rect 3480 10854 3532 10906
rect 3544 10854 3596 10906
rect 3608 10854 3660 10906
rect 3672 10854 3724 10906
rect 8478 10854 8530 10906
rect 8542 10854 8594 10906
rect 8606 10854 8658 10906
rect 8670 10854 8722 10906
rect 13475 10854 13527 10906
rect 13539 10854 13591 10906
rect 13603 10854 13655 10906
rect 13667 10854 13719 10906
rect 1584 10752 1636 10804
rect 2320 10752 2372 10804
rect 3976 10795 4028 10804
rect 3976 10761 3985 10795
rect 3985 10761 4019 10795
rect 4019 10761 4028 10795
rect 3976 10752 4028 10761
rect 4344 10752 4396 10804
rect 8208 10752 8260 10804
rect 9680 10752 9732 10804
rect 10784 10752 10836 10804
rect 12624 10752 12676 10804
rect 2688 10659 2740 10668
rect 2688 10625 2697 10659
rect 2697 10625 2731 10659
rect 2731 10625 2740 10659
rect 2688 10616 2740 10625
rect 2872 10548 2924 10600
rect 7840 10684 7892 10736
rect 5540 10616 5592 10668
rect 6000 10659 6052 10668
rect 6000 10625 6009 10659
rect 6009 10625 6043 10659
rect 6043 10625 6052 10659
rect 6000 10616 6052 10625
rect 7748 10616 7800 10668
rect 9128 10659 9180 10668
rect 9128 10625 9137 10659
rect 9137 10625 9171 10659
rect 9171 10625 9180 10659
rect 9128 10616 9180 10625
rect 12072 10684 12124 10736
rect 12992 10752 13044 10804
rect 13912 10752 13964 10804
rect 14188 10795 14240 10804
rect 14188 10761 14197 10795
rect 14197 10761 14231 10795
rect 14231 10761 14240 10795
rect 14188 10752 14240 10761
rect 10232 10616 10284 10668
rect 10508 10659 10560 10668
rect 10508 10625 10517 10659
rect 10517 10625 10551 10659
rect 10551 10625 10560 10659
rect 10508 10616 10560 10625
rect 11796 10616 11848 10668
rect 12256 10659 12308 10668
rect 12256 10625 12265 10659
rect 12265 10625 12299 10659
rect 12299 10625 12308 10659
rect 12256 10616 12308 10625
rect 3884 10480 3936 10532
rect 5540 10480 5592 10532
rect 3332 10455 3384 10464
rect 3332 10421 3341 10455
rect 3341 10421 3375 10455
rect 3375 10421 3384 10455
rect 3332 10412 3384 10421
rect 4896 10412 4948 10464
rect 6644 10480 6696 10532
rect 7932 10548 7984 10600
rect 8576 10548 8628 10600
rect 9220 10591 9272 10600
rect 9220 10557 9229 10591
rect 9229 10557 9263 10591
rect 9263 10557 9272 10591
rect 9220 10548 9272 10557
rect 11060 10548 11112 10600
rect 11428 10480 11480 10532
rect 12900 10480 12952 10532
rect 13360 10480 13412 10532
rect 5816 10455 5868 10464
rect 5816 10421 5825 10455
rect 5825 10421 5859 10455
rect 5859 10421 5868 10455
rect 6552 10455 6604 10464
rect 5816 10412 5868 10421
rect 6552 10421 6561 10455
rect 6561 10421 6595 10455
rect 6595 10421 6604 10455
rect 6552 10412 6604 10421
rect 7196 10455 7248 10464
rect 7196 10421 7205 10455
rect 7205 10421 7239 10455
rect 7239 10421 7248 10455
rect 7196 10412 7248 10421
rect 7748 10455 7800 10464
rect 7748 10421 7757 10455
rect 7757 10421 7791 10455
rect 7791 10421 7800 10455
rect 7748 10412 7800 10421
rect 8392 10412 8444 10464
rect 9128 10412 9180 10464
rect 9864 10455 9916 10464
rect 9864 10421 9873 10455
rect 9873 10421 9907 10455
rect 9907 10421 9916 10455
rect 9864 10412 9916 10421
rect 10048 10412 10100 10464
rect 10784 10412 10836 10464
rect 11336 10412 11388 10464
rect 12440 10412 12492 10464
rect 13176 10412 13228 10464
rect 14464 10455 14516 10464
rect 14464 10421 14473 10455
rect 14473 10421 14507 10455
rect 14507 10421 14516 10455
rect 14464 10412 14516 10421
rect 15108 10412 15160 10464
rect 5979 10310 6031 10362
rect 6043 10310 6095 10362
rect 6107 10310 6159 10362
rect 6171 10310 6223 10362
rect 10976 10310 11028 10362
rect 11040 10310 11092 10362
rect 11104 10310 11156 10362
rect 11168 10310 11220 10362
rect 3332 10208 3384 10260
rect 5724 10208 5776 10260
rect 7196 10208 7248 10260
rect 8392 10251 8444 10260
rect 8392 10217 8401 10251
rect 8401 10217 8435 10251
rect 8435 10217 8444 10251
rect 8392 10208 8444 10217
rect 8852 10208 8904 10260
rect 9864 10208 9916 10260
rect 11336 10208 11388 10260
rect 11428 10208 11480 10260
rect 13176 10208 13228 10260
rect 14464 10208 14516 10260
rect 15016 10208 15068 10260
rect 10508 10140 10560 10192
rect 1400 9979 1452 9988
rect 1400 9945 1409 9979
rect 1409 9945 1443 9979
rect 1443 9945 1452 9979
rect 1400 9936 1452 9945
rect 5632 10072 5684 10124
rect 7748 10072 7800 10124
rect 9220 10072 9272 10124
rect 9956 10072 10008 10124
rect 5540 10004 5592 10056
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 8944 10004 8996 10056
rect 11612 10140 11664 10192
rect 12256 10140 12308 10192
rect 13452 10140 13504 10192
rect 15292 10140 15344 10192
rect 11796 10072 11848 10124
rect 15108 10072 15160 10124
rect 5816 9936 5868 9988
rect 7288 9936 7340 9988
rect 7564 9936 7616 9988
rect 6920 9868 6972 9920
rect 10416 9936 10468 9988
rect 13360 10004 13412 10056
rect 12256 9868 12308 9920
rect 13268 9936 13320 9988
rect 13820 10004 13872 10056
rect 15660 9979 15712 9988
rect 15660 9945 15669 9979
rect 15669 9945 15703 9979
rect 15703 9945 15712 9979
rect 15660 9936 15712 9945
rect 12992 9911 13044 9920
rect 12992 9877 13001 9911
rect 13001 9877 13035 9911
rect 13035 9877 13044 9911
rect 14096 9911 14148 9920
rect 12992 9868 13044 9877
rect 14096 9877 14105 9911
rect 14105 9877 14139 9911
rect 14139 9877 14148 9911
rect 14096 9868 14148 9877
rect 14188 9868 14240 9920
rect 3480 9766 3532 9818
rect 3544 9766 3596 9818
rect 3608 9766 3660 9818
rect 3672 9766 3724 9818
rect 8478 9766 8530 9818
rect 8542 9766 8594 9818
rect 8606 9766 8658 9818
rect 8670 9766 8722 9818
rect 13475 9766 13527 9818
rect 13539 9766 13591 9818
rect 13603 9766 13655 9818
rect 13667 9766 13719 9818
rect 3884 9664 3936 9716
rect 5540 9664 5592 9716
rect 7196 9664 7248 9716
rect 9312 9664 9364 9716
rect 13820 9664 13872 9716
rect 8300 9596 8352 9648
rect 9036 9596 9088 9648
rect 9956 9639 10008 9648
rect 9956 9605 9965 9639
rect 9965 9605 9999 9639
rect 9999 9605 10008 9639
rect 9956 9596 10008 9605
rect 4160 9528 4212 9580
rect 5172 9571 5224 9580
rect 5172 9537 5181 9571
rect 5181 9537 5215 9571
rect 5215 9537 5224 9571
rect 5172 9528 5224 9537
rect 6000 9528 6052 9580
rect 6460 9528 6512 9580
rect 10784 9596 10836 9648
rect 12440 9596 12492 9648
rect 10508 9571 10560 9580
rect 5356 9460 5408 9512
rect 6276 9460 6328 9512
rect 6736 9460 6788 9512
rect 10508 9537 10517 9571
rect 10517 9537 10551 9571
rect 10551 9537 10560 9571
rect 10508 9528 10560 9537
rect 13268 9528 13320 9580
rect 13912 9528 13964 9580
rect 14096 9528 14148 9580
rect 9680 9460 9732 9512
rect 12808 9460 12860 9512
rect 12900 9460 12952 9512
rect 14188 9503 14240 9512
rect 3332 9324 3384 9376
rect 4988 9324 5040 9376
rect 7564 9435 7616 9444
rect 7564 9401 7582 9435
rect 7582 9401 7616 9435
rect 7564 9392 7616 9401
rect 9496 9392 9548 9444
rect 10784 9435 10836 9444
rect 10784 9401 10793 9435
rect 10793 9401 10827 9435
rect 10827 9401 10836 9435
rect 10784 9392 10836 9401
rect 5724 9367 5776 9376
rect 5724 9333 5733 9367
rect 5733 9333 5767 9367
rect 5767 9333 5776 9367
rect 5724 9324 5776 9333
rect 5816 9324 5868 9376
rect 7196 9324 7248 9376
rect 7472 9324 7524 9376
rect 9956 9324 10008 9376
rect 10324 9367 10376 9376
rect 10324 9333 10333 9367
rect 10333 9333 10367 9367
rect 10367 9333 10376 9367
rect 10324 9324 10376 9333
rect 10692 9324 10744 9376
rect 11612 9324 11664 9376
rect 12440 9367 12492 9376
rect 12440 9333 12449 9367
rect 12449 9333 12483 9367
rect 12483 9333 12492 9367
rect 12440 9324 12492 9333
rect 12808 9324 12860 9376
rect 14188 9469 14197 9503
rect 14197 9469 14231 9503
rect 14231 9469 14240 9503
rect 14188 9460 14240 9469
rect 13452 9367 13504 9376
rect 13452 9333 13461 9367
rect 13461 9333 13495 9367
rect 13495 9333 13504 9367
rect 13452 9324 13504 9333
rect 5979 9222 6031 9274
rect 6043 9222 6095 9274
rect 6107 9222 6159 9274
rect 6171 9222 6223 9274
rect 10976 9222 11028 9274
rect 11040 9222 11092 9274
rect 11104 9222 11156 9274
rect 11168 9222 11220 9274
rect 3332 9163 3384 9172
rect 3332 9129 3341 9163
rect 3341 9129 3375 9163
rect 3375 9129 3384 9163
rect 3332 9120 3384 9129
rect 1400 9095 1452 9104
rect 1400 9061 1409 9095
rect 1409 9061 1443 9095
rect 1443 9061 1452 9095
rect 1400 9052 1452 9061
rect 1584 9027 1636 9036
rect 1584 8993 1593 9027
rect 1593 8993 1627 9027
rect 1627 8993 1636 9027
rect 1584 8984 1636 8993
rect 6920 9120 6972 9172
rect 8760 9120 8812 9172
rect 9496 9163 9548 9172
rect 9496 9129 9505 9163
rect 9505 9129 9539 9163
rect 9539 9129 9548 9163
rect 9496 9120 9548 9129
rect 9772 9120 9824 9172
rect 10140 9120 10192 9172
rect 10416 9163 10468 9172
rect 10416 9129 10425 9163
rect 10425 9129 10459 9163
rect 10459 9129 10468 9163
rect 10416 9120 10468 9129
rect 7748 9052 7800 9104
rect 4160 9027 4212 9036
rect 4160 8993 4194 9027
rect 4194 8993 4212 9027
rect 4160 8984 4212 8993
rect 6460 8984 6512 9036
rect 8208 9027 8260 9036
rect 8208 8993 8217 9027
rect 8217 8993 8251 9027
rect 8251 8993 8260 9027
rect 8208 8984 8260 8993
rect 9404 8984 9456 9036
rect 7932 8959 7984 8968
rect 3792 8848 3844 8900
rect 2872 8780 2924 8832
rect 3056 8780 3108 8832
rect 6736 8891 6788 8900
rect 6736 8857 6745 8891
rect 6745 8857 6779 8891
rect 6779 8857 6788 8891
rect 6736 8848 6788 8857
rect 6460 8780 6512 8832
rect 7564 8823 7616 8832
rect 7564 8789 7573 8823
rect 7573 8789 7607 8823
rect 7607 8789 7616 8823
rect 7564 8780 7616 8789
rect 7932 8925 7941 8959
rect 7941 8925 7975 8959
rect 7975 8925 7984 8959
rect 7932 8916 7984 8925
rect 8116 8959 8168 8968
rect 8116 8925 8125 8959
rect 8125 8925 8159 8959
rect 8159 8925 8168 8959
rect 8116 8916 8168 8925
rect 8760 8959 8812 8968
rect 8760 8925 8769 8959
rect 8769 8925 8803 8959
rect 8803 8925 8812 8959
rect 8760 8916 8812 8925
rect 8944 8848 8996 8900
rect 9220 8848 9272 8900
rect 10600 8916 10652 8968
rect 12808 9120 12860 9172
rect 12992 9120 13044 9172
rect 14464 9120 14516 9172
rect 10784 9052 10836 9104
rect 15108 9052 15160 9104
rect 11336 8984 11388 9036
rect 12716 8984 12768 9036
rect 8852 8780 8904 8832
rect 9036 8780 9088 8832
rect 9956 8780 10008 8832
rect 11428 8780 11480 8832
rect 11796 8780 11848 8832
rect 11980 8780 12032 8832
rect 12532 8780 12584 8832
rect 12900 8780 12952 8832
rect 3480 8678 3532 8730
rect 3544 8678 3596 8730
rect 3608 8678 3660 8730
rect 3672 8678 3724 8730
rect 8478 8678 8530 8730
rect 8542 8678 8594 8730
rect 8606 8678 8658 8730
rect 8670 8678 8722 8730
rect 13475 8678 13527 8730
rect 13539 8678 13591 8730
rect 13603 8678 13655 8730
rect 13667 8678 13719 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 3792 8576 3844 8628
rect 4252 8440 4304 8492
rect 6276 8551 6328 8560
rect 6276 8517 6285 8551
rect 6285 8517 6319 8551
rect 6319 8517 6328 8551
rect 6276 8508 6328 8517
rect 8208 8576 8260 8628
rect 11336 8619 11388 8628
rect 9864 8508 9916 8560
rect 9956 8508 10008 8560
rect 11336 8585 11345 8619
rect 11345 8585 11379 8619
rect 11379 8585 11388 8619
rect 11336 8576 11388 8585
rect 11796 8576 11848 8628
rect 2964 8304 3016 8356
rect 4160 8372 4212 8424
rect 5172 8440 5224 8492
rect 5724 8440 5776 8492
rect 6460 8483 6512 8492
rect 6460 8449 6469 8483
rect 6469 8449 6503 8483
rect 6503 8449 6512 8483
rect 6460 8440 6512 8449
rect 9220 8440 9272 8492
rect 4252 8304 4304 8356
rect 4620 8304 4672 8356
rect 5632 8304 5684 8356
rect 6736 8415 6788 8424
rect 6736 8381 6770 8415
rect 6770 8381 6788 8415
rect 6736 8372 6788 8381
rect 7196 8372 7248 8424
rect 7472 8372 7524 8424
rect 8024 8372 8076 8424
rect 6920 8304 6972 8356
rect 7288 8304 7340 8356
rect 9772 8372 9824 8424
rect 4344 8279 4396 8288
rect 4344 8245 4353 8279
rect 4353 8245 4387 8279
rect 4387 8245 4396 8279
rect 4344 8236 4396 8245
rect 5080 8236 5132 8288
rect 5540 8279 5592 8288
rect 5540 8245 5549 8279
rect 5549 8245 5583 8279
rect 5583 8245 5592 8279
rect 5540 8236 5592 8245
rect 9496 8279 9548 8288
rect 9496 8245 9505 8279
rect 9505 8245 9539 8279
rect 9539 8245 9548 8279
rect 9496 8236 9548 8245
rect 9680 8236 9732 8288
rect 10600 8372 10652 8424
rect 10232 8347 10284 8356
rect 10232 8313 10266 8347
rect 10266 8313 10284 8347
rect 10232 8304 10284 8313
rect 13268 8576 13320 8628
rect 11980 8440 12032 8492
rect 12808 8372 12860 8424
rect 13452 8304 13504 8356
rect 14372 8304 14424 8356
rect 12808 8279 12860 8288
rect 12808 8245 12817 8279
rect 12817 8245 12851 8279
rect 12851 8245 12860 8279
rect 12808 8236 12860 8245
rect 5979 8134 6031 8186
rect 6043 8134 6095 8186
rect 6107 8134 6159 8186
rect 6171 8134 6223 8186
rect 10976 8134 11028 8186
rect 11040 8134 11092 8186
rect 11104 8134 11156 8186
rect 11168 8134 11220 8186
rect 1492 8075 1544 8084
rect 1492 8041 1501 8075
rect 1501 8041 1535 8075
rect 1535 8041 1544 8075
rect 1492 8032 1544 8041
rect 4344 8032 4396 8084
rect 4896 8032 4948 8084
rect 5448 8032 5500 8084
rect 7104 8032 7156 8084
rect 7564 8032 7616 8084
rect 8116 8032 8168 8084
rect 4344 7896 4396 7948
rect 4896 7939 4948 7948
rect 4896 7905 4905 7939
rect 4905 7905 4939 7939
rect 4939 7905 4948 7939
rect 4896 7896 4948 7905
rect 6184 7896 6236 7948
rect 6920 7896 6972 7948
rect 2780 7828 2832 7880
rect 4068 7828 4120 7880
rect 4528 7871 4580 7880
rect 4528 7837 4537 7871
rect 4537 7837 4571 7871
rect 4571 7837 4580 7871
rect 4528 7828 4580 7837
rect 4620 7871 4672 7880
rect 4620 7837 4629 7871
rect 4629 7837 4663 7871
rect 4663 7837 4672 7871
rect 4620 7828 4672 7837
rect 2964 7760 3016 7812
rect 7196 7964 7248 8016
rect 7472 7964 7524 8016
rect 8300 7964 8352 8016
rect 9496 8075 9548 8084
rect 9496 8041 9505 8075
rect 9505 8041 9539 8075
rect 9539 8041 9548 8075
rect 9496 8032 9548 8041
rect 12440 8032 12492 8084
rect 12808 8032 12860 8084
rect 13360 8075 13412 8084
rect 13360 8041 13369 8075
rect 13369 8041 13403 8075
rect 13403 8041 13412 8075
rect 13360 8032 13412 8041
rect 9036 7964 9088 8016
rect 9220 7896 9272 7948
rect 7288 7828 7340 7880
rect 7932 7828 7984 7880
rect 9312 7828 9364 7880
rect 9588 7871 9640 7880
rect 9588 7837 9597 7871
rect 9597 7837 9631 7871
rect 9631 7837 9640 7871
rect 9588 7828 9640 7837
rect 8116 7760 8168 7812
rect 8392 7760 8444 7812
rect 10324 7896 10376 7948
rect 10600 7896 10652 7948
rect 12900 8007 12952 8016
rect 10232 7871 10284 7880
rect 10232 7837 10241 7871
rect 10241 7837 10275 7871
rect 10275 7837 10284 7871
rect 10232 7828 10284 7837
rect 10416 7871 10468 7880
rect 10416 7837 10425 7871
rect 10425 7837 10459 7871
rect 10459 7837 10468 7871
rect 10416 7828 10468 7837
rect 11336 7828 11388 7880
rect 11980 7871 12032 7880
rect 11980 7837 11989 7871
rect 11989 7837 12023 7871
rect 12023 7837 12032 7871
rect 11980 7828 12032 7837
rect 12900 7973 12909 8007
rect 12909 7973 12943 8007
rect 12943 7973 12952 8007
rect 12900 7964 12952 7973
rect 9864 7760 9916 7812
rect 3240 7692 3292 7744
rect 5172 7692 5224 7744
rect 5816 7692 5868 7744
rect 7564 7692 7616 7744
rect 8208 7692 8260 7744
rect 8852 7692 8904 7744
rect 9956 7692 10008 7744
rect 12256 7692 12308 7744
rect 13084 7896 13136 7948
rect 13268 7828 13320 7880
rect 12716 7760 12768 7812
rect 14004 8032 14056 8084
rect 12992 7692 13044 7744
rect 3480 7590 3532 7642
rect 3544 7590 3596 7642
rect 3608 7590 3660 7642
rect 3672 7590 3724 7642
rect 8478 7590 8530 7642
rect 8542 7590 8594 7642
rect 8606 7590 8658 7642
rect 8670 7590 8722 7642
rect 13475 7590 13527 7642
rect 13539 7590 13591 7642
rect 13603 7590 13655 7642
rect 13667 7590 13719 7642
rect 2044 7488 2096 7540
rect 2320 7488 2372 7540
rect 2780 7488 2832 7540
rect 3240 7488 3292 7540
rect 4528 7488 4580 7540
rect 5540 7531 5592 7540
rect 5540 7497 5549 7531
rect 5549 7497 5583 7531
rect 5583 7497 5592 7531
rect 5540 7488 5592 7497
rect 5724 7488 5776 7540
rect 6276 7488 6328 7540
rect 7196 7488 7248 7540
rect 7656 7488 7708 7540
rect 7932 7488 7984 7540
rect 2872 7352 2924 7404
rect 8116 7420 8168 7472
rect 6184 7395 6236 7404
rect 6184 7361 6193 7395
rect 6193 7361 6227 7395
rect 6227 7361 6236 7395
rect 6184 7352 6236 7361
rect 6920 7352 6972 7404
rect 9864 7488 9916 7540
rect 10048 7488 10100 7540
rect 10324 7488 10376 7540
rect 10784 7488 10836 7540
rect 11520 7488 11572 7540
rect 9036 7395 9088 7404
rect 2964 7327 3016 7336
rect 2964 7293 2973 7327
rect 2973 7293 3007 7327
rect 3007 7293 3016 7327
rect 2964 7284 3016 7293
rect 4712 7284 4764 7336
rect 5540 7284 5592 7336
rect 7564 7284 7616 7336
rect 9036 7361 9045 7395
rect 9045 7361 9079 7395
rect 9079 7361 9088 7395
rect 9036 7352 9088 7361
rect 9680 7395 9732 7404
rect 9680 7361 9689 7395
rect 9689 7361 9723 7395
rect 9723 7361 9732 7395
rect 9680 7352 9732 7361
rect 11336 7352 11388 7404
rect 12072 7395 12124 7404
rect 12072 7361 12081 7395
rect 12081 7361 12115 7395
rect 12115 7361 12124 7395
rect 12072 7352 12124 7361
rect 12624 7352 12676 7404
rect 13268 7352 13320 7404
rect 8852 7327 8904 7336
rect 8852 7293 8861 7327
rect 8861 7293 8895 7327
rect 8895 7293 8904 7327
rect 8852 7284 8904 7293
rect 8944 7327 8996 7336
rect 8944 7293 8953 7327
rect 8953 7293 8987 7327
rect 8987 7293 8996 7327
rect 8944 7284 8996 7293
rect 3240 7259 3292 7268
rect 3240 7225 3274 7259
rect 3274 7225 3292 7259
rect 1492 7191 1544 7200
rect 1492 7157 1501 7191
rect 1501 7157 1535 7191
rect 1535 7157 1544 7191
rect 1492 7148 1544 7157
rect 3240 7216 3292 7225
rect 3424 7216 3476 7268
rect 5080 7216 5132 7268
rect 5172 7216 5224 7268
rect 2320 7191 2372 7200
rect 2320 7157 2329 7191
rect 2329 7157 2363 7191
rect 2363 7157 2372 7191
rect 2320 7148 2372 7157
rect 5264 7148 5316 7200
rect 5816 7148 5868 7200
rect 6460 7191 6512 7200
rect 6460 7157 6469 7191
rect 6469 7157 6503 7191
rect 6503 7157 6512 7191
rect 6460 7148 6512 7157
rect 6828 7216 6880 7268
rect 10508 7216 10560 7268
rect 11612 7284 11664 7336
rect 12164 7327 12216 7336
rect 12164 7293 12173 7327
rect 12173 7293 12207 7327
rect 12207 7293 12216 7327
rect 12164 7284 12216 7293
rect 12716 7216 12768 7268
rect 7656 7148 7708 7200
rect 10048 7148 10100 7200
rect 11336 7148 11388 7200
rect 12532 7191 12584 7200
rect 12532 7157 12541 7191
rect 12541 7157 12575 7191
rect 12575 7157 12584 7191
rect 12532 7148 12584 7157
rect 12624 7191 12676 7200
rect 12624 7157 12633 7191
rect 12633 7157 12667 7191
rect 12667 7157 12676 7191
rect 12624 7148 12676 7157
rect 15844 7148 15896 7200
rect 5979 7046 6031 7098
rect 6043 7046 6095 7098
rect 6107 7046 6159 7098
rect 6171 7046 6223 7098
rect 10976 7046 11028 7098
rect 11040 7046 11092 7098
rect 11104 7046 11156 7098
rect 11168 7046 11220 7098
rect 3332 6944 3384 6996
rect 7472 6944 7524 6996
rect 2504 6876 2556 6928
rect 3424 6919 3476 6928
rect 3424 6885 3433 6919
rect 3433 6885 3467 6919
rect 3467 6885 3476 6919
rect 3424 6876 3476 6885
rect 4068 6876 4120 6928
rect 5540 6876 5592 6928
rect 1768 6808 1820 6860
rect 1952 6808 2004 6860
rect 2688 6808 2740 6860
rect 5264 6808 5316 6860
rect 5724 6808 5776 6860
rect 1492 6647 1544 6656
rect 1492 6613 1501 6647
rect 1501 6613 1535 6647
rect 1535 6613 1544 6647
rect 1492 6604 1544 6613
rect 4896 6740 4948 6792
rect 3148 6672 3200 6724
rect 4528 6672 4580 6724
rect 2964 6604 3016 6656
rect 3240 6647 3292 6656
rect 3240 6613 3249 6647
rect 3249 6613 3283 6647
rect 3283 6613 3292 6647
rect 3240 6604 3292 6613
rect 4252 6647 4304 6656
rect 4252 6613 4261 6647
rect 4261 6613 4295 6647
rect 4295 6613 4304 6647
rect 4252 6604 4304 6613
rect 5264 6647 5316 6656
rect 5264 6613 5273 6647
rect 5273 6613 5307 6647
rect 5307 6613 5316 6647
rect 5264 6604 5316 6613
rect 5632 6672 5684 6724
rect 6276 6740 6328 6792
rect 8208 6944 8260 6996
rect 9036 6944 9088 6996
rect 10416 6944 10468 6996
rect 11336 6944 11388 6996
rect 7932 6876 7984 6928
rect 10692 6876 10744 6928
rect 9680 6808 9732 6860
rect 12532 6944 12584 6996
rect 6920 6740 6972 6792
rect 7472 6783 7524 6792
rect 6736 6715 6788 6724
rect 6736 6681 6745 6715
rect 6745 6681 6779 6715
rect 6779 6681 6788 6715
rect 6736 6672 6788 6681
rect 7472 6749 7481 6783
rect 7481 6749 7515 6783
rect 7515 6749 7524 6783
rect 7472 6740 7524 6749
rect 10232 6740 10284 6792
rect 10508 6715 10560 6724
rect 7012 6647 7064 6656
rect 7012 6613 7021 6647
rect 7021 6613 7055 6647
rect 7055 6613 7064 6647
rect 7012 6604 7064 6613
rect 10508 6681 10517 6715
rect 10517 6681 10551 6715
rect 10551 6681 10560 6715
rect 10508 6672 10560 6681
rect 10692 6740 10744 6792
rect 11336 6740 11388 6792
rect 12716 6808 12768 6860
rect 11244 6604 11296 6656
rect 11428 6647 11480 6656
rect 11428 6613 11437 6647
rect 11437 6613 11471 6647
rect 11471 6613 11480 6647
rect 11428 6604 11480 6613
rect 13084 6715 13136 6724
rect 13084 6681 13093 6715
rect 13093 6681 13127 6715
rect 13127 6681 13136 6715
rect 13084 6672 13136 6681
rect 3480 6502 3532 6554
rect 3544 6502 3596 6554
rect 3608 6502 3660 6554
rect 3672 6502 3724 6554
rect 8478 6502 8530 6554
rect 8542 6502 8594 6554
rect 8606 6502 8658 6554
rect 8670 6502 8722 6554
rect 13475 6502 13527 6554
rect 13539 6502 13591 6554
rect 13603 6502 13655 6554
rect 13667 6502 13719 6554
rect 1860 6400 1912 6452
rect 2688 6400 2740 6452
rect 3332 6400 3384 6452
rect 5264 6400 5316 6452
rect 5540 6400 5592 6452
rect 5816 6400 5868 6452
rect 6276 6400 6328 6452
rect 7012 6400 7064 6452
rect 8116 6400 8168 6452
rect 9128 6443 9180 6452
rect 9128 6409 9137 6443
rect 9137 6409 9171 6443
rect 9171 6409 9180 6443
rect 9128 6400 9180 6409
rect 10140 6400 10192 6452
rect 10600 6443 10652 6452
rect 10600 6409 10609 6443
rect 10609 6409 10643 6443
rect 10643 6409 10652 6443
rect 10600 6400 10652 6409
rect 11612 6400 11664 6452
rect 2964 6332 3016 6384
rect 9404 6332 9456 6384
rect 9588 6332 9640 6384
rect 11980 6332 12032 6384
rect 12716 6400 12768 6452
rect 13360 6400 13412 6452
rect 14096 6400 14148 6452
rect 14556 6400 14608 6452
rect 14740 6400 14792 6452
rect 4344 6307 4396 6316
rect 4344 6273 4353 6307
rect 4353 6273 4387 6307
rect 4387 6273 4396 6307
rect 4344 6264 4396 6273
rect 5172 6307 5224 6316
rect 5172 6273 5181 6307
rect 5181 6273 5215 6307
rect 5215 6273 5224 6307
rect 5172 6264 5224 6273
rect 5264 6264 5316 6316
rect 6552 6307 6604 6316
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 6920 6264 6972 6316
rect 9680 6264 9732 6316
rect 10508 6264 10560 6316
rect 11336 6264 11388 6316
rect 13268 6264 13320 6316
rect 3332 6196 3384 6248
rect 2228 6128 2280 6180
rect 2688 6171 2740 6180
rect 2688 6137 2706 6171
rect 2706 6137 2740 6171
rect 2688 6128 2740 6137
rect 5816 6196 5868 6248
rect 7012 6196 7064 6248
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 1952 6060 2004 6112
rect 3148 6060 3200 6112
rect 7288 6128 7340 6180
rect 7748 6128 7800 6180
rect 8024 6171 8076 6180
rect 8024 6137 8042 6171
rect 8042 6137 8076 6171
rect 8024 6128 8076 6137
rect 8208 6128 8260 6180
rect 9864 6196 9916 6248
rect 10324 6196 10376 6248
rect 10600 6196 10652 6248
rect 11612 6196 11664 6248
rect 12624 6196 12676 6248
rect 5632 6060 5684 6112
rect 6828 6060 6880 6112
rect 7380 6060 7432 6112
rect 7656 6060 7708 6112
rect 9036 6060 9088 6112
rect 9312 6060 9364 6112
rect 12348 6128 12400 6180
rect 9772 6060 9824 6112
rect 10140 6060 10192 6112
rect 10692 6060 10744 6112
rect 10876 6060 10928 6112
rect 11796 6060 11848 6112
rect 15384 6103 15436 6112
rect 15384 6069 15393 6103
rect 15393 6069 15427 6103
rect 15427 6069 15436 6103
rect 15384 6060 15436 6069
rect 5979 5958 6031 6010
rect 6043 5958 6095 6010
rect 6107 5958 6159 6010
rect 6171 5958 6223 6010
rect 10976 5958 11028 6010
rect 11040 5958 11092 6010
rect 11104 5958 11156 6010
rect 11168 5958 11220 6010
rect 1768 5899 1820 5908
rect 1768 5865 1777 5899
rect 1777 5865 1811 5899
rect 1811 5865 1820 5899
rect 1768 5856 1820 5865
rect 4252 5899 4304 5908
rect 4252 5865 4261 5899
rect 4261 5865 4295 5899
rect 4295 5865 4304 5899
rect 4252 5856 4304 5865
rect 1584 5788 1636 5840
rect 2136 5720 2188 5772
rect 4344 5788 4396 5840
rect 5632 5856 5684 5908
rect 6828 5788 6880 5840
rect 7472 5856 7524 5908
rect 9588 5856 9640 5908
rect 9864 5856 9916 5908
rect 11704 5856 11756 5908
rect 12256 5856 12308 5908
rect 12348 5856 12400 5908
rect 12900 5856 12952 5908
rect 15752 5856 15804 5908
rect 9312 5788 9364 5840
rect 3424 5720 3476 5772
rect 2412 5695 2464 5704
rect 2412 5661 2421 5695
rect 2421 5661 2455 5695
rect 2455 5661 2464 5695
rect 2412 5652 2464 5661
rect 2688 5652 2740 5704
rect 4160 5652 4212 5704
rect 4528 5720 4580 5772
rect 4896 5763 4948 5772
rect 4896 5729 4905 5763
rect 4905 5729 4939 5763
rect 4939 5729 4948 5763
rect 4896 5720 4948 5729
rect 6920 5720 6972 5772
rect 7472 5720 7524 5772
rect 8116 5720 8168 5772
rect 8944 5720 8996 5772
rect 9772 5720 9824 5772
rect 3884 5584 3936 5636
rect 4528 5584 4580 5636
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 2872 5559 2924 5568
rect 2872 5525 2881 5559
rect 2881 5525 2915 5559
rect 2915 5525 2924 5559
rect 2872 5516 2924 5525
rect 3332 5516 3384 5568
rect 6736 5652 6788 5704
rect 8024 5652 8076 5704
rect 7012 5584 7064 5636
rect 8852 5584 8904 5636
rect 9220 5584 9272 5636
rect 9404 5584 9456 5636
rect 6000 5516 6052 5568
rect 6368 5516 6420 5568
rect 6644 5516 6696 5568
rect 6920 5559 6972 5568
rect 6920 5525 6929 5559
rect 6929 5525 6963 5559
rect 6963 5525 6972 5559
rect 6920 5516 6972 5525
rect 7748 5559 7800 5568
rect 7748 5525 7757 5559
rect 7757 5525 7791 5559
rect 7791 5525 7800 5559
rect 7748 5516 7800 5525
rect 8944 5559 8996 5568
rect 8944 5525 8953 5559
rect 8953 5525 8987 5559
rect 8987 5525 8996 5559
rect 8944 5516 8996 5525
rect 9312 5559 9364 5568
rect 9312 5525 9321 5559
rect 9321 5525 9355 5559
rect 9355 5525 9364 5559
rect 9312 5516 9364 5525
rect 9588 5559 9640 5568
rect 9588 5525 9597 5559
rect 9597 5525 9631 5559
rect 9631 5525 9640 5559
rect 9588 5516 9640 5525
rect 9772 5516 9824 5568
rect 10324 5788 10376 5840
rect 10324 5695 10376 5704
rect 10324 5661 10333 5695
rect 10333 5661 10367 5695
rect 10367 5661 10376 5695
rect 10324 5652 10376 5661
rect 10140 5584 10192 5636
rect 10232 5584 10284 5636
rect 12808 5788 12860 5840
rect 14372 5831 14424 5840
rect 11612 5720 11664 5772
rect 14372 5797 14381 5831
rect 14381 5797 14415 5831
rect 14415 5797 14424 5831
rect 14372 5788 14424 5797
rect 15660 5831 15712 5840
rect 15660 5797 15669 5831
rect 15669 5797 15703 5831
rect 15703 5797 15712 5831
rect 15660 5788 15712 5797
rect 13360 5763 13412 5772
rect 11980 5652 12032 5704
rect 13360 5729 13369 5763
rect 13369 5729 13403 5763
rect 13403 5729 13412 5763
rect 13360 5720 13412 5729
rect 14648 5720 14700 5772
rect 14924 5720 14976 5772
rect 15476 5763 15528 5772
rect 15476 5729 15485 5763
rect 15485 5729 15519 5763
rect 15519 5729 15528 5763
rect 15476 5720 15528 5729
rect 12440 5695 12492 5704
rect 12440 5661 12449 5695
rect 12449 5661 12483 5695
rect 12483 5661 12492 5695
rect 12440 5652 12492 5661
rect 12808 5652 12860 5704
rect 13268 5695 13320 5704
rect 13268 5661 13277 5695
rect 13277 5661 13311 5695
rect 13311 5661 13320 5695
rect 13268 5652 13320 5661
rect 15568 5652 15620 5704
rect 13176 5584 13228 5636
rect 15292 5584 15344 5636
rect 10600 5559 10652 5568
rect 10600 5525 10609 5559
rect 10609 5525 10643 5559
rect 10643 5525 10652 5559
rect 10600 5516 10652 5525
rect 10968 5516 11020 5568
rect 11336 5516 11388 5568
rect 11520 5516 11572 5568
rect 11980 5559 12032 5568
rect 11980 5525 11989 5559
rect 11989 5525 12023 5559
rect 12023 5525 12032 5559
rect 11980 5516 12032 5525
rect 12164 5516 12216 5568
rect 13820 5559 13872 5568
rect 13820 5525 13829 5559
rect 13829 5525 13863 5559
rect 13863 5525 13872 5559
rect 13820 5516 13872 5525
rect 13912 5516 13964 5568
rect 15200 5559 15252 5568
rect 15200 5525 15209 5559
rect 15209 5525 15243 5559
rect 15243 5525 15252 5559
rect 15200 5516 15252 5525
rect 3480 5414 3532 5466
rect 3544 5414 3596 5466
rect 3608 5414 3660 5466
rect 3672 5414 3724 5466
rect 8478 5414 8530 5466
rect 8542 5414 8594 5466
rect 8606 5414 8658 5466
rect 8670 5414 8722 5466
rect 13475 5414 13527 5466
rect 13539 5414 13591 5466
rect 13603 5414 13655 5466
rect 13667 5414 13719 5466
rect 2412 5312 2464 5364
rect 4160 5312 4212 5364
rect 5264 5355 5316 5364
rect 5264 5321 5273 5355
rect 5273 5321 5307 5355
rect 5307 5321 5316 5355
rect 5264 5312 5316 5321
rect 6552 5312 6604 5364
rect 6828 5312 6880 5364
rect 1400 5287 1452 5296
rect 1400 5253 1409 5287
rect 1409 5253 1443 5287
rect 1443 5253 1452 5287
rect 1400 5244 1452 5253
rect 2136 5244 2188 5296
rect 2688 5176 2740 5228
rect 2872 5176 2924 5228
rect 3240 5219 3292 5228
rect 3240 5185 3249 5219
rect 3249 5185 3283 5219
rect 3283 5185 3292 5219
rect 3240 5176 3292 5185
rect 3332 5176 3384 5228
rect 1492 5108 1544 5160
rect 2964 5151 3016 5160
rect 2964 5117 2973 5151
rect 2973 5117 3007 5151
rect 3007 5117 3016 5151
rect 2964 5108 3016 5117
rect 2044 5015 2096 5024
rect 2044 4981 2053 5015
rect 2053 4981 2087 5015
rect 2087 4981 2096 5015
rect 2044 4972 2096 4981
rect 2136 5015 2188 5024
rect 2136 4981 2145 5015
rect 2145 4981 2179 5015
rect 2179 4981 2188 5015
rect 2136 4972 2188 4981
rect 3332 4972 3384 5024
rect 6092 5219 6144 5228
rect 6092 5185 6101 5219
rect 6101 5185 6135 5219
rect 6135 5185 6144 5219
rect 6092 5176 6144 5185
rect 6552 5176 6604 5228
rect 6920 5219 6972 5228
rect 6920 5185 6929 5219
rect 6929 5185 6963 5219
rect 6963 5185 6972 5219
rect 6920 5176 6972 5185
rect 7840 5312 7892 5364
rect 8944 5312 8996 5364
rect 11060 5355 11112 5364
rect 11060 5321 11069 5355
rect 11069 5321 11103 5355
rect 11103 5321 11112 5355
rect 11060 5312 11112 5321
rect 13176 5312 13228 5364
rect 8024 5244 8076 5296
rect 9956 5244 10008 5296
rect 10232 5244 10284 5296
rect 9680 5219 9732 5228
rect 9680 5185 9689 5219
rect 9689 5185 9723 5219
rect 9723 5185 9732 5219
rect 9680 5176 9732 5185
rect 4160 5151 4212 5160
rect 4160 5117 4194 5151
rect 4194 5117 4212 5151
rect 3700 5083 3752 5092
rect 3700 5049 3709 5083
rect 3709 5049 3743 5083
rect 3743 5049 3752 5083
rect 3700 5040 3752 5049
rect 4160 5108 4212 5117
rect 4528 5108 4580 5160
rect 3976 5040 4028 5092
rect 6736 5108 6788 5160
rect 7748 5108 7800 5160
rect 9772 5108 9824 5160
rect 10508 5151 10560 5160
rect 10508 5117 10517 5151
rect 10517 5117 10551 5151
rect 10551 5117 10560 5151
rect 10508 5108 10560 5117
rect 6184 5040 6236 5092
rect 6460 5040 6512 5092
rect 6920 5040 6972 5092
rect 7196 5040 7248 5092
rect 7472 5040 7524 5092
rect 8852 5040 8904 5092
rect 11612 5040 11664 5092
rect 15476 5312 15528 5364
rect 12072 5108 12124 5160
rect 13176 5040 13228 5092
rect 15292 5108 15344 5160
rect 5356 5015 5408 5024
rect 5356 4981 5365 5015
rect 5365 4981 5399 5015
rect 5399 4981 5408 5015
rect 5540 5015 5592 5024
rect 5356 4972 5408 4981
rect 5540 4981 5549 5015
rect 5549 4981 5583 5015
rect 5583 4981 5592 5015
rect 5540 4972 5592 4981
rect 6276 4972 6328 5024
rect 7012 4972 7064 5024
rect 7380 4972 7432 5024
rect 7748 5015 7800 5024
rect 7748 4981 7757 5015
rect 7757 4981 7791 5015
rect 7791 4981 7800 5015
rect 8116 5015 8168 5024
rect 7748 4972 7800 4981
rect 8116 4981 8125 5015
rect 8125 4981 8159 5015
rect 8159 4981 8168 5015
rect 8116 4972 8168 4981
rect 8576 4972 8628 5024
rect 9220 4972 9272 5024
rect 9312 4972 9364 5024
rect 10416 5015 10468 5024
rect 10416 4981 10425 5015
rect 10425 4981 10459 5015
rect 10459 4981 10468 5015
rect 10416 4972 10468 4981
rect 11336 5015 11388 5024
rect 11336 4981 11345 5015
rect 11345 4981 11379 5015
rect 11379 4981 11388 5015
rect 11336 4972 11388 4981
rect 11704 5015 11756 5024
rect 11704 4981 11713 5015
rect 11713 4981 11747 5015
rect 11747 4981 11756 5015
rect 11704 4972 11756 4981
rect 11796 4972 11848 5024
rect 14924 5015 14976 5024
rect 14924 4981 14933 5015
rect 14933 4981 14967 5015
rect 14967 4981 14976 5015
rect 14924 4972 14976 4981
rect 15016 4972 15068 5024
rect 5979 4870 6031 4922
rect 6043 4870 6095 4922
rect 6107 4870 6159 4922
rect 6171 4870 6223 4922
rect 10976 4870 11028 4922
rect 11040 4870 11092 4922
rect 11104 4870 11156 4922
rect 11168 4870 11220 4922
rect 2044 4811 2096 4820
rect 2044 4777 2053 4811
rect 2053 4777 2087 4811
rect 2087 4777 2096 4811
rect 2044 4768 2096 4777
rect 2136 4768 2188 4820
rect 3700 4768 3752 4820
rect 3884 4811 3936 4820
rect 3884 4777 3893 4811
rect 3893 4777 3927 4811
rect 3927 4777 3936 4811
rect 3884 4768 3936 4777
rect 7196 4811 7248 4820
rect 3792 4700 3844 4752
rect 1676 4675 1728 4684
rect 1676 4641 1685 4675
rect 1685 4641 1719 4675
rect 1719 4641 1728 4675
rect 1676 4632 1728 4641
rect 2136 4632 2188 4684
rect 3148 4632 3200 4684
rect 4712 4700 4764 4752
rect 5724 4700 5776 4752
rect 7196 4777 7205 4811
rect 7205 4777 7239 4811
rect 7239 4777 7248 4811
rect 7196 4768 7248 4777
rect 7380 4811 7432 4820
rect 7380 4777 7389 4811
rect 7389 4777 7423 4811
rect 7423 4777 7432 4811
rect 7380 4768 7432 4777
rect 7656 4768 7708 4820
rect 4252 4675 4304 4684
rect 4252 4641 4261 4675
rect 4261 4641 4295 4675
rect 4295 4641 4304 4675
rect 4252 4632 4304 4641
rect 4804 4632 4856 4684
rect 5080 4632 5132 4684
rect 5264 4632 5316 4684
rect 5356 4632 5408 4684
rect 5632 4632 5684 4684
rect 5816 4675 5868 4684
rect 5816 4641 5825 4675
rect 5825 4641 5859 4675
rect 5859 4641 5868 4675
rect 5816 4632 5868 4641
rect 6460 4632 6512 4684
rect 7932 4768 7984 4820
rect 10048 4768 10100 4820
rect 12072 4768 12124 4820
rect 13176 4811 13228 4820
rect 13176 4777 13185 4811
rect 13185 4777 13219 4811
rect 13219 4777 13228 4811
rect 13176 4768 13228 4777
rect 14924 4768 14976 4820
rect 15844 4768 15896 4820
rect 9312 4743 9364 4752
rect 3056 4564 3108 4616
rect 4068 4564 4120 4616
rect 4160 4564 4212 4616
rect 7196 4632 7248 4684
rect 8576 4675 8628 4684
rect 8576 4641 8585 4675
rect 8585 4641 8619 4675
rect 8619 4641 8628 4675
rect 8576 4632 8628 4641
rect 9312 4709 9321 4743
rect 9321 4709 9355 4743
rect 9355 4709 9364 4743
rect 9312 4700 9364 4709
rect 9220 4632 9272 4684
rect 7104 4564 7156 4616
rect 8024 4607 8076 4616
rect 8024 4573 8033 4607
rect 8033 4573 8067 4607
rect 8067 4573 8076 4607
rect 8024 4564 8076 4573
rect 8668 4607 8720 4616
rect 8668 4573 8677 4607
rect 8677 4573 8711 4607
rect 8711 4573 8720 4607
rect 8668 4564 8720 4573
rect 8852 4607 8904 4616
rect 8852 4573 8861 4607
rect 8861 4573 8895 4607
rect 8895 4573 8904 4607
rect 8852 4564 8904 4573
rect 4620 4496 4672 4548
rect 5540 4496 5592 4548
rect 6828 4539 6880 4548
rect 1492 4471 1544 4480
rect 1492 4437 1501 4471
rect 1501 4437 1535 4471
rect 1535 4437 1544 4471
rect 1492 4428 1544 4437
rect 1768 4471 1820 4480
rect 1768 4437 1777 4471
rect 1777 4437 1811 4471
rect 1811 4437 1820 4471
rect 1768 4428 1820 4437
rect 4344 4428 4396 4480
rect 4988 4471 5040 4480
rect 4988 4437 4997 4471
rect 4997 4437 5031 4471
rect 5031 4437 5040 4471
rect 4988 4428 5040 4437
rect 6276 4428 6328 4480
rect 6828 4505 6837 4539
rect 6837 4505 6871 4539
rect 6871 4505 6880 4539
rect 6828 4496 6880 4505
rect 8300 4496 8352 4548
rect 10784 4700 10836 4752
rect 11796 4700 11848 4752
rect 14556 4700 14608 4752
rect 14740 4743 14792 4752
rect 14740 4709 14749 4743
rect 14749 4709 14783 4743
rect 14783 4709 14792 4743
rect 14740 4700 14792 4709
rect 15292 4700 15344 4752
rect 12072 4675 12124 4684
rect 12072 4641 12106 4675
rect 12106 4641 12124 4675
rect 12072 4632 12124 4641
rect 14372 4632 14424 4684
rect 15752 4632 15804 4684
rect 16488 4632 16540 4684
rect 14188 4564 14240 4616
rect 10692 4496 10744 4548
rect 7104 4428 7156 4480
rect 8208 4471 8260 4480
rect 8208 4437 8217 4471
rect 8217 4437 8251 4471
rect 8251 4437 8260 4471
rect 8208 4428 8260 4437
rect 9680 4428 9732 4480
rect 10324 4471 10376 4480
rect 10324 4437 10333 4471
rect 10333 4437 10367 4471
rect 10367 4437 10376 4471
rect 10324 4428 10376 4437
rect 12440 4428 12492 4480
rect 14004 4428 14056 4480
rect 14372 4471 14424 4480
rect 14372 4437 14381 4471
rect 14381 4437 14415 4471
rect 14415 4437 14424 4471
rect 14372 4428 14424 4437
rect 14648 4428 14700 4480
rect 3480 4326 3532 4378
rect 3544 4326 3596 4378
rect 3608 4326 3660 4378
rect 3672 4326 3724 4378
rect 8478 4326 8530 4378
rect 8542 4326 8594 4378
rect 8606 4326 8658 4378
rect 8670 4326 8722 4378
rect 13475 4326 13527 4378
rect 13539 4326 13591 4378
rect 13603 4326 13655 4378
rect 13667 4326 13719 4378
rect 3056 4267 3108 4276
rect 3056 4233 3065 4267
rect 3065 4233 3099 4267
rect 3099 4233 3108 4267
rect 3056 4224 3108 4233
rect 4068 4224 4120 4276
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 4804 4224 4856 4276
rect 4712 4156 4764 4208
rect 7748 4224 7800 4276
rect 8024 4224 8076 4276
rect 7840 4156 7892 4208
rect 1768 4020 1820 4072
rect 1860 4020 1912 4072
rect 2320 4020 2372 4072
rect 2504 4020 2556 4072
rect 4344 4020 4396 4072
rect 3240 3952 3292 4004
rect 4160 3995 4212 4004
rect 4160 3961 4178 3995
rect 4178 3961 4212 3995
rect 4528 4088 4580 4140
rect 4988 4020 5040 4072
rect 8208 4088 8260 4140
rect 10048 4224 10100 4276
rect 10324 4156 10376 4208
rect 9680 4088 9732 4140
rect 10784 4156 10836 4208
rect 11520 4224 11572 4276
rect 14924 4224 14976 4276
rect 15108 4267 15160 4276
rect 15108 4233 15117 4267
rect 15117 4233 15151 4267
rect 15151 4233 15160 4267
rect 15108 4224 15160 4233
rect 11244 4156 11296 4208
rect 6184 4020 6236 4072
rect 6552 4020 6604 4072
rect 7564 4020 7616 4072
rect 8852 4020 8904 4072
rect 9404 4020 9456 4072
rect 10416 4020 10468 4072
rect 10876 4020 10928 4072
rect 11152 4063 11204 4072
rect 11152 4029 11161 4063
rect 11161 4029 11195 4063
rect 11195 4029 11204 4063
rect 11152 4020 11204 4029
rect 12072 4156 12124 4208
rect 12256 4088 12308 4140
rect 13176 4156 13228 4208
rect 11520 4020 11572 4072
rect 11888 4063 11940 4072
rect 11888 4029 11897 4063
rect 11897 4029 11931 4063
rect 11931 4029 11940 4063
rect 11888 4020 11940 4029
rect 13084 4088 13136 4140
rect 13728 4088 13780 4140
rect 14924 4088 14976 4140
rect 14004 4063 14056 4072
rect 4160 3952 4212 3961
rect 5632 3952 5684 4004
rect 7104 3952 7156 4004
rect 10968 3952 11020 4004
rect 12072 3952 12124 4004
rect 12532 3952 12584 4004
rect 1584 3884 1636 3936
rect 2320 3884 2372 3936
rect 2596 3927 2648 3936
rect 2596 3893 2605 3927
rect 2605 3893 2639 3927
rect 2639 3893 2648 3927
rect 2596 3884 2648 3893
rect 3976 3884 4028 3936
rect 5540 3927 5592 3936
rect 5540 3893 5549 3927
rect 5549 3893 5583 3927
rect 5583 3893 5592 3927
rect 5540 3884 5592 3893
rect 7656 3884 7708 3936
rect 7840 3927 7892 3936
rect 7840 3893 7849 3927
rect 7849 3893 7883 3927
rect 7883 3893 7892 3927
rect 7840 3884 7892 3893
rect 7932 3884 7984 3936
rect 9588 3884 9640 3936
rect 9772 3884 9824 3936
rect 10140 3927 10192 3936
rect 10140 3893 10149 3927
rect 10149 3893 10183 3927
rect 10183 3893 10192 3927
rect 10508 3927 10560 3936
rect 10140 3884 10192 3893
rect 10508 3893 10517 3927
rect 10517 3893 10551 3927
rect 10551 3893 10560 3927
rect 10508 3884 10560 3893
rect 10876 3884 10928 3936
rect 11520 3884 11572 3936
rect 11796 3884 11848 3936
rect 12164 3884 12216 3936
rect 13360 3952 13412 4004
rect 12900 3884 12952 3936
rect 13268 3884 13320 3936
rect 14004 4029 14013 4063
rect 14013 4029 14047 4063
rect 14047 4029 14056 4063
rect 14004 4020 14056 4029
rect 14372 4020 14424 4072
rect 15016 4020 15068 4072
rect 14280 3952 14332 4004
rect 14924 3995 14976 4004
rect 14924 3961 14933 3995
rect 14933 3961 14967 3995
rect 14967 3961 14976 3995
rect 14924 3952 14976 3961
rect 15568 4063 15620 4072
rect 15568 4029 15577 4063
rect 15577 4029 15611 4063
rect 15611 4029 15620 4063
rect 15568 4020 15620 4029
rect 15384 3952 15436 4004
rect 16120 3884 16172 3936
rect 5979 3782 6031 3834
rect 6043 3782 6095 3834
rect 6107 3782 6159 3834
rect 6171 3782 6223 3834
rect 10976 3782 11028 3834
rect 11040 3782 11092 3834
rect 11104 3782 11156 3834
rect 11168 3782 11220 3834
rect 1492 3612 1544 3664
rect 1952 3655 2004 3664
rect 1952 3621 1961 3655
rect 1961 3621 1995 3655
rect 1995 3621 2004 3655
rect 1952 3612 2004 3621
rect 2044 3476 2096 3528
rect 4160 3680 4212 3732
rect 4528 3680 4580 3732
rect 3884 3612 3936 3664
rect 6736 3680 6788 3732
rect 8944 3723 8996 3732
rect 6276 3612 6328 3664
rect 8944 3689 8953 3723
rect 8953 3689 8987 3723
rect 8987 3689 8996 3723
rect 8944 3680 8996 3689
rect 9772 3723 9824 3732
rect 9772 3689 9781 3723
rect 9781 3689 9815 3723
rect 9815 3689 9824 3723
rect 9772 3680 9824 3689
rect 9864 3723 9916 3732
rect 9864 3689 9873 3723
rect 9873 3689 9907 3723
rect 9907 3689 9916 3723
rect 9864 3680 9916 3689
rect 10876 3680 10928 3732
rect 4528 3544 4580 3596
rect 5816 3544 5868 3596
rect 5908 3544 5960 3596
rect 4712 3476 4764 3528
rect 1492 3383 1544 3392
rect 1492 3349 1501 3383
rect 1501 3349 1535 3383
rect 1535 3349 1544 3383
rect 1492 3340 1544 3349
rect 2780 3340 2832 3392
rect 3056 3340 3108 3392
rect 4068 3340 4120 3392
rect 6460 3476 6512 3528
rect 6920 3587 6972 3596
rect 6920 3553 6929 3587
rect 6929 3553 6963 3587
rect 6963 3553 6972 3587
rect 6920 3544 6972 3553
rect 7288 3544 7340 3596
rect 8300 3544 8352 3596
rect 9128 3544 9180 3596
rect 9496 3612 9548 3664
rect 10600 3612 10652 3664
rect 12716 3680 12768 3732
rect 13084 3680 13136 3732
rect 15292 3680 15344 3732
rect 12348 3612 12400 3664
rect 12624 3612 12676 3664
rect 14648 3655 14700 3664
rect 14648 3621 14657 3655
rect 14657 3621 14691 3655
rect 14691 3621 14700 3655
rect 14648 3612 14700 3621
rect 15016 3655 15068 3664
rect 15016 3621 15025 3655
rect 15025 3621 15059 3655
rect 15059 3621 15068 3655
rect 15016 3612 15068 3621
rect 15200 3612 15252 3664
rect 11244 3587 11296 3596
rect 11244 3553 11253 3587
rect 11253 3553 11287 3587
rect 11287 3553 11296 3587
rect 11244 3544 11296 3553
rect 11520 3544 11572 3596
rect 11980 3544 12032 3596
rect 12808 3587 12860 3596
rect 12808 3553 12817 3587
rect 12817 3553 12851 3587
rect 12851 3553 12860 3587
rect 12808 3544 12860 3553
rect 12992 3544 13044 3596
rect 13728 3587 13780 3596
rect 6276 3408 6328 3460
rect 6000 3340 6052 3392
rect 7288 3383 7340 3392
rect 7288 3349 7297 3383
rect 7297 3349 7331 3383
rect 7331 3349 7340 3383
rect 7288 3340 7340 3349
rect 8944 3476 8996 3528
rect 9772 3476 9824 3528
rect 9956 3519 10008 3528
rect 9956 3485 9965 3519
rect 9965 3485 9999 3519
rect 9999 3485 10008 3519
rect 9956 3476 10008 3485
rect 10324 3476 10376 3528
rect 10784 3476 10836 3528
rect 12624 3519 12676 3528
rect 12624 3485 12633 3519
rect 12633 3485 12667 3519
rect 12667 3485 12676 3519
rect 12624 3476 12676 3485
rect 13728 3553 13737 3587
rect 13737 3553 13771 3587
rect 13771 3553 13780 3587
rect 13728 3544 13780 3553
rect 13912 3587 13964 3596
rect 13912 3553 13921 3587
rect 13921 3553 13955 3587
rect 13955 3553 13964 3587
rect 13912 3544 13964 3553
rect 13820 3476 13872 3528
rect 9220 3408 9272 3460
rect 7840 3340 7892 3392
rect 9128 3383 9180 3392
rect 9128 3349 9137 3383
rect 9137 3349 9171 3383
rect 9171 3349 9180 3383
rect 9128 3340 9180 3349
rect 9404 3383 9456 3392
rect 9404 3349 9413 3383
rect 9413 3349 9447 3383
rect 9447 3349 9456 3383
rect 9404 3340 9456 3349
rect 9588 3340 9640 3392
rect 10600 3383 10652 3392
rect 10600 3349 10609 3383
rect 10609 3349 10643 3383
rect 10643 3349 10652 3383
rect 10600 3340 10652 3349
rect 10876 3383 10928 3392
rect 10876 3349 10885 3383
rect 10885 3349 10919 3383
rect 10919 3349 10928 3383
rect 10876 3340 10928 3349
rect 11244 3408 11296 3460
rect 12256 3408 12308 3460
rect 12348 3408 12400 3460
rect 13360 3340 13412 3392
rect 14096 3383 14148 3392
rect 14096 3349 14105 3383
rect 14105 3349 14139 3383
rect 14139 3349 14148 3383
rect 14096 3340 14148 3349
rect 3480 3238 3532 3290
rect 3544 3238 3596 3290
rect 3608 3238 3660 3290
rect 3672 3238 3724 3290
rect 8478 3238 8530 3290
rect 8542 3238 8594 3290
rect 8606 3238 8658 3290
rect 8670 3238 8722 3290
rect 13475 3238 13527 3290
rect 13539 3238 13591 3290
rect 13603 3238 13655 3290
rect 13667 3238 13719 3290
rect 4252 3136 4304 3188
rect 5540 3179 5592 3188
rect 5540 3145 5549 3179
rect 5549 3145 5583 3179
rect 5583 3145 5592 3179
rect 5540 3136 5592 3145
rect 8300 3179 8352 3188
rect 8300 3145 8309 3179
rect 8309 3145 8343 3179
rect 8343 3145 8352 3179
rect 8300 3136 8352 3145
rect 1400 3068 1452 3120
rect 2228 3068 2280 3120
rect 5816 3068 5868 3120
rect 1860 3000 1912 3052
rect 2688 3000 2740 3052
rect 4528 3000 4580 3052
rect 6000 3043 6052 3052
rect 6000 3009 6009 3043
rect 6009 3009 6043 3043
rect 6043 3009 6052 3043
rect 6000 3000 6052 3009
rect 6368 3068 6420 3120
rect 9680 3136 9732 3188
rect 11888 3068 11940 3120
rect 11980 3111 12032 3120
rect 11980 3077 11989 3111
rect 11989 3077 12023 3111
rect 12023 3077 12032 3111
rect 11980 3068 12032 3077
rect 14188 3136 14240 3188
rect 14464 3179 14516 3188
rect 14464 3145 14473 3179
rect 14473 3145 14507 3179
rect 14507 3145 14516 3179
rect 14464 3136 14516 3145
rect 1584 2975 1636 2984
rect 1584 2941 1593 2975
rect 1593 2941 1627 2975
rect 1627 2941 1636 2975
rect 1584 2932 1636 2941
rect 2320 2975 2372 2984
rect 2320 2941 2329 2975
rect 2329 2941 2363 2975
rect 2363 2941 2372 2975
rect 2320 2932 2372 2941
rect 2596 2932 2648 2984
rect 3332 2932 3384 2984
rect 4344 2932 4396 2984
rect 4436 2932 4488 2984
rect 5908 2932 5960 2984
rect 7840 2932 7892 2984
rect 572 2864 624 2916
rect 1032 2796 1084 2848
rect 3792 2864 3844 2916
rect 3516 2796 3568 2848
rect 4712 2864 4764 2916
rect 4804 2839 4856 2848
rect 4804 2805 4813 2839
rect 4813 2805 4847 2839
rect 4847 2805 4856 2839
rect 4804 2796 4856 2805
rect 5264 2839 5316 2848
rect 5264 2805 5273 2839
rect 5273 2805 5307 2839
rect 5307 2805 5316 2839
rect 5264 2796 5316 2805
rect 5540 2864 5592 2916
rect 8484 2932 8536 2984
rect 9128 2932 9180 2984
rect 9772 2932 9824 2984
rect 6644 2796 6696 2848
rect 9036 2864 9088 2916
rect 10232 2864 10284 2916
rect 9956 2796 10008 2848
rect 10600 2796 10652 2848
rect 10784 2864 10836 2916
rect 11612 2932 11664 2984
rect 11704 2932 11756 2984
rect 12532 2864 12584 2916
rect 13452 2932 13504 2984
rect 14740 2932 14792 2984
rect 14004 2864 14056 2916
rect 15476 2864 15528 2916
rect 11888 2796 11940 2848
rect 12808 2839 12860 2848
rect 12808 2805 12817 2839
rect 12817 2805 12851 2839
rect 12851 2805 12860 2839
rect 12808 2796 12860 2805
rect 14740 2839 14792 2848
rect 14740 2805 14749 2839
rect 14749 2805 14783 2839
rect 14783 2805 14792 2839
rect 14740 2796 14792 2805
rect 5979 2694 6031 2746
rect 6043 2694 6095 2746
rect 6107 2694 6159 2746
rect 6171 2694 6223 2746
rect 10976 2694 11028 2746
rect 11040 2694 11092 2746
rect 11104 2694 11156 2746
rect 11168 2694 11220 2746
rect 3516 2635 3568 2644
rect 3516 2601 3525 2635
rect 3525 2601 3559 2635
rect 3559 2601 3568 2635
rect 3516 2592 3568 2601
rect 3792 2592 3844 2644
rect 4344 2592 4396 2644
rect 5264 2592 5316 2644
rect 5632 2592 5684 2644
rect 5816 2592 5868 2644
rect 6736 2592 6788 2644
rect 7196 2592 7248 2644
rect 9220 2635 9272 2644
rect 2136 2456 2188 2508
rect 3148 2456 3200 2508
rect 2044 2431 2096 2440
rect 2044 2397 2053 2431
rect 2053 2397 2087 2431
rect 2087 2397 2096 2431
rect 2044 2388 2096 2397
rect 4804 2524 4856 2576
rect 4068 2499 4120 2508
rect 4068 2465 4077 2499
rect 4077 2465 4111 2499
rect 4111 2465 4120 2499
rect 4068 2456 4120 2465
rect 5540 2456 5592 2508
rect 7288 2524 7340 2576
rect 9220 2601 9229 2635
rect 9229 2601 9263 2635
rect 9263 2601 9272 2635
rect 9220 2592 9272 2601
rect 11336 2592 11388 2644
rect 12624 2592 12676 2644
rect 12808 2592 12860 2644
rect 13360 2635 13412 2644
rect 13360 2601 13369 2635
rect 13369 2601 13403 2635
rect 13403 2601 13412 2635
rect 14188 2635 14240 2644
rect 13360 2592 13412 2601
rect 14188 2601 14197 2635
rect 14197 2601 14231 2635
rect 14231 2601 14240 2635
rect 14188 2592 14240 2601
rect 6276 2456 6328 2508
rect 4620 2388 4672 2440
rect 4988 2431 5040 2440
rect 4988 2397 4997 2431
rect 4997 2397 5031 2431
rect 5031 2397 5040 2431
rect 4988 2388 5040 2397
rect 6368 2388 6420 2440
rect 204 2320 256 2372
rect 4804 2320 4856 2372
rect 4160 2252 4212 2304
rect 4344 2252 4396 2304
rect 5632 2320 5684 2372
rect 8484 2524 8536 2576
rect 8852 2456 8904 2508
rect 9036 2456 9088 2508
rect 9404 2524 9456 2576
rect 13176 2524 13228 2576
rect 14740 2524 14792 2576
rect 10876 2456 10928 2508
rect 7656 2431 7708 2440
rect 7656 2397 7665 2431
rect 7665 2397 7699 2431
rect 7699 2397 7708 2431
rect 7656 2388 7708 2397
rect 8300 2388 8352 2440
rect 10600 2431 10652 2440
rect 10600 2397 10609 2431
rect 10609 2397 10643 2431
rect 10643 2397 10652 2431
rect 10600 2388 10652 2397
rect 10784 2388 10836 2440
rect 11336 2431 11388 2440
rect 11336 2397 11345 2431
rect 11345 2397 11379 2431
rect 11379 2397 11388 2431
rect 11336 2388 11388 2397
rect 11980 2456 12032 2508
rect 12716 2456 12768 2508
rect 14096 2456 14148 2508
rect 14832 2499 14884 2508
rect 14832 2465 14841 2499
rect 14841 2465 14875 2499
rect 14875 2465 14884 2499
rect 14832 2456 14884 2465
rect 15476 2499 15528 2508
rect 15476 2465 15485 2499
rect 15485 2465 15519 2499
rect 15519 2465 15528 2499
rect 15476 2456 15528 2465
rect 12624 2431 12676 2440
rect 12624 2397 12633 2431
rect 12633 2397 12667 2431
rect 12667 2397 12676 2431
rect 12624 2388 12676 2397
rect 11796 2320 11848 2372
rect 12440 2320 12492 2372
rect 12900 2363 12952 2372
rect 12900 2329 12909 2363
rect 12909 2329 12943 2363
rect 12943 2329 12952 2363
rect 12900 2320 12952 2329
rect 14004 2388 14056 2440
rect 15108 2388 15160 2440
rect 14280 2320 14332 2372
rect 6736 2252 6788 2304
rect 7104 2252 7156 2304
rect 9312 2252 9364 2304
rect 12256 2252 12308 2304
rect 16948 2252 17000 2304
rect 3480 2150 3532 2202
rect 3544 2150 3596 2202
rect 3608 2150 3660 2202
rect 3672 2150 3724 2202
rect 8478 2150 8530 2202
rect 8542 2150 8594 2202
rect 8606 2150 8658 2202
rect 8670 2150 8722 2202
rect 13475 2150 13527 2202
rect 13539 2150 13591 2202
rect 13603 2150 13655 2202
rect 13667 2150 13719 2202
rect 4988 2048 5040 2100
rect 6552 2048 6604 2100
rect 4160 1980 4212 2032
rect 12624 2048 12676 2100
rect 4068 1912 4120 1964
rect 14648 1980 14700 2032
rect 3608 1844 3660 1896
rect 5356 1844 5408 1896
rect 11888 1844 11940 1896
rect 13820 1844 13872 1896
rect 6000 1436 6052 1488
rect 7656 1436 7708 1488
rect 5172 1368 5224 1420
rect 6736 1368 6788 1420
<< metal2 >>
rect 202 19200 258 20000
rect 570 19200 626 20000
rect 938 19200 994 20000
rect 1398 19200 1454 20000
rect 1766 19200 1822 20000
rect 2226 19200 2282 20000
rect 2594 19200 2650 20000
rect 2962 19544 3018 19553
rect 2962 19479 3018 19488
rect 216 15366 244 19200
rect 584 17270 612 19200
rect 952 17338 980 19200
rect 1412 17354 1440 19200
rect 940 17332 992 17338
rect 1412 17326 1532 17354
rect 940 17274 992 17280
rect 1504 17270 1532 17326
rect 572 17264 624 17270
rect 572 17206 624 17212
rect 1492 17264 1544 17270
rect 1492 17206 1544 17212
rect 1780 17202 1808 19200
rect 1858 17640 1914 17649
rect 1858 17575 1914 17584
rect 1768 17196 1820 17202
rect 1768 17138 1820 17144
rect 1676 17060 1728 17066
rect 1676 17002 1728 17008
rect 1400 16720 1452 16726
rect 1398 16688 1400 16697
rect 1452 16688 1454 16697
rect 1398 16623 1454 16632
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1490 15736 1546 15745
rect 1490 15671 1492 15680
rect 1544 15671 1546 15680
rect 1492 15642 1544 15648
rect 1596 15434 1624 16594
rect 1584 15428 1636 15434
rect 1584 15370 1636 15376
rect 204 15360 256 15366
rect 204 15302 256 15308
rect 1584 14884 1636 14890
rect 1584 14826 1636 14832
rect 1492 14816 1544 14822
rect 1490 14784 1492 14793
rect 1544 14784 1546 14793
rect 1490 14719 1546 14728
rect 1596 14074 1624 14826
rect 1688 14618 1716 17002
rect 1872 16794 1900 17575
rect 2240 17270 2268 19200
rect 2228 17264 2280 17270
rect 2228 17206 2280 17212
rect 2502 17096 2558 17105
rect 2136 17060 2188 17066
rect 2136 17002 2188 17008
rect 2228 17060 2280 17066
rect 2502 17031 2558 17040
rect 2228 17002 2280 17008
rect 2148 16794 2176 17002
rect 1860 16788 1912 16794
rect 1860 16730 1912 16736
rect 2136 16788 2188 16794
rect 2136 16730 2188 16736
rect 1952 16652 2004 16658
rect 1952 16594 2004 16600
rect 1964 15706 1992 16594
rect 2044 16040 2096 16046
rect 2044 15982 2096 15988
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 1676 14612 1728 14618
rect 1676 14554 1728 14560
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 2056 14006 2084 15982
rect 2134 15736 2190 15745
rect 2134 15671 2190 15680
rect 2148 15570 2176 15671
rect 2136 15564 2188 15570
rect 2136 15506 2188 15512
rect 2240 15162 2268 17002
rect 2412 16652 2464 16658
rect 2412 16594 2464 16600
rect 2424 16454 2452 16594
rect 2412 16448 2464 16454
rect 2412 16390 2464 16396
rect 2228 15156 2280 15162
rect 2228 15098 2280 15104
rect 2136 14816 2188 14822
rect 2136 14758 2188 14764
rect 2044 14000 2096 14006
rect 1950 13968 2006 13977
rect 2044 13942 2096 13948
rect 1950 13903 2006 13912
rect 1964 13870 1992 13903
rect 1400 13864 1452 13870
rect 1398 13832 1400 13841
rect 1952 13864 2004 13870
rect 1452 13832 1454 13841
rect 1952 13806 2004 13812
rect 1398 13767 1454 13776
rect 1676 13796 1728 13802
rect 1676 13738 1728 13744
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 1400 12912 1452 12918
rect 1398 12880 1400 12889
rect 1452 12880 1454 12889
rect 1398 12815 1454 12824
rect 1596 12782 1624 13126
rect 1688 12986 1716 13738
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 1584 12776 1636 12782
rect 1584 12718 1636 12724
rect 1860 12300 1912 12306
rect 1860 12242 1912 12248
rect 1492 12096 1544 12102
rect 1492 12038 1544 12044
rect 1504 11937 1532 12038
rect 1490 11928 1546 11937
rect 1490 11863 1546 11872
rect 1872 11354 1900 12242
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1584 11212 1636 11218
rect 1584 11154 1636 11160
rect 1400 11076 1452 11082
rect 1400 11018 1452 11024
rect 1412 10985 1440 11018
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 1596 10810 1624 11154
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1398 10024 1454 10033
rect 1398 9959 1400 9968
rect 1452 9959 1454 9968
rect 1400 9930 1452 9936
rect 1400 9104 1452 9110
rect 1398 9072 1400 9081
rect 1452 9072 1454 9081
rect 1398 9007 1454 9016
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1596 8634 1624 8978
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1490 8120 1546 8129
rect 1490 8055 1492 8064
rect 1544 8055 1546 8064
rect 1492 8026 1544 8032
rect 2056 7546 2084 13942
rect 2148 13394 2176 14758
rect 2136 13388 2188 13394
rect 2136 13330 2188 13336
rect 2424 12646 2452 16390
rect 2516 15570 2544 17031
rect 2608 16726 2636 19200
rect 2688 17060 2740 17066
rect 2688 17002 2740 17008
rect 2872 17060 2924 17066
rect 2872 17002 2924 17008
rect 2596 16720 2648 16726
rect 2596 16662 2648 16668
rect 2700 16250 2728 17002
rect 2780 16516 2832 16522
rect 2780 16458 2832 16464
rect 2792 16250 2820 16458
rect 2688 16244 2740 16250
rect 2688 16186 2740 16192
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 2884 15910 2912 17002
rect 2976 16182 3004 19479
rect 3054 19200 3110 20000
rect 3422 19200 3478 20000
rect 3882 19200 3938 20000
rect 4250 19200 4306 20000
rect 4618 19200 4674 20000
rect 5078 19200 5134 20000
rect 5446 19200 5502 20000
rect 5906 19200 5962 20000
rect 6274 19200 6330 20000
rect 6734 19200 6790 20000
rect 7102 19200 7158 20000
rect 7562 19200 7618 20000
rect 7930 19200 7986 20000
rect 8390 19200 8446 20000
rect 8758 19200 8814 20000
rect 9126 19200 9182 20000
rect 9586 19200 9642 20000
rect 9954 19200 10010 20000
rect 10414 19200 10470 20000
rect 10782 19200 10838 20000
rect 11242 19200 11298 20000
rect 11610 19200 11666 20000
rect 12070 19200 12126 20000
rect 12438 19200 12494 20000
rect 12898 19200 12954 20000
rect 13266 19200 13322 20000
rect 13634 19200 13690 20000
rect 14094 19200 14150 20000
rect 14462 19200 14518 20000
rect 14922 19200 14978 20000
rect 15290 19200 15346 20000
rect 15750 19200 15806 20000
rect 16118 19200 16174 20000
rect 16578 19200 16634 20000
rect 16946 19200 17002 20000
rect 3068 16726 3096 19200
rect 3146 18592 3202 18601
rect 3146 18527 3202 18536
rect 3056 16720 3108 16726
rect 3056 16662 3108 16668
rect 2964 16176 3016 16182
rect 2964 16118 3016 16124
rect 2964 16040 3016 16046
rect 2962 16008 2964 16017
rect 3016 16008 3018 16017
rect 2962 15943 3018 15952
rect 2596 15904 2648 15910
rect 2872 15904 2924 15910
rect 2648 15864 2820 15892
rect 2596 15846 2648 15852
rect 2504 15564 2556 15570
rect 2792 15552 2820 15864
rect 2872 15846 2924 15852
rect 3160 15638 3188 18527
rect 3436 17626 3464 19200
rect 3344 17598 3464 17626
rect 3344 16726 3372 17598
rect 3454 17436 3750 17456
rect 3510 17434 3534 17436
rect 3590 17434 3614 17436
rect 3670 17434 3694 17436
rect 3532 17382 3534 17434
rect 3596 17382 3608 17434
rect 3670 17382 3672 17434
rect 3510 17380 3534 17382
rect 3590 17380 3614 17382
rect 3670 17380 3694 17382
rect 3454 17360 3750 17380
rect 3896 16726 3924 19200
rect 3976 17604 4028 17610
rect 3976 17546 4028 17552
rect 3988 17134 4016 17546
rect 3976 17128 4028 17134
rect 3976 17070 4028 17076
rect 4264 16726 4292 19200
rect 4344 17536 4396 17542
rect 4344 17478 4396 17484
rect 4356 17066 4384 17478
rect 4632 17270 4660 19200
rect 5092 17270 5120 19200
rect 5460 17270 5488 19200
rect 5920 17270 5948 19200
rect 6288 17270 6316 19200
rect 6748 17270 6776 19200
rect 7116 17338 7144 19200
rect 7472 17536 7524 17542
rect 7472 17478 7524 17484
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 4620 17264 4672 17270
rect 4620 17206 4672 17212
rect 5080 17264 5132 17270
rect 5080 17206 5132 17212
rect 5448 17264 5500 17270
rect 5448 17206 5500 17212
rect 5908 17264 5960 17270
rect 5908 17206 5960 17212
rect 6276 17264 6328 17270
rect 6276 17206 6328 17212
rect 6736 17264 6788 17270
rect 6736 17206 6788 17212
rect 4344 17060 4396 17066
rect 4344 17002 4396 17008
rect 4804 17060 4856 17066
rect 4804 17002 4856 17008
rect 5080 17060 5132 17066
rect 5080 17002 5132 17008
rect 5632 17060 5684 17066
rect 5632 17002 5684 17008
rect 5816 17060 5868 17066
rect 5816 17002 5868 17008
rect 6736 17060 6788 17066
rect 6736 17002 6788 17008
rect 7104 17060 7156 17066
rect 7104 17002 7156 17008
rect 3332 16720 3384 16726
rect 3332 16662 3384 16668
rect 3884 16720 3936 16726
rect 3884 16662 3936 16668
rect 4252 16720 4304 16726
rect 4252 16662 4304 16668
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 3792 16652 3844 16658
rect 3792 16594 3844 16600
rect 3976 16652 4028 16658
rect 3976 16594 4028 16600
rect 3252 16250 3280 16594
rect 3454 16348 3750 16368
rect 3510 16346 3534 16348
rect 3590 16346 3614 16348
rect 3670 16346 3694 16348
rect 3532 16294 3534 16346
rect 3596 16294 3608 16346
rect 3670 16294 3672 16346
rect 3510 16292 3534 16294
rect 3590 16292 3614 16294
rect 3670 16292 3694 16294
rect 3454 16272 3750 16292
rect 3804 16250 3832 16594
rect 3988 16250 4016 16594
rect 4816 16250 4844 17002
rect 5092 16794 5120 17002
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5080 16788 5132 16794
rect 5080 16730 5132 16736
rect 5460 16658 5488 16934
rect 5540 16720 5592 16726
rect 5540 16662 5592 16668
rect 4896 16652 4948 16658
rect 4896 16594 4948 16600
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 3240 16244 3292 16250
rect 3240 16186 3292 16192
rect 3792 16244 3844 16250
rect 3792 16186 3844 16192
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 4804 16244 4856 16250
rect 4804 16186 4856 16192
rect 4160 16176 4212 16182
rect 4160 16118 4212 16124
rect 3240 16108 3292 16114
rect 3240 16050 3292 16056
rect 3976 16108 4028 16114
rect 3976 16050 4028 16056
rect 3148 15632 3200 15638
rect 3148 15574 3200 15580
rect 2792 15524 2912 15552
rect 2504 15506 2556 15512
rect 2778 15464 2834 15473
rect 2778 15399 2834 15408
rect 2792 15366 2820 15399
rect 2780 15360 2832 15366
rect 2780 15302 2832 15308
rect 2884 15162 2912 15524
rect 2872 15156 2924 15162
rect 2872 15098 2924 15104
rect 2780 15020 2832 15026
rect 2780 14962 2832 14968
rect 2596 14816 2648 14822
rect 2792 14793 2820 14962
rect 2596 14758 2648 14764
rect 2778 14784 2834 14793
rect 2608 14074 2636 14758
rect 2778 14719 2834 14728
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 2688 14476 2740 14482
rect 2688 14418 2740 14424
rect 2596 14068 2648 14074
rect 2596 14010 2648 14016
rect 2596 13728 2648 13734
rect 2596 13670 2648 13676
rect 2608 13530 2636 13670
rect 2596 13524 2648 13530
rect 2596 13466 2648 13472
rect 2700 13394 2728 14418
rect 2792 13938 2820 14554
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2884 13530 2912 15098
rect 2964 15088 3016 15094
rect 2964 15030 3016 15036
rect 2976 14822 3004 15030
rect 3148 15020 3200 15026
rect 3148 14962 3200 14968
rect 3160 14929 3188 14962
rect 3146 14920 3202 14929
rect 3146 14855 3202 14864
rect 2964 14816 3016 14822
rect 2964 14758 3016 14764
rect 3160 14006 3188 14855
rect 3148 14000 3200 14006
rect 3148 13942 3200 13948
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2688 13388 2740 13394
rect 2688 13330 2740 13336
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 3160 12986 3188 13262
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 2412 12640 2464 12646
rect 2412 12582 2464 12588
rect 2688 12640 2740 12646
rect 2688 12582 2740 12588
rect 2320 12300 2372 12306
rect 2320 12242 2372 12248
rect 2332 11558 2360 12242
rect 2700 12102 2728 12582
rect 2792 12374 2820 12718
rect 2884 12646 2912 12854
rect 2872 12640 2924 12646
rect 2872 12582 2924 12588
rect 2780 12368 2832 12374
rect 2780 12310 2832 12316
rect 2688 12096 2740 12102
rect 2688 12038 2740 12044
rect 2792 11830 2820 12310
rect 2780 11824 2832 11830
rect 2780 11766 2832 11772
rect 2792 11694 2820 11766
rect 2688 11688 2740 11694
rect 2688 11630 2740 11636
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2332 11286 2360 11494
rect 2320 11280 2372 11286
rect 2320 11222 2372 11228
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2332 10810 2360 11086
rect 2320 10804 2372 10810
rect 2320 10746 2372 10752
rect 2700 10674 2728 11630
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 3160 11150 3188 11494
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 2872 11008 2924 11014
rect 2872 10950 2924 10956
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 2884 10606 2912 10950
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 2872 8832 2924 8838
rect 3056 8832 3108 8838
rect 2872 8774 2924 8780
rect 2976 8792 3056 8820
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2792 7546 2820 7822
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 2320 7540 2372 7546
rect 2320 7482 2372 7488
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 1492 7200 1544 7206
rect 1490 7168 1492 7177
rect 1544 7168 1546 7177
rect 1490 7103 1546 7112
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1504 6225 1532 6598
rect 1490 6216 1546 6225
rect 1490 6151 1546 6160
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1596 5846 1624 6054
rect 1780 5914 1808 6802
rect 1860 6452 1912 6458
rect 1860 6394 1912 6400
rect 1768 5908 1820 5914
rect 1768 5850 1820 5856
rect 1584 5840 1636 5846
rect 1584 5782 1636 5788
rect 1492 5568 1544 5574
rect 1492 5510 1544 5516
rect 1400 5296 1452 5302
rect 1398 5264 1400 5273
rect 1452 5264 1454 5273
rect 1398 5199 1454 5208
rect 1504 5166 1532 5510
rect 1492 5160 1544 5166
rect 1492 5102 1544 5108
rect 1676 4684 1728 4690
rect 1676 4626 1728 4632
rect 1492 4480 1544 4486
rect 1492 4422 1544 4428
rect 1398 4312 1454 4321
rect 1398 4247 1454 4256
rect 1412 4146 1440 4247
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1504 3670 1532 4422
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1492 3664 1544 3670
rect 1492 3606 1544 3612
rect 1492 3392 1544 3398
rect 1490 3360 1492 3369
rect 1544 3360 1546 3369
rect 1490 3295 1546 3304
rect 1400 3120 1452 3126
rect 1400 3062 1452 3068
rect 572 2916 624 2922
rect 572 2858 624 2864
rect 204 2372 256 2378
rect 204 2314 256 2320
rect 216 800 244 2314
rect 584 800 612 2858
rect 1032 2848 1084 2854
rect 1032 2790 1084 2796
rect 1044 800 1072 2790
rect 1412 800 1440 3062
rect 1596 2990 1624 3878
rect 1584 2984 1636 2990
rect 1688 2961 1716 4626
rect 1768 4480 1820 4486
rect 1768 4422 1820 4428
rect 1780 4078 1808 4422
rect 1872 4078 1900 6394
rect 1964 6118 1992 6802
rect 1952 6112 2004 6118
rect 1952 6054 2004 6060
rect 2056 5930 2084 7482
rect 2332 7206 2360 7482
rect 2884 7410 2912 8774
rect 2976 8362 3004 8792
rect 3056 8774 3108 8780
rect 2964 8356 3016 8362
rect 2964 8298 3016 8304
rect 2976 7818 3004 8298
rect 2964 7812 3016 7818
rect 2964 7754 3016 7760
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2976 7342 3004 7754
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 2320 7200 2372 7206
rect 2320 7142 2372 7148
rect 2228 6180 2280 6186
rect 2228 6122 2280 6128
rect 1964 5902 2084 5930
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1860 4072 1912 4078
rect 1860 4014 1912 4020
rect 1964 3670 1992 5902
rect 2136 5772 2188 5778
rect 2136 5714 2188 5720
rect 2148 5302 2176 5714
rect 2136 5296 2188 5302
rect 2136 5238 2188 5244
rect 2044 5024 2096 5030
rect 2044 4966 2096 4972
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 2056 4826 2084 4966
rect 2148 4826 2176 4966
rect 2044 4820 2096 4826
rect 2044 4762 2096 4768
rect 2136 4820 2188 4826
rect 2136 4762 2188 4768
rect 2240 4729 2268 6122
rect 2226 4720 2282 4729
rect 2136 4684 2188 4690
rect 2188 4664 2226 4672
rect 2188 4655 2282 4664
rect 2188 4644 2268 4655
rect 2136 4626 2188 4632
rect 1952 3664 2004 3670
rect 1952 3606 2004 3612
rect 2044 3528 2096 3534
rect 2044 3470 2096 3476
rect 1860 3052 1912 3058
rect 1860 2994 1912 3000
rect 1584 2926 1636 2932
rect 1674 2952 1730 2961
rect 1674 2887 1730 2896
rect 1872 800 1900 2994
rect 2056 2446 2084 3470
rect 2148 2514 2176 4626
rect 2240 4595 2268 4644
rect 2332 4078 2360 7142
rect 2504 6928 2556 6934
rect 2504 6870 2556 6876
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2424 5370 2452 5646
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 2516 4078 2544 6870
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 2700 6458 2728 6802
rect 2976 6662 3004 7278
rect 3160 6730 3188 11086
rect 3252 7834 3280 16050
rect 3424 16040 3476 16046
rect 3424 15982 3476 15988
rect 3436 15910 3464 15982
rect 3988 15910 4016 16050
rect 3424 15904 3476 15910
rect 3424 15846 3476 15852
rect 3976 15904 4028 15910
rect 3976 15846 4028 15852
rect 3330 15600 3386 15609
rect 3330 15535 3386 15544
rect 3344 15366 3372 15535
rect 3332 15360 3384 15366
rect 3332 15302 3384 15308
rect 3454 15260 3750 15280
rect 3510 15258 3534 15260
rect 3590 15258 3614 15260
rect 3670 15258 3694 15260
rect 3532 15206 3534 15258
rect 3596 15206 3608 15258
rect 3670 15206 3672 15258
rect 3510 15204 3534 15206
rect 3590 15204 3614 15206
rect 3670 15204 3694 15206
rect 3454 15184 3750 15204
rect 3792 15088 3844 15094
rect 3792 15030 3844 15036
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 3712 14618 3740 14758
rect 3700 14612 3752 14618
rect 3700 14554 3752 14560
rect 3804 14414 3832 15030
rect 3884 15020 3936 15026
rect 3884 14962 3936 14968
rect 3896 14550 3924 14962
rect 3884 14544 3936 14550
rect 3884 14486 3936 14492
rect 3792 14408 3844 14414
rect 3792 14350 3844 14356
rect 3454 14172 3750 14192
rect 3510 14170 3534 14172
rect 3590 14170 3614 14172
rect 3670 14170 3694 14172
rect 3532 14118 3534 14170
rect 3596 14118 3608 14170
rect 3670 14118 3672 14170
rect 3510 14116 3534 14118
rect 3590 14116 3614 14118
rect 3670 14116 3694 14118
rect 3454 14096 3750 14116
rect 3424 13728 3476 13734
rect 3988 13716 4016 15846
rect 4172 15366 4200 16118
rect 4264 16017 4292 16186
rect 4250 16008 4306 16017
rect 4250 15943 4306 15952
rect 4344 15904 4396 15910
rect 4344 15846 4396 15852
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 4080 15065 4108 15098
rect 4066 15056 4122 15065
rect 4066 14991 4122 15000
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 4080 14074 4108 14758
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 4068 13728 4120 13734
rect 3988 13688 4068 13716
rect 3424 13670 3476 13676
rect 4068 13670 4120 13676
rect 3436 13530 3464 13670
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 3884 13524 3936 13530
rect 3884 13466 3936 13472
rect 3454 13084 3750 13104
rect 3510 13082 3534 13084
rect 3590 13082 3614 13084
rect 3670 13082 3694 13084
rect 3532 13030 3534 13082
rect 3596 13030 3608 13082
rect 3670 13030 3672 13082
rect 3510 13028 3534 13030
rect 3590 13028 3614 13030
rect 3670 13028 3694 13030
rect 3454 13008 3750 13028
rect 3424 12708 3476 12714
rect 3424 12650 3476 12656
rect 3436 12442 3464 12650
rect 3424 12436 3476 12442
rect 3424 12378 3476 12384
rect 3454 11996 3750 12016
rect 3510 11994 3534 11996
rect 3590 11994 3614 11996
rect 3670 11994 3694 11996
rect 3532 11942 3534 11994
rect 3596 11942 3608 11994
rect 3670 11942 3672 11994
rect 3510 11940 3534 11942
rect 3590 11940 3614 11942
rect 3670 11940 3694 11942
rect 3454 11920 3750 11940
rect 3332 11892 3384 11898
rect 3332 11834 3384 11840
rect 3344 11286 3372 11834
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3332 11280 3384 11286
rect 3332 11222 3384 11228
rect 3804 11082 3832 11698
rect 3896 11642 3924 13466
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 3988 12442 4016 12922
rect 3976 12436 4028 12442
rect 3976 12378 4028 12384
rect 4080 11937 4108 13670
rect 4356 12850 4384 15846
rect 4908 15434 4936 16594
rect 5080 15904 5132 15910
rect 5080 15846 5132 15852
rect 5092 15706 5120 15846
rect 5080 15700 5132 15706
rect 5080 15642 5132 15648
rect 4896 15428 4948 15434
rect 4896 15370 4948 15376
rect 4620 15360 4672 15366
rect 4620 15302 4672 15308
rect 4528 14884 4580 14890
rect 4528 14826 4580 14832
rect 4540 14793 4568 14826
rect 4526 14784 4582 14793
rect 4526 14719 4582 14728
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 4448 13802 4476 14010
rect 4436 13796 4488 13802
rect 4436 13738 4488 13744
rect 4528 13728 4580 13734
rect 4528 13670 4580 13676
rect 4540 13258 4568 13670
rect 4528 13252 4580 13258
rect 4528 13194 4580 13200
rect 4344 12844 4396 12850
rect 4344 12786 4396 12792
rect 4160 12708 4212 12714
rect 4160 12650 4212 12656
rect 4066 11928 4122 11937
rect 4066 11863 4122 11872
rect 3896 11614 4016 11642
rect 4172 11626 4200 12650
rect 4356 11898 4384 12786
rect 4436 12640 4488 12646
rect 4436 12582 4488 12588
rect 4448 11898 4476 12582
rect 4344 11892 4396 11898
rect 4344 11834 4396 11840
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 3896 11354 3924 11494
rect 3988 11370 4016 11614
rect 4160 11620 4212 11626
rect 4160 11562 4212 11568
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 3884 11348 3936 11354
rect 3988 11342 4108 11370
rect 4264 11354 4292 11494
rect 3884 11290 3936 11296
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 3792 11076 3844 11082
rect 3792 11018 3844 11024
rect 3454 10908 3750 10928
rect 3510 10906 3534 10908
rect 3590 10906 3614 10908
rect 3670 10906 3694 10908
rect 3532 10854 3534 10906
rect 3596 10854 3608 10906
rect 3670 10854 3672 10906
rect 3510 10852 3534 10854
rect 3590 10852 3614 10854
rect 3670 10852 3694 10854
rect 3454 10832 3750 10852
rect 3988 10810 4016 11154
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 3884 10532 3936 10538
rect 3884 10474 3936 10480
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3344 10266 3372 10406
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3454 9820 3750 9840
rect 3510 9818 3534 9820
rect 3590 9818 3614 9820
rect 3670 9818 3694 9820
rect 3532 9766 3534 9818
rect 3596 9766 3608 9818
rect 3670 9766 3672 9818
rect 3510 9764 3534 9766
rect 3590 9764 3614 9766
rect 3670 9764 3694 9766
rect 3454 9744 3750 9764
rect 3896 9722 3924 10474
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3344 9178 3372 9318
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3792 8900 3844 8906
rect 3792 8842 3844 8848
rect 3454 8732 3750 8752
rect 3510 8730 3534 8732
rect 3590 8730 3614 8732
rect 3670 8730 3694 8732
rect 3532 8678 3534 8730
rect 3596 8678 3608 8730
rect 3670 8678 3672 8730
rect 3510 8676 3534 8678
rect 3590 8676 3614 8678
rect 3670 8676 3694 8678
rect 3454 8656 3750 8676
rect 3804 8634 3832 8842
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3252 7806 3372 7834
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 3252 7546 3280 7686
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 3148 6724 3200 6730
rect 3148 6666 3200 6672
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 2688 6180 2740 6186
rect 2688 6122 2740 6128
rect 2700 5710 2728 6122
rect 2688 5704 2740 5710
rect 2688 5646 2740 5652
rect 2700 5234 2728 5646
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2884 5234 2912 5510
rect 2688 5228 2740 5234
rect 2688 5170 2740 5176
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 2976 5166 3004 6326
rect 3160 6118 3188 6666
rect 3252 6662 3280 7210
rect 3344 7002 3372 7806
rect 3454 7644 3750 7664
rect 3510 7642 3534 7644
rect 3590 7642 3614 7644
rect 3670 7642 3694 7644
rect 3532 7590 3534 7642
rect 3596 7590 3608 7642
rect 3670 7590 3672 7642
rect 3510 7588 3534 7590
rect 3590 7588 3614 7590
rect 3670 7588 3694 7590
rect 3454 7568 3750 7588
rect 3424 7268 3476 7274
rect 3424 7210 3476 7216
rect 3332 6996 3384 7002
rect 3332 6938 3384 6944
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 2964 5160 3016 5166
rect 2964 5102 3016 5108
rect 3160 4690 3188 6054
rect 3252 5234 3280 6598
rect 3344 6458 3372 6938
rect 3436 6934 3464 7210
rect 3424 6928 3476 6934
rect 3424 6870 3476 6876
rect 3454 6556 3750 6576
rect 3510 6554 3534 6556
rect 3590 6554 3614 6556
rect 3670 6554 3694 6556
rect 3532 6502 3534 6554
rect 3596 6502 3608 6554
rect 3670 6502 3672 6554
rect 3510 6500 3534 6502
rect 3590 6500 3614 6502
rect 3670 6500 3694 6502
rect 3454 6480 3750 6500
rect 3332 6452 3384 6458
rect 3384 6412 3464 6440
rect 3332 6394 3384 6400
rect 3332 6248 3384 6254
rect 3332 6190 3384 6196
rect 3344 5574 3372 6190
rect 3436 5778 3464 6412
rect 3424 5772 3476 5778
rect 3896 5760 3924 9658
rect 4080 7886 4108 11342
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4356 10810 4384 11494
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 4172 9042 4200 9522
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 4172 8430 4200 8978
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4160 8424 4212 8430
rect 4160 8366 4212 8372
rect 4264 8362 4292 8434
rect 4252 8356 4304 8362
rect 4252 8298 4304 8304
rect 4344 8288 4396 8294
rect 4344 8230 4396 8236
rect 4356 8090 4384 8230
rect 4344 8084 4396 8090
rect 4344 8026 4396 8032
rect 4540 7970 4568 13194
rect 4632 12434 4660 15302
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 4724 13938 4752 14418
rect 4804 14000 4856 14006
rect 4804 13942 4856 13948
rect 4712 13932 4764 13938
rect 4712 13874 4764 13880
rect 4724 13326 4752 13874
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4724 12986 4752 13262
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4816 12442 4844 13942
rect 4804 12436 4856 12442
rect 4632 12406 4752 12434
rect 4620 8356 4672 8362
rect 4620 8298 4672 8304
rect 4356 7954 4568 7970
rect 4344 7948 4568 7954
rect 4396 7942 4568 7948
rect 4344 7890 4396 7896
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 4080 6934 4108 7822
rect 4068 6928 4120 6934
rect 4068 6870 4120 6876
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 4264 5914 4292 6598
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 3424 5714 3476 5720
rect 3804 5732 3924 5760
rect 3332 5568 3384 5574
rect 3332 5510 3384 5516
rect 3344 5234 3372 5510
rect 3454 5468 3750 5488
rect 3510 5466 3534 5468
rect 3590 5466 3614 5468
rect 3670 5466 3694 5468
rect 3532 5414 3534 5466
rect 3596 5414 3608 5466
rect 3670 5414 3672 5466
rect 3510 5412 3534 5414
rect 3590 5412 3614 5414
rect 3670 5412 3694 5414
rect 3454 5392 3750 5412
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3700 5092 3752 5098
rect 3700 5034 3752 5040
rect 3332 5024 3384 5030
rect 3332 4966 3384 4972
rect 3148 4684 3200 4690
rect 3148 4626 3200 4632
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 3068 4282 3096 4558
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 2320 4072 2372 4078
rect 2320 4014 2372 4020
rect 2504 4072 2556 4078
rect 2504 4014 2556 4020
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 2228 3120 2280 3126
rect 2228 3062 2280 3068
rect 2136 2508 2188 2514
rect 2136 2450 2188 2456
rect 2044 2440 2096 2446
rect 2044 2382 2096 2388
rect 2240 800 2268 3062
rect 2332 2990 2360 3878
rect 2608 2990 2636 3878
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 2688 3052 2740 3058
rect 2688 2994 2740 3000
rect 2320 2984 2372 2990
rect 2320 2926 2372 2932
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 2700 800 2728 2994
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1398 0 1454 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2686 0 2742 800
rect 2792 513 2820 3334
rect 3068 800 3096 3334
rect 3160 2514 3188 4626
rect 3240 4004 3292 4010
rect 3240 3946 3292 3952
rect 3252 2774 3280 3946
rect 3344 2990 3372 4966
rect 3712 4826 3740 5034
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3712 4593 3740 4762
rect 3804 4758 3832 5732
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 3884 5636 3936 5642
rect 3884 5578 3936 5584
rect 3896 4826 3924 5578
rect 4172 5370 4200 5646
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4160 5160 4212 5166
rect 4080 5120 4160 5148
rect 3976 5092 4028 5098
rect 3976 5034 4028 5040
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 3792 4752 3844 4758
rect 3792 4694 3844 4700
rect 3698 4584 3754 4593
rect 3698 4519 3754 4528
rect 3454 4380 3750 4400
rect 3510 4378 3534 4380
rect 3590 4378 3614 4380
rect 3670 4378 3694 4380
rect 3532 4326 3534 4378
rect 3596 4326 3608 4378
rect 3670 4326 3672 4378
rect 3510 4324 3534 4326
rect 3590 4324 3614 4326
rect 3670 4324 3694 4326
rect 3454 4304 3750 4324
rect 3988 4298 4016 5034
rect 4080 4622 4108 5120
rect 4160 5102 4212 5108
rect 4264 4865 4292 5850
rect 4356 5846 4384 6258
rect 4344 5840 4396 5846
rect 4344 5782 4396 5788
rect 4250 4856 4306 4865
rect 4250 4791 4306 4800
rect 4252 4684 4304 4690
rect 4252 4626 4304 4632
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 3896 4282 4108 4298
rect 3896 4276 4120 4282
rect 3896 4270 4068 4276
rect 3896 3670 3924 4270
rect 4068 4218 4120 4224
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 3884 3664 3936 3670
rect 3884 3606 3936 3612
rect 3454 3292 3750 3312
rect 3510 3290 3534 3292
rect 3590 3290 3614 3292
rect 3670 3290 3694 3292
rect 3532 3238 3534 3290
rect 3596 3238 3608 3290
rect 3670 3238 3672 3290
rect 3510 3236 3534 3238
rect 3590 3236 3614 3238
rect 3670 3236 3694 3238
rect 3454 3216 3750 3236
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 3792 2916 3844 2922
rect 3792 2858 3844 2864
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 3252 2746 3372 2774
rect 3148 2508 3200 2514
rect 3148 2450 3200 2456
rect 3344 1442 3372 2746
rect 3528 2650 3556 2790
rect 3804 2650 3832 2858
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 3454 2204 3750 2224
rect 3510 2202 3534 2204
rect 3590 2202 3614 2204
rect 3670 2202 3694 2204
rect 3532 2150 3534 2202
rect 3596 2150 3608 2202
rect 3670 2150 3672 2202
rect 3510 2148 3534 2150
rect 3590 2148 3614 2150
rect 3670 2148 3694 2150
rect 3454 2128 3750 2148
rect 3608 1896 3660 1902
rect 3608 1838 3660 1844
rect 3620 1465 3648 1838
rect 3606 1456 3662 1465
rect 3344 1414 3556 1442
rect 3528 800 3556 1414
rect 3606 1391 3662 1400
rect 3988 800 4016 3878
rect 4080 3398 4108 4218
rect 4172 4010 4200 4558
rect 4160 4004 4212 4010
rect 4160 3946 4212 3952
rect 4172 3738 4200 3946
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 4264 3194 4292 4626
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4356 4078 4384 4422
rect 4344 4072 4396 4078
rect 4344 4014 4396 4020
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 4448 2990 4476 7942
rect 4632 7886 4660 8298
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4540 7546 4568 7822
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4724 7342 4752 12406
rect 4804 12378 4856 12384
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4816 11898 4844 12038
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 4908 10470 4936 15370
rect 5552 15366 5580 16662
rect 5644 16250 5672 17002
rect 5828 16250 5856 17002
rect 5953 16892 6249 16912
rect 6009 16890 6033 16892
rect 6089 16890 6113 16892
rect 6169 16890 6193 16892
rect 6031 16838 6033 16890
rect 6095 16838 6107 16890
rect 6169 16838 6171 16890
rect 6009 16836 6033 16838
rect 6089 16836 6113 16838
rect 6169 16836 6193 16838
rect 5953 16816 6249 16836
rect 6644 16720 6696 16726
rect 6644 16662 6696 16668
rect 6656 16522 6684 16662
rect 6644 16516 6696 16522
rect 6644 16458 6696 16464
rect 6368 16448 6420 16454
rect 6368 16390 6420 16396
rect 5632 16244 5684 16250
rect 5632 16186 5684 16192
rect 5816 16244 5868 16250
rect 5816 16186 5868 16192
rect 5724 16040 5776 16046
rect 5724 15982 5776 15988
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 5264 14884 5316 14890
rect 5264 14826 5316 14832
rect 4988 14816 5040 14822
rect 4988 14758 5040 14764
rect 5000 14414 5028 14758
rect 4988 14408 5040 14414
rect 4988 14350 5040 14356
rect 5276 14346 5304 14826
rect 5540 14476 5592 14482
rect 5540 14418 5592 14424
rect 5264 14340 5316 14346
rect 5264 14282 5316 14288
rect 5448 14340 5500 14346
rect 5448 14282 5500 14288
rect 4988 14068 5040 14074
rect 4988 14010 5040 14016
rect 5000 12434 5028 14010
rect 5460 13938 5488 14282
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5552 13802 5580 14418
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5448 13728 5500 13734
rect 5500 13676 5580 13682
rect 5448 13670 5580 13676
rect 5460 13654 5580 13670
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 5000 12406 5120 12434
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4908 8090 4936 10406
rect 5092 9674 5120 12406
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 5184 11762 5212 12038
rect 5172 11756 5224 11762
rect 5172 11698 5224 11704
rect 5276 11626 5304 13330
rect 5552 12918 5580 13654
rect 5540 12912 5592 12918
rect 5540 12854 5592 12860
rect 5644 12730 5672 15846
rect 5736 14890 5764 15982
rect 5816 15904 5868 15910
rect 5816 15846 5868 15852
rect 5828 15745 5856 15846
rect 5953 15804 6249 15824
rect 6009 15802 6033 15804
rect 6089 15802 6113 15804
rect 6169 15802 6193 15804
rect 6031 15750 6033 15802
rect 6095 15750 6107 15802
rect 6169 15750 6171 15802
rect 6009 15748 6033 15750
rect 6089 15748 6113 15750
rect 6169 15748 6193 15750
rect 5814 15736 5870 15745
rect 5953 15728 6249 15748
rect 5814 15671 5870 15680
rect 6092 15564 6144 15570
rect 6092 15506 6144 15512
rect 6276 15564 6328 15570
rect 6380 15552 6408 16390
rect 6460 16244 6512 16250
rect 6460 16186 6512 16192
rect 6472 15570 6500 16186
rect 6656 16114 6684 16458
rect 6748 16182 6776 17002
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 7024 16250 7052 16390
rect 7116 16250 7144 17002
rect 7012 16244 7064 16250
rect 7012 16186 7064 16192
rect 7104 16244 7156 16250
rect 7104 16186 7156 16192
rect 6736 16176 6788 16182
rect 6736 16118 6788 16124
rect 6644 16108 6696 16114
rect 6644 16050 6696 16056
rect 7288 15972 7340 15978
rect 7288 15914 7340 15920
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7208 15706 7236 15846
rect 7300 15706 7328 15914
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7288 15700 7340 15706
rect 7288 15642 7340 15648
rect 6328 15524 6408 15552
rect 6276 15506 6328 15512
rect 6104 15026 6132 15506
rect 6380 15162 6408 15524
rect 6460 15564 6512 15570
rect 6460 15506 6512 15512
rect 6828 15564 6880 15570
rect 6828 15506 6880 15512
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 6368 15156 6420 15162
rect 6368 15098 6420 15104
rect 6276 15088 6328 15094
rect 6276 15030 6328 15036
rect 6092 15020 6144 15026
rect 6092 14962 6144 14968
rect 5724 14884 5776 14890
rect 5724 14826 5776 14832
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 5828 14532 5856 14758
rect 5953 14716 6249 14736
rect 6009 14714 6033 14716
rect 6089 14714 6113 14716
rect 6169 14714 6193 14716
rect 6031 14662 6033 14714
rect 6095 14662 6107 14714
rect 6169 14662 6171 14714
rect 6009 14660 6033 14662
rect 6089 14660 6113 14662
rect 6169 14660 6193 14662
rect 5953 14640 6249 14660
rect 5828 14504 5948 14532
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5736 12986 5764 13806
rect 5920 13802 5948 14504
rect 5908 13796 5960 13802
rect 5908 13738 5960 13744
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5828 13530 5856 13670
rect 5953 13628 6249 13648
rect 6009 13626 6033 13628
rect 6089 13626 6113 13628
rect 6169 13626 6193 13628
rect 6031 13574 6033 13626
rect 6095 13574 6107 13626
rect 6169 13574 6171 13626
rect 6009 13572 6033 13574
rect 6089 13572 6113 13574
rect 6169 13572 6193 13574
rect 5953 13552 6249 13572
rect 5816 13524 5868 13530
rect 5816 13466 5868 13472
rect 5814 13424 5870 13433
rect 5814 13359 5816 13368
rect 5868 13359 5870 13368
rect 5816 13330 5868 13336
rect 6184 13320 6236 13326
rect 6288 13308 6316 15030
rect 6380 14618 6408 15098
rect 6642 14920 6698 14929
rect 6460 14884 6512 14890
rect 6642 14855 6644 14864
rect 6460 14826 6512 14832
rect 6696 14855 6698 14864
rect 6644 14826 6696 14832
rect 6368 14612 6420 14618
rect 6368 14554 6420 14560
rect 6368 14476 6420 14482
rect 6368 14418 6420 14424
rect 6236 13280 6316 13308
rect 6184 13262 6236 13268
rect 5998 13016 6054 13025
rect 5724 12980 5776 12986
rect 5998 12951 6054 12960
rect 5724 12922 5776 12928
rect 6012 12850 6040 12951
rect 6196 12850 6224 13262
rect 6276 12912 6328 12918
rect 6380 12889 6408 14418
rect 6276 12854 6328 12860
rect 6366 12880 6422 12889
rect 6000 12844 6052 12850
rect 6000 12786 6052 12792
rect 6184 12844 6236 12850
rect 6184 12786 6236 12792
rect 5816 12776 5868 12782
rect 5460 12702 5672 12730
rect 5814 12744 5816 12753
rect 5868 12744 5870 12753
rect 5460 12322 5488 12702
rect 5814 12679 5870 12688
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5552 12442 5580 12582
rect 5953 12540 6249 12560
rect 6009 12538 6033 12540
rect 6089 12538 6113 12540
rect 6169 12538 6193 12540
rect 6031 12486 6033 12538
rect 6095 12486 6107 12538
rect 6169 12486 6171 12538
rect 6009 12484 6033 12486
rect 6089 12484 6113 12486
rect 6169 12484 6193 12486
rect 5722 12472 5778 12481
rect 5540 12436 5592 12442
rect 5953 12464 6249 12484
rect 5722 12407 5778 12416
rect 5540 12378 5592 12384
rect 5460 12306 5580 12322
rect 5460 12300 5592 12306
rect 5460 12294 5540 12300
rect 5540 12242 5592 12248
rect 5356 12164 5408 12170
rect 5356 12106 5408 12112
rect 5368 11762 5396 12106
rect 5540 11824 5592 11830
rect 5540 11766 5592 11772
rect 5356 11756 5408 11762
rect 5356 11698 5408 11704
rect 5264 11620 5316 11626
rect 5264 11562 5316 11568
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5460 11354 5488 11494
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5552 11218 5580 11766
rect 5736 11694 5764 12407
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 6196 12084 6224 12242
rect 6288 12238 6316 12854
rect 6366 12815 6422 12824
rect 6380 12782 6408 12815
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 6472 12434 6500 14826
rect 6748 14618 6776 15438
rect 6840 15162 6868 15506
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 7024 15076 7052 15642
rect 7104 15088 7156 15094
rect 7024 15048 7104 15076
rect 7104 15030 7156 15036
rect 7116 14958 7144 15030
rect 7288 15020 7340 15026
rect 7288 14962 7340 14968
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 7104 14952 7156 14958
rect 7104 14894 7156 14900
rect 6840 14822 6868 14894
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 6736 14612 6788 14618
rect 6736 14554 6788 14560
rect 6564 13190 6592 14554
rect 6736 14476 6788 14482
rect 6736 14418 6788 14424
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 6642 14376 6698 14385
rect 6642 14311 6698 14320
rect 6656 13870 6684 14311
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 6656 13530 6684 13806
rect 6644 13524 6696 13530
rect 6644 13466 6696 13472
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 6644 13184 6696 13190
rect 6644 13126 6696 13132
rect 6656 12753 6684 13126
rect 6642 12744 6698 12753
rect 6642 12679 6698 12688
rect 6380 12406 6500 12434
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 6276 12096 6328 12102
rect 5814 12064 5870 12073
rect 6196 12056 6276 12084
rect 6380 12073 6408 12406
rect 6656 12322 6684 12679
rect 6460 12300 6512 12306
rect 6460 12242 6512 12248
rect 6564 12294 6684 12322
rect 6276 12038 6328 12044
rect 6366 12064 6422 12073
rect 5814 11999 5870 12008
rect 5724 11688 5776 11694
rect 5724 11630 5776 11636
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5552 10674 5580 11154
rect 5540 10668 5592 10674
rect 5592 10628 5672 10656
rect 5540 10610 5592 10616
rect 5540 10532 5592 10538
rect 5540 10474 5592 10480
rect 5552 10062 5580 10474
rect 5644 10130 5672 10628
rect 5736 10266 5764 11154
rect 5828 10470 5856 11999
rect 5953 11452 6249 11472
rect 6009 11450 6033 11452
rect 6089 11450 6113 11452
rect 6169 11450 6193 11452
rect 6031 11398 6033 11450
rect 6095 11398 6107 11450
rect 6169 11398 6171 11450
rect 6009 11396 6033 11398
rect 6089 11396 6113 11398
rect 6169 11396 6193 11398
rect 5953 11376 6249 11396
rect 6288 11286 6316 12038
rect 6366 11999 6422 12008
rect 6366 11928 6422 11937
rect 6366 11863 6422 11872
rect 6380 11694 6408 11863
rect 6472 11762 6500 12242
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6368 11688 6420 11694
rect 6368 11630 6420 11636
rect 6276 11280 6328 11286
rect 6276 11222 6328 11228
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 6012 10674 6040 11086
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5953 10364 6249 10384
rect 6009 10362 6033 10364
rect 6089 10362 6113 10364
rect 6169 10362 6193 10364
rect 6031 10310 6033 10362
rect 6095 10310 6107 10362
rect 6169 10310 6171 10362
rect 6009 10308 6033 10310
rect 6089 10308 6113 10310
rect 6169 10308 6193 10310
rect 5953 10288 6249 10308
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5552 9722 5580 9998
rect 5816 9988 5868 9994
rect 5816 9930 5868 9936
rect 5000 9646 5120 9674
rect 5540 9716 5592 9722
rect 5540 9658 5592 9664
rect 5828 9674 5856 9930
rect 5828 9646 6040 9674
rect 5000 9382 5028 9646
rect 6012 9586 6040 9646
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 4988 9376 5040 9382
rect 4986 9344 4988 9353
rect 5040 9344 5042 9353
rect 4986 9279 5042 9288
rect 4896 8084 4948 8090
rect 4896 8026 4948 8032
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4908 6798 4936 7890
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4528 6724 4580 6730
rect 4528 6666 4580 6672
rect 4540 5778 4568 6666
rect 4908 5778 4936 6734
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 5000 5658 5028 9279
rect 5184 8498 5212 9522
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 6276 9512 6328 9518
rect 6276 9454 6328 9460
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 5092 7857 5120 8230
rect 5078 7848 5134 7857
rect 5078 7783 5134 7792
rect 5092 7274 5120 7783
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 5184 7274 5212 7686
rect 5080 7268 5132 7274
rect 5080 7210 5132 7216
rect 5172 7268 5224 7274
rect 5172 7210 5224 7216
rect 5184 6322 5212 7210
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 5276 6866 5304 7142
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5276 6458 5304 6598
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 5172 6316 5224 6322
rect 4528 5636 4580 5642
rect 4528 5578 4580 5584
rect 4908 5630 5028 5658
rect 5092 6276 5172 6304
rect 4540 5166 4568 5578
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 4712 4752 4764 4758
rect 4712 4694 4764 4700
rect 4620 4548 4672 4554
rect 4620 4490 4672 4496
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 4540 3738 4568 4082
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 4540 3602 4568 3674
rect 4528 3596 4580 3602
rect 4528 3538 4580 3544
rect 4540 3058 4568 3538
rect 4528 3052 4580 3058
rect 4528 2994 4580 3000
rect 4344 2984 4396 2990
rect 4344 2926 4396 2932
rect 4436 2984 4488 2990
rect 4436 2926 4488 2932
rect 4356 2650 4384 2926
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 4066 2544 4122 2553
rect 4066 2479 4068 2488
rect 4120 2479 4122 2488
rect 4068 2450 4120 2456
rect 4632 2446 4660 4490
rect 4724 4214 4752 4694
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4816 4282 4844 4626
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 4712 4208 4764 4214
rect 4712 4150 4764 4156
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 4724 2922 4752 3470
rect 4712 2916 4764 2922
rect 4712 2858 4764 2864
rect 4804 2848 4856 2854
rect 4908 2836 4936 5630
rect 5092 4690 5120 6276
rect 5172 6258 5224 6264
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5276 5370 5304 6258
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 5368 5250 5396 9454
rect 5724 9376 5776 9382
rect 5816 9376 5868 9382
rect 5724 9318 5776 9324
rect 5814 9344 5816 9353
rect 5868 9344 5870 9353
rect 5736 8498 5764 9318
rect 5814 9279 5870 9288
rect 5953 9276 6249 9296
rect 6009 9274 6033 9276
rect 6089 9274 6113 9276
rect 6169 9274 6193 9276
rect 6031 9222 6033 9274
rect 6095 9222 6107 9274
rect 6169 9222 6171 9274
rect 6009 9220 6033 9222
rect 6089 9220 6113 9222
rect 6169 9220 6193 9222
rect 5953 9200 6249 9220
rect 6288 8566 6316 9454
rect 6276 8560 6328 8566
rect 6276 8502 6328 8508
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 5276 5222 5396 5250
rect 5460 6882 5488 8026
rect 5552 7546 5580 8230
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5540 7336 5592 7342
rect 5538 7304 5540 7313
rect 5592 7304 5594 7313
rect 5538 7239 5594 7248
rect 5540 6928 5592 6934
rect 5460 6876 5540 6882
rect 5460 6870 5592 6876
rect 5460 6854 5580 6870
rect 5276 4690 5304 5222
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5368 4690 5396 4966
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 4988 4480 5040 4486
rect 4988 4422 5040 4428
rect 5000 4078 5028 4422
rect 4988 4072 5040 4078
rect 4988 4014 5040 4020
rect 4856 2808 4936 2836
rect 5264 2848 5316 2854
rect 4804 2790 4856 2796
rect 5264 2790 5316 2796
rect 4816 2582 4844 2790
rect 5276 2650 5304 2790
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 4804 2576 4856 2582
rect 4804 2518 4856 2524
rect 4620 2440 4672 2446
rect 4066 2408 4122 2417
rect 4620 2382 4672 2388
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 4066 2343 4122 2352
rect 4804 2372 4856 2378
rect 4080 1970 4108 2343
rect 4804 2314 4856 2320
rect 4160 2304 4212 2310
rect 4160 2246 4212 2252
rect 4344 2304 4396 2310
rect 4344 2246 4396 2252
rect 4172 2038 4200 2246
rect 4160 2032 4212 2038
rect 4160 1974 4212 1980
rect 4068 1964 4120 1970
rect 4068 1906 4120 1912
rect 4356 800 4384 2246
rect 4816 800 4844 2314
rect 5000 2106 5028 2382
rect 4988 2100 5040 2106
rect 4988 2042 5040 2048
rect 5368 1902 5396 4626
rect 5460 2825 5488 6854
rect 5644 6730 5672 8298
rect 5953 8188 6249 8208
rect 6009 8186 6033 8188
rect 6089 8186 6113 8188
rect 6169 8186 6193 8188
rect 6031 8134 6033 8186
rect 6095 8134 6107 8186
rect 6169 8134 6171 8186
rect 6009 8132 6033 8134
rect 6089 8132 6113 8134
rect 6169 8132 6193 8134
rect 5953 8112 6249 8132
rect 6184 7948 6236 7954
rect 6184 7890 6236 7896
rect 5816 7744 5868 7750
rect 5816 7686 5868 7692
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5736 6866 5764 7482
rect 5828 7206 5856 7686
rect 6196 7410 6224 7890
rect 6288 7546 6316 8502
rect 6276 7540 6328 7546
rect 6276 7482 6328 7488
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 5816 7200 5868 7206
rect 6196 7188 6224 7346
rect 6196 7160 6316 7188
rect 5816 7142 5868 7148
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5632 6724 5684 6730
rect 5632 6666 5684 6672
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5552 5114 5580 6394
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 5644 5914 5672 6054
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5630 5128 5686 5137
rect 5552 5086 5630 5114
rect 5630 5063 5686 5072
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5552 4554 5580 4966
rect 5644 4690 5672 5063
rect 5736 4758 5764 6802
rect 5828 6458 5856 7142
rect 5953 7100 6249 7120
rect 6009 7098 6033 7100
rect 6089 7098 6113 7100
rect 6169 7098 6193 7100
rect 6031 7046 6033 7098
rect 6095 7046 6107 7098
rect 6169 7046 6171 7098
rect 6009 7044 6033 7046
rect 6089 7044 6113 7046
rect 6169 7044 6193 7046
rect 5953 7024 6249 7044
rect 6288 6798 6316 7160
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 5724 4752 5776 4758
rect 5724 4694 5776 4700
rect 5828 4690 5856 6190
rect 5953 6012 6249 6032
rect 6009 6010 6033 6012
rect 6089 6010 6113 6012
rect 6169 6010 6193 6012
rect 6031 5958 6033 6010
rect 6095 5958 6107 6010
rect 6169 5958 6171 6010
rect 6009 5956 6033 5958
rect 6089 5956 6113 5958
rect 6169 5956 6193 5958
rect 5953 5936 6249 5956
rect 6000 5568 6052 5574
rect 6000 5510 6052 5516
rect 6012 5216 6040 5510
rect 6182 5400 6238 5409
rect 6182 5335 6238 5344
rect 6092 5228 6144 5234
rect 6012 5188 6092 5216
rect 6092 5170 6144 5176
rect 6196 5098 6224 5335
rect 6288 5114 6316 6394
rect 6380 5574 6408 11630
rect 6460 11620 6512 11626
rect 6460 11562 6512 11568
rect 6472 9586 6500 11562
rect 6564 11506 6592 12294
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6656 11626 6684 12174
rect 6644 11620 6696 11626
rect 6644 11562 6696 11568
rect 6564 11478 6684 11506
rect 6656 10538 6684 11478
rect 6644 10532 6696 10538
rect 6644 10474 6696 10480
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6460 9580 6512 9586
rect 6460 9522 6512 9528
rect 6472 9042 6500 9522
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6472 8498 6500 8774
rect 6460 8492 6512 8498
rect 6460 8434 6512 8440
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6368 5568 6420 5574
rect 6368 5510 6420 5516
rect 6184 5092 6236 5098
rect 6288 5086 6408 5114
rect 6472 5098 6500 7142
rect 6564 6322 6592 10406
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6656 5692 6684 10474
rect 6748 9518 6776 14418
rect 6828 13932 6880 13938
rect 6828 13874 6880 13880
rect 6840 13530 6868 13874
rect 7208 13852 7236 14418
rect 7300 14414 7328 14962
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7300 14074 7328 14350
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7208 13824 7328 13852
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6840 12918 6868 13466
rect 6932 13433 6960 13670
rect 7300 13462 7328 13824
rect 7288 13456 7340 13462
rect 6918 13424 6974 13433
rect 6974 13382 7052 13410
rect 7288 13398 7340 13404
rect 6918 13359 6974 13368
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 6828 12708 6880 12714
rect 6828 12650 6880 12656
rect 6840 11218 6868 12650
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6932 11150 6960 11562
rect 7024 11200 7052 13382
rect 7300 12730 7328 13398
rect 7392 13394 7420 17274
rect 7484 16250 7512 17478
rect 7576 17134 7604 19200
rect 7748 17604 7800 17610
rect 7748 17546 7800 17552
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7656 17060 7708 17066
rect 7656 17002 7708 17008
rect 7472 16244 7524 16250
rect 7472 16186 7524 16192
rect 7668 16114 7696 17002
rect 7760 16250 7788 17546
rect 7840 17264 7892 17270
rect 7944 17252 7972 19200
rect 8404 17626 8432 19200
rect 7892 17224 7972 17252
rect 8312 17598 8432 17626
rect 8772 17626 8800 19200
rect 8772 17598 8892 17626
rect 7840 17206 7892 17212
rect 8024 17060 8076 17066
rect 8024 17002 8076 17008
rect 8116 17060 8168 17066
rect 8116 17002 8168 17008
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 8036 16182 8064 17002
rect 8128 16794 8156 17002
rect 8208 16992 8260 16998
rect 8208 16934 8260 16940
rect 8116 16788 8168 16794
rect 8116 16730 8168 16736
rect 8024 16176 8076 16182
rect 8024 16118 8076 16124
rect 7656 16108 7708 16114
rect 7656 16050 7708 16056
rect 7472 16040 7524 16046
rect 7472 15982 7524 15988
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 7484 15706 7512 15982
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7484 14074 7512 15642
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 7760 15162 7788 15438
rect 7852 15366 7880 15982
rect 7932 15972 7984 15978
rect 7932 15914 7984 15920
rect 7944 15434 7972 15914
rect 7932 15428 7984 15434
rect 7932 15370 7984 15376
rect 7840 15360 7892 15366
rect 7840 15302 7892 15308
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 7472 14068 7524 14074
rect 7472 14010 7524 14016
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 7576 13190 7604 14758
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7378 13016 7434 13025
rect 7378 12951 7434 12960
rect 7116 12702 7328 12730
rect 7116 12646 7144 12702
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7116 11354 7144 12038
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 7024 11172 7144 11200
rect 6920 11144 6972 11150
rect 6972 11104 7052 11132
rect 6920 11086 6972 11092
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6932 9926 6960 10950
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6736 9512 6788 9518
rect 6736 9454 6788 9460
rect 6932 9178 6960 9862
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 6736 8900 6788 8906
rect 6736 8842 6788 8848
rect 6748 8430 6776 8842
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6826 7984 6882 7993
rect 6932 7954 6960 8298
rect 6826 7919 6882 7928
rect 6920 7948 6972 7954
rect 6840 7274 6868 7919
rect 6920 7890 6972 7896
rect 6932 7410 6960 7890
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6828 7268 6880 7274
rect 6828 7210 6880 7216
rect 6932 6798 6960 7346
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6736 6724 6788 6730
rect 6736 6666 6788 6672
rect 6748 6633 6776 6666
rect 7024 6662 7052 11104
rect 7116 11014 7144 11172
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7208 10554 7236 12702
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7300 11354 7328 12582
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7116 10526 7236 10554
rect 7116 10146 7144 10526
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 7208 10266 7236 10406
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7116 10118 7236 10146
rect 7208 9722 7236 10118
rect 7300 9994 7328 11018
rect 7288 9988 7340 9994
rect 7288 9930 7340 9936
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 7208 9382 7236 9658
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 7102 8120 7158 8129
rect 7102 8055 7104 8064
rect 7156 8055 7158 8064
rect 7104 8026 7156 8032
rect 7208 8022 7236 8366
rect 7288 8356 7340 8362
rect 7288 8298 7340 8304
rect 7196 8016 7248 8022
rect 7300 7993 7328 8298
rect 7196 7958 7248 7964
rect 7286 7984 7342 7993
rect 7286 7919 7342 7928
rect 7300 7886 7328 7919
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7196 7540 7248 7546
rect 7116 7500 7196 7528
rect 7012 6656 7064 6662
rect 6734 6624 6790 6633
rect 7012 6598 7064 6604
rect 6734 6559 6790 6568
rect 7024 6458 7052 6598
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6840 5846 6868 6054
rect 6828 5840 6880 5846
rect 6828 5782 6880 5788
rect 6736 5704 6788 5710
rect 6656 5664 6736 5692
rect 6736 5646 6788 5652
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6550 5400 6606 5409
rect 6550 5335 6552 5344
rect 6604 5335 6606 5344
rect 6552 5306 6604 5312
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6184 5034 6236 5040
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 5953 4924 6249 4944
rect 6009 4922 6033 4924
rect 6089 4922 6113 4924
rect 6169 4922 6193 4924
rect 6031 4870 6033 4922
rect 6095 4870 6107 4922
rect 6169 4870 6171 4922
rect 6009 4868 6033 4870
rect 6089 4868 6113 4870
rect 6169 4868 6193 4870
rect 5953 4848 6249 4868
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 6288 4570 6316 4966
rect 5540 4548 5592 4554
rect 5540 4490 5592 4496
rect 6196 4542 6316 4570
rect 6196 4078 6224 4542
rect 6276 4480 6328 4486
rect 6276 4422 6328 4428
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5552 3194 5580 3878
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 5446 2816 5502 2825
rect 5446 2751 5502 2760
rect 5552 2514 5580 2858
rect 5644 2650 5672 3946
rect 5953 3836 6249 3856
rect 6009 3834 6033 3836
rect 6089 3834 6113 3836
rect 6169 3834 6193 3836
rect 6031 3782 6033 3834
rect 6095 3782 6107 3834
rect 6169 3782 6171 3834
rect 6009 3780 6033 3782
rect 6089 3780 6113 3782
rect 6169 3780 6193 3782
rect 5953 3760 6249 3780
rect 6288 3670 6316 4422
rect 6276 3664 6328 3670
rect 6276 3606 6328 3612
rect 5816 3596 5868 3602
rect 5816 3538 5868 3544
rect 5908 3596 5960 3602
rect 5908 3538 5960 3544
rect 5828 3126 5856 3538
rect 5816 3120 5868 3126
rect 5816 3062 5868 3068
rect 5920 2990 5948 3538
rect 6276 3460 6328 3466
rect 6380 3448 6408 5086
rect 6460 5092 6512 5098
rect 6460 5034 6512 5040
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6472 3924 6500 4626
rect 6564 4078 6592 5170
rect 6656 4978 6684 5510
rect 6748 5166 6776 5646
rect 6840 5370 6868 5782
rect 6932 5778 6960 6258
rect 7024 6254 7052 6394
rect 7012 6248 7064 6254
rect 7012 6190 7064 6196
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 7012 5636 7064 5642
rect 7012 5578 7064 5584
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 6932 5234 6960 5510
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6920 5092 6972 5098
rect 6920 5034 6972 5040
rect 6656 4950 6776 4978
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6472 3896 6592 3924
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 6328 3420 6408 3448
rect 6276 3402 6328 3408
rect 6000 3392 6052 3398
rect 6000 3334 6052 3340
rect 6012 3058 6040 3334
rect 6368 3120 6420 3126
rect 6274 3088 6330 3097
rect 6000 3052 6052 3058
rect 6368 3062 6420 3068
rect 6274 3023 6330 3032
rect 6000 2994 6052 3000
rect 5908 2984 5960 2990
rect 5908 2926 5960 2932
rect 5814 2816 5870 2825
rect 5814 2751 5870 2760
rect 5828 2650 5856 2751
rect 5953 2748 6249 2768
rect 6009 2746 6033 2748
rect 6089 2746 6113 2748
rect 6169 2746 6193 2748
rect 6031 2694 6033 2746
rect 6095 2694 6107 2746
rect 6169 2694 6171 2746
rect 6009 2692 6033 2694
rect 6089 2692 6113 2694
rect 6169 2692 6193 2694
rect 5953 2672 6249 2692
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 6288 2514 6316 3023
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 6276 2508 6328 2514
rect 6276 2450 6328 2456
rect 6380 2446 6408 3062
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 5632 2372 5684 2378
rect 5632 2314 5684 2320
rect 5356 1896 5408 1902
rect 5356 1838 5408 1844
rect 5172 1420 5224 1426
rect 5172 1362 5224 1368
rect 5184 800 5212 1362
rect 5644 800 5672 2314
rect 6000 1488 6052 1494
rect 6000 1430 6052 1436
rect 6012 800 6040 1430
rect 6472 800 6500 3470
rect 6564 2106 6592 3896
rect 6642 3768 6698 3777
rect 6748 3738 6776 4950
rect 6828 4548 6880 4554
rect 6828 4490 6880 4496
rect 6642 3703 6698 3712
rect 6736 3732 6788 3738
rect 6656 2854 6684 3703
rect 6736 3674 6788 3680
rect 6644 2848 6696 2854
rect 6644 2790 6696 2796
rect 6748 2650 6776 3674
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 6736 2304 6788 2310
rect 6736 2246 6788 2252
rect 6552 2100 6604 2106
rect 6552 2042 6604 2048
rect 6748 1426 6776 2246
rect 6736 1420 6788 1426
rect 6736 1362 6788 1368
rect 6840 800 6868 4490
rect 6932 3602 6960 5034
rect 7024 5030 7052 5578
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 7116 4622 7144 7500
rect 7196 7482 7248 7488
rect 7288 6180 7340 6186
rect 7288 6122 7340 6128
rect 7194 5264 7250 5273
rect 7194 5199 7250 5208
rect 7208 5098 7236 5199
rect 7196 5092 7248 5098
rect 7196 5034 7248 5040
rect 7208 4826 7236 5034
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 7116 4010 7144 4422
rect 7104 4004 7156 4010
rect 7104 3946 7156 3952
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 6932 2292 6960 3538
rect 7208 2650 7236 4626
rect 7300 3602 7328 6122
rect 7392 6118 7420 12951
rect 7576 12714 7604 13126
rect 7852 12986 7880 15302
rect 8220 14618 8248 16934
rect 8312 16794 8340 17598
rect 8452 17436 8748 17456
rect 8508 17434 8532 17436
rect 8588 17434 8612 17436
rect 8668 17434 8692 17436
rect 8530 17382 8532 17434
rect 8594 17382 8606 17434
rect 8668 17382 8670 17434
rect 8508 17380 8532 17382
rect 8588 17380 8612 17382
rect 8668 17380 8692 17382
rect 8452 17360 8748 17380
rect 8864 17134 8892 17598
rect 9140 17202 9168 19200
rect 9220 17264 9272 17270
rect 9220 17206 9272 17212
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 8852 17128 8904 17134
rect 8852 17070 8904 17076
rect 9128 17060 9180 17066
rect 9128 17002 9180 17008
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 8944 16652 8996 16658
rect 8944 16594 8996 16600
rect 8312 16250 8340 16594
rect 8852 16516 8904 16522
rect 8852 16458 8904 16464
rect 8452 16348 8748 16368
rect 8508 16346 8532 16348
rect 8588 16346 8612 16348
rect 8668 16346 8692 16348
rect 8530 16294 8532 16346
rect 8594 16294 8606 16346
rect 8668 16294 8670 16346
rect 8508 16292 8532 16294
rect 8588 16292 8612 16294
rect 8668 16292 8692 16294
rect 8452 16272 8748 16292
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8864 16114 8892 16458
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 8312 15706 8340 15982
rect 8760 15972 8812 15978
rect 8760 15914 8812 15920
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 8772 15570 8800 15914
rect 8956 15586 8984 16594
rect 9140 16590 9168 17002
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8760 15564 8812 15570
rect 8760 15506 8812 15512
rect 8864 15558 8984 15586
rect 8312 15162 8340 15506
rect 8452 15260 8748 15280
rect 8508 15258 8532 15260
rect 8588 15258 8612 15260
rect 8668 15258 8692 15260
rect 8530 15206 8532 15258
rect 8594 15206 8606 15258
rect 8668 15206 8670 15258
rect 8508 15204 8532 15206
rect 8588 15204 8612 15206
rect 8668 15204 8692 15206
rect 8452 15184 8748 15204
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8760 14952 8812 14958
rect 8864 14940 8892 15558
rect 8944 15496 8996 15502
rect 8944 15438 8996 15444
rect 8956 14958 8984 15438
rect 8812 14912 8892 14940
rect 8944 14952 8996 14958
rect 8760 14894 8812 14900
rect 8944 14894 8996 14900
rect 8772 14618 8800 14894
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 8208 14612 8260 14618
rect 8208 14554 8260 14560
rect 8760 14612 8812 14618
rect 8760 14554 8812 14560
rect 8024 14408 8076 14414
rect 8022 14376 8024 14385
rect 8076 14376 8078 14385
rect 8022 14311 8078 14320
rect 8220 13734 8248 14554
rect 8300 14544 8352 14550
rect 8300 14486 8352 14492
rect 8312 13852 8340 14486
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 8452 14172 8748 14192
rect 8508 14170 8532 14172
rect 8588 14170 8612 14172
rect 8668 14170 8692 14172
rect 8530 14118 8532 14170
rect 8594 14118 8606 14170
rect 8668 14118 8670 14170
rect 8508 14116 8532 14118
rect 8588 14116 8612 14118
rect 8668 14116 8692 14118
rect 8452 14096 8748 14116
rect 8864 14074 8892 14350
rect 8852 14068 8904 14074
rect 8852 14010 8904 14016
rect 8392 13864 8444 13870
rect 8312 13824 8392 13852
rect 8392 13806 8444 13812
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 8220 13546 8248 13670
rect 8220 13530 8340 13546
rect 8956 13530 8984 14758
rect 9048 14414 9076 15642
rect 9140 15162 9168 16526
rect 9232 15910 9260 17206
rect 9600 17048 9628 19200
rect 9772 17060 9824 17066
rect 9600 17020 9772 17048
rect 9600 16250 9628 17020
rect 9772 17002 9824 17008
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9588 16244 9640 16250
rect 9588 16186 9640 16192
rect 9772 15972 9824 15978
rect 9772 15914 9824 15920
rect 9220 15904 9272 15910
rect 9220 15846 9272 15852
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9128 15156 9180 15162
rect 9128 15098 9180 15104
rect 9140 14550 9168 15098
rect 9128 14544 9180 14550
rect 9128 14486 9180 14492
rect 9036 14408 9088 14414
rect 9036 14350 9088 14356
rect 9128 14340 9180 14346
rect 9128 14282 9180 14288
rect 9140 13977 9168 14282
rect 9126 13968 9182 13977
rect 9126 13903 9182 13912
rect 9232 13802 9260 15846
rect 9416 15706 9444 15846
rect 9404 15700 9456 15706
rect 9404 15642 9456 15648
rect 9312 15564 9364 15570
rect 9312 15506 9364 15512
rect 9324 15065 9352 15506
rect 9588 15088 9640 15094
rect 9310 15056 9366 15065
rect 9310 14991 9366 15000
rect 9586 15056 9588 15065
rect 9680 15088 9732 15094
rect 9640 15056 9642 15065
rect 9680 15030 9732 15036
rect 9586 14991 9642 15000
rect 9312 14952 9364 14958
rect 9312 14894 9364 14900
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 9220 13796 9272 13802
rect 9220 13738 9272 13744
rect 8220 13524 8352 13530
rect 8220 13518 8300 13524
rect 8300 13466 8352 13472
rect 8944 13524 8996 13530
rect 8944 13466 8996 13472
rect 8208 13456 8260 13462
rect 8206 13424 8208 13433
rect 8260 13424 8262 13433
rect 8206 13359 8262 13368
rect 8452 13084 8748 13104
rect 8508 13082 8532 13084
rect 8588 13082 8612 13084
rect 8668 13082 8692 13084
rect 8530 13030 8532 13082
rect 8594 13030 8606 13082
rect 8668 13030 8670 13082
rect 8508 13028 8532 13030
rect 8588 13028 8612 13030
rect 8668 13028 8692 13030
rect 8452 13008 8748 13028
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7564 12708 7616 12714
rect 7564 12650 7616 12656
rect 7748 12708 7800 12714
rect 7748 12650 7800 12656
rect 7656 12436 7708 12442
rect 7760 12434 7788 12650
rect 7852 12646 7880 12922
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 8956 12442 8984 12718
rect 8944 12436 8996 12442
rect 7760 12406 7972 12434
rect 7656 12378 7708 12384
rect 7668 11354 7696 12378
rect 7748 12368 7800 12374
rect 7748 12310 7800 12316
rect 7760 11558 7788 12310
rect 7944 11694 7972 12406
rect 8944 12378 8996 12384
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 8944 12300 8996 12306
rect 8996 12260 9076 12288
rect 8944 12242 8996 12248
rect 8312 11778 8340 12242
rect 8452 11996 8748 12016
rect 8508 11994 8532 11996
rect 8588 11994 8612 11996
rect 8668 11994 8692 11996
rect 8530 11942 8532 11994
rect 8594 11942 8606 11994
rect 8668 11942 8670 11994
rect 8508 11940 8532 11942
rect 8588 11940 8612 11942
rect 8668 11940 8692 11942
rect 8452 11920 8748 11940
rect 8208 11756 8260 11762
rect 8312 11750 8432 11778
rect 8208 11698 8260 11704
rect 7932 11688 7984 11694
rect 7932 11630 7984 11636
rect 8116 11688 8168 11694
rect 8116 11630 8168 11636
rect 7748 11552 7800 11558
rect 7932 11552 7984 11558
rect 7748 11494 7800 11500
rect 7852 11512 7932 11540
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 7564 9988 7616 9994
rect 7564 9930 7616 9936
rect 7576 9450 7604 9930
rect 7564 9444 7616 9450
rect 7564 9386 7616 9392
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7484 8430 7512 9318
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7576 8090 7604 8774
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7472 8016 7524 8022
rect 7472 7958 7524 7964
rect 7484 7002 7512 7958
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7576 7342 7604 7686
rect 7668 7546 7696 11290
rect 7760 11150 7788 11494
rect 7748 11144 7800 11150
rect 7748 11086 7800 11092
rect 7852 10742 7880 11512
rect 7932 11494 7984 11500
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 7932 11008 7984 11014
rect 7932 10950 7984 10956
rect 7840 10736 7892 10742
rect 7840 10678 7892 10684
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 7760 10470 7788 10610
rect 7944 10606 7972 10950
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 7760 10130 7788 10406
rect 7838 10160 7894 10169
rect 7748 10124 7800 10130
rect 7838 10095 7894 10104
rect 7748 10066 7800 10072
rect 7760 9110 7788 10066
rect 7748 9104 7800 9110
rect 7748 9046 7800 9052
rect 7852 8650 7880 10095
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 7760 8622 7880 8650
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7654 7304 7710 7313
rect 7654 7239 7710 7248
rect 7668 7206 7696 7239
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7484 5914 7512 6734
rect 7760 6186 7788 8622
rect 7944 7886 7972 8910
rect 8036 8430 8064 11154
rect 8128 10169 8156 11630
rect 8220 11082 8248 11698
rect 8404 11558 8432 11750
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 8208 11076 8260 11082
rect 8208 11018 8260 11024
rect 8208 10804 8260 10810
rect 8312 10792 8340 11494
rect 8852 11212 8904 11218
rect 8852 11154 8904 11160
rect 8452 10908 8748 10928
rect 8508 10906 8532 10908
rect 8588 10906 8612 10908
rect 8668 10906 8692 10908
rect 8530 10854 8532 10906
rect 8594 10854 8606 10906
rect 8668 10854 8670 10906
rect 8508 10852 8532 10854
rect 8588 10852 8612 10854
rect 8668 10852 8692 10854
rect 8452 10832 8748 10852
rect 8260 10764 8340 10792
rect 8208 10746 8260 10752
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8404 10266 8432 10406
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8114 10160 8170 10169
rect 8114 10095 8170 10104
rect 8588 10062 8616 10542
rect 8864 10266 8892 11154
rect 8944 11144 8996 11150
rect 8944 11086 8996 11092
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 8956 10062 8984 11086
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 8452 9820 8748 9840
rect 8508 9818 8532 9820
rect 8588 9818 8612 9820
rect 8668 9818 8692 9820
rect 8530 9766 8532 9818
rect 8594 9766 8606 9818
rect 8668 9766 8670 9818
rect 8508 9764 8532 9766
rect 8588 9764 8612 9766
rect 8668 9764 8692 9766
rect 8452 9744 8748 9764
rect 9048 9654 9076 12260
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9140 11014 9168 12174
rect 9232 11558 9260 13738
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 9140 10674 9168 10950
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 9036 9648 9088 9654
rect 9036 9590 9088 9596
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 8024 8424 8076 8430
rect 8024 8366 8076 8372
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 7944 7546 7972 7822
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 7944 6934 7972 7482
rect 7932 6928 7984 6934
rect 7932 6870 7984 6876
rect 8036 6304 8064 8366
rect 8128 8090 8156 8910
rect 8220 8634 8248 8978
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 8116 8084 8168 8090
rect 8116 8026 8168 8032
rect 8312 8022 8340 9590
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 8772 8974 8800 9114
rect 8760 8968 8812 8974
rect 8758 8936 8760 8945
rect 8812 8936 8814 8945
rect 8758 8871 8814 8880
rect 8944 8900 8996 8906
rect 8944 8842 8996 8848
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 8452 8732 8748 8752
rect 8508 8730 8532 8732
rect 8588 8730 8612 8732
rect 8668 8730 8692 8732
rect 8530 8678 8532 8730
rect 8594 8678 8606 8730
rect 8668 8678 8670 8730
rect 8508 8676 8532 8678
rect 8588 8676 8612 8678
rect 8668 8676 8692 8678
rect 8452 8656 8748 8676
rect 8300 8016 8352 8022
rect 8300 7958 8352 7964
rect 8864 7857 8892 8774
rect 8390 7848 8446 7857
rect 8116 7812 8168 7818
rect 8390 7783 8392 7792
rect 8116 7754 8168 7760
rect 8444 7783 8446 7792
rect 8850 7848 8906 7857
rect 8850 7783 8906 7792
rect 8392 7754 8444 7760
rect 8128 7478 8156 7754
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8852 7744 8904 7750
rect 8852 7686 8904 7692
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 8220 7002 8248 7686
rect 8452 7644 8748 7664
rect 8508 7642 8532 7644
rect 8588 7642 8612 7644
rect 8668 7642 8692 7644
rect 8530 7590 8532 7642
rect 8594 7590 8606 7642
rect 8668 7590 8670 7642
rect 8508 7588 8532 7590
rect 8588 7588 8612 7590
rect 8668 7588 8692 7590
rect 8452 7568 8748 7588
rect 8864 7342 8892 7686
rect 8956 7342 8984 8842
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 9048 8022 9076 8774
rect 9036 8016 9088 8022
rect 9036 7958 9088 7964
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 8942 7168 8998 7177
rect 8942 7103 8998 7112
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 7944 6276 8064 6304
rect 7748 6180 7800 6186
rect 7748 6122 7800 6128
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 7472 5772 7524 5778
rect 7472 5714 7524 5720
rect 7484 5098 7512 5714
rect 7472 5092 7524 5098
rect 7472 5034 7524 5040
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7392 4826 7420 4966
rect 7668 4826 7696 6054
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7760 5166 7788 5510
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7760 4282 7788 4966
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7852 4214 7880 5306
rect 7944 4826 7972 6276
rect 8024 6180 8076 6186
rect 8024 6122 8076 6128
rect 8036 5710 8064 6122
rect 8128 5778 8156 6394
rect 8220 6186 8248 6938
rect 8452 6556 8748 6576
rect 8508 6554 8532 6556
rect 8588 6554 8612 6556
rect 8668 6554 8692 6556
rect 8530 6502 8532 6554
rect 8594 6502 8606 6554
rect 8668 6502 8670 6554
rect 8508 6500 8532 6502
rect 8588 6500 8612 6502
rect 8668 6500 8692 6502
rect 8452 6480 8748 6500
rect 8208 6180 8260 6186
rect 8208 6122 8260 6128
rect 8956 5778 8984 7103
rect 9048 7002 9076 7346
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 9140 6458 9168 10406
rect 9232 10130 9260 10542
rect 9220 10124 9272 10130
rect 9220 10066 9272 10072
rect 9324 9722 9352 14894
rect 9600 14822 9628 14894
rect 9496 14816 9548 14822
rect 9496 14758 9548 14764
rect 9588 14816 9640 14822
rect 9588 14758 9640 14764
rect 9508 14634 9536 14758
rect 9416 14618 9536 14634
rect 9404 14612 9536 14618
rect 9456 14606 9536 14612
rect 9404 14554 9456 14560
rect 9404 13728 9456 13734
rect 9404 13670 9456 13676
rect 9416 13530 9444 13670
rect 9404 13524 9456 13530
rect 9404 13466 9456 13472
rect 9312 9716 9364 9722
rect 9312 9658 9364 9664
rect 9220 8900 9272 8906
rect 9220 8842 9272 8848
rect 9232 8498 9260 8842
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9232 7993 9260 8434
rect 9218 7984 9274 7993
rect 9218 7919 9220 7928
rect 9272 7919 9274 7928
rect 9220 7890 9272 7896
rect 9232 7859 9260 7890
rect 9324 7886 9352 9658
rect 9416 9042 9444 13466
rect 9508 9450 9536 14606
rect 9692 14550 9720 15030
rect 9784 14958 9812 15914
rect 9876 15570 9904 16934
rect 9968 16658 9996 19200
rect 10428 16810 10456 19200
rect 10508 17128 10560 17134
rect 10508 17070 10560 17076
rect 10796 17082 10824 19200
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 11072 17105 11100 17138
rect 11058 17096 11114 17105
rect 10336 16782 10456 16810
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 10048 16448 10100 16454
rect 10048 16390 10100 16396
rect 9956 15972 10008 15978
rect 9956 15914 10008 15920
rect 9968 15706 9996 15914
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9864 15564 9916 15570
rect 9864 15506 9916 15512
rect 9862 15328 9918 15337
rect 9862 15263 9918 15272
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 9680 14544 9732 14550
rect 9680 14486 9732 14492
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 9600 13530 9628 14282
rect 9588 13524 9640 13530
rect 9588 13466 9640 13472
rect 9784 13410 9812 14894
rect 9876 14618 9904 15263
rect 9954 14920 10010 14929
rect 9954 14855 10010 14864
rect 9968 14618 9996 14855
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9876 14006 9904 14350
rect 9864 14000 9916 14006
rect 9864 13942 9916 13948
rect 9692 13382 9812 13410
rect 9692 11898 9720 13382
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9784 12986 9812 13262
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 10060 12374 10088 16390
rect 10336 16250 10364 16782
rect 10416 16652 10468 16658
rect 10416 16594 10468 16600
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 10140 15360 10192 15366
rect 10140 15302 10192 15308
rect 10152 15201 10180 15302
rect 10138 15192 10194 15201
rect 10138 15127 10194 15136
rect 10244 14958 10272 16050
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 10336 15706 10364 15846
rect 10324 15700 10376 15706
rect 10324 15642 10376 15648
rect 10232 14952 10284 14958
rect 10232 14894 10284 14900
rect 10140 14884 10192 14890
rect 10140 14826 10192 14832
rect 10152 14385 10180 14826
rect 10428 14618 10456 16594
rect 10520 16454 10548 17070
rect 10796 17054 10916 17082
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10508 16448 10560 16454
rect 10508 16390 10560 16396
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10520 15502 10548 16390
rect 10704 15706 10732 16390
rect 10796 16114 10824 16934
rect 10888 16250 10916 17054
rect 11058 17031 11114 17040
rect 11256 16980 11284 19200
rect 11520 16992 11572 16998
rect 11256 16952 11468 16980
rect 10950 16892 11246 16912
rect 11006 16890 11030 16892
rect 11086 16890 11110 16892
rect 11166 16890 11190 16892
rect 11028 16838 11030 16890
rect 11092 16838 11104 16890
rect 11166 16838 11168 16890
rect 11006 16836 11030 16838
rect 11086 16836 11110 16838
rect 11166 16836 11190 16838
rect 10950 16816 11246 16836
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 11152 16448 11204 16454
rect 11152 16390 11204 16396
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 10600 15428 10652 15434
rect 10600 15370 10652 15376
rect 10506 15192 10562 15201
rect 10506 15127 10562 15136
rect 10232 14612 10284 14618
rect 10232 14554 10284 14560
rect 10416 14612 10468 14618
rect 10416 14554 10468 14560
rect 10138 14376 10194 14385
rect 10138 14311 10194 14320
rect 10244 14090 10272 14554
rect 10244 14062 10364 14090
rect 10230 13832 10286 13841
rect 10230 13767 10286 13776
rect 10244 13190 10272 13767
rect 10232 13184 10284 13190
rect 10232 13126 10284 13132
rect 10232 12912 10284 12918
rect 10230 12880 10232 12889
rect 10284 12880 10286 12889
rect 10230 12815 10286 12824
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 10048 12368 10100 12374
rect 10048 12310 10100 12316
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9692 11801 9720 11834
rect 9678 11792 9734 11801
rect 9678 11727 9734 11736
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9600 11218 9628 11494
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9692 10810 9720 11086
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 9508 9178 9536 9386
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 9218 7712 9274 7721
rect 9218 7647 9274 7656
rect 9232 7313 9260 7647
rect 9218 7304 9274 7313
rect 9218 7239 9274 7248
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 9034 6352 9090 6361
rect 9034 6287 9090 6296
rect 9048 6118 9076 6287
rect 9036 6112 9088 6118
rect 9036 6054 9088 6060
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 8944 5772 8996 5778
rect 8944 5714 8996 5720
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 8036 5302 8064 5646
rect 8852 5636 8904 5642
rect 8852 5578 8904 5584
rect 8452 5468 8748 5488
rect 8508 5466 8532 5468
rect 8588 5466 8612 5468
rect 8668 5466 8692 5468
rect 8530 5414 8532 5466
rect 8594 5414 8606 5466
rect 8668 5414 8670 5466
rect 8508 5412 8532 5414
rect 8588 5412 8612 5414
rect 8668 5412 8692 5414
rect 8452 5392 8748 5412
rect 8864 5352 8892 5578
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 8956 5370 8984 5510
rect 8680 5324 8892 5352
rect 8944 5364 8996 5370
rect 8024 5296 8076 5302
rect 8024 5238 8076 5244
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 8036 4622 8064 5238
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 8576 5024 8628 5030
rect 8576 4966 8628 4972
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 8036 4282 8064 4558
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 7840 4208 7892 4214
rect 7892 4168 7972 4196
rect 8128 4185 8156 4966
rect 8588 4729 8616 4966
rect 8574 4720 8630 4729
rect 8574 4655 8576 4664
rect 8628 4655 8630 4664
rect 8576 4626 8628 4632
rect 8680 4622 8708 5324
rect 8944 5306 8996 5312
rect 8852 5092 8904 5098
rect 8852 5034 8904 5040
rect 8864 4622 8892 5034
rect 8668 4616 8720 4622
rect 8666 4584 8668 4593
rect 8852 4616 8904 4622
rect 8720 4584 8722 4593
rect 8300 4548 8352 4554
rect 8904 4576 8984 4604
rect 8852 4558 8904 4564
rect 8666 4519 8722 4528
rect 8300 4490 8352 4496
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 7840 4150 7892 4156
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7300 2582 7328 3334
rect 7576 2774 7604 4014
rect 7944 3942 7972 4168
rect 8114 4176 8170 4185
rect 8220 4146 8248 4422
rect 8114 4111 8170 4120
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 7392 2746 7604 2774
rect 7668 2774 7696 3878
rect 7852 3398 7880 3878
rect 8312 3720 8340 4490
rect 8452 4380 8748 4400
rect 8508 4378 8532 4380
rect 8588 4378 8612 4380
rect 8668 4378 8692 4380
rect 8530 4326 8532 4378
rect 8594 4326 8606 4378
rect 8668 4326 8670 4378
rect 8508 4324 8532 4326
rect 8588 4324 8612 4326
rect 8668 4324 8692 4326
rect 8452 4304 8748 4324
rect 8852 4072 8904 4078
rect 8852 4014 8904 4020
rect 8128 3692 8340 3720
rect 7840 3392 7892 3398
rect 7840 3334 7892 3340
rect 7852 2990 7880 3334
rect 7840 2984 7892 2990
rect 7840 2926 7892 2932
rect 7668 2746 7788 2774
rect 7288 2576 7340 2582
rect 7288 2518 7340 2524
rect 7104 2304 7156 2310
rect 6932 2264 7104 2292
rect 7104 2246 7156 2252
rect 7392 1034 7420 2746
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 7668 1494 7696 2382
rect 7656 1488 7708 1494
rect 7656 1430 7708 1436
rect 7300 1006 7420 1034
rect 7300 800 7328 1006
rect 7760 800 7788 2746
rect 8128 800 8156 3692
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8312 3194 8340 3538
rect 8452 3292 8748 3312
rect 8508 3290 8532 3292
rect 8588 3290 8612 3292
rect 8668 3290 8692 3292
rect 8530 3238 8532 3290
rect 8594 3238 8606 3290
rect 8668 3238 8670 3290
rect 8508 3236 8532 3238
rect 8588 3236 8612 3238
rect 8668 3236 8692 3238
rect 8452 3216 8748 3236
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8312 2446 8340 3130
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 8496 2582 8524 2926
rect 8484 2576 8536 2582
rect 8484 2518 8536 2524
rect 8864 2514 8892 4014
rect 8956 3738 8984 4576
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 8956 3097 8984 3470
rect 8942 3088 8998 3097
rect 8942 3023 8998 3032
rect 9048 2922 9076 6054
rect 9140 3602 9168 6394
rect 9232 5642 9260 7239
rect 9416 6474 9444 8978
rect 9692 8294 9720 9454
rect 9784 9178 9812 11630
rect 10060 11354 10088 12310
rect 10152 11830 10180 12582
rect 10244 11898 10272 12582
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 10140 11824 10192 11830
rect 10140 11766 10192 11772
rect 10230 11792 10286 11801
rect 10336 11778 10364 14062
rect 10416 13796 10468 13802
rect 10416 13738 10468 13744
rect 10428 13530 10456 13738
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 10428 13326 10456 13466
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10520 13161 10548 15127
rect 10612 14929 10640 15370
rect 10598 14920 10654 14929
rect 10598 14855 10654 14864
rect 10600 14476 10652 14482
rect 10600 14418 10652 14424
rect 10612 14074 10640 14418
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 10600 13388 10652 13394
rect 10600 13330 10652 13336
rect 10506 13152 10562 13161
rect 10506 13087 10562 13096
rect 10612 12646 10640 13330
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10612 12442 10640 12582
rect 10416 12436 10468 12442
rect 10416 12378 10468 12384
rect 10600 12436 10652 12442
rect 10704 12434 10732 15642
rect 10784 15564 10836 15570
rect 10784 15506 10836 15512
rect 10796 14414 10824 15506
rect 10888 15162 10916 16186
rect 11072 16114 11100 16390
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 11164 16046 11192 16390
rect 11152 16040 11204 16046
rect 11152 15982 11204 15988
rect 11336 15904 11388 15910
rect 11336 15846 11388 15852
rect 10950 15804 11246 15824
rect 11006 15802 11030 15804
rect 11086 15802 11110 15804
rect 11166 15802 11190 15804
rect 11028 15750 11030 15802
rect 11092 15750 11104 15802
rect 11166 15750 11168 15802
rect 11006 15748 11030 15750
rect 11086 15748 11110 15750
rect 11166 15748 11190 15750
rect 10950 15728 11246 15748
rect 11348 15638 11376 15846
rect 11336 15632 11388 15638
rect 11336 15574 11388 15580
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 11440 14958 11468 16952
rect 11520 16934 11572 16940
rect 11532 15858 11560 16934
rect 11624 15978 11652 19200
rect 11796 17060 11848 17066
rect 11796 17002 11848 17008
rect 11980 17060 12032 17066
rect 11980 17002 12032 17008
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11716 16182 11744 16594
rect 11704 16176 11756 16182
rect 11704 16118 11756 16124
rect 11704 16040 11756 16046
rect 11808 15994 11836 17002
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11756 15988 11836 15994
rect 11704 15982 11836 15988
rect 11612 15972 11664 15978
rect 11716 15966 11836 15982
rect 11612 15914 11664 15920
rect 11704 15904 11756 15910
rect 11532 15830 11652 15858
rect 11704 15846 11756 15852
rect 11518 15736 11574 15745
rect 11518 15671 11574 15680
rect 11532 15337 11560 15671
rect 11518 15328 11574 15337
rect 11518 15263 11574 15272
rect 11428 14952 11480 14958
rect 11428 14894 11480 14900
rect 10950 14716 11246 14736
rect 11006 14714 11030 14716
rect 11086 14714 11110 14716
rect 11166 14714 11190 14716
rect 11028 14662 11030 14714
rect 11092 14662 11104 14714
rect 11166 14662 11168 14714
rect 11006 14660 11030 14662
rect 11086 14660 11110 14662
rect 11166 14660 11190 14662
rect 10950 14640 11246 14660
rect 10876 14476 10928 14482
rect 10928 14436 11376 14464
rect 10876 14418 10928 14424
rect 10784 14408 10836 14414
rect 10836 14356 10916 14362
rect 10784 14350 10916 14356
rect 10796 14334 10916 14350
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10796 13530 10824 14214
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 10704 12406 10824 12434
rect 10600 12378 10652 12384
rect 10428 12238 10456 12378
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10796 12102 10824 12406
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10336 11750 10732 11778
rect 10230 11727 10232 11736
rect 10284 11727 10286 11736
rect 10232 11698 10284 11704
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 10060 10470 10088 11154
rect 10140 11076 10192 11082
rect 10140 11018 10192 11024
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 9876 10266 9904 10406
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9968 9654 9996 10066
rect 9956 9648 10008 9654
rect 9956 9590 10008 9596
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9968 8838 9996 9318
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9864 8560 9916 8566
rect 9864 8502 9916 8508
rect 9956 8560 10008 8566
rect 9956 8502 10008 8508
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9496 8288 9548 8294
rect 9496 8230 9548 8236
rect 9680 8288 9732 8294
rect 9680 8230 9732 8236
rect 9508 8090 9536 8230
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9600 7177 9628 7822
rect 9692 7410 9720 8230
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9586 7168 9642 7177
rect 9586 7103 9642 7112
rect 9692 6866 9720 7346
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9408 6446 9444 6474
rect 9408 6390 9436 6446
rect 9404 6384 9456 6390
rect 9588 6384 9640 6390
rect 9404 6326 9456 6332
rect 9586 6352 9588 6361
rect 9640 6352 9642 6361
rect 9586 6287 9642 6296
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 9324 5846 9352 6054
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 9312 5840 9364 5846
rect 9312 5782 9364 5788
rect 9220 5636 9272 5642
rect 9220 5578 9272 5584
rect 9404 5636 9456 5642
rect 9404 5578 9456 5584
rect 9312 5568 9364 5574
rect 9218 5536 9274 5545
rect 9274 5516 9312 5522
rect 9274 5510 9364 5516
rect 9274 5494 9352 5510
rect 9218 5471 9274 5480
rect 9232 5030 9260 5471
rect 9416 5137 9444 5578
rect 9600 5574 9628 5850
rect 9588 5568 9640 5574
rect 9692 5545 9720 6258
rect 9784 6118 9812 8366
rect 9876 7818 9904 8502
rect 9864 7812 9916 7818
rect 9864 7754 9916 7760
rect 9968 7750 9996 8502
rect 9956 7744 10008 7750
rect 9956 7686 10008 7692
rect 10060 7546 10088 10406
rect 10152 9178 10180 11018
rect 10244 10674 10272 11698
rect 10704 11626 10732 11750
rect 10508 11620 10560 11626
rect 10508 11562 10560 11568
rect 10692 11620 10744 11626
rect 10692 11562 10744 11568
rect 10520 11354 10548 11562
rect 10508 11348 10560 11354
rect 10508 11290 10560 11296
rect 10324 11076 10376 11082
rect 10324 11018 10376 11024
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10244 8480 10272 10610
rect 10336 9382 10364 11018
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 10520 10198 10548 10610
rect 10508 10192 10560 10198
rect 10508 10134 10560 10140
rect 10416 9988 10468 9994
rect 10416 9930 10468 9936
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10152 8452 10272 8480
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 9876 6254 9904 7482
rect 10048 7200 10100 7206
rect 10048 7142 10100 7148
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9772 6112 9824 6118
rect 9824 6072 9996 6100
rect 9772 6054 9824 6060
rect 9770 5944 9826 5953
rect 9770 5879 9826 5888
rect 9864 5908 9916 5914
rect 9784 5778 9812 5879
rect 9864 5850 9916 5856
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9772 5568 9824 5574
rect 9588 5510 9640 5516
rect 9678 5536 9734 5545
rect 9600 5273 9628 5510
rect 9772 5510 9824 5516
rect 9678 5471 9734 5480
rect 9586 5264 9642 5273
rect 9692 5234 9720 5471
rect 9784 5409 9812 5510
rect 9770 5400 9826 5409
rect 9770 5335 9826 5344
rect 9770 5264 9826 5273
rect 9586 5199 9642 5208
rect 9680 5228 9732 5234
rect 9770 5199 9826 5208
rect 9680 5170 9732 5176
rect 9402 5128 9458 5137
rect 9402 5063 9458 5072
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9324 4758 9352 4966
rect 9312 4752 9364 4758
rect 9312 4694 9364 4700
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 9232 3466 9260 4626
rect 9310 4584 9366 4593
rect 9692 4570 9720 5170
rect 9784 5166 9812 5199
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9692 4542 9812 4570
rect 9310 4519 9366 4528
rect 9220 3460 9272 3466
rect 9220 3402 9272 3408
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 9140 2990 9168 3334
rect 9128 2984 9180 2990
rect 9128 2926 9180 2932
rect 9218 2952 9274 2961
rect 9036 2916 9088 2922
rect 9218 2887 9274 2896
rect 9036 2858 9088 2864
rect 9232 2650 9260 2887
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 8852 2508 8904 2514
rect 9036 2508 9088 2514
rect 8852 2450 8904 2456
rect 8956 2468 9036 2496
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 8452 2204 8748 2224
rect 8508 2202 8532 2204
rect 8588 2202 8612 2204
rect 8668 2202 8692 2204
rect 8530 2150 8532 2202
rect 8594 2150 8606 2202
rect 8668 2150 8670 2202
rect 8508 2148 8532 2150
rect 8588 2148 8612 2150
rect 8668 2148 8692 2150
rect 8452 2128 8748 2148
rect 8864 1850 8892 2450
rect 8588 1822 8892 1850
rect 8588 800 8616 1822
rect 8956 800 8984 2468
rect 9036 2450 9088 2456
rect 9324 2310 9352 4519
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9692 4146 9720 4422
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 9404 4072 9456 4078
rect 9784 4026 9812 4542
rect 9404 4014 9456 4020
rect 9416 3777 9444 4014
rect 9692 3998 9812 4026
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9402 3768 9458 3777
rect 9402 3703 9458 3712
rect 9496 3664 9548 3670
rect 9496 3606 9548 3612
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9416 2582 9444 3334
rect 9404 2576 9456 2582
rect 9404 2518 9456 2524
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 9508 1034 9536 3606
rect 9600 3398 9628 3878
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9692 3194 9720 3998
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9784 3738 9812 3878
rect 9876 3738 9904 5850
rect 9968 5302 9996 6072
rect 10060 5930 10088 7142
rect 10152 6458 10180 8452
rect 10232 8356 10284 8362
rect 10232 8298 10284 8304
rect 10244 7886 10272 8298
rect 10336 8129 10364 9318
rect 10428 9178 10456 9930
rect 10520 9586 10548 10134
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10704 9382 10732 11562
rect 10796 11558 10824 12038
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10796 11082 10824 11494
rect 10784 11076 10836 11082
rect 10784 11018 10836 11024
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10796 10470 10824 10746
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10796 9654 10824 10406
rect 10784 9648 10836 9654
rect 10784 9590 10836 9596
rect 10784 9444 10836 9450
rect 10784 9386 10836 9392
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10612 8430 10640 8910
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10322 8120 10378 8129
rect 10322 8055 10378 8064
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 10600 7948 10652 7954
rect 10600 7890 10652 7896
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 10244 6798 10272 7822
rect 10336 7546 10364 7890
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10428 7002 10456 7822
rect 10508 7268 10560 7274
rect 10508 7210 10560 7216
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10520 6730 10548 7210
rect 10508 6724 10560 6730
rect 10508 6666 10560 6672
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10152 6118 10180 6394
rect 10520 6322 10548 6666
rect 10612 6458 10640 7890
rect 10704 6934 10732 9318
rect 10796 9110 10824 9386
rect 10784 9104 10836 9110
rect 10784 9046 10836 9052
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 10692 6928 10744 6934
rect 10690 6896 10692 6905
rect 10744 6896 10746 6905
rect 10690 6831 10746 6840
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 10140 6112 10192 6118
rect 10138 6080 10140 6089
rect 10192 6080 10194 6089
rect 10138 6015 10194 6024
rect 10336 5930 10364 6190
rect 10506 6080 10562 6089
rect 10506 6015 10562 6024
rect 10060 5902 10272 5930
rect 10336 5902 10456 5930
rect 9956 5296 10008 5302
rect 9956 5238 10008 5244
rect 10060 4826 10088 5902
rect 10244 5828 10272 5902
rect 10324 5840 10376 5846
rect 10244 5800 10324 5828
rect 10324 5782 10376 5788
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10140 5636 10192 5642
rect 10140 5578 10192 5584
rect 10232 5636 10284 5642
rect 10232 5578 10284 5584
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 10060 4282 10088 4762
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 10152 3942 10180 5578
rect 10244 5302 10272 5578
rect 10232 5296 10284 5302
rect 10232 5238 10284 5244
rect 10336 4486 10364 5646
rect 10428 5030 10456 5902
rect 10520 5166 10548 6015
rect 10612 5930 10640 6190
rect 10704 6118 10732 6734
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10612 5902 10732 5930
rect 10600 5568 10652 5574
rect 10600 5510 10652 5516
rect 10508 5160 10560 5166
rect 10508 5102 10560 5108
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 10506 4992 10562 5001
rect 10506 4927 10562 4936
rect 10324 4480 10376 4486
rect 10324 4422 10376 4428
rect 10336 4214 10364 4422
rect 10324 4208 10376 4214
rect 10324 4150 10376 4156
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 10336 3534 10364 4150
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 9784 3233 9812 3470
rect 9770 3224 9826 3233
rect 9680 3188 9732 3194
rect 9770 3159 9826 3168
rect 9680 3130 9732 3136
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 9416 1006 9536 1034
rect 9416 800 9444 1006
rect 9784 800 9812 2926
rect 9968 2854 9996 3470
rect 10428 3369 10456 4014
rect 10520 3942 10548 4927
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10612 3670 10640 5510
rect 10704 5001 10732 5902
rect 10690 4992 10746 5001
rect 10690 4927 10746 4936
rect 10796 4842 10824 7482
rect 10888 6118 10916 14334
rect 10950 13628 11246 13648
rect 11006 13626 11030 13628
rect 11086 13626 11110 13628
rect 11166 13626 11190 13628
rect 11028 13574 11030 13626
rect 11092 13574 11104 13626
rect 11166 13574 11168 13626
rect 11006 13572 11030 13574
rect 11086 13572 11110 13574
rect 11166 13572 11190 13574
rect 10950 13552 11246 13572
rect 11348 12714 11376 14436
rect 11440 14006 11468 14894
rect 11624 14822 11652 15830
rect 11716 15706 11744 15846
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11716 15162 11744 15438
rect 11808 15366 11836 15966
rect 11796 15360 11848 15366
rect 11796 15302 11848 15308
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 11612 14816 11664 14822
rect 11612 14758 11664 14764
rect 11716 14550 11744 15098
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 11704 14544 11756 14550
rect 11704 14486 11756 14492
rect 11520 14476 11572 14482
rect 11520 14418 11572 14424
rect 11428 14000 11480 14006
rect 11428 13942 11480 13948
rect 11532 13870 11560 14418
rect 11520 13864 11572 13870
rect 11808 13841 11836 14758
rect 11520 13806 11572 13812
rect 11794 13832 11850 13841
rect 11794 13767 11850 13776
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11808 13569 11836 13670
rect 11794 13560 11850 13569
rect 11440 13518 11744 13546
rect 11440 13462 11468 13518
rect 11428 13456 11480 13462
rect 11428 13398 11480 13404
rect 11520 13456 11572 13462
rect 11520 13398 11572 13404
rect 11532 12918 11560 13398
rect 11716 12986 11744 13518
rect 11900 13530 11928 16730
rect 11992 16250 12020 17002
rect 12084 16454 12112 19200
rect 12164 17264 12216 17270
rect 12164 17206 12216 17212
rect 12176 16726 12204 17206
rect 12256 17128 12308 17134
rect 12308 17076 12388 17082
rect 12256 17070 12388 17076
rect 12268 17054 12388 17070
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 12164 16720 12216 16726
rect 12164 16662 12216 16668
rect 12072 16448 12124 16454
rect 12072 16390 12124 16396
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 11992 15094 12020 16186
rect 12072 15904 12124 15910
rect 12072 15846 12124 15852
rect 11980 15088 12032 15094
rect 11980 15030 12032 15036
rect 11980 14816 12032 14822
rect 11980 14758 12032 14764
rect 11794 13495 11850 13504
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11520 12912 11572 12918
rect 11520 12854 11572 12860
rect 11428 12776 11480 12782
rect 11428 12718 11480 12724
rect 11520 12776 11572 12782
rect 11520 12718 11572 12724
rect 11612 12776 11664 12782
rect 11612 12718 11664 12724
rect 11702 12744 11758 12753
rect 11336 12708 11388 12714
rect 11336 12650 11388 12656
rect 10950 12540 11246 12560
rect 11006 12538 11030 12540
rect 11086 12538 11110 12540
rect 11166 12538 11190 12540
rect 11028 12486 11030 12538
rect 11092 12486 11104 12538
rect 11166 12486 11168 12538
rect 11006 12484 11030 12486
rect 11086 12484 11110 12486
rect 11166 12484 11190 12486
rect 10950 12464 11246 12484
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 11072 11694 11100 12038
rect 11256 11830 11284 12174
rect 11244 11824 11296 11830
rect 11244 11766 11296 11772
rect 11060 11688 11112 11694
rect 11348 11676 11376 12650
rect 11440 12102 11468 12718
rect 11532 12306 11560 12718
rect 11624 12442 11652 12718
rect 11702 12679 11758 12688
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11428 12096 11480 12102
rect 11428 12038 11480 12044
rect 11532 11762 11560 12242
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 11428 11688 11480 11694
rect 11348 11648 11428 11676
rect 11060 11630 11112 11636
rect 11428 11630 11480 11636
rect 10950 11452 11246 11472
rect 11006 11450 11030 11452
rect 11086 11450 11110 11452
rect 11166 11450 11190 11452
rect 11028 11398 11030 11450
rect 11092 11398 11104 11450
rect 11166 11398 11168 11450
rect 11006 11396 11030 11398
rect 11086 11396 11110 11398
rect 11166 11396 11190 11398
rect 10950 11376 11246 11396
rect 11058 11248 11114 11257
rect 11058 11183 11114 11192
rect 11520 11212 11572 11218
rect 11072 10606 11100 11183
rect 11520 11154 11572 11160
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 11428 10532 11480 10538
rect 11428 10474 11480 10480
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 10950 10364 11246 10384
rect 11006 10362 11030 10364
rect 11086 10362 11110 10364
rect 11166 10362 11190 10364
rect 11028 10310 11030 10362
rect 11092 10310 11104 10362
rect 11166 10310 11168 10362
rect 11006 10308 11030 10310
rect 11086 10308 11110 10310
rect 11166 10308 11190 10310
rect 10950 10288 11246 10308
rect 11348 10266 11376 10406
rect 11440 10266 11468 10474
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 11428 10260 11480 10266
rect 11428 10202 11480 10208
rect 10950 9276 11246 9296
rect 11006 9274 11030 9276
rect 11086 9274 11110 9276
rect 11166 9274 11190 9276
rect 11028 9222 11030 9274
rect 11092 9222 11104 9274
rect 11166 9222 11168 9274
rect 11006 9220 11030 9222
rect 11086 9220 11110 9222
rect 11166 9220 11190 9222
rect 10950 9200 11246 9220
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 11348 8634 11376 8978
rect 11428 8832 11480 8838
rect 11428 8774 11480 8780
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 10950 8188 11246 8208
rect 11006 8186 11030 8188
rect 11086 8186 11110 8188
rect 11166 8186 11190 8188
rect 11028 8134 11030 8186
rect 11092 8134 11104 8186
rect 11166 8134 11168 8186
rect 11006 8132 11030 8134
rect 11086 8132 11110 8134
rect 11166 8132 11190 8134
rect 10950 8112 11246 8132
rect 11348 7886 11376 8570
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 11348 7206 11376 7346
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 10950 7100 11246 7120
rect 11006 7098 11030 7100
rect 11086 7098 11110 7100
rect 11166 7098 11190 7100
rect 11028 7046 11030 7098
rect 11092 7046 11104 7098
rect 11166 7046 11168 7098
rect 11006 7044 11030 7046
rect 11086 7044 11110 7046
rect 11166 7044 11190 7046
rect 10950 7024 11246 7044
rect 11348 7002 11376 7142
rect 11336 6996 11388 7002
rect 11336 6938 11388 6944
rect 11348 6798 11376 6938
rect 11336 6792 11388 6798
rect 11242 6760 11298 6769
rect 11336 6734 11388 6740
rect 11440 6746 11468 8774
rect 11532 7546 11560 11154
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 11624 10198 11652 10950
rect 11612 10192 11664 10198
rect 11612 10134 11664 10140
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11624 7993 11652 9318
rect 11610 7984 11666 7993
rect 11610 7919 11666 7928
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 11624 7342 11652 7919
rect 11612 7336 11664 7342
rect 11612 7278 11664 7284
rect 11242 6695 11298 6704
rect 11256 6662 11284 6695
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11348 6322 11376 6734
rect 11440 6718 11560 6746
rect 11428 6656 11480 6662
rect 11426 6624 11428 6633
rect 11480 6624 11482 6633
rect 11426 6559 11482 6568
rect 11336 6316 11388 6322
rect 11336 6258 11388 6264
rect 11440 6202 11468 6559
rect 11348 6174 11468 6202
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10888 5896 10916 6054
rect 10950 6012 11246 6032
rect 11006 6010 11030 6012
rect 11086 6010 11110 6012
rect 11166 6010 11190 6012
rect 11028 5958 11030 6010
rect 11092 5958 11104 6010
rect 11166 5958 11168 6010
rect 11006 5956 11030 5958
rect 11086 5956 11110 5958
rect 11166 5956 11190 5958
rect 10950 5936 11246 5956
rect 10888 5868 11008 5896
rect 10980 5574 11008 5868
rect 11348 5574 11376 6174
rect 11532 5760 11560 6718
rect 11624 6458 11652 7278
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11624 6254 11652 6394
rect 11612 6248 11664 6254
rect 11612 6190 11664 6196
rect 11716 5914 11744 12679
rect 11808 11830 11836 13262
rect 11900 13190 11928 13466
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11796 11824 11848 11830
rect 11796 11766 11848 11772
rect 11808 11082 11836 11766
rect 11900 11150 11928 12922
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 11808 10674 11836 11018
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11808 10130 11836 10610
rect 11796 10124 11848 10130
rect 11796 10066 11848 10072
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11808 8634 11836 8774
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11900 6610 11928 11086
rect 11992 9674 12020 14758
rect 12084 13274 12112 15846
rect 12176 14822 12204 16662
rect 12164 14816 12216 14822
rect 12164 14758 12216 14764
rect 12162 14512 12218 14521
rect 12162 14447 12164 14456
rect 12216 14447 12218 14456
rect 12164 14418 12216 14424
rect 12164 13728 12216 13734
rect 12164 13670 12216 13676
rect 12176 13530 12204 13670
rect 12164 13524 12216 13530
rect 12164 13466 12216 13472
rect 12268 13462 12296 16934
rect 12360 13938 12388 17054
rect 12452 15586 12480 19200
rect 12624 17332 12676 17338
rect 12624 17274 12676 17280
rect 12532 16720 12584 16726
rect 12532 16662 12584 16668
rect 12544 16153 12572 16662
rect 12530 16144 12586 16153
rect 12530 16079 12586 16088
rect 12532 15972 12584 15978
rect 12532 15914 12584 15920
rect 12544 15706 12572 15914
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12452 15558 12572 15586
rect 12440 15496 12492 15502
rect 12440 15438 12492 15444
rect 12452 15162 12480 15438
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12438 14920 12494 14929
rect 12438 14855 12494 14864
rect 12452 14822 12480 14855
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12544 14550 12572 15558
rect 12636 14906 12664 17274
rect 12912 17066 12940 19200
rect 13280 17134 13308 19200
rect 13648 17626 13676 19200
rect 13648 17598 13860 17626
rect 13449 17436 13745 17456
rect 13505 17434 13529 17436
rect 13585 17434 13609 17436
rect 13665 17434 13689 17436
rect 13527 17382 13529 17434
rect 13591 17382 13603 17434
rect 13665 17382 13667 17434
rect 13505 17380 13529 17382
rect 13585 17380 13609 17382
rect 13665 17380 13689 17382
rect 13449 17360 13745 17380
rect 13268 17128 13320 17134
rect 13268 17070 13320 17076
rect 12900 17060 12952 17066
rect 12900 17002 12952 17008
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 12728 15094 12756 16934
rect 12808 15972 12860 15978
rect 12808 15914 12860 15920
rect 12716 15088 12768 15094
rect 12716 15030 12768 15036
rect 12716 14952 12768 14958
rect 12636 14900 12716 14906
rect 12636 14894 12768 14900
rect 12636 14878 12756 14894
rect 12532 14544 12584 14550
rect 12532 14486 12584 14492
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 12452 13802 12480 14418
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12728 14226 12756 14878
rect 12820 14482 12848 15914
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 12912 15065 12940 15506
rect 13004 15434 13032 16934
rect 13176 16448 13228 16454
rect 13176 16390 13228 16396
rect 13188 15570 13216 16390
rect 13280 16250 13308 17070
rect 13832 16998 13860 17598
rect 13912 17332 13964 17338
rect 13964 17292 14044 17320
rect 13912 17274 13964 17280
rect 13912 17196 13964 17202
rect 13912 17138 13964 17144
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13924 16794 13952 17138
rect 13912 16788 13964 16794
rect 13912 16730 13964 16736
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13268 16244 13320 16250
rect 13268 16186 13320 16192
rect 13372 16046 13400 16390
rect 13449 16348 13745 16368
rect 13505 16346 13529 16348
rect 13585 16346 13609 16348
rect 13665 16346 13689 16348
rect 13527 16294 13529 16346
rect 13591 16294 13603 16346
rect 13665 16294 13667 16346
rect 13505 16292 13529 16294
rect 13585 16292 13609 16294
rect 13665 16292 13689 16294
rect 13449 16272 13745 16292
rect 13360 16040 13412 16046
rect 13360 15982 13412 15988
rect 13832 15910 13860 16594
rect 13924 16046 13952 16730
rect 13912 16040 13964 16046
rect 13912 15982 13964 15988
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 13728 15700 13780 15706
rect 13728 15642 13780 15648
rect 13268 15632 13320 15638
rect 13268 15574 13320 15580
rect 13176 15564 13228 15570
rect 13176 15506 13228 15512
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 12992 15428 13044 15434
rect 12992 15370 13044 15376
rect 13096 15162 13124 15438
rect 13084 15156 13136 15162
rect 13084 15098 13136 15104
rect 12898 15056 12954 15065
rect 13174 15056 13230 15065
rect 12898 14991 12954 15000
rect 13084 15020 13136 15026
rect 13280 15026 13308 15574
rect 13740 15348 13768 15642
rect 13832 15502 13860 15846
rect 14016 15706 14044 17292
rect 14108 16980 14136 19200
rect 14280 17264 14332 17270
rect 14280 17206 14332 17212
rect 14188 16992 14240 16998
rect 14108 16952 14188 16980
rect 14004 15700 14056 15706
rect 14004 15642 14056 15648
rect 14004 15564 14056 15570
rect 14004 15506 14056 15512
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13912 15360 13964 15366
rect 13740 15320 13860 15348
rect 13449 15260 13745 15280
rect 13505 15258 13529 15260
rect 13585 15258 13609 15260
rect 13665 15258 13689 15260
rect 13527 15206 13529 15258
rect 13591 15206 13603 15258
rect 13665 15206 13667 15258
rect 13505 15204 13529 15206
rect 13585 15204 13609 15206
rect 13665 15204 13689 15206
rect 13449 15184 13745 15204
rect 13174 14991 13230 15000
rect 13268 15020 13320 15026
rect 13084 14962 13136 14968
rect 12898 14920 12954 14929
rect 12898 14855 12954 14864
rect 12808 14476 12860 14482
rect 12808 14418 12860 14424
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 12440 13796 12492 13802
rect 12440 13738 12492 13744
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12256 13456 12308 13462
rect 12452 13433 12480 13466
rect 12256 13398 12308 13404
rect 12438 13424 12494 13433
rect 12084 13246 12204 13274
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 12084 10742 12112 13126
rect 12176 11218 12204 13246
rect 12268 12753 12296 13398
rect 12438 13359 12494 13368
rect 12346 13152 12402 13161
rect 12346 13087 12402 13096
rect 12254 12744 12310 12753
rect 12254 12679 12310 12688
rect 12164 11212 12216 11218
rect 12164 11154 12216 11160
rect 12072 10736 12124 10742
rect 12124 10696 12204 10724
rect 12072 10678 12124 10684
rect 11992 9646 12112 9674
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 11992 8498 12020 8774
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 11992 7886 12020 8434
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 12084 7410 12112 9646
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 11808 6582 11928 6610
rect 11808 6118 11836 6582
rect 12084 6474 12112 7346
rect 12176 7342 12204 10696
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12268 10198 12296 10610
rect 12256 10192 12308 10198
rect 12256 10134 12308 10140
rect 12256 9920 12308 9926
rect 12256 9862 12308 9868
rect 12268 7750 12296 9862
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12164 7336 12216 7342
rect 12164 7278 12216 7284
rect 12268 7188 12296 7686
rect 11900 6446 12112 6474
rect 12176 7160 12296 7188
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11612 5772 11664 5778
rect 11532 5732 11612 5760
rect 11612 5714 11664 5720
rect 10968 5568 11020 5574
rect 11336 5568 11388 5574
rect 10968 5510 11020 5516
rect 11058 5536 11114 5545
rect 10980 5012 11008 5510
rect 11336 5510 11388 5516
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11058 5471 11114 5480
rect 11072 5370 11100 5471
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 10704 4814 10824 4842
rect 10888 4984 11008 5012
rect 11336 5024 11388 5030
rect 10704 4554 10732 4814
rect 10888 4808 10916 4984
rect 11336 4966 11388 4972
rect 10950 4924 11246 4944
rect 11006 4922 11030 4924
rect 11086 4922 11110 4924
rect 11166 4922 11190 4924
rect 11028 4870 11030 4922
rect 11092 4870 11104 4922
rect 11166 4870 11168 4922
rect 11006 4868 11030 4870
rect 11086 4868 11110 4870
rect 11166 4868 11190 4870
rect 10950 4848 11246 4868
rect 11348 4808 11376 4966
rect 10888 4780 11008 4808
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 10692 4548 10744 4554
rect 10692 4490 10744 4496
rect 10796 4214 10824 4694
rect 10784 4208 10836 4214
rect 10784 4150 10836 4156
rect 10876 4072 10928 4078
rect 10704 4032 10876 4060
rect 10600 3664 10652 3670
rect 10600 3606 10652 3612
rect 10600 3392 10652 3398
rect 10414 3360 10470 3369
rect 10600 3334 10652 3340
rect 10414 3295 10470 3304
rect 10612 2961 10640 3334
rect 10598 2952 10654 2961
rect 10232 2916 10284 2922
rect 10598 2887 10654 2896
rect 10232 2858 10284 2864
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 10244 800 10272 2858
rect 10600 2848 10652 2854
rect 10600 2790 10652 2796
rect 10612 2446 10640 2790
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10704 800 10732 4032
rect 10876 4014 10928 4020
rect 10980 4010 11008 4780
rect 11164 4780 11376 4808
rect 11164 4078 11192 4780
rect 11532 4282 11560 5510
rect 11716 5409 11744 5850
rect 11702 5400 11758 5409
rect 11702 5335 11758 5344
rect 11808 5273 11836 6054
rect 11794 5264 11850 5273
rect 11794 5199 11850 5208
rect 11612 5092 11664 5098
rect 11612 5034 11664 5040
rect 11520 4276 11572 4282
rect 11520 4218 11572 4224
rect 11244 4208 11296 4214
rect 11244 4150 11296 4156
rect 11152 4072 11204 4078
rect 11152 4014 11204 4020
rect 10968 4004 11020 4010
rect 10968 3946 11020 3952
rect 10876 3936 10928 3942
rect 11256 3924 11284 4150
rect 11520 4072 11572 4078
rect 11520 4014 11572 4020
rect 11532 3942 11560 4014
rect 11520 3936 11572 3942
rect 11256 3896 11376 3924
rect 10876 3878 10928 3884
rect 10888 3738 10916 3878
rect 10950 3836 11246 3856
rect 11006 3834 11030 3836
rect 11086 3834 11110 3836
rect 11166 3834 11190 3836
rect 11028 3782 11030 3834
rect 11092 3782 11104 3834
rect 11166 3782 11168 3834
rect 11006 3780 11030 3782
rect 11086 3780 11110 3782
rect 11166 3780 11190 3782
rect 10950 3760 11246 3780
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 10796 2922 10824 3470
rect 11256 3466 11284 3538
rect 11244 3460 11296 3466
rect 11244 3402 11296 3408
rect 10876 3392 10928 3398
rect 10876 3334 10928 3340
rect 10784 2916 10836 2922
rect 10784 2858 10836 2864
rect 10796 2446 10824 2858
rect 10888 2514 10916 3334
rect 10950 2748 11246 2768
rect 11006 2746 11030 2748
rect 11086 2746 11110 2748
rect 11166 2746 11190 2748
rect 11028 2694 11030 2746
rect 11092 2694 11104 2746
rect 11166 2694 11168 2746
rect 11006 2692 11030 2694
rect 11086 2692 11110 2694
rect 11166 2692 11190 2694
rect 10950 2672 11246 2692
rect 11348 2650 11376 3896
rect 11520 3878 11572 3884
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 11426 3496 11482 3505
rect 11426 3431 11482 3440
rect 11336 2644 11388 2650
rect 11336 2586 11388 2592
rect 11334 2544 11390 2553
rect 10876 2508 10928 2514
rect 11334 2479 11390 2488
rect 10876 2450 10928 2456
rect 11348 2446 11376 2479
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 11336 2440 11388 2446
rect 11336 2382 11388 2388
rect 11440 1442 11468 3431
rect 11072 1414 11468 1442
rect 11072 800 11100 1414
rect 11532 800 11560 3538
rect 11624 2990 11652 5034
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11716 2990 11744 4966
rect 11808 4758 11836 4966
rect 11796 4752 11848 4758
rect 11796 4694 11848 4700
rect 11900 4078 11928 6446
rect 11980 6384 12032 6390
rect 11980 6326 12032 6332
rect 11992 5710 12020 6326
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 12176 5574 12204 7160
rect 12360 6440 12388 13087
rect 12544 12782 12572 13806
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12544 10554 12572 11494
rect 12636 10810 12664 14214
rect 12728 14198 12848 14226
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12728 12850 12756 13262
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12728 12442 12756 12786
rect 12716 12436 12768 12442
rect 12716 12378 12768 12384
rect 12820 12322 12848 14198
rect 12912 13190 12940 14855
rect 12992 14544 13044 14550
rect 12992 14486 13044 14492
rect 13004 13326 13032 14486
rect 13096 14482 13124 14962
rect 13084 14476 13136 14482
rect 13084 14418 13136 14424
rect 13096 14278 13124 14418
rect 13084 14272 13136 14278
rect 13084 14214 13136 14220
rect 13096 13938 13124 14214
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 13188 13818 13216 14991
rect 13268 14962 13320 14968
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 13360 14952 13412 14958
rect 13360 14894 13412 14900
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13280 14006 13308 14758
rect 13372 14074 13400 14894
rect 13740 14550 13768 14962
rect 13728 14544 13780 14550
rect 13728 14486 13780 14492
rect 13449 14172 13745 14192
rect 13505 14170 13529 14172
rect 13585 14170 13609 14172
rect 13665 14170 13689 14172
rect 13527 14118 13529 14170
rect 13591 14118 13603 14170
rect 13665 14118 13667 14170
rect 13505 14116 13529 14118
rect 13585 14116 13609 14118
rect 13665 14116 13689 14118
rect 13449 14096 13745 14116
rect 13360 14068 13412 14074
rect 13832 14056 13860 15320
rect 13912 15302 13964 15308
rect 13360 14010 13412 14016
rect 13740 14028 13860 14056
rect 13268 14000 13320 14006
rect 13268 13942 13320 13948
rect 13084 13796 13136 13802
rect 13188 13790 13308 13818
rect 13084 13738 13136 13744
rect 13096 13326 13124 13738
rect 13280 13326 13308 13790
rect 13544 13796 13596 13802
rect 13544 13738 13596 13744
rect 13556 13530 13584 13738
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 13648 13530 13676 13670
rect 13740 13569 13768 14028
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13726 13560 13782 13569
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13636 13524 13688 13530
rect 13726 13495 13782 13504
rect 13636 13466 13688 13472
rect 13360 13388 13412 13394
rect 13360 13330 13412 13336
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 12900 13184 12952 13190
rect 13084 13184 13136 13190
rect 12900 13126 12952 13132
rect 12990 13152 13046 13161
rect 13084 13126 13136 13132
rect 12990 13087 13046 13096
rect 12898 13016 12954 13025
rect 12898 12951 12900 12960
rect 12952 12951 12954 12960
rect 12900 12922 12952 12928
rect 13004 12730 13032 13087
rect 12912 12714 13032 12730
rect 12900 12708 13032 12714
rect 12952 12702 13032 12708
rect 12900 12650 12952 12656
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 12728 12294 12848 12322
rect 12728 11558 12756 12294
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12544 10526 12664 10554
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12452 9654 12480 10406
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12452 8090 12480 9318
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12438 7304 12494 7313
rect 12544 7290 12572 8774
rect 12636 7410 12664 10526
rect 12820 9518 12848 12174
rect 12900 11280 12952 11286
rect 13004 11257 13032 12582
rect 12900 11222 12952 11228
rect 12990 11248 13046 11257
rect 12912 10690 12940 11222
rect 12990 11183 13046 11192
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 13004 10810 13032 11086
rect 12992 10804 13044 10810
rect 12992 10746 13044 10752
rect 12912 10662 13032 10690
rect 12900 10532 12952 10538
rect 12900 10474 12952 10480
rect 12912 9518 12940 10474
rect 13004 9926 13032 10662
rect 12992 9920 13044 9926
rect 12992 9862 13044 9868
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12900 9512 12952 9518
rect 12900 9454 12952 9460
rect 12808 9376 12860 9382
rect 13004 9330 13032 9862
rect 12860 9324 13032 9330
rect 12808 9318 13032 9324
rect 12820 9302 13032 9318
rect 13004 9178 13032 9302
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12728 7936 12756 8978
rect 12820 8430 12848 9114
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12808 8424 12860 8430
rect 12808 8366 12860 8372
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12820 8090 12848 8230
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 12912 8022 12940 8774
rect 13096 8072 13124 13126
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 13188 10266 13216 10406
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 13004 8044 13124 8072
rect 12900 8016 12952 8022
rect 12900 7958 12952 7964
rect 12728 7908 12848 7936
rect 12716 7812 12768 7818
rect 12716 7754 12768 7760
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 12494 7262 12572 7290
rect 12728 7274 12756 7754
rect 12716 7268 12768 7274
rect 12438 7239 12494 7248
rect 12268 6412 12388 6440
rect 12268 5914 12296 6412
rect 12346 6352 12402 6361
rect 12346 6287 12402 6296
rect 12360 6186 12388 6287
rect 12348 6180 12400 6186
rect 12348 6122 12400 6128
rect 12256 5908 12308 5914
rect 12256 5850 12308 5856
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 12164 5568 12216 5574
rect 12164 5510 12216 5516
rect 11888 4072 11940 4078
rect 11888 4014 11940 4020
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11886 3904 11942 3913
rect 11612 2984 11664 2990
rect 11612 2926 11664 2932
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 11808 2378 11836 3878
rect 11886 3839 11942 3848
rect 11900 3482 11928 3839
rect 11992 3602 12020 5510
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 12084 4826 12112 5102
rect 12072 4820 12124 4826
rect 12072 4762 12124 4768
rect 12072 4684 12124 4690
rect 12072 4626 12124 4632
rect 12084 4214 12112 4626
rect 12072 4208 12124 4214
rect 12072 4150 12124 4156
rect 12072 4004 12124 4010
rect 12072 3946 12124 3952
rect 11980 3596 12032 3602
rect 11980 3538 12032 3544
rect 11900 3454 12020 3482
rect 11886 3360 11942 3369
rect 11886 3295 11942 3304
rect 11900 3126 11928 3295
rect 11992 3126 12020 3454
rect 11888 3120 11940 3126
rect 11888 3062 11940 3068
rect 11980 3120 12032 3126
rect 11980 3062 12032 3068
rect 11886 2952 11942 2961
rect 11886 2887 11942 2896
rect 11900 2854 11928 2887
rect 11888 2848 11940 2854
rect 11888 2790 11940 2796
rect 11992 2514 12020 3062
rect 12084 2961 12112 3946
rect 12176 3942 12204 5510
rect 12268 4146 12296 5850
rect 12256 4140 12308 4146
rect 12256 4082 12308 4088
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 12176 3346 12204 3878
rect 12268 3466 12296 4082
rect 12360 3913 12388 5850
rect 12452 5710 12480 7239
rect 12716 7210 12768 7216
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12544 7002 12572 7142
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12636 6361 12664 7142
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 12728 6458 12756 6802
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12622 6352 12678 6361
rect 12622 6287 12678 6296
rect 12624 6248 12676 6254
rect 12624 6190 12676 6196
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 12346 3904 12402 3913
rect 12346 3839 12402 3848
rect 12360 3670 12388 3701
rect 12348 3664 12400 3670
rect 12346 3632 12348 3641
rect 12400 3632 12402 3641
rect 12452 3618 12480 4422
rect 12636 4321 12664 6190
rect 12820 5846 12848 7908
rect 13004 7834 13032 8044
rect 13084 7948 13136 7954
rect 13084 7890 13136 7896
rect 12912 7806 13032 7834
rect 12912 6769 12940 7806
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 12898 6760 12954 6769
rect 12898 6695 12954 6704
rect 12912 5914 12940 6695
rect 12900 5908 12952 5914
rect 12900 5850 12952 5856
rect 12808 5840 12860 5846
rect 12728 5800 12808 5828
rect 12622 4312 12678 4321
rect 12622 4247 12678 4256
rect 12622 4176 12678 4185
rect 12622 4111 12678 4120
rect 12532 4004 12584 4010
rect 12532 3946 12584 3952
rect 12402 3590 12480 3618
rect 12346 3567 12402 3576
rect 12256 3460 12308 3466
rect 12256 3402 12308 3408
rect 12348 3460 12400 3466
rect 12348 3402 12400 3408
rect 12176 3318 12296 3346
rect 12070 2952 12126 2961
rect 12070 2887 12126 2896
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 11796 2372 11848 2378
rect 11796 2314 11848 2320
rect 12268 2310 12296 3318
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 11888 1896 11940 1902
rect 11888 1838 11940 1844
rect 11900 800 11928 1838
rect 12360 800 12388 3402
rect 12544 3108 12572 3946
rect 12636 3670 12664 4111
rect 12728 3738 12756 5800
rect 12808 5782 12860 5788
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 12624 3664 12676 3670
rect 12624 3606 12676 3612
rect 12820 3602 12848 5646
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12624 3528 12676 3534
rect 12624 3470 12676 3476
rect 12452 3080 12572 3108
rect 12452 2378 12480 3080
rect 12532 2916 12584 2922
rect 12636 2904 12664 3470
rect 12584 2876 12664 2904
rect 12532 2858 12584 2864
rect 12544 2428 12572 2858
rect 12808 2848 12860 2854
rect 12808 2790 12860 2796
rect 12622 2680 12678 2689
rect 12820 2650 12848 2790
rect 12622 2615 12624 2624
rect 12676 2615 12678 2624
rect 12808 2644 12860 2650
rect 12624 2586 12676 2592
rect 12808 2586 12860 2592
rect 12716 2508 12768 2514
rect 12716 2450 12768 2456
rect 12624 2440 12676 2446
rect 12544 2400 12624 2428
rect 12624 2382 12676 2388
rect 12440 2372 12492 2378
rect 12440 2314 12492 2320
rect 12636 2106 12664 2382
rect 12624 2100 12676 2106
rect 12624 2042 12676 2048
rect 12728 800 12756 2450
rect 12912 2378 12940 3878
rect 13004 3602 13032 7686
rect 13096 6730 13124 7890
rect 13084 6724 13136 6730
rect 13084 6666 13136 6672
rect 13188 6610 13216 10202
rect 13280 9994 13308 13262
rect 13372 12850 13400 13330
rect 13648 13258 13676 13466
rect 13636 13252 13688 13258
rect 13636 13194 13688 13200
rect 13449 13084 13745 13104
rect 13505 13082 13529 13084
rect 13585 13082 13609 13084
rect 13665 13082 13689 13084
rect 13527 13030 13529 13082
rect 13591 13030 13603 13082
rect 13665 13030 13667 13082
rect 13505 13028 13529 13030
rect 13585 13028 13609 13030
rect 13665 13028 13689 13030
rect 13449 13008 13745 13028
rect 13832 12986 13860 13806
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 13449 11996 13745 12016
rect 13505 11994 13529 11996
rect 13585 11994 13609 11996
rect 13665 11994 13689 11996
rect 13527 11942 13529 11994
rect 13591 11942 13603 11994
rect 13665 11942 13667 11994
rect 13505 11940 13529 11942
rect 13585 11940 13609 11942
rect 13665 11940 13689 11942
rect 13449 11920 13745 11940
rect 13924 10962 13952 15302
rect 14016 14074 14044 15506
rect 14108 15162 14136 16952
rect 14188 16934 14240 16940
rect 14188 16584 14240 16590
rect 14188 16526 14240 16532
rect 14200 15978 14228 16526
rect 14188 15972 14240 15978
rect 14188 15914 14240 15920
rect 14292 15586 14320 17206
rect 14476 16658 14504 19200
rect 14832 17332 14884 17338
rect 14832 17274 14884 17280
rect 14556 17128 14608 17134
rect 14556 17070 14608 17076
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 14372 15904 14424 15910
rect 14372 15846 14424 15852
rect 14200 15558 14320 15586
rect 14096 15156 14148 15162
rect 14096 15098 14148 15104
rect 14004 14068 14056 14074
rect 14004 14010 14056 14016
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 14016 12374 14044 13466
rect 14200 12714 14228 15558
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 14292 15094 14320 15438
rect 14280 15088 14332 15094
rect 14280 15030 14332 15036
rect 14384 14906 14412 15846
rect 14292 14878 14412 14906
rect 14188 12708 14240 12714
rect 14188 12650 14240 12656
rect 14004 12368 14056 12374
rect 14004 12310 14056 12316
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 13924 10934 14044 10962
rect 13449 10908 13745 10928
rect 13505 10906 13529 10908
rect 13585 10906 13609 10908
rect 13665 10906 13689 10908
rect 13527 10854 13529 10906
rect 13591 10854 13603 10906
rect 13665 10854 13667 10906
rect 13505 10852 13529 10854
rect 13585 10852 13609 10854
rect 13665 10852 13689 10854
rect 13449 10832 13745 10852
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 13360 10532 13412 10538
rect 13360 10474 13412 10480
rect 13372 10062 13400 10474
rect 13452 10192 13504 10198
rect 13450 10160 13452 10169
rect 13504 10160 13506 10169
rect 13450 10095 13506 10104
rect 13360 10056 13412 10062
rect 13360 9998 13412 10004
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13268 9988 13320 9994
rect 13268 9930 13320 9936
rect 13372 9874 13400 9998
rect 13280 9846 13400 9874
rect 13280 9586 13308 9846
rect 13449 9820 13745 9840
rect 13505 9818 13529 9820
rect 13585 9818 13609 9820
rect 13665 9818 13689 9820
rect 13527 9766 13529 9818
rect 13591 9766 13603 9818
rect 13665 9766 13667 9818
rect 13505 9764 13529 9766
rect 13585 9764 13609 9766
rect 13665 9764 13689 9766
rect 13449 9744 13745 9764
rect 13832 9722 13860 9998
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 13924 9586 13952 10746
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13912 9580 13964 9586
rect 13912 9522 13964 9528
rect 13280 8634 13308 9522
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13464 8820 13492 9318
rect 13372 8792 13492 8820
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13280 7886 13308 8570
rect 13372 8090 13400 8792
rect 13449 8732 13745 8752
rect 13505 8730 13529 8732
rect 13585 8730 13609 8732
rect 13665 8730 13689 8732
rect 13527 8678 13529 8730
rect 13591 8678 13603 8730
rect 13665 8678 13667 8730
rect 13505 8676 13529 8678
rect 13585 8676 13609 8678
rect 13665 8676 13689 8678
rect 13449 8656 13745 8676
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13464 7732 13492 8298
rect 14016 8090 14044 10934
rect 14200 10810 14228 11154
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 14108 9586 14136 9862
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14200 9518 14228 9862
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 14004 8084 14056 8090
rect 14004 8026 14056 8032
rect 13372 7704 13492 7732
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 13096 6582 13216 6610
rect 13096 4146 13124 6582
rect 13280 6322 13308 7346
rect 13372 6458 13400 7704
rect 13449 7644 13745 7664
rect 13505 7642 13529 7644
rect 13585 7642 13609 7644
rect 13665 7642 13689 7644
rect 13527 7590 13529 7642
rect 13591 7590 13603 7642
rect 13665 7590 13667 7642
rect 13505 7588 13529 7590
rect 13585 7588 13609 7590
rect 13665 7588 13689 7590
rect 13449 7568 13745 7588
rect 13449 6556 13745 6576
rect 13505 6554 13529 6556
rect 13585 6554 13609 6556
rect 13665 6554 13689 6556
rect 13527 6502 13529 6554
rect 13591 6502 13603 6554
rect 13665 6502 13667 6554
rect 13505 6500 13529 6502
rect 13585 6500 13609 6502
rect 13665 6500 13689 6502
rect 13449 6480 13745 6500
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 13268 6316 13320 6322
rect 13268 6258 13320 6264
rect 13360 5772 13412 5778
rect 13360 5714 13412 5720
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 13176 5636 13228 5642
rect 13176 5578 13228 5584
rect 13188 5370 13216 5578
rect 13176 5364 13228 5370
rect 13176 5306 13228 5312
rect 13176 5092 13228 5098
rect 13176 5034 13228 5040
rect 13188 4826 13216 5034
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 13188 4214 13216 4762
rect 13176 4208 13228 4214
rect 13176 4150 13228 4156
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 13280 3942 13308 5646
rect 13372 4010 13400 5714
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13912 5568 13964 5574
rect 13912 5510 13964 5516
rect 13449 5468 13745 5488
rect 13505 5466 13529 5468
rect 13585 5466 13609 5468
rect 13665 5466 13689 5468
rect 13527 5414 13529 5466
rect 13591 5414 13603 5466
rect 13665 5414 13667 5466
rect 13505 5412 13529 5414
rect 13585 5412 13609 5414
rect 13665 5412 13689 5414
rect 13449 5392 13745 5412
rect 13449 4380 13745 4400
rect 13505 4378 13529 4380
rect 13585 4378 13609 4380
rect 13665 4378 13689 4380
rect 13527 4326 13529 4378
rect 13591 4326 13603 4378
rect 13665 4326 13667 4378
rect 13505 4324 13529 4326
rect 13585 4324 13609 4326
rect 13665 4324 13689 4326
rect 13449 4304 13745 4324
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13360 4004 13412 4010
rect 13360 3946 13412 3952
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 13096 3233 13124 3674
rect 13740 3602 13768 4082
rect 13728 3596 13780 3602
rect 13728 3538 13780 3544
rect 13832 3534 13860 5510
rect 13924 3602 13952 5510
rect 14004 4480 14056 4486
rect 14004 4422 14056 4428
rect 14016 4078 14044 4422
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 13820 3528 13872 3534
rect 14108 3482 14136 6394
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 13820 3470 13872 3476
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13082 3224 13138 3233
rect 13082 3159 13138 3168
rect 13372 2650 13400 3334
rect 13449 3292 13745 3312
rect 13505 3290 13529 3292
rect 13585 3290 13609 3292
rect 13665 3290 13689 3292
rect 13527 3238 13529 3290
rect 13591 3238 13603 3290
rect 13665 3238 13667 3290
rect 13505 3236 13529 3238
rect 13585 3236 13609 3238
rect 13665 3236 13689 3238
rect 13449 3216 13745 3236
rect 13452 2984 13504 2990
rect 13452 2926 13504 2932
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 13176 2576 13228 2582
rect 13464 2530 13492 2926
rect 13176 2518 13228 2524
rect 12900 2372 12952 2378
rect 12900 2314 12952 2320
rect 13188 800 13216 2518
rect 13372 2502 13492 2530
rect 13372 1952 13400 2502
rect 13449 2204 13745 2224
rect 13505 2202 13529 2204
rect 13585 2202 13609 2204
rect 13665 2202 13689 2204
rect 13527 2150 13529 2202
rect 13591 2150 13603 2202
rect 13665 2150 13667 2202
rect 13505 2148 13529 2150
rect 13585 2148 13609 2150
rect 13665 2148 13689 2150
rect 13449 2128 13745 2148
rect 13372 1924 13584 1952
rect 13556 800 13584 1924
rect 13832 1902 13860 3470
rect 14016 3454 14136 3482
rect 14016 2922 14044 3454
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 14004 2916 14056 2922
rect 14004 2858 14056 2864
rect 14108 2514 14136 3334
rect 14200 3194 14228 4558
rect 14292 4010 14320 14878
rect 14476 14550 14504 16594
rect 14568 15473 14596 17070
rect 14648 16788 14700 16794
rect 14648 16730 14700 16736
rect 14554 15464 14610 15473
rect 14554 15399 14610 15408
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14568 14618 14596 14758
rect 14556 14612 14608 14618
rect 14556 14554 14608 14560
rect 14464 14544 14516 14550
rect 14464 14486 14516 14492
rect 14554 14376 14610 14385
rect 14554 14311 14610 14320
rect 14568 13938 14596 14311
rect 14556 13932 14608 13938
rect 14556 13874 14608 13880
rect 14370 13560 14426 13569
rect 14370 13495 14426 13504
rect 14384 13462 14412 13495
rect 14372 13456 14424 13462
rect 14372 13398 14424 13404
rect 14372 12980 14424 12986
rect 14372 12922 14424 12928
rect 14384 8362 14412 12922
rect 14556 12368 14608 12374
rect 14556 12310 14608 12316
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14476 10266 14504 10406
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 14372 8356 14424 8362
rect 14372 8298 14424 8304
rect 14372 5840 14424 5846
rect 14372 5782 14424 5788
rect 14384 4690 14412 5782
rect 14372 4684 14424 4690
rect 14372 4626 14424 4632
rect 14372 4480 14424 4486
rect 14372 4422 14424 4428
rect 14384 4078 14412 4422
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14280 4004 14332 4010
rect 14280 3946 14332 3952
rect 14476 3194 14504 9114
rect 14568 6458 14596 12310
rect 14660 11354 14688 16730
rect 14740 16652 14792 16658
rect 14740 16594 14792 16600
rect 14752 15609 14780 16594
rect 14738 15600 14794 15609
rect 14738 15535 14794 15544
rect 14740 15020 14792 15026
rect 14740 14962 14792 14968
rect 14752 13530 14780 14962
rect 14844 14226 14872 17274
rect 14936 16046 14964 19200
rect 15016 17332 15068 17338
rect 15016 17274 15068 17280
rect 14924 16040 14976 16046
rect 14924 15982 14976 15988
rect 14936 14414 14964 15982
rect 15028 15910 15056 17274
rect 15304 17082 15332 19200
rect 15304 17054 15700 17082
rect 15292 16992 15344 16998
rect 15292 16934 15344 16940
rect 15304 16658 15332 16934
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15304 16538 15332 16594
rect 15304 16510 15424 16538
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 15016 15904 15068 15910
rect 15016 15846 15068 15852
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 15028 14906 15056 15506
rect 15108 15496 15160 15502
rect 15108 15438 15160 15444
rect 15120 15026 15148 15438
rect 15108 15020 15160 15026
rect 15108 14962 15160 14968
rect 15028 14878 15148 14906
rect 14924 14408 14976 14414
rect 14924 14350 14976 14356
rect 14844 14198 15056 14226
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 14740 13184 14792 13190
rect 14844 13172 14872 14010
rect 14792 13144 14872 13172
rect 14740 13126 14792 13132
rect 14752 12889 14780 13126
rect 14738 12880 14794 12889
rect 14738 12815 14794 12824
rect 14648 11348 14700 11354
rect 14648 11290 14700 11296
rect 14752 6458 14780 12815
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 14568 4758 14596 6394
rect 14648 5772 14700 5778
rect 14648 5714 14700 5720
rect 14556 4752 14608 4758
rect 14556 4694 14608 4700
rect 14660 4570 14688 5714
rect 14752 4758 14780 6394
rect 14740 4752 14792 4758
rect 14740 4694 14792 4700
rect 14660 4542 14780 4570
rect 14648 4480 14700 4486
rect 14648 4422 14700 4428
rect 14660 3670 14688 4422
rect 14648 3664 14700 3670
rect 14568 3624 14648 3652
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 14464 3188 14516 3194
rect 14464 3130 14516 3136
rect 14200 3074 14228 3130
rect 14200 3046 14320 3074
rect 14186 2952 14242 2961
rect 14186 2887 14242 2896
rect 14200 2650 14228 2887
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 14096 2508 14148 2514
rect 14096 2450 14148 2456
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 13820 1896 13872 1902
rect 13820 1838 13872 1844
rect 14016 800 14044 2382
rect 14292 2378 14320 3046
rect 14280 2372 14332 2378
rect 14280 2314 14332 2320
rect 14568 2258 14596 3624
rect 14648 3606 14700 3612
rect 14752 2990 14780 4542
rect 14740 2984 14792 2990
rect 14476 2230 14596 2258
rect 14660 2944 14740 2972
rect 14476 800 14504 2230
rect 14660 2038 14688 2944
rect 14740 2926 14792 2932
rect 14740 2848 14792 2854
rect 14740 2790 14792 2796
rect 14752 2582 14780 2790
rect 14740 2576 14792 2582
rect 14740 2518 14792 2524
rect 14844 2514 14872 12718
rect 14924 12300 14976 12306
rect 14924 12242 14976 12248
rect 14936 5778 14964 12242
rect 15028 10266 15056 14198
rect 15120 14074 15148 14878
rect 15212 14550 15240 16390
rect 15292 15972 15344 15978
rect 15292 15914 15344 15920
rect 15304 15745 15332 15914
rect 15290 15736 15346 15745
rect 15290 15671 15346 15680
rect 15292 15360 15344 15366
rect 15292 15302 15344 15308
rect 15304 15026 15332 15302
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 15396 14906 15424 16510
rect 15304 14878 15424 14906
rect 15200 14544 15252 14550
rect 15200 14486 15252 14492
rect 15200 14340 15252 14346
rect 15200 14282 15252 14288
rect 15108 14068 15160 14074
rect 15108 14010 15160 14016
rect 15108 13796 15160 13802
rect 15108 13738 15160 13744
rect 15120 13530 15148 13738
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 15212 12918 15240 14282
rect 15304 13394 15332 14878
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15396 13530 15424 14418
rect 15384 13524 15436 13530
rect 15384 13466 15436 13472
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15200 12912 15252 12918
rect 15200 12854 15252 12860
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 15120 12306 15148 12718
rect 15108 12300 15160 12306
rect 15108 12242 15160 12248
rect 15108 10464 15160 10470
rect 15108 10406 15160 10412
rect 15016 10260 15068 10266
rect 15016 10202 15068 10208
rect 15120 10130 15148 10406
rect 15304 10198 15332 13330
rect 15488 12850 15516 16594
rect 15672 15638 15700 17054
rect 15764 16250 15792 19200
rect 16132 18034 16160 19200
rect 16040 18006 16160 18034
rect 16040 16522 16068 18006
rect 16118 17912 16174 17921
rect 16118 17847 16174 17856
rect 16028 16516 16080 16522
rect 16028 16458 16080 16464
rect 15752 16244 15804 16250
rect 15752 16186 15804 16192
rect 15660 15632 15712 15638
rect 15660 15574 15712 15580
rect 16132 15162 16160 17847
rect 16120 15156 16172 15162
rect 16120 15098 16172 15104
rect 16592 14482 16620 19200
rect 16960 16794 16988 19200
rect 16948 16788 17000 16794
rect 16948 16730 17000 16736
rect 16580 14476 16632 14482
rect 16580 14418 16632 14424
rect 15658 13968 15714 13977
rect 15658 13903 15714 13912
rect 15568 13796 15620 13802
rect 15568 13738 15620 13744
rect 15580 13530 15608 13738
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 15672 13394 15700 13903
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 15672 12986 15700 13330
rect 15660 12980 15712 12986
rect 15660 12922 15712 12928
rect 15476 12844 15528 12850
rect 15476 12786 15528 12792
rect 15292 10192 15344 10198
rect 15292 10134 15344 10140
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 15120 9110 15148 10066
rect 15660 9988 15712 9994
rect 15660 9930 15712 9936
rect 15672 9897 15700 9930
rect 15658 9888 15714 9897
rect 15658 9823 15714 9832
rect 15108 9104 15160 9110
rect 15108 9046 15160 9052
rect 14924 5772 14976 5778
rect 14924 5714 14976 5720
rect 14924 5024 14976 5030
rect 14924 4966 14976 4972
rect 15016 5024 15068 5030
rect 15016 4966 15068 4972
rect 14936 4826 14964 4966
rect 14924 4820 14976 4826
rect 14924 4762 14976 4768
rect 15028 4298 15056 4966
rect 14936 4282 15056 4298
rect 15120 4282 15148 9046
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 15292 5636 15344 5642
rect 15292 5578 15344 5584
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 14924 4276 15056 4282
rect 14976 4270 15056 4276
rect 15108 4276 15160 4282
rect 14924 4218 14976 4224
rect 15108 4218 15160 4224
rect 14936 4146 15148 4162
rect 14924 4140 15148 4146
rect 14976 4134 15148 4140
rect 14924 4082 14976 4088
rect 15016 4072 15068 4078
rect 15016 4014 15068 4020
rect 14924 4004 14976 4010
rect 14924 3946 14976 3952
rect 14832 2508 14884 2514
rect 14832 2450 14884 2456
rect 14648 2032 14700 2038
rect 14936 2009 14964 3946
rect 15028 3670 15056 4014
rect 15016 3664 15068 3670
rect 15016 3606 15068 3612
rect 14648 1974 14700 1980
rect 14922 2000 14978 2009
rect 14922 1935 14978 1944
rect 15028 1850 15056 3606
rect 15120 2446 15148 4134
rect 15212 3670 15240 5510
rect 15304 5166 15332 5578
rect 15292 5160 15344 5166
rect 15292 5102 15344 5108
rect 15292 4752 15344 4758
rect 15292 4694 15344 4700
rect 15304 3738 15332 4694
rect 15396 4010 15424 6054
rect 15658 5944 15714 5953
rect 15658 5879 15714 5888
rect 15752 5908 15804 5914
rect 15672 5846 15700 5879
rect 15752 5850 15804 5856
rect 15660 5840 15712 5846
rect 15660 5782 15712 5788
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 15488 5370 15516 5714
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 15476 5364 15528 5370
rect 15476 5306 15528 5312
rect 15580 4078 15608 5646
rect 15764 4690 15792 5850
rect 15856 4826 15884 7142
rect 15844 4820 15896 4826
rect 15844 4762 15896 4768
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 16488 4684 16540 4690
rect 16488 4626 16540 4632
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 15384 4004 15436 4010
rect 15384 3946 15436 3952
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 15200 3664 15252 3670
rect 15200 3606 15252 3612
rect 15212 2774 15240 3606
rect 15476 2916 15528 2922
rect 15476 2858 15528 2864
rect 15212 2746 15332 2774
rect 15108 2440 15160 2446
rect 15108 2382 15160 2388
rect 14844 1822 15056 1850
rect 14844 800 14872 1822
rect 15304 800 15332 2746
rect 15488 2514 15516 2858
rect 15580 2774 15608 4014
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 15580 2746 15700 2774
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 15672 800 15700 2746
rect 16132 800 16160 3878
rect 16500 800 16528 4626
rect 16948 2304 17000 2310
rect 16948 2246 17000 2252
rect 16960 800 16988 2246
rect 2778 504 2834 513
rect 2778 439 2834 448
rect 3054 0 3110 800
rect 3514 0 3570 800
rect 3974 0 4030 800
rect 4342 0 4398 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5630 0 5686 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7286 0 7342 800
rect 7746 0 7802 800
rect 8114 0 8170 800
rect 8574 0 8630 800
rect 8942 0 8998 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10230 0 10286 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11518 0 11574 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 13174 0 13230 800
rect 13542 0 13598 800
rect 14002 0 14058 800
rect 14462 0 14518 800
rect 14830 0 14886 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 16486 0 16542 800
rect 16946 0 17002 800
<< via2 >>
rect 2962 19488 3018 19544
rect 1858 17584 1914 17640
rect 1398 16668 1400 16688
rect 1400 16668 1452 16688
rect 1452 16668 1454 16688
rect 1398 16632 1454 16668
rect 1490 15700 1546 15736
rect 1490 15680 1492 15700
rect 1492 15680 1544 15700
rect 1544 15680 1546 15700
rect 1490 14764 1492 14784
rect 1492 14764 1544 14784
rect 1544 14764 1546 14784
rect 1490 14728 1546 14764
rect 2502 17040 2558 17096
rect 2134 15680 2190 15736
rect 1950 13912 2006 13968
rect 1398 13812 1400 13832
rect 1400 13812 1452 13832
rect 1452 13812 1454 13832
rect 1398 13776 1454 13812
rect 1398 12860 1400 12880
rect 1400 12860 1452 12880
rect 1452 12860 1454 12880
rect 1398 12824 1454 12860
rect 1490 11872 1546 11928
rect 1398 10920 1454 10976
rect 1398 9988 1454 10024
rect 1398 9968 1400 9988
rect 1400 9968 1452 9988
rect 1452 9968 1454 9988
rect 1398 9052 1400 9072
rect 1400 9052 1452 9072
rect 1452 9052 1454 9072
rect 1398 9016 1454 9052
rect 1490 8084 1546 8120
rect 1490 8064 1492 8084
rect 1492 8064 1544 8084
rect 1544 8064 1546 8084
rect 3146 18536 3202 18592
rect 2962 15988 2964 16008
rect 2964 15988 3016 16008
rect 3016 15988 3018 16008
rect 2962 15952 3018 15988
rect 3454 17434 3510 17436
rect 3534 17434 3590 17436
rect 3614 17434 3670 17436
rect 3694 17434 3750 17436
rect 3454 17382 3480 17434
rect 3480 17382 3510 17434
rect 3534 17382 3544 17434
rect 3544 17382 3590 17434
rect 3614 17382 3660 17434
rect 3660 17382 3670 17434
rect 3694 17382 3724 17434
rect 3724 17382 3750 17434
rect 3454 17380 3510 17382
rect 3534 17380 3590 17382
rect 3614 17380 3670 17382
rect 3694 17380 3750 17382
rect 3454 16346 3510 16348
rect 3534 16346 3590 16348
rect 3614 16346 3670 16348
rect 3694 16346 3750 16348
rect 3454 16294 3480 16346
rect 3480 16294 3510 16346
rect 3534 16294 3544 16346
rect 3544 16294 3590 16346
rect 3614 16294 3660 16346
rect 3660 16294 3670 16346
rect 3694 16294 3724 16346
rect 3724 16294 3750 16346
rect 3454 16292 3510 16294
rect 3534 16292 3590 16294
rect 3614 16292 3670 16294
rect 3694 16292 3750 16294
rect 2778 15408 2834 15464
rect 2778 14728 2834 14784
rect 3146 14864 3202 14920
rect 1490 7148 1492 7168
rect 1492 7148 1544 7168
rect 1544 7148 1546 7168
rect 1490 7112 1546 7148
rect 1490 6160 1546 6216
rect 1398 5244 1400 5264
rect 1400 5244 1452 5264
rect 1452 5244 1454 5264
rect 1398 5208 1454 5244
rect 1398 4256 1454 4312
rect 1490 3340 1492 3360
rect 1492 3340 1544 3360
rect 1544 3340 1546 3360
rect 1490 3304 1546 3340
rect 2226 4664 2282 4720
rect 1674 2896 1730 2952
rect 3330 15544 3386 15600
rect 3454 15258 3510 15260
rect 3534 15258 3590 15260
rect 3614 15258 3670 15260
rect 3694 15258 3750 15260
rect 3454 15206 3480 15258
rect 3480 15206 3510 15258
rect 3534 15206 3544 15258
rect 3544 15206 3590 15258
rect 3614 15206 3660 15258
rect 3660 15206 3670 15258
rect 3694 15206 3724 15258
rect 3724 15206 3750 15258
rect 3454 15204 3510 15206
rect 3534 15204 3590 15206
rect 3614 15204 3670 15206
rect 3694 15204 3750 15206
rect 3454 14170 3510 14172
rect 3534 14170 3590 14172
rect 3614 14170 3670 14172
rect 3694 14170 3750 14172
rect 3454 14118 3480 14170
rect 3480 14118 3510 14170
rect 3534 14118 3544 14170
rect 3544 14118 3590 14170
rect 3614 14118 3660 14170
rect 3660 14118 3670 14170
rect 3694 14118 3724 14170
rect 3724 14118 3750 14170
rect 3454 14116 3510 14118
rect 3534 14116 3590 14118
rect 3614 14116 3670 14118
rect 3694 14116 3750 14118
rect 4250 15952 4306 16008
rect 4066 15000 4122 15056
rect 3454 13082 3510 13084
rect 3534 13082 3590 13084
rect 3614 13082 3670 13084
rect 3694 13082 3750 13084
rect 3454 13030 3480 13082
rect 3480 13030 3510 13082
rect 3534 13030 3544 13082
rect 3544 13030 3590 13082
rect 3614 13030 3660 13082
rect 3660 13030 3670 13082
rect 3694 13030 3724 13082
rect 3724 13030 3750 13082
rect 3454 13028 3510 13030
rect 3534 13028 3590 13030
rect 3614 13028 3670 13030
rect 3694 13028 3750 13030
rect 3454 11994 3510 11996
rect 3534 11994 3590 11996
rect 3614 11994 3670 11996
rect 3694 11994 3750 11996
rect 3454 11942 3480 11994
rect 3480 11942 3510 11994
rect 3534 11942 3544 11994
rect 3544 11942 3590 11994
rect 3614 11942 3660 11994
rect 3660 11942 3670 11994
rect 3694 11942 3724 11994
rect 3724 11942 3750 11994
rect 3454 11940 3510 11942
rect 3534 11940 3590 11942
rect 3614 11940 3670 11942
rect 3694 11940 3750 11942
rect 4526 14728 4582 14784
rect 4066 11872 4122 11928
rect 3454 10906 3510 10908
rect 3534 10906 3590 10908
rect 3614 10906 3670 10908
rect 3694 10906 3750 10908
rect 3454 10854 3480 10906
rect 3480 10854 3510 10906
rect 3534 10854 3544 10906
rect 3544 10854 3590 10906
rect 3614 10854 3660 10906
rect 3660 10854 3670 10906
rect 3694 10854 3724 10906
rect 3724 10854 3750 10906
rect 3454 10852 3510 10854
rect 3534 10852 3590 10854
rect 3614 10852 3670 10854
rect 3694 10852 3750 10854
rect 3454 9818 3510 9820
rect 3534 9818 3590 9820
rect 3614 9818 3670 9820
rect 3694 9818 3750 9820
rect 3454 9766 3480 9818
rect 3480 9766 3510 9818
rect 3534 9766 3544 9818
rect 3544 9766 3590 9818
rect 3614 9766 3660 9818
rect 3660 9766 3670 9818
rect 3694 9766 3724 9818
rect 3724 9766 3750 9818
rect 3454 9764 3510 9766
rect 3534 9764 3590 9766
rect 3614 9764 3670 9766
rect 3694 9764 3750 9766
rect 3454 8730 3510 8732
rect 3534 8730 3590 8732
rect 3614 8730 3670 8732
rect 3694 8730 3750 8732
rect 3454 8678 3480 8730
rect 3480 8678 3510 8730
rect 3534 8678 3544 8730
rect 3544 8678 3590 8730
rect 3614 8678 3660 8730
rect 3660 8678 3670 8730
rect 3694 8678 3724 8730
rect 3724 8678 3750 8730
rect 3454 8676 3510 8678
rect 3534 8676 3590 8678
rect 3614 8676 3670 8678
rect 3694 8676 3750 8678
rect 3454 7642 3510 7644
rect 3534 7642 3590 7644
rect 3614 7642 3670 7644
rect 3694 7642 3750 7644
rect 3454 7590 3480 7642
rect 3480 7590 3510 7642
rect 3534 7590 3544 7642
rect 3544 7590 3590 7642
rect 3614 7590 3660 7642
rect 3660 7590 3670 7642
rect 3694 7590 3724 7642
rect 3724 7590 3750 7642
rect 3454 7588 3510 7590
rect 3534 7588 3590 7590
rect 3614 7588 3670 7590
rect 3694 7588 3750 7590
rect 3454 6554 3510 6556
rect 3534 6554 3590 6556
rect 3614 6554 3670 6556
rect 3694 6554 3750 6556
rect 3454 6502 3480 6554
rect 3480 6502 3510 6554
rect 3534 6502 3544 6554
rect 3544 6502 3590 6554
rect 3614 6502 3660 6554
rect 3660 6502 3670 6554
rect 3694 6502 3724 6554
rect 3724 6502 3750 6554
rect 3454 6500 3510 6502
rect 3534 6500 3590 6502
rect 3614 6500 3670 6502
rect 3694 6500 3750 6502
rect 3454 5466 3510 5468
rect 3534 5466 3590 5468
rect 3614 5466 3670 5468
rect 3694 5466 3750 5468
rect 3454 5414 3480 5466
rect 3480 5414 3510 5466
rect 3534 5414 3544 5466
rect 3544 5414 3590 5466
rect 3614 5414 3660 5466
rect 3660 5414 3670 5466
rect 3694 5414 3724 5466
rect 3724 5414 3750 5466
rect 3454 5412 3510 5414
rect 3534 5412 3590 5414
rect 3614 5412 3670 5414
rect 3694 5412 3750 5414
rect 3698 4528 3754 4584
rect 3454 4378 3510 4380
rect 3534 4378 3590 4380
rect 3614 4378 3670 4380
rect 3694 4378 3750 4380
rect 3454 4326 3480 4378
rect 3480 4326 3510 4378
rect 3534 4326 3544 4378
rect 3544 4326 3590 4378
rect 3614 4326 3660 4378
rect 3660 4326 3670 4378
rect 3694 4326 3724 4378
rect 3724 4326 3750 4378
rect 3454 4324 3510 4326
rect 3534 4324 3590 4326
rect 3614 4324 3670 4326
rect 3694 4324 3750 4326
rect 4250 4800 4306 4856
rect 3454 3290 3510 3292
rect 3534 3290 3590 3292
rect 3614 3290 3670 3292
rect 3694 3290 3750 3292
rect 3454 3238 3480 3290
rect 3480 3238 3510 3290
rect 3534 3238 3544 3290
rect 3544 3238 3590 3290
rect 3614 3238 3660 3290
rect 3660 3238 3670 3290
rect 3694 3238 3724 3290
rect 3724 3238 3750 3290
rect 3454 3236 3510 3238
rect 3534 3236 3590 3238
rect 3614 3236 3670 3238
rect 3694 3236 3750 3238
rect 3454 2202 3510 2204
rect 3534 2202 3590 2204
rect 3614 2202 3670 2204
rect 3694 2202 3750 2204
rect 3454 2150 3480 2202
rect 3480 2150 3510 2202
rect 3534 2150 3544 2202
rect 3544 2150 3590 2202
rect 3614 2150 3660 2202
rect 3660 2150 3670 2202
rect 3694 2150 3724 2202
rect 3724 2150 3750 2202
rect 3454 2148 3510 2150
rect 3534 2148 3590 2150
rect 3614 2148 3670 2150
rect 3694 2148 3750 2150
rect 3606 1400 3662 1456
rect 5953 16890 6009 16892
rect 6033 16890 6089 16892
rect 6113 16890 6169 16892
rect 6193 16890 6249 16892
rect 5953 16838 5979 16890
rect 5979 16838 6009 16890
rect 6033 16838 6043 16890
rect 6043 16838 6089 16890
rect 6113 16838 6159 16890
rect 6159 16838 6169 16890
rect 6193 16838 6223 16890
rect 6223 16838 6249 16890
rect 5953 16836 6009 16838
rect 6033 16836 6089 16838
rect 6113 16836 6169 16838
rect 6193 16836 6249 16838
rect 5953 15802 6009 15804
rect 6033 15802 6089 15804
rect 6113 15802 6169 15804
rect 6193 15802 6249 15804
rect 5953 15750 5979 15802
rect 5979 15750 6009 15802
rect 6033 15750 6043 15802
rect 6043 15750 6089 15802
rect 6113 15750 6159 15802
rect 6159 15750 6169 15802
rect 6193 15750 6223 15802
rect 6223 15750 6249 15802
rect 5953 15748 6009 15750
rect 6033 15748 6089 15750
rect 6113 15748 6169 15750
rect 6193 15748 6249 15750
rect 5814 15680 5870 15736
rect 5953 14714 6009 14716
rect 6033 14714 6089 14716
rect 6113 14714 6169 14716
rect 6193 14714 6249 14716
rect 5953 14662 5979 14714
rect 5979 14662 6009 14714
rect 6033 14662 6043 14714
rect 6043 14662 6089 14714
rect 6113 14662 6159 14714
rect 6159 14662 6169 14714
rect 6193 14662 6223 14714
rect 6223 14662 6249 14714
rect 5953 14660 6009 14662
rect 6033 14660 6089 14662
rect 6113 14660 6169 14662
rect 6193 14660 6249 14662
rect 5953 13626 6009 13628
rect 6033 13626 6089 13628
rect 6113 13626 6169 13628
rect 6193 13626 6249 13628
rect 5953 13574 5979 13626
rect 5979 13574 6009 13626
rect 6033 13574 6043 13626
rect 6043 13574 6089 13626
rect 6113 13574 6159 13626
rect 6159 13574 6169 13626
rect 6193 13574 6223 13626
rect 6223 13574 6249 13626
rect 5953 13572 6009 13574
rect 6033 13572 6089 13574
rect 6113 13572 6169 13574
rect 6193 13572 6249 13574
rect 5814 13388 5870 13424
rect 5814 13368 5816 13388
rect 5816 13368 5868 13388
rect 5868 13368 5870 13388
rect 6642 14884 6698 14920
rect 6642 14864 6644 14884
rect 6644 14864 6696 14884
rect 6696 14864 6698 14884
rect 5998 12960 6054 13016
rect 5814 12724 5816 12744
rect 5816 12724 5868 12744
rect 5868 12724 5870 12744
rect 5814 12688 5870 12724
rect 5953 12538 6009 12540
rect 6033 12538 6089 12540
rect 6113 12538 6169 12540
rect 6193 12538 6249 12540
rect 5953 12486 5979 12538
rect 5979 12486 6009 12538
rect 6033 12486 6043 12538
rect 6043 12486 6089 12538
rect 6113 12486 6159 12538
rect 6159 12486 6169 12538
rect 6193 12486 6223 12538
rect 6223 12486 6249 12538
rect 5953 12484 6009 12486
rect 6033 12484 6089 12486
rect 6113 12484 6169 12486
rect 6193 12484 6249 12486
rect 5722 12416 5778 12472
rect 6366 12824 6422 12880
rect 6642 14320 6698 14376
rect 6642 12688 6698 12744
rect 5814 12008 5870 12064
rect 5953 11450 6009 11452
rect 6033 11450 6089 11452
rect 6113 11450 6169 11452
rect 6193 11450 6249 11452
rect 5953 11398 5979 11450
rect 5979 11398 6009 11450
rect 6033 11398 6043 11450
rect 6043 11398 6089 11450
rect 6113 11398 6159 11450
rect 6159 11398 6169 11450
rect 6193 11398 6223 11450
rect 6223 11398 6249 11450
rect 5953 11396 6009 11398
rect 6033 11396 6089 11398
rect 6113 11396 6169 11398
rect 6193 11396 6249 11398
rect 6366 12008 6422 12064
rect 6366 11872 6422 11928
rect 5953 10362 6009 10364
rect 6033 10362 6089 10364
rect 6113 10362 6169 10364
rect 6193 10362 6249 10364
rect 5953 10310 5979 10362
rect 5979 10310 6009 10362
rect 6033 10310 6043 10362
rect 6043 10310 6089 10362
rect 6113 10310 6159 10362
rect 6159 10310 6169 10362
rect 6193 10310 6223 10362
rect 6223 10310 6249 10362
rect 5953 10308 6009 10310
rect 6033 10308 6089 10310
rect 6113 10308 6169 10310
rect 6193 10308 6249 10310
rect 4986 9324 4988 9344
rect 4988 9324 5040 9344
rect 5040 9324 5042 9344
rect 4986 9288 5042 9324
rect 5078 7792 5134 7848
rect 4066 2508 4122 2544
rect 4066 2488 4068 2508
rect 4068 2488 4120 2508
rect 4120 2488 4122 2508
rect 5814 9324 5816 9344
rect 5816 9324 5868 9344
rect 5868 9324 5870 9344
rect 5814 9288 5870 9324
rect 5953 9274 6009 9276
rect 6033 9274 6089 9276
rect 6113 9274 6169 9276
rect 6193 9274 6249 9276
rect 5953 9222 5979 9274
rect 5979 9222 6009 9274
rect 6033 9222 6043 9274
rect 6043 9222 6089 9274
rect 6113 9222 6159 9274
rect 6159 9222 6169 9274
rect 6193 9222 6223 9274
rect 6223 9222 6249 9274
rect 5953 9220 6009 9222
rect 6033 9220 6089 9222
rect 6113 9220 6169 9222
rect 6193 9220 6249 9222
rect 5538 7284 5540 7304
rect 5540 7284 5592 7304
rect 5592 7284 5594 7304
rect 5538 7248 5594 7284
rect 4066 2352 4122 2408
rect 5953 8186 6009 8188
rect 6033 8186 6089 8188
rect 6113 8186 6169 8188
rect 6193 8186 6249 8188
rect 5953 8134 5979 8186
rect 5979 8134 6009 8186
rect 6033 8134 6043 8186
rect 6043 8134 6089 8186
rect 6113 8134 6159 8186
rect 6159 8134 6169 8186
rect 6193 8134 6223 8186
rect 6223 8134 6249 8186
rect 5953 8132 6009 8134
rect 6033 8132 6089 8134
rect 6113 8132 6169 8134
rect 6193 8132 6249 8134
rect 5630 5072 5686 5128
rect 5953 7098 6009 7100
rect 6033 7098 6089 7100
rect 6113 7098 6169 7100
rect 6193 7098 6249 7100
rect 5953 7046 5979 7098
rect 5979 7046 6009 7098
rect 6033 7046 6043 7098
rect 6043 7046 6089 7098
rect 6113 7046 6159 7098
rect 6159 7046 6169 7098
rect 6193 7046 6223 7098
rect 6223 7046 6249 7098
rect 5953 7044 6009 7046
rect 6033 7044 6089 7046
rect 6113 7044 6169 7046
rect 6193 7044 6249 7046
rect 5953 6010 6009 6012
rect 6033 6010 6089 6012
rect 6113 6010 6169 6012
rect 6193 6010 6249 6012
rect 5953 5958 5979 6010
rect 5979 5958 6009 6010
rect 6033 5958 6043 6010
rect 6043 5958 6089 6010
rect 6113 5958 6159 6010
rect 6159 5958 6169 6010
rect 6193 5958 6223 6010
rect 6223 5958 6249 6010
rect 5953 5956 6009 5958
rect 6033 5956 6089 5958
rect 6113 5956 6169 5958
rect 6193 5956 6249 5958
rect 6182 5344 6238 5400
rect 6918 13368 6974 13424
rect 7378 12960 7434 13016
rect 6826 7928 6882 7984
rect 7102 8084 7158 8120
rect 7102 8064 7104 8084
rect 7104 8064 7156 8084
rect 7156 8064 7158 8084
rect 7286 7928 7342 7984
rect 6734 6568 6790 6624
rect 6550 5364 6606 5400
rect 6550 5344 6552 5364
rect 6552 5344 6604 5364
rect 6604 5344 6606 5364
rect 5953 4922 6009 4924
rect 6033 4922 6089 4924
rect 6113 4922 6169 4924
rect 6193 4922 6249 4924
rect 5953 4870 5979 4922
rect 5979 4870 6009 4922
rect 6033 4870 6043 4922
rect 6043 4870 6089 4922
rect 6113 4870 6159 4922
rect 6159 4870 6169 4922
rect 6193 4870 6223 4922
rect 6223 4870 6249 4922
rect 5953 4868 6009 4870
rect 6033 4868 6089 4870
rect 6113 4868 6169 4870
rect 6193 4868 6249 4870
rect 5446 2760 5502 2816
rect 5953 3834 6009 3836
rect 6033 3834 6089 3836
rect 6113 3834 6169 3836
rect 6193 3834 6249 3836
rect 5953 3782 5979 3834
rect 5979 3782 6009 3834
rect 6033 3782 6043 3834
rect 6043 3782 6089 3834
rect 6113 3782 6159 3834
rect 6159 3782 6169 3834
rect 6193 3782 6223 3834
rect 6223 3782 6249 3834
rect 5953 3780 6009 3782
rect 6033 3780 6089 3782
rect 6113 3780 6169 3782
rect 6193 3780 6249 3782
rect 6274 3032 6330 3088
rect 5814 2760 5870 2816
rect 5953 2746 6009 2748
rect 6033 2746 6089 2748
rect 6113 2746 6169 2748
rect 6193 2746 6249 2748
rect 5953 2694 5979 2746
rect 5979 2694 6009 2746
rect 6033 2694 6043 2746
rect 6043 2694 6089 2746
rect 6113 2694 6159 2746
rect 6159 2694 6169 2746
rect 6193 2694 6223 2746
rect 6223 2694 6249 2746
rect 5953 2692 6009 2694
rect 6033 2692 6089 2694
rect 6113 2692 6169 2694
rect 6193 2692 6249 2694
rect 6642 3712 6698 3768
rect 7194 5208 7250 5264
rect 8452 17434 8508 17436
rect 8532 17434 8588 17436
rect 8612 17434 8668 17436
rect 8692 17434 8748 17436
rect 8452 17382 8478 17434
rect 8478 17382 8508 17434
rect 8532 17382 8542 17434
rect 8542 17382 8588 17434
rect 8612 17382 8658 17434
rect 8658 17382 8668 17434
rect 8692 17382 8722 17434
rect 8722 17382 8748 17434
rect 8452 17380 8508 17382
rect 8532 17380 8588 17382
rect 8612 17380 8668 17382
rect 8692 17380 8748 17382
rect 8452 16346 8508 16348
rect 8532 16346 8588 16348
rect 8612 16346 8668 16348
rect 8692 16346 8748 16348
rect 8452 16294 8478 16346
rect 8478 16294 8508 16346
rect 8532 16294 8542 16346
rect 8542 16294 8588 16346
rect 8612 16294 8658 16346
rect 8658 16294 8668 16346
rect 8692 16294 8722 16346
rect 8722 16294 8748 16346
rect 8452 16292 8508 16294
rect 8532 16292 8588 16294
rect 8612 16292 8668 16294
rect 8692 16292 8748 16294
rect 8452 15258 8508 15260
rect 8532 15258 8588 15260
rect 8612 15258 8668 15260
rect 8692 15258 8748 15260
rect 8452 15206 8478 15258
rect 8478 15206 8508 15258
rect 8532 15206 8542 15258
rect 8542 15206 8588 15258
rect 8612 15206 8658 15258
rect 8658 15206 8668 15258
rect 8692 15206 8722 15258
rect 8722 15206 8748 15258
rect 8452 15204 8508 15206
rect 8532 15204 8588 15206
rect 8612 15204 8668 15206
rect 8692 15204 8748 15206
rect 8022 14356 8024 14376
rect 8024 14356 8076 14376
rect 8076 14356 8078 14376
rect 8022 14320 8078 14356
rect 8452 14170 8508 14172
rect 8532 14170 8588 14172
rect 8612 14170 8668 14172
rect 8692 14170 8748 14172
rect 8452 14118 8478 14170
rect 8478 14118 8508 14170
rect 8532 14118 8542 14170
rect 8542 14118 8588 14170
rect 8612 14118 8658 14170
rect 8658 14118 8668 14170
rect 8692 14118 8722 14170
rect 8722 14118 8748 14170
rect 8452 14116 8508 14118
rect 8532 14116 8588 14118
rect 8612 14116 8668 14118
rect 8692 14116 8748 14118
rect 9126 13912 9182 13968
rect 9310 15000 9366 15056
rect 9586 15036 9588 15056
rect 9588 15036 9640 15056
rect 9640 15036 9642 15056
rect 9586 15000 9642 15036
rect 8206 13404 8208 13424
rect 8208 13404 8260 13424
rect 8260 13404 8262 13424
rect 8206 13368 8262 13404
rect 8452 13082 8508 13084
rect 8532 13082 8588 13084
rect 8612 13082 8668 13084
rect 8692 13082 8748 13084
rect 8452 13030 8478 13082
rect 8478 13030 8508 13082
rect 8532 13030 8542 13082
rect 8542 13030 8588 13082
rect 8612 13030 8658 13082
rect 8658 13030 8668 13082
rect 8692 13030 8722 13082
rect 8722 13030 8748 13082
rect 8452 13028 8508 13030
rect 8532 13028 8588 13030
rect 8612 13028 8668 13030
rect 8692 13028 8748 13030
rect 8452 11994 8508 11996
rect 8532 11994 8588 11996
rect 8612 11994 8668 11996
rect 8692 11994 8748 11996
rect 8452 11942 8478 11994
rect 8478 11942 8508 11994
rect 8532 11942 8542 11994
rect 8542 11942 8588 11994
rect 8612 11942 8658 11994
rect 8658 11942 8668 11994
rect 8692 11942 8722 11994
rect 8722 11942 8748 11994
rect 8452 11940 8508 11942
rect 8532 11940 8588 11942
rect 8612 11940 8668 11942
rect 8692 11940 8748 11942
rect 7838 10104 7894 10160
rect 7654 7248 7710 7304
rect 8452 10906 8508 10908
rect 8532 10906 8588 10908
rect 8612 10906 8668 10908
rect 8692 10906 8748 10908
rect 8452 10854 8478 10906
rect 8478 10854 8508 10906
rect 8532 10854 8542 10906
rect 8542 10854 8588 10906
rect 8612 10854 8658 10906
rect 8658 10854 8668 10906
rect 8692 10854 8722 10906
rect 8722 10854 8748 10906
rect 8452 10852 8508 10854
rect 8532 10852 8588 10854
rect 8612 10852 8668 10854
rect 8692 10852 8748 10854
rect 8114 10104 8170 10160
rect 8452 9818 8508 9820
rect 8532 9818 8588 9820
rect 8612 9818 8668 9820
rect 8692 9818 8748 9820
rect 8452 9766 8478 9818
rect 8478 9766 8508 9818
rect 8532 9766 8542 9818
rect 8542 9766 8588 9818
rect 8612 9766 8658 9818
rect 8658 9766 8668 9818
rect 8692 9766 8722 9818
rect 8722 9766 8748 9818
rect 8452 9764 8508 9766
rect 8532 9764 8588 9766
rect 8612 9764 8668 9766
rect 8692 9764 8748 9766
rect 8758 8916 8760 8936
rect 8760 8916 8812 8936
rect 8812 8916 8814 8936
rect 8758 8880 8814 8916
rect 8452 8730 8508 8732
rect 8532 8730 8588 8732
rect 8612 8730 8668 8732
rect 8692 8730 8748 8732
rect 8452 8678 8478 8730
rect 8478 8678 8508 8730
rect 8532 8678 8542 8730
rect 8542 8678 8588 8730
rect 8612 8678 8658 8730
rect 8658 8678 8668 8730
rect 8692 8678 8722 8730
rect 8722 8678 8748 8730
rect 8452 8676 8508 8678
rect 8532 8676 8588 8678
rect 8612 8676 8668 8678
rect 8692 8676 8748 8678
rect 8390 7812 8446 7848
rect 8390 7792 8392 7812
rect 8392 7792 8444 7812
rect 8444 7792 8446 7812
rect 8850 7792 8906 7848
rect 8452 7642 8508 7644
rect 8532 7642 8588 7644
rect 8612 7642 8668 7644
rect 8692 7642 8748 7644
rect 8452 7590 8478 7642
rect 8478 7590 8508 7642
rect 8532 7590 8542 7642
rect 8542 7590 8588 7642
rect 8612 7590 8658 7642
rect 8658 7590 8668 7642
rect 8692 7590 8722 7642
rect 8722 7590 8748 7642
rect 8452 7588 8508 7590
rect 8532 7588 8588 7590
rect 8612 7588 8668 7590
rect 8692 7588 8748 7590
rect 8942 7112 8998 7168
rect 8452 6554 8508 6556
rect 8532 6554 8588 6556
rect 8612 6554 8668 6556
rect 8692 6554 8748 6556
rect 8452 6502 8478 6554
rect 8478 6502 8508 6554
rect 8532 6502 8542 6554
rect 8542 6502 8588 6554
rect 8612 6502 8658 6554
rect 8658 6502 8668 6554
rect 8692 6502 8722 6554
rect 8722 6502 8748 6554
rect 8452 6500 8508 6502
rect 8532 6500 8588 6502
rect 8612 6500 8668 6502
rect 8692 6500 8748 6502
rect 9218 7948 9274 7984
rect 9218 7928 9220 7948
rect 9220 7928 9272 7948
rect 9272 7928 9274 7948
rect 9862 15272 9918 15328
rect 9954 14864 10010 14920
rect 10138 15136 10194 15192
rect 11058 17040 11114 17096
rect 10950 16890 11006 16892
rect 11030 16890 11086 16892
rect 11110 16890 11166 16892
rect 11190 16890 11246 16892
rect 10950 16838 10976 16890
rect 10976 16838 11006 16890
rect 11030 16838 11040 16890
rect 11040 16838 11086 16890
rect 11110 16838 11156 16890
rect 11156 16838 11166 16890
rect 11190 16838 11220 16890
rect 11220 16838 11246 16890
rect 10950 16836 11006 16838
rect 11030 16836 11086 16838
rect 11110 16836 11166 16838
rect 11190 16836 11246 16838
rect 10506 15136 10562 15192
rect 10138 14320 10194 14376
rect 10230 13776 10286 13832
rect 10230 12860 10232 12880
rect 10232 12860 10284 12880
rect 10284 12860 10286 12880
rect 10230 12824 10286 12860
rect 9678 11736 9734 11792
rect 9218 7656 9274 7712
rect 9218 7248 9274 7304
rect 9034 6296 9090 6352
rect 8452 5466 8508 5468
rect 8532 5466 8588 5468
rect 8612 5466 8668 5468
rect 8692 5466 8748 5468
rect 8452 5414 8478 5466
rect 8478 5414 8508 5466
rect 8532 5414 8542 5466
rect 8542 5414 8588 5466
rect 8612 5414 8658 5466
rect 8658 5414 8668 5466
rect 8692 5414 8722 5466
rect 8722 5414 8748 5466
rect 8452 5412 8508 5414
rect 8532 5412 8588 5414
rect 8612 5412 8668 5414
rect 8692 5412 8748 5414
rect 8574 4684 8630 4720
rect 8574 4664 8576 4684
rect 8576 4664 8628 4684
rect 8628 4664 8630 4684
rect 8666 4564 8668 4584
rect 8668 4564 8720 4584
rect 8720 4564 8722 4584
rect 8666 4528 8722 4564
rect 8114 4120 8170 4176
rect 8452 4378 8508 4380
rect 8532 4378 8588 4380
rect 8612 4378 8668 4380
rect 8692 4378 8748 4380
rect 8452 4326 8478 4378
rect 8478 4326 8508 4378
rect 8532 4326 8542 4378
rect 8542 4326 8588 4378
rect 8612 4326 8658 4378
rect 8658 4326 8668 4378
rect 8692 4326 8722 4378
rect 8722 4326 8748 4378
rect 8452 4324 8508 4326
rect 8532 4324 8588 4326
rect 8612 4324 8668 4326
rect 8692 4324 8748 4326
rect 8452 3290 8508 3292
rect 8532 3290 8588 3292
rect 8612 3290 8668 3292
rect 8692 3290 8748 3292
rect 8452 3238 8478 3290
rect 8478 3238 8508 3290
rect 8532 3238 8542 3290
rect 8542 3238 8588 3290
rect 8612 3238 8658 3290
rect 8658 3238 8668 3290
rect 8692 3238 8722 3290
rect 8722 3238 8748 3290
rect 8452 3236 8508 3238
rect 8532 3236 8588 3238
rect 8612 3236 8668 3238
rect 8692 3236 8748 3238
rect 8942 3032 8998 3088
rect 10230 11756 10286 11792
rect 10230 11736 10232 11756
rect 10232 11736 10284 11756
rect 10284 11736 10286 11756
rect 10598 14864 10654 14920
rect 10506 13096 10562 13152
rect 10950 15802 11006 15804
rect 11030 15802 11086 15804
rect 11110 15802 11166 15804
rect 11190 15802 11246 15804
rect 10950 15750 10976 15802
rect 10976 15750 11006 15802
rect 11030 15750 11040 15802
rect 11040 15750 11086 15802
rect 11110 15750 11156 15802
rect 11156 15750 11166 15802
rect 11190 15750 11220 15802
rect 11220 15750 11246 15802
rect 10950 15748 11006 15750
rect 11030 15748 11086 15750
rect 11110 15748 11166 15750
rect 11190 15748 11246 15750
rect 11518 15680 11574 15736
rect 11518 15272 11574 15328
rect 10950 14714 11006 14716
rect 11030 14714 11086 14716
rect 11110 14714 11166 14716
rect 11190 14714 11246 14716
rect 10950 14662 10976 14714
rect 10976 14662 11006 14714
rect 11030 14662 11040 14714
rect 11040 14662 11086 14714
rect 11110 14662 11156 14714
rect 11156 14662 11166 14714
rect 11190 14662 11220 14714
rect 11220 14662 11246 14714
rect 10950 14660 11006 14662
rect 11030 14660 11086 14662
rect 11110 14660 11166 14662
rect 11190 14660 11246 14662
rect 9586 7112 9642 7168
rect 9586 6332 9588 6352
rect 9588 6332 9640 6352
rect 9640 6332 9642 6352
rect 9586 6296 9642 6332
rect 9218 5480 9274 5536
rect 9770 5888 9826 5944
rect 9678 5480 9734 5536
rect 9586 5208 9642 5264
rect 9770 5344 9826 5400
rect 9770 5208 9826 5264
rect 9402 5072 9458 5128
rect 9310 4528 9366 4584
rect 9218 2896 9274 2952
rect 8452 2202 8508 2204
rect 8532 2202 8588 2204
rect 8612 2202 8668 2204
rect 8692 2202 8748 2204
rect 8452 2150 8478 2202
rect 8478 2150 8508 2202
rect 8532 2150 8542 2202
rect 8542 2150 8588 2202
rect 8612 2150 8658 2202
rect 8658 2150 8668 2202
rect 8692 2150 8722 2202
rect 8722 2150 8748 2202
rect 8452 2148 8508 2150
rect 8532 2148 8588 2150
rect 8612 2148 8668 2150
rect 8692 2148 8748 2150
rect 9402 3712 9458 3768
rect 10322 8064 10378 8120
rect 10690 6876 10692 6896
rect 10692 6876 10744 6896
rect 10744 6876 10746 6896
rect 10690 6840 10746 6876
rect 10138 6060 10140 6080
rect 10140 6060 10192 6080
rect 10192 6060 10194 6080
rect 10138 6024 10194 6060
rect 10506 6024 10562 6080
rect 10506 4936 10562 4992
rect 9770 3168 9826 3224
rect 10690 4936 10746 4992
rect 10950 13626 11006 13628
rect 11030 13626 11086 13628
rect 11110 13626 11166 13628
rect 11190 13626 11246 13628
rect 10950 13574 10976 13626
rect 10976 13574 11006 13626
rect 11030 13574 11040 13626
rect 11040 13574 11086 13626
rect 11110 13574 11156 13626
rect 11156 13574 11166 13626
rect 11190 13574 11220 13626
rect 11220 13574 11246 13626
rect 10950 13572 11006 13574
rect 11030 13572 11086 13574
rect 11110 13572 11166 13574
rect 11190 13572 11246 13574
rect 11794 13776 11850 13832
rect 11794 13504 11850 13560
rect 10950 12538 11006 12540
rect 11030 12538 11086 12540
rect 11110 12538 11166 12540
rect 11190 12538 11246 12540
rect 10950 12486 10976 12538
rect 10976 12486 11006 12538
rect 11030 12486 11040 12538
rect 11040 12486 11086 12538
rect 11110 12486 11156 12538
rect 11156 12486 11166 12538
rect 11190 12486 11220 12538
rect 11220 12486 11246 12538
rect 10950 12484 11006 12486
rect 11030 12484 11086 12486
rect 11110 12484 11166 12486
rect 11190 12484 11246 12486
rect 11702 12688 11758 12744
rect 10950 11450 11006 11452
rect 11030 11450 11086 11452
rect 11110 11450 11166 11452
rect 11190 11450 11246 11452
rect 10950 11398 10976 11450
rect 10976 11398 11006 11450
rect 11030 11398 11040 11450
rect 11040 11398 11086 11450
rect 11110 11398 11156 11450
rect 11156 11398 11166 11450
rect 11190 11398 11220 11450
rect 11220 11398 11246 11450
rect 10950 11396 11006 11398
rect 11030 11396 11086 11398
rect 11110 11396 11166 11398
rect 11190 11396 11246 11398
rect 11058 11192 11114 11248
rect 10950 10362 11006 10364
rect 11030 10362 11086 10364
rect 11110 10362 11166 10364
rect 11190 10362 11246 10364
rect 10950 10310 10976 10362
rect 10976 10310 11006 10362
rect 11030 10310 11040 10362
rect 11040 10310 11086 10362
rect 11110 10310 11156 10362
rect 11156 10310 11166 10362
rect 11190 10310 11220 10362
rect 11220 10310 11246 10362
rect 10950 10308 11006 10310
rect 11030 10308 11086 10310
rect 11110 10308 11166 10310
rect 11190 10308 11246 10310
rect 10950 9274 11006 9276
rect 11030 9274 11086 9276
rect 11110 9274 11166 9276
rect 11190 9274 11246 9276
rect 10950 9222 10976 9274
rect 10976 9222 11006 9274
rect 11030 9222 11040 9274
rect 11040 9222 11086 9274
rect 11110 9222 11156 9274
rect 11156 9222 11166 9274
rect 11190 9222 11220 9274
rect 11220 9222 11246 9274
rect 10950 9220 11006 9222
rect 11030 9220 11086 9222
rect 11110 9220 11166 9222
rect 11190 9220 11246 9222
rect 10950 8186 11006 8188
rect 11030 8186 11086 8188
rect 11110 8186 11166 8188
rect 11190 8186 11246 8188
rect 10950 8134 10976 8186
rect 10976 8134 11006 8186
rect 11030 8134 11040 8186
rect 11040 8134 11086 8186
rect 11110 8134 11156 8186
rect 11156 8134 11166 8186
rect 11190 8134 11220 8186
rect 11220 8134 11246 8186
rect 10950 8132 11006 8134
rect 11030 8132 11086 8134
rect 11110 8132 11166 8134
rect 11190 8132 11246 8134
rect 10950 7098 11006 7100
rect 11030 7098 11086 7100
rect 11110 7098 11166 7100
rect 11190 7098 11246 7100
rect 10950 7046 10976 7098
rect 10976 7046 11006 7098
rect 11030 7046 11040 7098
rect 11040 7046 11086 7098
rect 11110 7046 11156 7098
rect 11156 7046 11166 7098
rect 11190 7046 11220 7098
rect 11220 7046 11246 7098
rect 10950 7044 11006 7046
rect 11030 7044 11086 7046
rect 11110 7044 11166 7046
rect 11190 7044 11246 7046
rect 11242 6704 11298 6760
rect 11610 7928 11666 7984
rect 11426 6604 11428 6624
rect 11428 6604 11480 6624
rect 11480 6604 11482 6624
rect 11426 6568 11482 6604
rect 10950 6010 11006 6012
rect 11030 6010 11086 6012
rect 11110 6010 11166 6012
rect 11190 6010 11246 6012
rect 10950 5958 10976 6010
rect 10976 5958 11006 6010
rect 11030 5958 11040 6010
rect 11040 5958 11086 6010
rect 11110 5958 11156 6010
rect 11156 5958 11166 6010
rect 11190 5958 11220 6010
rect 11220 5958 11246 6010
rect 10950 5956 11006 5958
rect 11030 5956 11086 5958
rect 11110 5956 11166 5958
rect 11190 5956 11246 5958
rect 12162 14476 12218 14512
rect 12162 14456 12164 14476
rect 12164 14456 12216 14476
rect 12216 14456 12218 14476
rect 12530 16088 12586 16144
rect 12438 14864 12494 14920
rect 13449 17434 13505 17436
rect 13529 17434 13585 17436
rect 13609 17434 13665 17436
rect 13689 17434 13745 17436
rect 13449 17382 13475 17434
rect 13475 17382 13505 17434
rect 13529 17382 13539 17434
rect 13539 17382 13585 17434
rect 13609 17382 13655 17434
rect 13655 17382 13665 17434
rect 13689 17382 13719 17434
rect 13719 17382 13745 17434
rect 13449 17380 13505 17382
rect 13529 17380 13585 17382
rect 13609 17380 13665 17382
rect 13689 17380 13745 17382
rect 13449 16346 13505 16348
rect 13529 16346 13585 16348
rect 13609 16346 13665 16348
rect 13689 16346 13745 16348
rect 13449 16294 13475 16346
rect 13475 16294 13505 16346
rect 13529 16294 13539 16346
rect 13539 16294 13585 16346
rect 13609 16294 13655 16346
rect 13655 16294 13665 16346
rect 13689 16294 13719 16346
rect 13719 16294 13745 16346
rect 13449 16292 13505 16294
rect 13529 16292 13585 16294
rect 13609 16292 13665 16294
rect 13689 16292 13745 16294
rect 12898 15000 12954 15056
rect 13174 15000 13230 15056
rect 13449 15258 13505 15260
rect 13529 15258 13585 15260
rect 13609 15258 13665 15260
rect 13689 15258 13745 15260
rect 13449 15206 13475 15258
rect 13475 15206 13505 15258
rect 13529 15206 13539 15258
rect 13539 15206 13585 15258
rect 13609 15206 13655 15258
rect 13655 15206 13665 15258
rect 13689 15206 13719 15258
rect 13719 15206 13745 15258
rect 13449 15204 13505 15206
rect 13529 15204 13585 15206
rect 13609 15204 13665 15206
rect 13689 15204 13745 15206
rect 12898 14864 12954 14920
rect 12438 13368 12494 13424
rect 12346 13096 12402 13152
rect 12254 12688 12310 12744
rect 11058 5480 11114 5536
rect 10950 4922 11006 4924
rect 11030 4922 11086 4924
rect 11110 4922 11166 4924
rect 11190 4922 11246 4924
rect 10950 4870 10976 4922
rect 10976 4870 11006 4922
rect 11030 4870 11040 4922
rect 11040 4870 11086 4922
rect 11110 4870 11156 4922
rect 11156 4870 11166 4922
rect 11190 4870 11220 4922
rect 11220 4870 11246 4922
rect 10950 4868 11006 4870
rect 11030 4868 11086 4870
rect 11110 4868 11166 4870
rect 11190 4868 11246 4870
rect 10414 3304 10470 3360
rect 10598 2896 10654 2952
rect 11702 5344 11758 5400
rect 11794 5208 11850 5264
rect 10950 3834 11006 3836
rect 11030 3834 11086 3836
rect 11110 3834 11166 3836
rect 11190 3834 11246 3836
rect 10950 3782 10976 3834
rect 10976 3782 11006 3834
rect 11030 3782 11040 3834
rect 11040 3782 11086 3834
rect 11110 3782 11156 3834
rect 11156 3782 11166 3834
rect 11190 3782 11220 3834
rect 11220 3782 11246 3834
rect 10950 3780 11006 3782
rect 11030 3780 11086 3782
rect 11110 3780 11166 3782
rect 11190 3780 11246 3782
rect 10950 2746 11006 2748
rect 11030 2746 11086 2748
rect 11110 2746 11166 2748
rect 11190 2746 11246 2748
rect 10950 2694 10976 2746
rect 10976 2694 11006 2746
rect 11030 2694 11040 2746
rect 11040 2694 11086 2746
rect 11110 2694 11156 2746
rect 11156 2694 11166 2746
rect 11190 2694 11220 2746
rect 11220 2694 11246 2746
rect 10950 2692 11006 2694
rect 11030 2692 11086 2694
rect 11110 2692 11166 2694
rect 11190 2692 11246 2694
rect 11426 3440 11482 3496
rect 11334 2488 11390 2544
rect 13449 14170 13505 14172
rect 13529 14170 13585 14172
rect 13609 14170 13665 14172
rect 13689 14170 13745 14172
rect 13449 14118 13475 14170
rect 13475 14118 13505 14170
rect 13529 14118 13539 14170
rect 13539 14118 13585 14170
rect 13609 14118 13655 14170
rect 13655 14118 13665 14170
rect 13689 14118 13719 14170
rect 13719 14118 13745 14170
rect 13449 14116 13505 14118
rect 13529 14116 13585 14118
rect 13609 14116 13665 14118
rect 13689 14116 13745 14118
rect 13726 13504 13782 13560
rect 12990 13096 13046 13152
rect 12898 12980 12954 13016
rect 12898 12960 12900 12980
rect 12900 12960 12952 12980
rect 12952 12960 12954 12980
rect 12438 7248 12494 7304
rect 12990 11192 13046 11248
rect 12346 6296 12402 6352
rect 11886 3848 11942 3904
rect 11886 3304 11942 3360
rect 11886 2896 11942 2952
rect 12622 6296 12678 6352
rect 12346 3848 12402 3904
rect 12346 3612 12348 3632
rect 12348 3612 12400 3632
rect 12400 3612 12402 3632
rect 12898 6704 12954 6760
rect 12622 4256 12678 4312
rect 12622 4120 12678 4176
rect 12346 3576 12402 3612
rect 12070 2896 12126 2952
rect 12622 2644 12678 2680
rect 12622 2624 12624 2644
rect 12624 2624 12676 2644
rect 12676 2624 12678 2644
rect 13449 13082 13505 13084
rect 13529 13082 13585 13084
rect 13609 13082 13665 13084
rect 13689 13082 13745 13084
rect 13449 13030 13475 13082
rect 13475 13030 13505 13082
rect 13529 13030 13539 13082
rect 13539 13030 13585 13082
rect 13609 13030 13655 13082
rect 13655 13030 13665 13082
rect 13689 13030 13719 13082
rect 13719 13030 13745 13082
rect 13449 13028 13505 13030
rect 13529 13028 13585 13030
rect 13609 13028 13665 13030
rect 13689 13028 13745 13030
rect 13449 11994 13505 11996
rect 13529 11994 13585 11996
rect 13609 11994 13665 11996
rect 13689 11994 13745 11996
rect 13449 11942 13475 11994
rect 13475 11942 13505 11994
rect 13529 11942 13539 11994
rect 13539 11942 13585 11994
rect 13609 11942 13655 11994
rect 13655 11942 13665 11994
rect 13689 11942 13719 11994
rect 13719 11942 13745 11994
rect 13449 11940 13505 11942
rect 13529 11940 13585 11942
rect 13609 11940 13665 11942
rect 13689 11940 13745 11942
rect 13449 10906 13505 10908
rect 13529 10906 13585 10908
rect 13609 10906 13665 10908
rect 13689 10906 13745 10908
rect 13449 10854 13475 10906
rect 13475 10854 13505 10906
rect 13529 10854 13539 10906
rect 13539 10854 13585 10906
rect 13609 10854 13655 10906
rect 13655 10854 13665 10906
rect 13689 10854 13719 10906
rect 13719 10854 13745 10906
rect 13449 10852 13505 10854
rect 13529 10852 13585 10854
rect 13609 10852 13665 10854
rect 13689 10852 13745 10854
rect 13450 10140 13452 10160
rect 13452 10140 13504 10160
rect 13504 10140 13506 10160
rect 13450 10104 13506 10140
rect 13449 9818 13505 9820
rect 13529 9818 13585 9820
rect 13609 9818 13665 9820
rect 13689 9818 13745 9820
rect 13449 9766 13475 9818
rect 13475 9766 13505 9818
rect 13529 9766 13539 9818
rect 13539 9766 13585 9818
rect 13609 9766 13655 9818
rect 13655 9766 13665 9818
rect 13689 9766 13719 9818
rect 13719 9766 13745 9818
rect 13449 9764 13505 9766
rect 13529 9764 13585 9766
rect 13609 9764 13665 9766
rect 13689 9764 13745 9766
rect 13449 8730 13505 8732
rect 13529 8730 13585 8732
rect 13609 8730 13665 8732
rect 13689 8730 13745 8732
rect 13449 8678 13475 8730
rect 13475 8678 13505 8730
rect 13529 8678 13539 8730
rect 13539 8678 13585 8730
rect 13609 8678 13655 8730
rect 13655 8678 13665 8730
rect 13689 8678 13719 8730
rect 13719 8678 13745 8730
rect 13449 8676 13505 8678
rect 13529 8676 13585 8678
rect 13609 8676 13665 8678
rect 13689 8676 13745 8678
rect 13449 7642 13505 7644
rect 13529 7642 13585 7644
rect 13609 7642 13665 7644
rect 13689 7642 13745 7644
rect 13449 7590 13475 7642
rect 13475 7590 13505 7642
rect 13529 7590 13539 7642
rect 13539 7590 13585 7642
rect 13609 7590 13655 7642
rect 13655 7590 13665 7642
rect 13689 7590 13719 7642
rect 13719 7590 13745 7642
rect 13449 7588 13505 7590
rect 13529 7588 13585 7590
rect 13609 7588 13665 7590
rect 13689 7588 13745 7590
rect 13449 6554 13505 6556
rect 13529 6554 13585 6556
rect 13609 6554 13665 6556
rect 13689 6554 13745 6556
rect 13449 6502 13475 6554
rect 13475 6502 13505 6554
rect 13529 6502 13539 6554
rect 13539 6502 13585 6554
rect 13609 6502 13655 6554
rect 13655 6502 13665 6554
rect 13689 6502 13719 6554
rect 13719 6502 13745 6554
rect 13449 6500 13505 6502
rect 13529 6500 13585 6502
rect 13609 6500 13665 6502
rect 13689 6500 13745 6502
rect 13449 5466 13505 5468
rect 13529 5466 13585 5468
rect 13609 5466 13665 5468
rect 13689 5466 13745 5468
rect 13449 5414 13475 5466
rect 13475 5414 13505 5466
rect 13529 5414 13539 5466
rect 13539 5414 13585 5466
rect 13609 5414 13655 5466
rect 13655 5414 13665 5466
rect 13689 5414 13719 5466
rect 13719 5414 13745 5466
rect 13449 5412 13505 5414
rect 13529 5412 13585 5414
rect 13609 5412 13665 5414
rect 13689 5412 13745 5414
rect 13449 4378 13505 4380
rect 13529 4378 13585 4380
rect 13609 4378 13665 4380
rect 13689 4378 13745 4380
rect 13449 4326 13475 4378
rect 13475 4326 13505 4378
rect 13529 4326 13539 4378
rect 13539 4326 13585 4378
rect 13609 4326 13655 4378
rect 13655 4326 13665 4378
rect 13689 4326 13719 4378
rect 13719 4326 13745 4378
rect 13449 4324 13505 4326
rect 13529 4324 13585 4326
rect 13609 4324 13665 4326
rect 13689 4324 13745 4326
rect 13082 3168 13138 3224
rect 13449 3290 13505 3292
rect 13529 3290 13585 3292
rect 13609 3290 13665 3292
rect 13689 3290 13745 3292
rect 13449 3238 13475 3290
rect 13475 3238 13505 3290
rect 13529 3238 13539 3290
rect 13539 3238 13585 3290
rect 13609 3238 13655 3290
rect 13655 3238 13665 3290
rect 13689 3238 13719 3290
rect 13719 3238 13745 3290
rect 13449 3236 13505 3238
rect 13529 3236 13585 3238
rect 13609 3236 13665 3238
rect 13689 3236 13745 3238
rect 13449 2202 13505 2204
rect 13529 2202 13585 2204
rect 13609 2202 13665 2204
rect 13689 2202 13745 2204
rect 13449 2150 13475 2202
rect 13475 2150 13505 2202
rect 13529 2150 13539 2202
rect 13539 2150 13585 2202
rect 13609 2150 13655 2202
rect 13655 2150 13665 2202
rect 13689 2150 13719 2202
rect 13719 2150 13745 2202
rect 13449 2148 13505 2150
rect 13529 2148 13585 2150
rect 13609 2148 13665 2150
rect 13689 2148 13745 2150
rect 14554 15408 14610 15464
rect 14554 14320 14610 14376
rect 14370 13504 14426 13560
rect 14738 15544 14794 15600
rect 14738 12824 14794 12880
rect 14186 2896 14242 2952
rect 15290 15680 15346 15736
rect 16118 17856 16174 17912
rect 15658 13912 15714 13968
rect 15658 9832 15714 9888
rect 14922 1944 14978 2000
rect 15658 5888 15714 5944
rect 2778 448 2834 504
<< metal3 >>
rect 0 19546 800 19576
rect 2957 19546 3023 19549
rect 0 19544 3023 19546
rect 0 19488 2962 19544
rect 3018 19488 3023 19544
rect 0 19486 3023 19488
rect 0 19456 800 19486
rect 2957 19483 3023 19486
rect 0 18594 800 18624
rect 3141 18594 3207 18597
rect 0 18592 3207 18594
rect 0 18536 3146 18592
rect 3202 18536 3207 18592
rect 0 18534 3207 18536
rect 0 18504 800 18534
rect 3141 18531 3207 18534
rect 16113 17914 16179 17917
rect 16400 17914 17200 17944
rect 16113 17912 17200 17914
rect 16113 17856 16118 17912
rect 16174 17856 17200 17912
rect 16113 17854 17200 17856
rect 16113 17851 16179 17854
rect 16400 17824 17200 17854
rect 0 17642 800 17672
rect 1853 17642 1919 17645
rect 0 17640 1919 17642
rect 0 17584 1858 17640
rect 1914 17584 1919 17640
rect 0 17582 1919 17584
rect 0 17552 800 17582
rect 1853 17579 1919 17582
rect 3442 17440 3762 17441
rect 3442 17376 3450 17440
rect 3514 17376 3530 17440
rect 3594 17376 3610 17440
rect 3674 17376 3690 17440
rect 3754 17376 3762 17440
rect 3442 17375 3762 17376
rect 8440 17440 8760 17441
rect 8440 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8760 17440
rect 8440 17375 8760 17376
rect 13437 17440 13757 17441
rect 13437 17376 13445 17440
rect 13509 17376 13525 17440
rect 13589 17376 13605 17440
rect 13669 17376 13685 17440
rect 13749 17376 13757 17440
rect 13437 17375 13757 17376
rect 2497 17098 2563 17101
rect 11053 17098 11119 17101
rect 2497 17096 11119 17098
rect 2497 17040 2502 17096
rect 2558 17040 11058 17096
rect 11114 17040 11119 17096
rect 2497 17038 11119 17040
rect 2497 17035 2563 17038
rect 11053 17035 11119 17038
rect 5941 16896 6261 16897
rect 5941 16832 5949 16896
rect 6013 16832 6029 16896
rect 6093 16832 6109 16896
rect 6173 16832 6189 16896
rect 6253 16832 6261 16896
rect 5941 16831 6261 16832
rect 10938 16896 11258 16897
rect 10938 16832 10946 16896
rect 11010 16832 11026 16896
rect 11090 16832 11106 16896
rect 11170 16832 11186 16896
rect 11250 16832 11258 16896
rect 10938 16831 11258 16832
rect 0 16690 800 16720
rect 1393 16690 1459 16693
rect 0 16688 1459 16690
rect 0 16632 1398 16688
rect 1454 16632 1459 16688
rect 0 16630 1459 16632
rect 0 16600 800 16630
rect 1393 16627 1459 16630
rect 3442 16352 3762 16353
rect 3442 16288 3450 16352
rect 3514 16288 3530 16352
rect 3594 16288 3610 16352
rect 3674 16288 3690 16352
rect 3754 16288 3762 16352
rect 3442 16287 3762 16288
rect 8440 16352 8760 16353
rect 8440 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8760 16352
rect 8440 16287 8760 16288
rect 13437 16352 13757 16353
rect 13437 16288 13445 16352
rect 13509 16288 13525 16352
rect 13589 16288 13605 16352
rect 13669 16288 13685 16352
rect 13749 16288 13757 16352
rect 13437 16287 13757 16288
rect 12525 16146 12591 16149
rect 12750 16146 12756 16148
rect 12525 16144 12756 16146
rect 12525 16088 12530 16144
rect 12586 16088 12756 16144
rect 12525 16086 12756 16088
rect 12525 16083 12591 16086
rect 12750 16084 12756 16086
rect 12820 16084 12826 16148
rect 2957 16010 3023 16013
rect 4245 16010 4311 16013
rect 2957 16008 4311 16010
rect 2957 15952 2962 16008
rect 3018 15952 4250 16008
rect 4306 15952 4311 16008
rect 2957 15950 4311 15952
rect 2957 15947 3023 15950
rect 4245 15947 4311 15950
rect 5941 15808 6261 15809
rect 0 15738 800 15768
rect 5941 15744 5949 15808
rect 6013 15744 6029 15808
rect 6093 15744 6109 15808
rect 6173 15744 6189 15808
rect 6253 15744 6261 15808
rect 5941 15743 6261 15744
rect 10938 15808 11258 15809
rect 10938 15744 10946 15808
rect 11010 15744 11026 15808
rect 11090 15744 11106 15808
rect 11170 15744 11186 15808
rect 11250 15744 11258 15808
rect 10938 15743 11258 15744
rect 1485 15738 1551 15741
rect 0 15736 1551 15738
rect 0 15680 1490 15736
rect 1546 15680 1551 15736
rect 0 15678 1551 15680
rect 0 15648 800 15678
rect 1485 15675 1551 15678
rect 2129 15738 2195 15741
rect 5809 15738 5875 15741
rect 2129 15736 5875 15738
rect 2129 15680 2134 15736
rect 2190 15680 5814 15736
rect 5870 15680 5875 15736
rect 2129 15678 5875 15680
rect 2129 15675 2195 15678
rect 5809 15675 5875 15678
rect 11513 15738 11579 15741
rect 15285 15738 15351 15741
rect 11513 15736 15351 15738
rect 11513 15680 11518 15736
rect 11574 15680 15290 15736
rect 15346 15680 15351 15736
rect 11513 15678 15351 15680
rect 11513 15675 11579 15678
rect 15285 15675 15351 15678
rect 3325 15602 3391 15605
rect 14733 15602 14799 15605
rect 3325 15600 14799 15602
rect 3325 15544 3330 15600
rect 3386 15544 14738 15600
rect 14794 15544 14799 15600
rect 3325 15542 14799 15544
rect 3325 15539 3391 15542
rect 14733 15539 14799 15542
rect 2773 15466 2839 15469
rect 14549 15466 14615 15469
rect 2773 15464 14615 15466
rect 2773 15408 2778 15464
rect 2834 15408 14554 15464
rect 14610 15408 14615 15464
rect 2773 15406 14615 15408
rect 2773 15403 2839 15406
rect 14549 15403 14615 15406
rect 9857 15330 9923 15333
rect 11513 15330 11579 15333
rect 9857 15328 11579 15330
rect 9857 15272 9862 15328
rect 9918 15272 11518 15328
rect 11574 15272 11579 15328
rect 9857 15270 11579 15272
rect 9857 15267 9923 15270
rect 11513 15267 11579 15270
rect 3442 15264 3762 15265
rect 3442 15200 3450 15264
rect 3514 15200 3530 15264
rect 3594 15200 3610 15264
rect 3674 15200 3690 15264
rect 3754 15200 3762 15264
rect 3442 15199 3762 15200
rect 8440 15264 8760 15265
rect 8440 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8760 15264
rect 8440 15199 8760 15200
rect 13437 15264 13757 15265
rect 13437 15200 13445 15264
rect 13509 15200 13525 15264
rect 13589 15200 13605 15264
rect 13669 15200 13685 15264
rect 13749 15200 13757 15264
rect 13437 15199 13757 15200
rect 10133 15194 10199 15197
rect 10501 15194 10567 15197
rect 10133 15192 10567 15194
rect 10133 15136 10138 15192
rect 10194 15136 10506 15192
rect 10562 15136 10567 15192
rect 10133 15134 10567 15136
rect 10133 15131 10199 15134
rect 10501 15131 10567 15134
rect 4061 15058 4127 15061
rect 9305 15058 9371 15061
rect 9581 15058 9647 15061
rect 12893 15058 12959 15061
rect 13169 15058 13235 15061
rect 4061 15056 9506 15058
rect 4061 15000 4066 15056
rect 4122 15000 9310 15056
rect 9366 15000 9506 15056
rect 4061 14998 9506 15000
rect 4061 14995 4127 14998
rect 9305 14995 9371 14998
rect 3141 14922 3207 14925
rect 6637 14922 6703 14925
rect 3141 14920 6703 14922
rect 3141 14864 3146 14920
rect 3202 14864 6642 14920
rect 6698 14864 6703 14920
rect 3141 14862 6703 14864
rect 9446 14922 9506 14998
rect 9581 15056 13235 15058
rect 9581 15000 9586 15056
rect 9642 15000 12898 15056
rect 12954 15000 13174 15056
rect 13230 15000 13235 15056
rect 9581 14998 13235 15000
rect 9581 14995 9647 14998
rect 12893 14995 12959 14998
rect 13169 14995 13235 14998
rect 9949 14922 10015 14925
rect 9446 14920 10015 14922
rect 9446 14864 9954 14920
rect 10010 14864 10015 14920
rect 9446 14862 10015 14864
rect 3141 14859 3207 14862
rect 6637 14859 6703 14862
rect 9949 14859 10015 14862
rect 10593 14922 10659 14925
rect 12433 14922 12499 14925
rect 12893 14922 12959 14925
rect 10593 14920 12959 14922
rect 10593 14864 10598 14920
rect 10654 14864 12438 14920
rect 12494 14864 12898 14920
rect 12954 14864 12959 14920
rect 10593 14862 12959 14864
rect 10593 14859 10659 14862
rect 12433 14859 12499 14862
rect 12893 14859 12959 14862
rect 0 14786 800 14816
rect 1485 14786 1551 14789
rect 0 14784 1551 14786
rect 0 14728 1490 14784
rect 1546 14728 1551 14784
rect 0 14726 1551 14728
rect 0 14696 800 14726
rect 1485 14723 1551 14726
rect 2773 14786 2839 14789
rect 4521 14786 4587 14789
rect 2773 14784 4587 14786
rect 2773 14728 2778 14784
rect 2834 14728 4526 14784
rect 4582 14728 4587 14784
rect 2773 14726 4587 14728
rect 2773 14723 2839 14726
rect 4521 14723 4587 14726
rect 5941 14720 6261 14721
rect 5941 14656 5949 14720
rect 6013 14656 6029 14720
rect 6093 14656 6109 14720
rect 6173 14656 6189 14720
rect 6253 14656 6261 14720
rect 5941 14655 6261 14656
rect 10938 14720 11258 14721
rect 10938 14656 10946 14720
rect 11010 14656 11026 14720
rect 11090 14656 11106 14720
rect 11170 14656 11186 14720
rect 11250 14656 11258 14720
rect 10938 14655 11258 14656
rect 12157 14514 12223 14517
rect 9630 14512 12223 14514
rect 9630 14456 12162 14512
rect 12218 14456 12223 14512
rect 9630 14454 12223 14456
rect 6637 14378 6703 14381
rect 8017 14378 8083 14381
rect 9630 14378 9690 14454
rect 12157 14451 12223 14454
rect 6637 14376 9690 14378
rect 6637 14320 6642 14376
rect 6698 14320 8022 14376
rect 8078 14320 9690 14376
rect 6637 14318 9690 14320
rect 10133 14378 10199 14381
rect 14549 14378 14615 14381
rect 10133 14376 14615 14378
rect 10133 14320 10138 14376
rect 10194 14320 14554 14376
rect 14610 14320 14615 14376
rect 10133 14318 14615 14320
rect 6637 14315 6703 14318
rect 8017 14315 8083 14318
rect 10133 14315 10199 14318
rect 14549 14315 14615 14318
rect 3442 14176 3762 14177
rect 3442 14112 3450 14176
rect 3514 14112 3530 14176
rect 3594 14112 3610 14176
rect 3674 14112 3690 14176
rect 3754 14112 3762 14176
rect 3442 14111 3762 14112
rect 8440 14176 8760 14177
rect 8440 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8760 14176
rect 8440 14111 8760 14112
rect 13437 14176 13757 14177
rect 13437 14112 13445 14176
rect 13509 14112 13525 14176
rect 13589 14112 13605 14176
rect 13669 14112 13685 14176
rect 13749 14112 13757 14176
rect 13437 14111 13757 14112
rect 1945 13970 2011 13973
rect 9121 13970 9187 13973
rect 1945 13968 9187 13970
rect 1945 13912 1950 13968
rect 2006 13912 9126 13968
rect 9182 13912 9187 13968
rect 1945 13910 9187 13912
rect 1945 13907 2011 13910
rect 9121 13907 9187 13910
rect 15653 13970 15719 13973
rect 16400 13970 17200 14000
rect 15653 13968 17200 13970
rect 15653 13912 15658 13968
rect 15714 13912 17200 13968
rect 15653 13910 17200 13912
rect 15653 13907 15719 13910
rect 16400 13880 17200 13910
rect 0 13834 800 13864
rect 1393 13834 1459 13837
rect 0 13832 1459 13834
rect 0 13776 1398 13832
rect 1454 13776 1459 13832
rect 0 13774 1459 13776
rect 0 13744 800 13774
rect 1393 13771 1459 13774
rect 10225 13834 10291 13837
rect 11789 13834 11855 13837
rect 10225 13832 11855 13834
rect 10225 13776 10230 13832
rect 10286 13776 11794 13832
rect 11850 13776 11855 13832
rect 10225 13774 11855 13776
rect 10225 13771 10291 13774
rect 11789 13771 11855 13774
rect 5941 13632 6261 13633
rect 5941 13568 5949 13632
rect 6013 13568 6029 13632
rect 6093 13568 6109 13632
rect 6173 13568 6189 13632
rect 6253 13568 6261 13632
rect 5941 13567 6261 13568
rect 10938 13632 11258 13633
rect 10938 13568 10946 13632
rect 11010 13568 11026 13632
rect 11090 13568 11106 13632
rect 11170 13568 11186 13632
rect 11250 13568 11258 13632
rect 10938 13567 11258 13568
rect 11789 13562 11855 13565
rect 13721 13562 13787 13565
rect 14365 13562 14431 13565
rect 11789 13560 14431 13562
rect 11789 13504 11794 13560
rect 11850 13504 13726 13560
rect 13782 13504 14370 13560
rect 14426 13504 14431 13560
rect 11789 13502 14431 13504
rect 11789 13499 11855 13502
rect 13721 13499 13787 13502
rect 14365 13499 14431 13502
rect 5809 13426 5875 13429
rect 6913 13426 6979 13429
rect 5809 13424 6979 13426
rect 5809 13368 5814 13424
rect 5870 13368 6918 13424
rect 6974 13368 6979 13424
rect 5809 13366 6979 13368
rect 5809 13363 5875 13366
rect 6913 13363 6979 13366
rect 8201 13426 8267 13429
rect 12433 13426 12499 13429
rect 8201 13424 12499 13426
rect 8201 13368 8206 13424
rect 8262 13368 12438 13424
rect 12494 13368 12499 13424
rect 8201 13366 12499 13368
rect 8201 13363 8267 13366
rect 12433 13363 12499 13366
rect 10501 13154 10567 13157
rect 12341 13154 12407 13157
rect 12985 13154 13051 13157
rect 10501 13152 13051 13154
rect 10501 13096 10506 13152
rect 10562 13096 12346 13152
rect 12402 13096 12990 13152
rect 13046 13096 13051 13152
rect 10501 13094 13051 13096
rect 10501 13091 10567 13094
rect 12341 13091 12407 13094
rect 12985 13091 13051 13094
rect 3442 13088 3762 13089
rect 3442 13024 3450 13088
rect 3514 13024 3530 13088
rect 3594 13024 3610 13088
rect 3674 13024 3690 13088
rect 3754 13024 3762 13088
rect 3442 13023 3762 13024
rect 8440 13088 8760 13089
rect 8440 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8760 13088
rect 8440 13023 8760 13024
rect 13437 13088 13757 13089
rect 13437 13024 13445 13088
rect 13509 13024 13525 13088
rect 13589 13024 13605 13088
rect 13669 13024 13685 13088
rect 13749 13024 13757 13088
rect 13437 13023 13757 13024
rect 5993 13018 6059 13021
rect 7373 13018 7439 13021
rect 5993 13016 7439 13018
rect 5993 12960 5998 13016
rect 6054 12960 7378 13016
rect 7434 12960 7439 13016
rect 5993 12958 7439 12960
rect 5993 12955 6059 12958
rect 7373 12955 7439 12958
rect 12750 12956 12756 13020
rect 12820 13018 12826 13020
rect 12893 13018 12959 13021
rect 12820 13016 12959 13018
rect 12820 12960 12898 13016
rect 12954 12960 12959 13016
rect 12820 12958 12959 12960
rect 12820 12956 12826 12958
rect 12893 12955 12959 12958
rect 0 12882 800 12912
rect 1393 12882 1459 12885
rect 6361 12882 6427 12885
rect 0 12880 1459 12882
rect 0 12824 1398 12880
rect 1454 12824 1459 12880
rect 0 12822 1459 12824
rect 0 12792 800 12822
rect 1393 12819 1459 12822
rect 5582 12880 6427 12882
rect 5582 12824 6366 12880
rect 6422 12824 6427 12880
rect 5582 12822 6427 12824
rect 5582 12474 5642 12822
rect 6361 12819 6427 12822
rect 10225 12882 10291 12885
rect 14733 12882 14799 12885
rect 10225 12880 14799 12882
rect 10225 12824 10230 12880
rect 10286 12824 14738 12880
rect 14794 12824 14799 12880
rect 10225 12822 14799 12824
rect 10225 12819 10291 12822
rect 14733 12819 14799 12822
rect 5809 12746 5875 12749
rect 6637 12746 6703 12749
rect 5809 12744 6703 12746
rect 5809 12688 5814 12744
rect 5870 12688 6642 12744
rect 6698 12688 6703 12744
rect 5809 12686 6703 12688
rect 5809 12683 5875 12686
rect 6637 12683 6703 12686
rect 11697 12746 11763 12749
rect 12249 12746 12315 12749
rect 11697 12744 12315 12746
rect 11697 12688 11702 12744
rect 11758 12688 12254 12744
rect 12310 12688 12315 12744
rect 11697 12686 12315 12688
rect 11697 12683 11763 12686
rect 12249 12683 12315 12686
rect 5941 12544 6261 12545
rect 5941 12480 5949 12544
rect 6013 12480 6029 12544
rect 6093 12480 6109 12544
rect 6173 12480 6189 12544
rect 6253 12480 6261 12544
rect 5941 12479 6261 12480
rect 10938 12544 11258 12545
rect 10938 12480 10946 12544
rect 11010 12480 11026 12544
rect 11090 12480 11106 12544
rect 11170 12480 11186 12544
rect 11250 12480 11258 12544
rect 10938 12479 11258 12480
rect 5717 12474 5783 12477
rect 5582 12472 5783 12474
rect 5582 12416 5722 12472
rect 5778 12416 5783 12472
rect 5582 12414 5783 12416
rect 5717 12411 5783 12414
rect 5809 12066 5875 12069
rect 6361 12066 6427 12069
rect 5809 12064 6427 12066
rect 5809 12008 5814 12064
rect 5870 12008 6366 12064
rect 6422 12008 6427 12064
rect 5809 12006 6427 12008
rect 5809 12003 5875 12006
rect 6361 12003 6427 12006
rect 3442 12000 3762 12001
rect 0 11930 800 11960
rect 3442 11936 3450 12000
rect 3514 11936 3530 12000
rect 3594 11936 3610 12000
rect 3674 11936 3690 12000
rect 3754 11936 3762 12000
rect 3442 11935 3762 11936
rect 8440 12000 8760 12001
rect 8440 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8760 12000
rect 8440 11935 8760 11936
rect 13437 12000 13757 12001
rect 13437 11936 13445 12000
rect 13509 11936 13525 12000
rect 13589 11936 13605 12000
rect 13669 11936 13685 12000
rect 13749 11936 13757 12000
rect 13437 11935 13757 11936
rect 1485 11930 1551 11933
rect 0 11928 1551 11930
rect 0 11872 1490 11928
rect 1546 11872 1551 11928
rect 0 11870 1551 11872
rect 0 11840 800 11870
rect 1485 11867 1551 11870
rect 4061 11930 4127 11933
rect 6361 11930 6427 11933
rect 4061 11928 6427 11930
rect 4061 11872 4066 11928
rect 4122 11872 6366 11928
rect 6422 11872 6427 11928
rect 4061 11870 6427 11872
rect 4061 11867 4127 11870
rect 6361 11867 6427 11870
rect 9673 11794 9739 11797
rect 10225 11794 10291 11797
rect 9673 11792 10291 11794
rect 9673 11736 9678 11792
rect 9734 11736 10230 11792
rect 10286 11736 10291 11792
rect 9673 11734 10291 11736
rect 9673 11731 9739 11734
rect 10225 11731 10291 11734
rect 5941 11456 6261 11457
rect 5941 11392 5949 11456
rect 6013 11392 6029 11456
rect 6093 11392 6109 11456
rect 6173 11392 6189 11456
rect 6253 11392 6261 11456
rect 5941 11391 6261 11392
rect 10938 11456 11258 11457
rect 10938 11392 10946 11456
rect 11010 11392 11026 11456
rect 11090 11392 11106 11456
rect 11170 11392 11186 11456
rect 11250 11392 11258 11456
rect 10938 11391 11258 11392
rect 11053 11250 11119 11253
rect 12985 11250 13051 11253
rect 11053 11248 13051 11250
rect 11053 11192 11058 11248
rect 11114 11192 12990 11248
rect 13046 11192 13051 11248
rect 11053 11190 13051 11192
rect 11053 11187 11119 11190
rect 12985 11187 13051 11190
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 3442 10912 3762 10913
rect 3442 10848 3450 10912
rect 3514 10848 3530 10912
rect 3594 10848 3610 10912
rect 3674 10848 3690 10912
rect 3754 10848 3762 10912
rect 3442 10847 3762 10848
rect 8440 10912 8760 10913
rect 8440 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8760 10912
rect 8440 10847 8760 10848
rect 13437 10912 13757 10913
rect 13437 10848 13445 10912
rect 13509 10848 13525 10912
rect 13589 10848 13605 10912
rect 13669 10848 13685 10912
rect 13749 10848 13757 10912
rect 13437 10847 13757 10848
rect 5941 10368 6261 10369
rect 5941 10304 5949 10368
rect 6013 10304 6029 10368
rect 6093 10304 6109 10368
rect 6173 10304 6189 10368
rect 6253 10304 6261 10368
rect 5941 10303 6261 10304
rect 10938 10368 11258 10369
rect 10938 10304 10946 10368
rect 11010 10304 11026 10368
rect 11090 10304 11106 10368
rect 11170 10304 11186 10368
rect 11250 10304 11258 10368
rect 10938 10303 11258 10304
rect 7833 10162 7899 10165
rect 8109 10162 8175 10165
rect 13445 10162 13511 10165
rect 7833 10160 13511 10162
rect 7833 10104 7838 10160
rect 7894 10104 8114 10160
rect 8170 10104 13450 10160
rect 13506 10104 13511 10160
rect 7833 10102 13511 10104
rect 7833 10099 7899 10102
rect 8109 10099 8175 10102
rect 13445 10099 13511 10102
rect 0 10026 800 10056
rect 1393 10026 1459 10029
rect 0 10024 1459 10026
rect 0 9968 1398 10024
rect 1454 9968 1459 10024
rect 0 9966 1459 9968
rect 0 9936 800 9966
rect 1393 9963 1459 9966
rect 15653 9890 15719 9893
rect 16400 9890 17200 9920
rect 15653 9888 17200 9890
rect 15653 9832 15658 9888
rect 15714 9832 17200 9888
rect 15653 9830 17200 9832
rect 15653 9827 15719 9830
rect 3442 9824 3762 9825
rect 3442 9760 3450 9824
rect 3514 9760 3530 9824
rect 3594 9760 3610 9824
rect 3674 9760 3690 9824
rect 3754 9760 3762 9824
rect 3442 9759 3762 9760
rect 8440 9824 8760 9825
rect 8440 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8760 9824
rect 8440 9759 8760 9760
rect 13437 9824 13757 9825
rect 13437 9760 13445 9824
rect 13509 9760 13525 9824
rect 13589 9760 13605 9824
rect 13669 9760 13685 9824
rect 13749 9760 13757 9824
rect 16400 9800 17200 9830
rect 13437 9759 13757 9760
rect 4981 9346 5047 9349
rect 5809 9346 5875 9349
rect 4981 9344 5875 9346
rect 4981 9288 4986 9344
rect 5042 9288 5814 9344
rect 5870 9288 5875 9344
rect 4981 9286 5875 9288
rect 4981 9283 5047 9286
rect 5809 9283 5875 9286
rect 5941 9280 6261 9281
rect 5941 9216 5949 9280
rect 6013 9216 6029 9280
rect 6093 9216 6109 9280
rect 6173 9216 6189 9280
rect 6253 9216 6261 9280
rect 5941 9215 6261 9216
rect 10938 9280 11258 9281
rect 10938 9216 10946 9280
rect 11010 9216 11026 9280
rect 11090 9216 11106 9280
rect 11170 9216 11186 9280
rect 11250 9216 11258 9280
rect 10938 9215 11258 9216
rect 0 9074 800 9104
rect 1393 9074 1459 9077
rect 0 9072 1459 9074
rect 0 9016 1398 9072
rect 1454 9016 1459 9072
rect 0 9014 1459 9016
rect 0 8984 800 9014
rect 1393 9011 1459 9014
rect 8753 8938 8819 8941
rect 8886 8938 8892 8940
rect 8753 8936 8892 8938
rect 8753 8880 8758 8936
rect 8814 8880 8892 8936
rect 8753 8878 8892 8880
rect 8753 8875 8819 8878
rect 8886 8876 8892 8878
rect 8956 8876 8962 8940
rect 3442 8736 3762 8737
rect 3442 8672 3450 8736
rect 3514 8672 3530 8736
rect 3594 8672 3610 8736
rect 3674 8672 3690 8736
rect 3754 8672 3762 8736
rect 3442 8671 3762 8672
rect 8440 8736 8760 8737
rect 8440 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8760 8736
rect 8440 8671 8760 8672
rect 13437 8736 13757 8737
rect 13437 8672 13445 8736
rect 13509 8672 13525 8736
rect 13589 8672 13605 8736
rect 13669 8672 13685 8736
rect 13749 8672 13757 8736
rect 13437 8671 13757 8672
rect 5941 8192 6261 8193
rect 0 8122 800 8152
rect 5941 8128 5949 8192
rect 6013 8128 6029 8192
rect 6093 8128 6109 8192
rect 6173 8128 6189 8192
rect 6253 8128 6261 8192
rect 5941 8127 6261 8128
rect 10938 8192 11258 8193
rect 10938 8128 10946 8192
rect 11010 8128 11026 8192
rect 11090 8128 11106 8192
rect 11170 8128 11186 8192
rect 11250 8128 11258 8192
rect 10938 8127 11258 8128
rect 1485 8122 1551 8125
rect 0 8120 1551 8122
rect 0 8064 1490 8120
rect 1546 8064 1551 8120
rect 0 8062 1551 8064
rect 0 8032 800 8062
rect 1485 8059 1551 8062
rect 7097 8122 7163 8125
rect 7097 8120 9690 8122
rect 7097 8064 7102 8120
rect 7158 8064 9690 8120
rect 7097 8062 9690 8064
rect 7097 8059 7163 8062
rect 6821 7986 6887 7989
rect 7281 7986 7347 7989
rect 9213 7986 9279 7989
rect 6821 7984 9279 7986
rect 6821 7928 6826 7984
rect 6882 7928 7286 7984
rect 7342 7928 9218 7984
rect 9274 7928 9279 7984
rect 6821 7926 9279 7928
rect 9630 7986 9690 8062
rect 10317 8120 10383 8125
rect 10317 8064 10322 8120
rect 10378 8064 10383 8120
rect 10317 8059 10383 8064
rect 10320 7986 10380 8059
rect 11605 7986 11671 7989
rect 9630 7984 11671 7986
rect 9630 7928 11610 7984
rect 11666 7928 11671 7984
rect 9630 7926 11671 7928
rect 6821 7923 6887 7926
rect 7281 7923 7347 7926
rect 9213 7923 9279 7926
rect 11605 7923 11671 7926
rect 5073 7850 5139 7853
rect 8385 7850 8451 7853
rect 5073 7848 8451 7850
rect 5073 7792 5078 7848
rect 5134 7792 8390 7848
rect 8446 7792 8451 7848
rect 5073 7790 8451 7792
rect 5073 7787 5139 7790
rect 8385 7787 8451 7790
rect 8845 7850 8911 7853
rect 8845 7848 9276 7850
rect 8845 7792 8850 7848
rect 8906 7792 9276 7848
rect 8845 7790 9276 7792
rect 8845 7787 8911 7790
rect 9216 7717 9276 7790
rect 9213 7712 9279 7717
rect 9213 7656 9218 7712
rect 9274 7656 9279 7712
rect 9213 7651 9279 7656
rect 3442 7648 3762 7649
rect 3442 7584 3450 7648
rect 3514 7584 3530 7648
rect 3594 7584 3610 7648
rect 3674 7584 3690 7648
rect 3754 7584 3762 7648
rect 3442 7583 3762 7584
rect 8440 7648 8760 7649
rect 8440 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8760 7648
rect 8440 7583 8760 7584
rect 13437 7648 13757 7649
rect 13437 7584 13445 7648
rect 13509 7584 13525 7648
rect 13589 7584 13605 7648
rect 13669 7584 13685 7648
rect 13749 7584 13757 7648
rect 13437 7583 13757 7584
rect 5533 7306 5599 7309
rect 7649 7306 7715 7309
rect 5533 7304 7715 7306
rect 5533 7248 5538 7304
rect 5594 7248 7654 7304
rect 7710 7248 7715 7304
rect 5533 7246 7715 7248
rect 5533 7243 5599 7246
rect 7649 7243 7715 7246
rect 9213 7306 9279 7309
rect 12433 7306 12499 7309
rect 9213 7304 12499 7306
rect 9213 7248 9218 7304
rect 9274 7248 12438 7304
rect 12494 7248 12499 7304
rect 9213 7246 12499 7248
rect 9213 7243 9279 7246
rect 12433 7243 12499 7246
rect 0 7170 800 7200
rect 1485 7170 1551 7173
rect 0 7168 1551 7170
rect 0 7112 1490 7168
rect 1546 7112 1551 7168
rect 0 7110 1551 7112
rect 0 7080 800 7110
rect 1485 7107 1551 7110
rect 8937 7170 9003 7173
rect 9581 7170 9647 7173
rect 8937 7168 9647 7170
rect 8937 7112 8942 7168
rect 8998 7112 9586 7168
rect 9642 7112 9647 7168
rect 8937 7110 9647 7112
rect 8937 7107 9003 7110
rect 9581 7107 9647 7110
rect 5941 7104 6261 7105
rect 5941 7040 5949 7104
rect 6013 7040 6029 7104
rect 6093 7040 6109 7104
rect 6173 7040 6189 7104
rect 6253 7040 6261 7104
rect 5941 7039 6261 7040
rect 10938 7104 11258 7105
rect 10938 7040 10946 7104
rect 11010 7040 11026 7104
rect 11090 7040 11106 7104
rect 11170 7040 11186 7104
rect 11250 7040 11258 7104
rect 10938 7039 11258 7040
rect 10685 6898 10751 6901
rect 10685 6896 10794 6898
rect 10685 6840 10690 6896
rect 10746 6840 10794 6896
rect 10685 6835 10794 6840
rect 6729 6628 6795 6629
rect 6678 6564 6684 6628
rect 6748 6626 6795 6628
rect 10734 6626 10794 6835
rect 11237 6762 11303 6765
rect 12893 6762 12959 6765
rect 11237 6760 12959 6762
rect 11237 6704 11242 6760
rect 11298 6704 12898 6760
rect 12954 6704 12959 6760
rect 11237 6702 12959 6704
rect 11237 6699 11303 6702
rect 12893 6699 12959 6702
rect 11421 6626 11487 6629
rect 6748 6624 6840 6626
rect 6790 6568 6840 6624
rect 6748 6566 6840 6568
rect 10734 6624 11487 6626
rect 10734 6568 11426 6624
rect 11482 6568 11487 6624
rect 10734 6566 11487 6568
rect 6748 6564 6795 6566
rect 6729 6563 6795 6564
rect 11421 6563 11487 6566
rect 3442 6560 3762 6561
rect 3442 6496 3450 6560
rect 3514 6496 3530 6560
rect 3594 6496 3610 6560
rect 3674 6496 3690 6560
rect 3754 6496 3762 6560
rect 3442 6495 3762 6496
rect 8440 6560 8760 6561
rect 8440 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8760 6560
rect 8440 6495 8760 6496
rect 13437 6560 13757 6561
rect 13437 6496 13445 6560
rect 13509 6496 13525 6560
rect 13589 6496 13605 6560
rect 13669 6496 13685 6560
rect 13749 6496 13757 6560
rect 13437 6495 13757 6496
rect 9029 6354 9095 6357
rect 9581 6354 9647 6357
rect 9029 6352 9647 6354
rect 9029 6296 9034 6352
rect 9090 6296 9586 6352
rect 9642 6296 9647 6352
rect 9029 6294 9647 6296
rect 9029 6291 9095 6294
rect 9581 6291 9647 6294
rect 12341 6354 12407 6357
rect 12617 6354 12683 6357
rect 12341 6352 12683 6354
rect 12341 6296 12346 6352
rect 12402 6296 12622 6352
rect 12678 6296 12683 6352
rect 12341 6294 12683 6296
rect 12341 6291 12407 6294
rect 12617 6291 12683 6294
rect 0 6218 800 6248
rect 1485 6218 1551 6221
rect 0 6216 1551 6218
rect 0 6160 1490 6216
rect 1546 6160 1551 6216
rect 0 6158 1551 6160
rect 0 6128 800 6158
rect 1485 6155 1551 6158
rect 10133 6082 10199 6085
rect 10501 6082 10567 6085
rect 9814 6080 10567 6082
rect 9814 6024 10138 6080
rect 10194 6024 10506 6080
rect 10562 6024 10567 6080
rect 9814 6022 10567 6024
rect 5941 6016 6261 6017
rect 5941 5952 5949 6016
rect 6013 5952 6029 6016
rect 6093 5952 6109 6016
rect 6173 5952 6189 6016
rect 6253 5952 6261 6016
rect 5941 5951 6261 5952
rect 9814 5949 9874 6022
rect 10133 6019 10199 6022
rect 10501 6019 10567 6022
rect 10938 6016 11258 6017
rect 10938 5952 10946 6016
rect 11010 5952 11026 6016
rect 11090 5952 11106 6016
rect 11170 5952 11186 6016
rect 11250 5952 11258 6016
rect 10938 5951 11258 5952
rect 9765 5944 9874 5949
rect 9765 5888 9770 5944
rect 9826 5888 9874 5944
rect 9765 5886 9874 5888
rect 15653 5946 15719 5949
rect 16400 5946 17200 5976
rect 15653 5944 17200 5946
rect 15653 5888 15658 5944
rect 15714 5888 17200 5944
rect 15653 5886 17200 5888
rect 9765 5883 9831 5886
rect 15653 5883 15719 5886
rect 16400 5856 17200 5886
rect 8886 5476 8892 5540
rect 8956 5538 8962 5540
rect 9213 5538 9279 5541
rect 8956 5536 9279 5538
rect 8956 5480 9218 5536
rect 9274 5480 9279 5536
rect 8956 5478 9279 5480
rect 8956 5476 8962 5478
rect 9213 5475 9279 5478
rect 9673 5538 9739 5541
rect 11053 5538 11119 5541
rect 9673 5536 11119 5538
rect 9673 5480 9678 5536
rect 9734 5480 11058 5536
rect 11114 5480 11119 5536
rect 9673 5478 11119 5480
rect 9673 5475 9739 5478
rect 11053 5475 11119 5478
rect 3442 5472 3762 5473
rect 3442 5408 3450 5472
rect 3514 5408 3530 5472
rect 3594 5408 3610 5472
rect 3674 5408 3690 5472
rect 3754 5408 3762 5472
rect 3442 5407 3762 5408
rect 8440 5472 8760 5473
rect 8440 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8760 5472
rect 8440 5407 8760 5408
rect 13437 5472 13757 5473
rect 13437 5408 13445 5472
rect 13509 5408 13525 5472
rect 13589 5408 13605 5472
rect 13669 5408 13685 5472
rect 13749 5408 13757 5472
rect 13437 5407 13757 5408
rect 6177 5402 6243 5405
rect 6545 5402 6611 5405
rect 6177 5400 6611 5402
rect 6177 5344 6182 5400
rect 6238 5344 6550 5400
rect 6606 5344 6611 5400
rect 6177 5342 6611 5344
rect 6177 5339 6243 5342
rect 6545 5339 6611 5342
rect 9765 5402 9831 5405
rect 11462 5402 11468 5404
rect 9765 5400 11468 5402
rect 9765 5344 9770 5400
rect 9826 5344 11468 5400
rect 9765 5342 11468 5344
rect 9765 5339 9831 5342
rect 11462 5340 11468 5342
rect 11532 5402 11538 5404
rect 11697 5402 11763 5405
rect 11532 5400 11763 5402
rect 11532 5344 11702 5400
rect 11758 5344 11763 5400
rect 11532 5342 11763 5344
rect 11532 5340 11538 5342
rect 11697 5339 11763 5342
rect 0 5266 800 5296
rect 1393 5266 1459 5269
rect 0 5264 1459 5266
rect 0 5208 1398 5264
rect 1454 5208 1459 5264
rect 0 5206 1459 5208
rect 0 5176 800 5206
rect 1393 5203 1459 5206
rect 7189 5266 7255 5269
rect 9581 5266 9647 5269
rect 7189 5264 9647 5266
rect 7189 5208 7194 5264
rect 7250 5208 9586 5264
rect 9642 5208 9647 5264
rect 7189 5206 9647 5208
rect 7189 5203 7255 5206
rect 9581 5203 9647 5206
rect 9765 5266 9831 5269
rect 11789 5266 11855 5269
rect 9765 5264 11855 5266
rect 9765 5208 9770 5264
rect 9826 5208 11794 5264
rect 11850 5208 11855 5264
rect 9765 5206 11855 5208
rect 9765 5203 9831 5206
rect 11789 5203 11855 5206
rect 5625 5130 5691 5133
rect 9397 5130 9463 5133
rect 5625 5128 9463 5130
rect 5625 5072 5630 5128
rect 5686 5072 9402 5128
rect 9458 5072 9463 5128
rect 5625 5070 9463 5072
rect 5625 5067 5691 5070
rect 9397 5067 9463 5070
rect 10501 4994 10567 4997
rect 10685 4994 10751 4997
rect 10501 4992 10751 4994
rect 10501 4936 10506 4992
rect 10562 4936 10690 4992
rect 10746 4936 10751 4992
rect 10501 4934 10751 4936
rect 10501 4931 10567 4934
rect 10685 4931 10751 4934
rect 5941 4928 6261 4929
rect 5941 4864 5949 4928
rect 6013 4864 6029 4928
rect 6093 4864 6109 4928
rect 6173 4864 6189 4928
rect 6253 4864 6261 4928
rect 5941 4863 6261 4864
rect 10938 4928 11258 4929
rect 10938 4864 10946 4928
rect 11010 4864 11026 4928
rect 11090 4864 11106 4928
rect 11170 4864 11186 4928
rect 11250 4864 11258 4928
rect 10938 4863 11258 4864
rect 4102 4796 4108 4860
rect 4172 4858 4178 4860
rect 4245 4858 4311 4861
rect 4172 4856 4311 4858
rect 4172 4800 4250 4856
rect 4306 4800 4311 4856
rect 4172 4798 4311 4800
rect 4172 4796 4178 4798
rect 4245 4795 4311 4798
rect 2221 4722 2287 4725
rect 8569 4722 8635 4725
rect 2221 4720 8635 4722
rect 2221 4664 2226 4720
rect 2282 4664 8574 4720
rect 8630 4664 8635 4720
rect 2221 4662 8635 4664
rect 2221 4659 2287 4662
rect 8569 4659 8635 4662
rect 3693 4586 3759 4589
rect 8661 4586 8727 4589
rect 9305 4586 9371 4589
rect 3693 4584 9371 4586
rect 3693 4528 3698 4584
rect 3754 4528 8666 4584
rect 8722 4528 9310 4584
rect 9366 4528 9371 4584
rect 3693 4526 9371 4528
rect 3693 4523 3759 4526
rect 8661 4523 8727 4526
rect 9305 4523 9371 4526
rect 3442 4384 3762 4385
rect 0 4314 800 4344
rect 3442 4320 3450 4384
rect 3514 4320 3530 4384
rect 3594 4320 3610 4384
rect 3674 4320 3690 4384
rect 3754 4320 3762 4384
rect 3442 4319 3762 4320
rect 8440 4384 8760 4385
rect 8440 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8760 4384
rect 8440 4319 8760 4320
rect 13437 4384 13757 4385
rect 13437 4320 13445 4384
rect 13509 4320 13525 4384
rect 13589 4320 13605 4384
rect 13669 4320 13685 4384
rect 13749 4320 13757 4384
rect 13437 4319 13757 4320
rect 1393 4314 1459 4317
rect 12617 4316 12683 4317
rect 12566 4314 12572 4316
rect 0 4312 1459 4314
rect 0 4256 1398 4312
rect 1454 4256 1459 4312
rect 0 4254 1459 4256
rect 12526 4254 12572 4314
rect 12636 4312 12683 4316
rect 12678 4256 12683 4312
rect 0 4224 800 4254
rect 1393 4251 1459 4254
rect 12566 4252 12572 4254
rect 12636 4252 12683 4256
rect 12617 4251 12683 4252
rect 8109 4178 8175 4181
rect 12617 4178 12683 4181
rect 8109 4176 12683 4178
rect 8109 4120 8114 4176
rect 8170 4120 12622 4176
rect 12678 4120 12683 4176
rect 8109 4118 12683 4120
rect 8109 4115 8175 4118
rect 12617 4115 12683 4118
rect 11881 3906 11947 3909
rect 12341 3906 12407 3909
rect 11881 3904 12407 3906
rect 11881 3848 11886 3904
rect 11942 3848 12346 3904
rect 12402 3848 12407 3904
rect 11881 3846 12407 3848
rect 11881 3843 11947 3846
rect 12341 3843 12407 3846
rect 5941 3840 6261 3841
rect 5941 3776 5949 3840
rect 6013 3776 6029 3840
rect 6093 3776 6109 3840
rect 6173 3776 6189 3840
rect 6253 3776 6261 3840
rect 5941 3775 6261 3776
rect 10938 3840 11258 3841
rect 10938 3776 10946 3840
rect 11010 3776 11026 3840
rect 11090 3776 11106 3840
rect 11170 3776 11186 3840
rect 11250 3776 11258 3840
rect 10938 3775 11258 3776
rect 6637 3772 6703 3773
rect 6637 3770 6684 3772
rect 6556 3768 6684 3770
rect 6748 3770 6754 3772
rect 9397 3770 9463 3773
rect 6748 3768 9463 3770
rect 6556 3712 6642 3768
rect 6748 3712 9402 3768
rect 9458 3712 9463 3768
rect 6556 3710 6684 3712
rect 6637 3708 6684 3710
rect 6748 3710 9463 3712
rect 6748 3708 6754 3710
rect 6637 3707 6703 3708
rect 9397 3707 9463 3710
rect 12341 3634 12407 3637
rect 11838 3632 12407 3634
rect 11838 3576 12346 3632
rect 12402 3576 12407 3632
rect 11838 3574 12407 3576
rect 11421 3498 11487 3501
rect 11838 3498 11898 3574
rect 12341 3571 12407 3574
rect 11421 3496 11898 3498
rect 11421 3440 11426 3496
rect 11482 3440 11898 3496
rect 11421 3438 11898 3440
rect 11421 3435 11487 3438
rect 0 3362 800 3392
rect 1485 3362 1551 3365
rect 0 3360 1551 3362
rect 0 3304 1490 3360
rect 1546 3304 1551 3360
rect 0 3302 1551 3304
rect 0 3272 800 3302
rect 1485 3299 1551 3302
rect 10409 3362 10475 3365
rect 11881 3362 11947 3365
rect 10409 3360 11947 3362
rect 10409 3304 10414 3360
rect 10470 3304 11886 3360
rect 11942 3304 11947 3360
rect 10409 3302 11947 3304
rect 10409 3299 10475 3302
rect 11881 3299 11947 3302
rect 3442 3296 3762 3297
rect 3442 3232 3450 3296
rect 3514 3232 3530 3296
rect 3594 3232 3610 3296
rect 3674 3232 3690 3296
rect 3754 3232 3762 3296
rect 3442 3231 3762 3232
rect 8440 3296 8760 3297
rect 8440 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8760 3296
rect 8440 3231 8760 3232
rect 13437 3296 13757 3297
rect 13437 3232 13445 3296
rect 13509 3232 13525 3296
rect 13589 3232 13605 3296
rect 13669 3232 13685 3296
rect 13749 3232 13757 3296
rect 13437 3231 13757 3232
rect 9765 3226 9831 3229
rect 13077 3226 13143 3229
rect 9765 3224 13143 3226
rect 9765 3168 9770 3224
rect 9826 3168 13082 3224
rect 13138 3168 13143 3224
rect 9765 3166 13143 3168
rect 9765 3163 9831 3166
rect 13077 3163 13143 3166
rect 6269 3090 6335 3093
rect 8937 3090 9003 3093
rect 6269 3088 9003 3090
rect 6269 3032 6274 3088
rect 6330 3032 8942 3088
rect 8998 3032 9003 3088
rect 6269 3030 9003 3032
rect 6269 3027 6335 3030
rect 8937 3027 9003 3030
rect 1669 2954 1735 2957
rect 9213 2954 9279 2957
rect 1669 2952 9279 2954
rect 1669 2896 1674 2952
rect 1730 2896 9218 2952
rect 9274 2896 9279 2952
rect 1669 2894 9279 2896
rect 1669 2891 1735 2894
rect 9213 2891 9279 2894
rect 10593 2954 10659 2957
rect 11881 2954 11947 2957
rect 10593 2952 11947 2954
rect 10593 2896 10598 2952
rect 10654 2896 11886 2952
rect 11942 2896 11947 2952
rect 10593 2894 11947 2896
rect 10593 2891 10659 2894
rect 11881 2891 11947 2894
rect 12065 2954 12131 2957
rect 14181 2954 14247 2957
rect 12065 2952 14247 2954
rect 12065 2896 12070 2952
rect 12126 2896 14186 2952
rect 14242 2896 14247 2952
rect 12065 2894 14247 2896
rect 12065 2891 12131 2894
rect 14181 2891 14247 2894
rect 5441 2818 5507 2821
rect 5809 2818 5875 2821
rect 5441 2816 5875 2818
rect 5441 2760 5446 2816
rect 5502 2760 5814 2816
rect 5870 2760 5875 2816
rect 5441 2758 5875 2760
rect 5441 2755 5507 2758
rect 5809 2755 5875 2758
rect 5941 2752 6261 2753
rect 5941 2688 5949 2752
rect 6013 2688 6029 2752
rect 6093 2688 6109 2752
rect 6173 2688 6189 2752
rect 6253 2688 6261 2752
rect 5941 2687 6261 2688
rect 10938 2752 11258 2753
rect 10938 2688 10946 2752
rect 11010 2688 11026 2752
rect 11090 2688 11106 2752
rect 11170 2688 11186 2752
rect 11250 2688 11258 2752
rect 10938 2687 11258 2688
rect 12617 2684 12683 2685
rect 12566 2620 12572 2684
rect 12636 2682 12683 2684
rect 12636 2680 12728 2682
rect 12678 2624 12728 2680
rect 12636 2622 12728 2624
rect 12636 2620 12683 2622
rect 12617 2619 12683 2620
rect 4061 2548 4127 2549
rect 4061 2546 4108 2548
rect 4016 2544 4108 2546
rect 4016 2488 4066 2544
rect 4016 2486 4108 2488
rect 4061 2484 4108 2486
rect 4172 2484 4178 2548
rect 11329 2546 11395 2549
rect 11462 2546 11468 2548
rect 11329 2544 11468 2546
rect 11329 2488 11334 2544
rect 11390 2488 11468 2544
rect 11329 2486 11468 2488
rect 4061 2483 4127 2484
rect 11329 2483 11395 2486
rect 11462 2484 11468 2486
rect 11532 2484 11538 2548
rect 0 2410 800 2440
rect 4061 2410 4127 2413
rect 0 2408 4127 2410
rect 0 2352 4066 2408
rect 4122 2352 4127 2408
rect 0 2350 4127 2352
rect 0 2320 800 2350
rect 4061 2347 4127 2350
rect 3442 2208 3762 2209
rect 3442 2144 3450 2208
rect 3514 2144 3530 2208
rect 3594 2144 3610 2208
rect 3674 2144 3690 2208
rect 3754 2144 3762 2208
rect 3442 2143 3762 2144
rect 8440 2208 8760 2209
rect 8440 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8760 2208
rect 8440 2143 8760 2144
rect 13437 2208 13757 2209
rect 13437 2144 13445 2208
rect 13509 2144 13525 2208
rect 13589 2144 13605 2208
rect 13669 2144 13685 2208
rect 13749 2144 13757 2208
rect 13437 2143 13757 2144
rect 14917 2002 14983 2005
rect 16400 2002 17200 2032
rect 14917 2000 17200 2002
rect 14917 1944 14922 2000
rect 14978 1944 17200 2000
rect 14917 1942 17200 1944
rect 14917 1939 14983 1942
rect 16400 1912 17200 1942
rect 0 1458 800 1488
rect 3601 1458 3667 1461
rect 0 1456 3667 1458
rect 0 1400 3606 1456
rect 3662 1400 3667 1456
rect 0 1398 3667 1400
rect 0 1368 800 1398
rect 3601 1395 3667 1398
rect 0 506 800 536
rect 2773 506 2839 509
rect 0 504 2839 506
rect 0 448 2778 504
rect 2834 448 2839 504
rect 0 446 2839 448
rect 0 416 800 446
rect 2773 443 2839 446
<< via3 >>
rect 3450 17436 3514 17440
rect 3450 17380 3454 17436
rect 3454 17380 3510 17436
rect 3510 17380 3514 17436
rect 3450 17376 3514 17380
rect 3530 17436 3594 17440
rect 3530 17380 3534 17436
rect 3534 17380 3590 17436
rect 3590 17380 3594 17436
rect 3530 17376 3594 17380
rect 3610 17436 3674 17440
rect 3610 17380 3614 17436
rect 3614 17380 3670 17436
rect 3670 17380 3674 17436
rect 3610 17376 3674 17380
rect 3690 17436 3754 17440
rect 3690 17380 3694 17436
rect 3694 17380 3750 17436
rect 3750 17380 3754 17436
rect 3690 17376 3754 17380
rect 8448 17436 8512 17440
rect 8448 17380 8452 17436
rect 8452 17380 8508 17436
rect 8508 17380 8512 17436
rect 8448 17376 8512 17380
rect 8528 17436 8592 17440
rect 8528 17380 8532 17436
rect 8532 17380 8588 17436
rect 8588 17380 8592 17436
rect 8528 17376 8592 17380
rect 8608 17436 8672 17440
rect 8608 17380 8612 17436
rect 8612 17380 8668 17436
rect 8668 17380 8672 17436
rect 8608 17376 8672 17380
rect 8688 17436 8752 17440
rect 8688 17380 8692 17436
rect 8692 17380 8748 17436
rect 8748 17380 8752 17436
rect 8688 17376 8752 17380
rect 13445 17436 13509 17440
rect 13445 17380 13449 17436
rect 13449 17380 13505 17436
rect 13505 17380 13509 17436
rect 13445 17376 13509 17380
rect 13525 17436 13589 17440
rect 13525 17380 13529 17436
rect 13529 17380 13585 17436
rect 13585 17380 13589 17436
rect 13525 17376 13589 17380
rect 13605 17436 13669 17440
rect 13605 17380 13609 17436
rect 13609 17380 13665 17436
rect 13665 17380 13669 17436
rect 13605 17376 13669 17380
rect 13685 17436 13749 17440
rect 13685 17380 13689 17436
rect 13689 17380 13745 17436
rect 13745 17380 13749 17436
rect 13685 17376 13749 17380
rect 5949 16892 6013 16896
rect 5949 16836 5953 16892
rect 5953 16836 6009 16892
rect 6009 16836 6013 16892
rect 5949 16832 6013 16836
rect 6029 16892 6093 16896
rect 6029 16836 6033 16892
rect 6033 16836 6089 16892
rect 6089 16836 6093 16892
rect 6029 16832 6093 16836
rect 6109 16892 6173 16896
rect 6109 16836 6113 16892
rect 6113 16836 6169 16892
rect 6169 16836 6173 16892
rect 6109 16832 6173 16836
rect 6189 16892 6253 16896
rect 6189 16836 6193 16892
rect 6193 16836 6249 16892
rect 6249 16836 6253 16892
rect 6189 16832 6253 16836
rect 10946 16892 11010 16896
rect 10946 16836 10950 16892
rect 10950 16836 11006 16892
rect 11006 16836 11010 16892
rect 10946 16832 11010 16836
rect 11026 16892 11090 16896
rect 11026 16836 11030 16892
rect 11030 16836 11086 16892
rect 11086 16836 11090 16892
rect 11026 16832 11090 16836
rect 11106 16892 11170 16896
rect 11106 16836 11110 16892
rect 11110 16836 11166 16892
rect 11166 16836 11170 16892
rect 11106 16832 11170 16836
rect 11186 16892 11250 16896
rect 11186 16836 11190 16892
rect 11190 16836 11246 16892
rect 11246 16836 11250 16892
rect 11186 16832 11250 16836
rect 3450 16348 3514 16352
rect 3450 16292 3454 16348
rect 3454 16292 3510 16348
rect 3510 16292 3514 16348
rect 3450 16288 3514 16292
rect 3530 16348 3594 16352
rect 3530 16292 3534 16348
rect 3534 16292 3590 16348
rect 3590 16292 3594 16348
rect 3530 16288 3594 16292
rect 3610 16348 3674 16352
rect 3610 16292 3614 16348
rect 3614 16292 3670 16348
rect 3670 16292 3674 16348
rect 3610 16288 3674 16292
rect 3690 16348 3754 16352
rect 3690 16292 3694 16348
rect 3694 16292 3750 16348
rect 3750 16292 3754 16348
rect 3690 16288 3754 16292
rect 8448 16348 8512 16352
rect 8448 16292 8452 16348
rect 8452 16292 8508 16348
rect 8508 16292 8512 16348
rect 8448 16288 8512 16292
rect 8528 16348 8592 16352
rect 8528 16292 8532 16348
rect 8532 16292 8588 16348
rect 8588 16292 8592 16348
rect 8528 16288 8592 16292
rect 8608 16348 8672 16352
rect 8608 16292 8612 16348
rect 8612 16292 8668 16348
rect 8668 16292 8672 16348
rect 8608 16288 8672 16292
rect 8688 16348 8752 16352
rect 8688 16292 8692 16348
rect 8692 16292 8748 16348
rect 8748 16292 8752 16348
rect 8688 16288 8752 16292
rect 13445 16348 13509 16352
rect 13445 16292 13449 16348
rect 13449 16292 13505 16348
rect 13505 16292 13509 16348
rect 13445 16288 13509 16292
rect 13525 16348 13589 16352
rect 13525 16292 13529 16348
rect 13529 16292 13585 16348
rect 13585 16292 13589 16348
rect 13525 16288 13589 16292
rect 13605 16348 13669 16352
rect 13605 16292 13609 16348
rect 13609 16292 13665 16348
rect 13665 16292 13669 16348
rect 13605 16288 13669 16292
rect 13685 16348 13749 16352
rect 13685 16292 13689 16348
rect 13689 16292 13745 16348
rect 13745 16292 13749 16348
rect 13685 16288 13749 16292
rect 12756 16084 12820 16148
rect 5949 15804 6013 15808
rect 5949 15748 5953 15804
rect 5953 15748 6009 15804
rect 6009 15748 6013 15804
rect 5949 15744 6013 15748
rect 6029 15804 6093 15808
rect 6029 15748 6033 15804
rect 6033 15748 6089 15804
rect 6089 15748 6093 15804
rect 6029 15744 6093 15748
rect 6109 15804 6173 15808
rect 6109 15748 6113 15804
rect 6113 15748 6169 15804
rect 6169 15748 6173 15804
rect 6109 15744 6173 15748
rect 6189 15804 6253 15808
rect 6189 15748 6193 15804
rect 6193 15748 6249 15804
rect 6249 15748 6253 15804
rect 6189 15744 6253 15748
rect 10946 15804 11010 15808
rect 10946 15748 10950 15804
rect 10950 15748 11006 15804
rect 11006 15748 11010 15804
rect 10946 15744 11010 15748
rect 11026 15804 11090 15808
rect 11026 15748 11030 15804
rect 11030 15748 11086 15804
rect 11086 15748 11090 15804
rect 11026 15744 11090 15748
rect 11106 15804 11170 15808
rect 11106 15748 11110 15804
rect 11110 15748 11166 15804
rect 11166 15748 11170 15804
rect 11106 15744 11170 15748
rect 11186 15804 11250 15808
rect 11186 15748 11190 15804
rect 11190 15748 11246 15804
rect 11246 15748 11250 15804
rect 11186 15744 11250 15748
rect 3450 15260 3514 15264
rect 3450 15204 3454 15260
rect 3454 15204 3510 15260
rect 3510 15204 3514 15260
rect 3450 15200 3514 15204
rect 3530 15260 3594 15264
rect 3530 15204 3534 15260
rect 3534 15204 3590 15260
rect 3590 15204 3594 15260
rect 3530 15200 3594 15204
rect 3610 15260 3674 15264
rect 3610 15204 3614 15260
rect 3614 15204 3670 15260
rect 3670 15204 3674 15260
rect 3610 15200 3674 15204
rect 3690 15260 3754 15264
rect 3690 15204 3694 15260
rect 3694 15204 3750 15260
rect 3750 15204 3754 15260
rect 3690 15200 3754 15204
rect 8448 15260 8512 15264
rect 8448 15204 8452 15260
rect 8452 15204 8508 15260
rect 8508 15204 8512 15260
rect 8448 15200 8512 15204
rect 8528 15260 8592 15264
rect 8528 15204 8532 15260
rect 8532 15204 8588 15260
rect 8588 15204 8592 15260
rect 8528 15200 8592 15204
rect 8608 15260 8672 15264
rect 8608 15204 8612 15260
rect 8612 15204 8668 15260
rect 8668 15204 8672 15260
rect 8608 15200 8672 15204
rect 8688 15260 8752 15264
rect 8688 15204 8692 15260
rect 8692 15204 8748 15260
rect 8748 15204 8752 15260
rect 8688 15200 8752 15204
rect 13445 15260 13509 15264
rect 13445 15204 13449 15260
rect 13449 15204 13505 15260
rect 13505 15204 13509 15260
rect 13445 15200 13509 15204
rect 13525 15260 13589 15264
rect 13525 15204 13529 15260
rect 13529 15204 13585 15260
rect 13585 15204 13589 15260
rect 13525 15200 13589 15204
rect 13605 15260 13669 15264
rect 13605 15204 13609 15260
rect 13609 15204 13665 15260
rect 13665 15204 13669 15260
rect 13605 15200 13669 15204
rect 13685 15260 13749 15264
rect 13685 15204 13689 15260
rect 13689 15204 13745 15260
rect 13745 15204 13749 15260
rect 13685 15200 13749 15204
rect 5949 14716 6013 14720
rect 5949 14660 5953 14716
rect 5953 14660 6009 14716
rect 6009 14660 6013 14716
rect 5949 14656 6013 14660
rect 6029 14716 6093 14720
rect 6029 14660 6033 14716
rect 6033 14660 6089 14716
rect 6089 14660 6093 14716
rect 6029 14656 6093 14660
rect 6109 14716 6173 14720
rect 6109 14660 6113 14716
rect 6113 14660 6169 14716
rect 6169 14660 6173 14716
rect 6109 14656 6173 14660
rect 6189 14716 6253 14720
rect 6189 14660 6193 14716
rect 6193 14660 6249 14716
rect 6249 14660 6253 14716
rect 6189 14656 6253 14660
rect 10946 14716 11010 14720
rect 10946 14660 10950 14716
rect 10950 14660 11006 14716
rect 11006 14660 11010 14716
rect 10946 14656 11010 14660
rect 11026 14716 11090 14720
rect 11026 14660 11030 14716
rect 11030 14660 11086 14716
rect 11086 14660 11090 14716
rect 11026 14656 11090 14660
rect 11106 14716 11170 14720
rect 11106 14660 11110 14716
rect 11110 14660 11166 14716
rect 11166 14660 11170 14716
rect 11106 14656 11170 14660
rect 11186 14716 11250 14720
rect 11186 14660 11190 14716
rect 11190 14660 11246 14716
rect 11246 14660 11250 14716
rect 11186 14656 11250 14660
rect 3450 14172 3514 14176
rect 3450 14116 3454 14172
rect 3454 14116 3510 14172
rect 3510 14116 3514 14172
rect 3450 14112 3514 14116
rect 3530 14172 3594 14176
rect 3530 14116 3534 14172
rect 3534 14116 3590 14172
rect 3590 14116 3594 14172
rect 3530 14112 3594 14116
rect 3610 14172 3674 14176
rect 3610 14116 3614 14172
rect 3614 14116 3670 14172
rect 3670 14116 3674 14172
rect 3610 14112 3674 14116
rect 3690 14172 3754 14176
rect 3690 14116 3694 14172
rect 3694 14116 3750 14172
rect 3750 14116 3754 14172
rect 3690 14112 3754 14116
rect 8448 14172 8512 14176
rect 8448 14116 8452 14172
rect 8452 14116 8508 14172
rect 8508 14116 8512 14172
rect 8448 14112 8512 14116
rect 8528 14172 8592 14176
rect 8528 14116 8532 14172
rect 8532 14116 8588 14172
rect 8588 14116 8592 14172
rect 8528 14112 8592 14116
rect 8608 14172 8672 14176
rect 8608 14116 8612 14172
rect 8612 14116 8668 14172
rect 8668 14116 8672 14172
rect 8608 14112 8672 14116
rect 8688 14172 8752 14176
rect 8688 14116 8692 14172
rect 8692 14116 8748 14172
rect 8748 14116 8752 14172
rect 8688 14112 8752 14116
rect 13445 14172 13509 14176
rect 13445 14116 13449 14172
rect 13449 14116 13505 14172
rect 13505 14116 13509 14172
rect 13445 14112 13509 14116
rect 13525 14172 13589 14176
rect 13525 14116 13529 14172
rect 13529 14116 13585 14172
rect 13585 14116 13589 14172
rect 13525 14112 13589 14116
rect 13605 14172 13669 14176
rect 13605 14116 13609 14172
rect 13609 14116 13665 14172
rect 13665 14116 13669 14172
rect 13605 14112 13669 14116
rect 13685 14172 13749 14176
rect 13685 14116 13689 14172
rect 13689 14116 13745 14172
rect 13745 14116 13749 14172
rect 13685 14112 13749 14116
rect 5949 13628 6013 13632
rect 5949 13572 5953 13628
rect 5953 13572 6009 13628
rect 6009 13572 6013 13628
rect 5949 13568 6013 13572
rect 6029 13628 6093 13632
rect 6029 13572 6033 13628
rect 6033 13572 6089 13628
rect 6089 13572 6093 13628
rect 6029 13568 6093 13572
rect 6109 13628 6173 13632
rect 6109 13572 6113 13628
rect 6113 13572 6169 13628
rect 6169 13572 6173 13628
rect 6109 13568 6173 13572
rect 6189 13628 6253 13632
rect 6189 13572 6193 13628
rect 6193 13572 6249 13628
rect 6249 13572 6253 13628
rect 6189 13568 6253 13572
rect 10946 13628 11010 13632
rect 10946 13572 10950 13628
rect 10950 13572 11006 13628
rect 11006 13572 11010 13628
rect 10946 13568 11010 13572
rect 11026 13628 11090 13632
rect 11026 13572 11030 13628
rect 11030 13572 11086 13628
rect 11086 13572 11090 13628
rect 11026 13568 11090 13572
rect 11106 13628 11170 13632
rect 11106 13572 11110 13628
rect 11110 13572 11166 13628
rect 11166 13572 11170 13628
rect 11106 13568 11170 13572
rect 11186 13628 11250 13632
rect 11186 13572 11190 13628
rect 11190 13572 11246 13628
rect 11246 13572 11250 13628
rect 11186 13568 11250 13572
rect 3450 13084 3514 13088
rect 3450 13028 3454 13084
rect 3454 13028 3510 13084
rect 3510 13028 3514 13084
rect 3450 13024 3514 13028
rect 3530 13084 3594 13088
rect 3530 13028 3534 13084
rect 3534 13028 3590 13084
rect 3590 13028 3594 13084
rect 3530 13024 3594 13028
rect 3610 13084 3674 13088
rect 3610 13028 3614 13084
rect 3614 13028 3670 13084
rect 3670 13028 3674 13084
rect 3610 13024 3674 13028
rect 3690 13084 3754 13088
rect 3690 13028 3694 13084
rect 3694 13028 3750 13084
rect 3750 13028 3754 13084
rect 3690 13024 3754 13028
rect 8448 13084 8512 13088
rect 8448 13028 8452 13084
rect 8452 13028 8508 13084
rect 8508 13028 8512 13084
rect 8448 13024 8512 13028
rect 8528 13084 8592 13088
rect 8528 13028 8532 13084
rect 8532 13028 8588 13084
rect 8588 13028 8592 13084
rect 8528 13024 8592 13028
rect 8608 13084 8672 13088
rect 8608 13028 8612 13084
rect 8612 13028 8668 13084
rect 8668 13028 8672 13084
rect 8608 13024 8672 13028
rect 8688 13084 8752 13088
rect 8688 13028 8692 13084
rect 8692 13028 8748 13084
rect 8748 13028 8752 13084
rect 8688 13024 8752 13028
rect 13445 13084 13509 13088
rect 13445 13028 13449 13084
rect 13449 13028 13505 13084
rect 13505 13028 13509 13084
rect 13445 13024 13509 13028
rect 13525 13084 13589 13088
rect 13525 13028 13529 13084
rect 13529 13028 13585 13084
rect 13585 13028 13589 13084
rect 13525 13024 13589 13028
rect 13605 13084 13669 13088
rect 13605 13028 13609 13084
rect 13609 13028 13665 13084
rect 13665 13028 13669 13084
rect 13605 13024 13669 13028
rect 13685 13084 13749 13088
rect 13685 13028 13689 13084
rect 13689 13028 13745 13084
rect 13745 13028 13749 13084
rect 13685 13024 13749 13028
rect 12756 12956 12820 13020
rect 5949 12540 6013 12544
rect 5949 12484 5953 12540
rect 5953 12484 6009 12540
rect 6009 12484 6013 12540
rect 5949 12480 6013 12484
rect 6029 12540 6093 12544
rect 6029 12484 6033 12540
rect 6033 12484 6089 12540
rect 6089 12484 6093 12540
rect 6029 12480 6093 12484
rect 6109 12540 6173 12544
rect 6109 12484 6113 12540
rect 6113 12484 6169 12540
rect 6169 12484 6173 12540
rect 6109 12480 6173 12484
rect 6189 12540 6253 12544
rect 6189 12484 6193 12540
rect 6193 12484 6249 12540
rect 6249 12484 6253 12540
rect 6189 12480 6253 12484
rect 10946 12540 11010 12544
rect 10946 12484 10950 12540
rect 10950 12484 11006 12540
rect 11006 12484 11010 12540
rect 10946 12480 11010 12484
rect 11026 12540 11090 12544
rect 11026 12484 11030 12540
rect 11030 12484 11086 12540
rect 11086 12484 11090 12540
rect 11026 12480 11090 12484
rect 11106 12540 11170 12544
rect 11106 12484 11110 12540
rect 11110 12484 11166 12540
rect 11166 12484 11170 12540
rect 11106 12480 11170 12484
rect 11186 12540 11250 12544
rect 11186 12484 11190 12540
rect 11190 12484 11246 12540
rect 11246 12484 11250 12540
rect 11186 12480 11250 12484
rect 3450 11996 3514 12000
rect 3450 11940 3454 11996
rect 3454 11940 3510 11996
rect 3510 11940 3514 11996
rect 3450 11936 3514 11940
rect 3530 11996 3594 12000
rect 3530 11940 3534 11996
rect 3534 11940 3590 11996
rect 3590 11940 3594 11996
rect 3530 11936 3594 11940
rect 3610 11996 3674 12000
rect 3610 11940 3614 11996
rect 3614 11940 3670 11996
rect 3670 11940 3674 11996
rect 3610 11936 3674 11940
rect 3690 11996 3754 12000
rect 3690 11940 3694 11996
rect 3694 11940 3750 11996
rect 3750 11940 3754 11996
rect 3690 11936 3754 11940
rect 8448 11996 8512 12000
rect 8448 11940 8452 11996
rect 8452 11940 8508 11996
rect 8508 11940 8512 11996
rect 8448 11936 8512 11940
rect 8528 11996 8592 12000
rect 8528 11940 8532 11996
rect 8532 11940 8588 11996
rect 8588 11940 8592 11996
rect 8528 11936 8592 11940
rect 8608 11996 8672 12000
rect 8608 11940 8612 11996
rect 8612 11940 8668 11996
rect 8668 11940 8672 11996
rect 8608 11936 8672 11940
rect 8688 11996 8752 12000
rect 8688 11940 8692 11996
rect 8692 11940 8748 11996
rect 8748 11940 8752 11996
rect 8688 11936 8752 11940
rect 13445 11996 13509 12000
rect 13445 11940 13449 11996
rect 13449 11940 13505 11996
rect 13505 11940 13509 11996
rect 13445 11936 13509 11940
rect 13525 11996 13589 12000
rect 13525 11940 13529 11996
rect 13529 11940 13585 11996
rect 13585 11940 13589 11996
rect 13525 11936 13589 11940
rect 13605 11996 13669 12000
rect 13605 11940 13609 11996
rect 13609 11940 13665 11996
rect 13665 11940 13669 11996
rect 13605 11936 13669 11940
rect 13685 11996 13749 12000
rect 13685 11940 13689 11996
rect 13689 11940 13745 11996
rect 13745 11940 13749 11996
rect 13685 11936 13749 11940
rect 5949 11452 6013 11456
rect 5949 11396 5953 11452
rect 5953 11396 6009 11452
rect 6009 11396 6013 11452
rect 5949 11392 6013 11396
rect 6029 11452 6093 11456
rect 6029 11396 6033 11452
rect 6033 11396 6089 11452
rect 6089 11396 6093 11452
rect 6029 11392 6093 11396
rect 6109 11452 6173 11456
rect 6109 11396 6113 11452
rect 6113 11396 6169 11452
rect 6169 11396 6173 11452
rect 6109 11392 6173 11396
rect 6189 11452 6253 11456
rect 6189 11396 6193 11452
rect 6193 11396 6249 11452
rect 6249 11396 6253 11452
rect 6189 11392 6253 11396
rect 10946 11452 11010 11456
rect 10946 11396 10950 11452
rect 10950 11396 11006 11452
rect 11006 11396 11010 11452
rect 10946 11392 11010 11396
rect 11026 11452 11090 11456
rect 11026 11396 11030 11452
rect 11030 11396 11086 11452
rect 11086 11396 11090 11452
rect 11026 11392 11090 11396
rect 11106 11452 11170 11456
rect 11106 11396 11110 11452
rect 11110 11396 11166 11452
rect 11166 11396 11170 11452
rect 11106 11392 11170 11396
rect 11186 11452 11250 11456
rect 11186 11396 11190 11452
rect 11190 11396 11246 11452
rect 11246 11396 11250 11452
rect 11186 11392 11250 11396
rect 3450 10908 3514 10912
rect 3450 10852 3454 10908
rect 3454 10852 3510 10908
rect 3510 10852 3514 10908
rect 3450 10848 3514 10852
rect 3530 10908 3594 10912
rect 3530 10852 3534 10908
rect 3534 10852 3590 10908
rect 3590 10852 3594 10908
rect 3530 10848 3594 10852
rect 3610 10908 3674 10912
rect 3610 10852 3614 10908
rect 3614 10852 3670 10908
rect 3670 10852 3674 10908
rect 3610 10848 3674 10852
rect 3690 10908 3754 10912
rect 3690 10852 3694 10908
rect 3694 10852 3750 10908
rect 3750 10852 3754 10908
rect 3690 10848 3754 10852
rect 8448 10908 8512 10912
rect 8448 10852 8452 10908
rect 8452 10852 8508 10908
rect 8508 10852 8512 10908
rect 8448 10848 8512 10852
rect 8528 10908 8592 10912
rect 8528 10852 8532 10908
rect 8532 10852 8588 10908
rect 8588 10852 8592 10908
rect 8528 10848 8592 10852
rect 8608 10908 8672 10912
rect 8608 10852 8612 10908
rect 8612 10852 8668 10908
rect 8668 10852 8672 10908
rect 8608 10848 8672 10852
rect 8688 10908 8752 10912
rect 8688 10852 8692 10908
rect 8692 10852 8748 10908
rect 8748 10852 8752 10908
rect 8688 10848 8752 10852
rect 13445 10908 13509 10912
rect 13445 10852 13449 10908
rect 13449 10852 13505 10908
rect 13505 10852 13509 10908
rect 13445 10848 13509 10852
rect 13525 10908 13589 10912
rect 13525 10852 13529 10908
rect 13529 10852 13585 10908
rect 13585 10852 13589 10908
rect 13525 10848 13589 10852
rect 13605 10908 13669 10912
rect 13605 10852 13609 10908
rect 13609 10852 13665 10908
rect 13665 10852 13669 10908
rect 13605 10848 13669 10852
rect 13685 10908 13749 10912
rect 13685 10852 13689 10908
rect 13689 10852 13745 10908
rect 13745 10852 13749 10908
rect 13685 10848 13749 10852
rect 5949 10364 6013 10368
rect 5949 10308 5953 10364
rect 5953 10308 6009 10364
rect 6009 10308 6013 10364
rect 5949 10304 6013 10308
rect 6029 10364 6093 10368
rect 6029 10308 6033 10364
rect 6033 10308 6089 10364
rect 6089 10308 6093 10364
rect 6029 10304 6093 10308
rect 6109 10364 6173 10368
rect 6109 10308 6113 10364
rect 6113 10308 6169 10364
rect 6169 10308 6173 10364
rect 6109 10304 6173 10308
rect 6189 10364 6253 10368
rect 6189 10308 6193 10364
rect 6193 10308 6249 10364
rect 6249 10308 6253 10364
rect 6189 10304 6253 10308
rect 10946 10364 11010 10368
rect 10946 10308 10950 10364
rect 10950 10308 11006 10364
rect 11006 10308 11010 10364
rect 10946 10304 11010 10308
rect 11026 10364 11090 10368
rect 11026 10308 11030 10364
rect 11030 10308 11086 10364
rect 11086 10308 11090 10364
rect 11026 10304 11090 10308
rect 11106 10364 11170 10368
rect 11106 10308 11110 10364
rect 11110 10308 11166 10364
rect 11166 10308 11170 10364
rect 11106 10304 11170 10308
rect 11186 10364 11250 10368
rect 11186 10308 11190 10364
rect 11190 10308 11246 10364
rect 11246 10308 11250 10364
rect 11186 10304 11250 10308
rect 3450 9820 3514 9824
rect 3450 9764 3454 9820
rect 3454 9764 3510 9820
rect 3510 9764 3514 9820
rect 3450 9760 3514 9764
rect 3530 9820 3594 9824
rect 3530 9764 3534 9820
rect 3534 9764 3590 9820
rect 3590 9764 3594 9820
rect 3530 9760 3594 9764
rect 3610 9820 3674 9824
rect 3610 9764 3614 9820
rect 3614 9764 3670 9820
rect 3670 9764 3674 9820
rect 3610 9760 3674 9764
rect 3690 9820 3754 9824
rect 3690 9764 3694 9820
rect 3694 9764 3750 9820
rect 3750 9764 3754 9820
rect 3690 9760 3754 9764
rect 8448 9820 8512 9824
rect 8448 9764 8452 9820
rect 8452 9764 8508 9820
rect 8508 9764 8512 9820
rect 8448 9760 8512 9764
rect 8528 9820 8592 9824
rect 8528 9764 8532 9820
rect 8532 9764 8588 9820
rect 8588 9764 8592 9820
rect 8528 9760 8592 9764
rect 8608 9820 8672 9824
rect 8608 9764 8612 9820
rect 8612 9764 8668 9820
rect 8668 9764 8672 9820
rect 8608 9760 8672 9764
rect 8688 9820 8752 9824
rect 8688 9764 8692 9820
rect 8692 9764 8748 9820
rect 8748 9764 8752 9820
rect 8688 9760 8752 9764
rect 13445 9820 13509 9824
rect 13445 9764 13449 9820
rect 13449 9764 13505 9820
rect 13505 9764 13509 9820
rect 13445 9760 13509 9764
rect 13525 9820 13589 9824
rect 13525 9764 13529 9820
rect 13529 9764 13585 9820
rect 13585 9764 13589 9820
rect 13525 9760 13589 9764
rect 13605 9820 13669 9824
rect 13605 9764 13609 9820
rect 13609 9764 13665 9820
rect 13665 9764 13669 9820
rect 13605 9760 13669 9764
rect 13685 9820 13749 9824
rect 13685 9764 13689 9820
rect 13689 9764 13745 9820
rect 13745 9764 13749 9820
rect 13685 9760 13749 9764
rect 5949 9276 6013 9280
rect 5949 9220 5953 9276
rect 5953 9220 6009 9276
rect 6009 9220 6013 9276
rect 5949 9216 6013 9220
rect 6029 9276 6093 9280
rect 6029 9220 6033 9276
rect 6033 9220 6089 9276
rect 6089 9220 6093 9276
rect 6029 9216 6093 9220
rect 6109 9276 6173 9280
rect 6109 9220 6113 9276
rect 6113 9220 6169 9276
rect 6169 9220 6173 9276
rect 6109 9216 6173 9220
rect 6189 9276 6253 9280
rect 6189 9220 6193 9276
rect 6193 9220 6249 9276
rect 6249 9220 6253 9276
rect 6189 9216 6253 9220
rect 10946 9276 11010 9280
rect 10946 9220 10950 9276
rect 10950 9220 11006 9276
rect 11006 9220 11010 9276
rect 10946 9216 11010 9220
rect 11026 9276 11090 9280
rect 11026 9220 11030 9276
rect 11030 9220 11086 9276
rect 11086 9220 11090 9276
rect 11026 9216 11090 9220
rect 11106 9276 11170 9280
rect 11106 9220 11110 9276
rect 11110 9220 11166 9276
rect 11166 9220 11170 9276
rect 11106 9216 11170 9220
rect 11186 9276 11250 9280
rect 11186 9220 11190 9276
rect 11190 9220 11246 9276
rect 11246 9220 11250 9276
rect 11186 9216 11250 9220
rect 8892 8876 8956 8940
rect 3450 8732 3514 8736
rect 3450 8676 3454 8732
rect 3454 8676 3510 8732
rect 3510 8676 3514 8732
rect 3450 8672 3514 8676
rect 3530 8732 3594 8736
rect 3530 8676 3534 8732
rect 3534 8676 3590 8732
rect 3590 8676 3594 8732
rect 3530 8672 3594 8676
rect 3610 8732 3674 8736
rect 3610 8676 3614 8732
rect 3614 8676 3670 8732
rect 3670 8676 3674 8732
rect 3610 8672 3674 8676
rect 3690 8732 3754 8736
rect 3690 8676 3694 8732
rect 3694 8676 3750 8732
rect 3750 8676 3754 8732
rect 3690 8672 3754 8676
rect 8448 8732 8512 8736
rect 8448 8676 8452 8732
rect 8452 8676 8508 8732
rect 8508 8676 8512 8732
rect 8448 8672 8512 8676
rect 8528 8732 8592 8736
rect 8528 8676 8532 8732
rect 8532 8676 8588 8732
rect 8588 8676 8592 8732
rect 8528 8672 8592 8676
rect 8608 8732 8672 8736
rect 8608 8676 8612 8732
rect 8612 8676 8668 8732
rect 8668 8676 8672 8732
rect 8608 8672 8672 8676
rect 8688 8732 8752 8736
rect 8688 8676 8692 8732
rect 8692 8676 8748 8732
rect 8748 8676 8752 8732
rect 8688 8672 8752 8676
rect 13445 8732 13509 8736
rect 13445 8676 13449 8732
rect 13449 8676 13505 8732
rect 13505 8676 13509 8732
rect 13445 8672 13509 8676
rect 13525 8732 13589 8736
rect 13525 8676 13529 8732
rect 13529 8676 13585 8732
rect 13585 8676 13589 8732
rect 13525 8672 13589 8676
rect 13605 8732 13669 8736
rect 13605 8676 13609 8732
rect 13609 8676 13665 8732
rect 13665 8676 13669 8732
rect 13605 8672 13669 8676
rect 13685 8732 13749 8736
rect 13685 8676 13689 8732
rect 13689 8676 13745 8732
rect 13745 8676 13749 8732
rect 13685 8672 13749 8676
rect 5949 8188 6013 8192
rect 5949 8132 5953 8188
rect 5953 8132 6009 8188
rect 6009 8132 6013 8188
rect 5949 8128 6013 8132
rect 6029 8188 6093 8192
rect 6029 8132 6033 8188
rect 6033 8132 6089 8188
rect 6089 8132 6093 8188
rect 6029 8128 6093 8132
rect 6109 8188 6173 8192
rect 6109 8132 6113 8188
rect 6113 8132 6169 8188
rect 6169 8132 6173 8188
rect 6109 8128 6173 8132
rect 6189 8188 6253 8192
rect 6189 8132 6193 8188
rect 6193 8132 6249 8188
rect 6249 8132 6253 8188
rect 6189 8128 6253 8132
rect 10946 8188 11010 8192
rect 10946 8132 10950 8188
rect 10950 8132 11006 8188
rect 11006 8132 11010 8188
rect 10946 8128 11010 8132
rect 11026 8188 11090 8192
rect 11026 8132 11030 8188
rect 11030 8132 11086 8188
rect 11086 8132 11090 8188
rect 11026 8128 11090 8132
rect 11106 8188 11170 8192
rect 11106 8132 11110 8188
rect 11110 8132 11166 8188
rect 11166 8132 11170 8188
rect 11106 8128 11170 8132
rect 11186 8188 11250 8192
rect 11186 8132 11190 8188
rect 11190 8132 11246 8188
rect 11246 8132 11250 8188
rect 11186 8128 11250 8132
rect 3450 7644 3514 7648
rect 3450 7588 3454 7644
rect 3454 7588 3510 7644
rect 3510 7588 3514 7644
rect 3450 7584 3514 7588
rect 3530 7644 3594 7648
rect 3530 7588 3534 7644
rect 3534 7588 3590 7644
rect 3590 7588 3594 7644
rect 3530 7584 3594 7588
rect 3610 7644 3674 7648
rect 3610 7588 3614 7644
rect 3614 7588 3670 7644
rect 3670 7588 3674 7644
rect 3610 7584 3674 7588
rect 3690 7644 3754 7648
rect 3690 7588 3694 7644
rect 3694 7588 3750 7644
rect 3750 7588 3754 7644
rect 3690 7584 3754 7588
rect 8448 7644 8512 7648
rect 8448 7588 8452 7644
rect 8452 7588 8508 7644
rect 8508 7588 8512 7644
rect 8448 7584 8512 7588
rect 8528 7644 8592 7648
rect 8528 7588 8532 7644
rect 8532 7588 8588 7644
rect 8588 7588 8592 7644
rect 8528 7584 8592 7588
rect 8608 7644 8672 7648
rect 8608 7588 8612 7644
rect 8612 7588 8668 7644
rect 8668 7588 8672 7644
rect 8608 7584 8672 7588
rect 8688 7644 8752 7648
rect 8688 7588 8692 7644
rect 8692 7588 8748 7644
rect 8748 7588 8752 7644
rect 8688 7584 8752 7588
rect 13445 7644 13509 7648
rect 13445 7588 13449 7644
rect 13449 7588 13505 7644
rect 13505 7588 13509 7644
rect 13445 7584 13509 7588
rect 13525 7644 13589 7648
rect 13525 7588 13529 7644
rect 13529 7588 13585 7644
rect 13585 7588 13589 7644
rect 13525 7584 13589 7588
rect 13605 7644 13669 7648
rect 13605 7588 13609 7644
rect 13609 7588 13665 7644
rect 13665 7588 13669 7644
rect 13605 7584 13669 7588
rect 13685 7644 13749 7648
rect 13685 7588 13689 7644
rect 13689 7588 13745 7644
rect 13745 7588 13749 7644
rect 13685 7584 13749 7588
rect 5949 7100 6013 7104
rect 5949 7044 5953 7100
rect 5953 7044 6009 7100
rect 6009 7044 6013 7100
rect 5949 7040 6013 7044
rect 6029 7100 6093 7104
rect 6029 7044 6033 7100
rect 6033 7044 6089 7100
rect 6089 7044 6093 7100
rect 6029 7040 6093 7044
rect 6109 7100 6173 7104
rect 6109 7044 6113 7100
rect 6113 7044 6169 7100
rect 6169 7044 6173 7100
rect 6109 7040 6173 7044
rect 6189 7100 6253 7104
rect 6189 7044 6193 7100
rect 6193 7044 6249 7100
rect 6249 7044 6253 7100
rect 6189 7040 6253 7044
rect 10946 7100 11010 7104
rect 10946 7044 10950 7100
rect 10950 7044 11006 7100
rect 11006 7044 11010 7100
rect 10946 7040 11010 7044
rect 11026 7100 11090 7104
rect 11026 7044 11030 7100
rect 11030 7044 11086 7100
rect 11086 7044 11090 7100
rect 11026 7040 11090 7044
rect 11106 7100 11170 7104
rect 11106 7044 11110 7100
rect 11110 7044 11166 7100
rect 11166 7044 11170 7100
rect 11106 7040 11170 7044
rect 11186 7100 11250 7104
rect 11186 7044 11190 7100
rect 11190 7044 11246 7100
rect 11246 7044 11250 7100
rect 11186 7040 11250 7044
rect 6684 6624 6748 6628
rect 6684 6568 6734 6624
rect 6734 6568 6748 6624
rect 6684 6564 6748 6568
rect 3450 6556 3514 6560
rect 3450 6500 3454 6556
rect 3454 6500 3510 6556
rect 3510 6500 3514 6556
rect 3450 6496 3514 6500
rect 3530 6556 3594 6560
rect 3530 6500 3534 6556
rect 3534 6500 3590 6556
rect 3590 6500 3594 6556
rect 3530 6496 3594 6500
rect 3610 6556 3674 6560
rect 3610 6500 3614 6556
rect 3614 6500 3670 6556
rect 3670 6500 3674 6556
rect 3610 6496 3674 6500
rect 3690 6556 3754 6560
rect 3690 6500 3694 6556
rect 3694 6500 3750 6556
rect 3750 6500 3754 6556
rect 3690 6496 3754 6500
rect 8448 6556 8512 6560
rect 8448 6500 8452 6556
rect 8452 6500 8508 6556
rect 8508 6500 8512 6556
rect 8448 6496 8512 6500
rect 8528 6556 8592 6560
rect 8528 6500 8532 6556
rect 8532 6500 8588 6556
rect 8588 6500 8592 6556
rect 8528 6496 8592 6500
rect 8608 6556 8672 6560
rect 8608 6500 8612 6556
rect 8612 6500 8668 6556
rect 8668 6500 8672 6556
rect 8608 6496 8672 6500
rect 8688 6556 8752 6560
rect 8688 6500 8692 6556
rect 8692 6500 8748 6556
rect 8748 6500 8752 6556
rect 8688 6496 8752 6500
rect 13445 6556 13509 6560
rect 13445 6500 13449 6556
rect 13449 6500 13505 6556
rect 13505 6500 13509 6556
rect 13445 6496 13509 6500
rect 13525 6556 13589 6560
rect 13525 6500 13529 6556
rect 13529 6500 13585 6556
rect 13585 6500 13589 6556
rect 13525 6496 13589 6500
rect 13605 6556 13669 6560
rect 13605 6500 13609 6556
rect 13609 6500 13665 6556
rect 13665 6500 13669 6556
rect 13605 6496 13669 6500
rect 13685 6556 13749 6560
rect 13685 6500 13689 6556
rect 13689 6500 13745 6556
rect 13745 6500 13749 6556
rect 13685 6496 13749 6500
rect 5949 6012 6013 6016
rect 5949 5956 5953 6012
rect 5953 5956 6009 6012
rect 6009 5956 6013 6012
rect 5949 5952 6013 5956
rect 6029 6012 6093 6016
rect 6029 5956 6033 6012
rect 6033 5956 6089 6012
rect 6089 5956 6093 6012
rect 6029 5952 6093 5956
rect 6109 6012 6173 6016
rect 6109 5956 6113 6012
rect 6113 5956 6169 6012
rect 6169 5956 6173 6012
rect 6109 5952 6173 5956
rect 6189 6012 6253 6016
rect 6189 5956 6193 6012
rect 6193 5956 6249 6012
rect 6249 5956 6253 6012
rect 6189 5952 6253 5956
rect 10946 6012 11010 6016
rect 10946 5956 10950 6012
rect 10950 5956 11006 6012
rect 11006 5956 11010 6012
rect 10946 5952 11010 5956
rect 11026 6012 11090 6016
rect 11026 5956 11030 6012
rect 11030 5956 11086 6012
rect 11086 5956 11090 6012
rect 11026 5952 11090 5956
rect 11106 6012 11170 6016
rect 11106 5956 11110 6012
rect 11110 5956 11166 6012
rect 11166 5956 11170 6012
rect 11106 5952 11170 5956
rect 11186 6012 11250 6016
rect 11186 5956 11190 6012
rect 11190 5956 11246 6012
rect 11246 5956 11250 6012
rect 11186 5952 11250 5956
rect 8892 5476 8956 5540
rect 3450 5468 3514 5472
rect 3450 5412 3454 5468
rect 3454 5412 3510 5468
rect 3510 5412 3514 5468
rect 3450 5408 3514 5412
rect 3530 5468 3594 5472
rect 3530 5412 3534 5468
rect 3534 5412 3590 5468
rect 3590 5412 3594 5468
rect 3530 5408 3594 5412
rect 3610 5468 3674 5472
rect 3610 5412 3614 5468
rect 3614 5412 3670 5468
rect 3670 5412 3674 5468
rect 3610 5408 3674 5412
rect 3690 5468 3754 5472
rect 3690 5412 3694 5468
rect 3694 5412 3750 5468
rect 3750 5412 3754 5468
rect 3690 5408 3754 5412
rect 8448 5468 8512 5472
rect 8448 5412 8452 5468
rect 8452 5412 8508 5468
rect 8508 5412 8512 5468
rect 8448 5408 8512 5412
rect 8528 5468 8592 5472
rect 8528 5412 8532 5468
rect 8532 5412 8588 5468
rect 8588 5412 8592 5468
rect 8528 5408 8592 5412
rect 8608 5468 8672 5472
rect 8608 5412 8612 5468
rect 8612 5412 8668 5468
rect 8668 5412 8672 5468
rect 8608 5408 8672 5412
rect 8688 5468 8752 5472
rect 8688 5412 8692 5468
rect 8692 5412 8748 5468
rect 8748 5412 8752 5468
rect 8688 5408 8752 5412
rect 13445 5468 13509 5472
rect 13445 5412 13449 5468
rect 13449 5412 13505 5468
rect 13505 5412 13509 5468
rect 13445 5408 13509 5412
rect 13525 5468 13589 5472
rect 13525 5412 13529 5468
rect 13529 5412 13585 5468
rect 13585 5412 13589 5468
rect 13525 5408 13589 5412
rect 13605 5468 13669 5472
rect 13605 5412 13609 5468
rect 13609 5412 13665 5468
rect 13665 5412 13669 5468
rect 13605 5408 13669 5412
rect 13685 5468 13749 5472
rect 13685 5412 13689 5468
rect 13689 5412 13745 5468
rect 13745 5412 13749 5468
rect 13685 5408 13749 5412
rect 11468 5340 11532 5404
rect 5949 4924 6013 4928
rect 5949 4868 5953 4924
rect 5953 4868 6009 4924
rect 6009 4868 6013 4924
rect 5949 4864 6013 4868
rect 6029 4924 6093 4928
rect 6029 4868 6033 4924
rect 6033 4868 6089 4924
rect 6089 4868 6093 4924
rect 6029 4864 6093 4868
rect 6109 4924 6173 4928
rect 6109 4868 6113 4924
rect 6113 4868 6169 4924
rect 6169 4868 6173 4924
rect 6109 4864 6173 4868
rect 6189 4924 6253 4928
rect 6189 4868 6193 4924
rect 6193 4868 6249 4924
rect 6249 4868 6253 4924
rect 6189 4864 6253 4868
rect 10946 4924 11010 4928
rect 10946 4868 10950 4924
rect 10950 4868 11006 4924
rect 11006 4868 11010 4924
rect 10946 4864 11010 4868
rect 11026 4924 11090 4928
rect 11026 4868 11030 4924
rect 11030 4868 11086 4924
rect 11086 4868 11090 4924
rect 11026 4864 11090 4868
rect 11106 4924 11170 4928
rect 11106 4868 11110 4924
rect 11110 4868 11166 4924
rect 11166 4868 11170 4924
rect 11106 4864 11170 4868
rect 11186 4924 11250 4928
rect 11186 4868 11190 4924
rect 11190 4868 11246 4924
rect 11246 4868 11250 4924
rect 11186 4864 11250 4868
rect 4108 4796 4172 4860
rect 3450 4380 3514 4384
rect 3450 4324 3454 4380
rect 3454 4324 3510 4380
rect 3510 4324 3514 4380
rect 3450 4320 3514 4324
rect 3530 4380 3594 4384
rect 3530 4324 3534 4380
rect 3534 4324 3590 4380
rect 3590 4324 3594 4380
rect 3530 4320 3594 4324
rect 3610 4380 3674 4384
rect 3610 4324 3614 4380
rect 3614 4324 3670 4380
rect 3670 4324 3674 4380
rect 3610 4320 3674 4324
rect 3690 4380 3754 4384
rect 3690 4324 3694 4380
rect 3694 4324 3750 4380
rect 3750 4324 3754 4380
rect 3690 4320 3754 4324
rect 8448 4380 8512 4384
rect 8448 4324 8452 4380
rect 8452 4324 8508 4380
rect 8508 4324 8512 4380
rect 8448 4320 8512 4324
rect 8528 4380 8592 4384
rect 8528 4324 8532 4380
rect 8532 4324 8588 4380
rect 8588 4324 8592 4380
rect 8528 4320 8592 4324
rect 8608 4380 8672 4384
rect 8608 4324 8612 4380
rect 8612 4324 8668 4380
rect 8668 4324 8672 4380
rect 8608 4320 8672 4324
rect 8688 4380 8752 4384
rect 8688 4324 8692 4380
rect 8692 4324 8748 4380
rect 8748 4324 8752 4380
rect 8688 4320 8752 4324
rect 13445 4380 13509 4384
rect 13445 4324 13449 4380
rect 13449 4324 13505 4380
rect 13505 4324 13509 4380
rect 13445 4320 13509 4324
rect 13525 4380 13589 4384
rect 13525 4324 13529 4380
rect 13529 4324 13585 4380
rect 13585 4324 13589 4380
rect 13525 4320 13589 4324
rect 13605 4380 13669 4384
rect 13605 4324 13609 4380
rect 13609 4324 13665 4380
rect 13665 4324 13669 4380
rect 13605 4320 13669 4324
rect 13685 4380 13749 4384
rect 13685 4324 13689 4380
rect 13689 4324 13745 4380
rect 13745 4324 13749 4380
rect 13685 4320 13749 4324
rect 12572 4312 12636 4316
rect 12572 4256 12622 4312
rect 12622 4256 12636 4312
rect 12572 4252 12636 4256
rect 5949 3836 6013 3840
rect 5949 3780 5953 3836
rect 5953 3780 6009 3836
rect 6009 3780 6013 3836
rect 5949 3776 6013 3780
rect 6029 3836 6093 3840
rect 6029 3780 6033 3836
rect 6033 3780 6089 3836
rect 6089 3780 6093 3836
rect 6029 3776 6093 3780
rect 6109 3836 6173 3840
rect 6109 3780 6113 3836
rect 6113 3780 6169 3836
rect 6169 3780 6173 3836
rect 6109 3776 6173 3780
rect 6189 3836 6253 3840
rect 6189 3780 6193 3836
rect 6193 3780 6249 3836
rect 6249 3780 6253 3836
rect 6189 3776 6253 3780
rect 10946 3836 11010 3840
rect 10946 3780 10950 3836
rect 10950 3780 11006 3836
rect 11006 3780 11010 3836
rect 10946 3776 11010 3780
rect 11026 3836 11090 3840
rect 11026 3780 11030 3836
rect 11030 3780 11086 3836
rect 11086 3780 11090 3836
rect 11026 3776 11090 3780
rect 11106 3836 11170 3840
rect 11106 3780 11110 3836
rect 11110 3780 11166 3836
rect 11166 3780 11170 3836
rect 11106 3776 11170 3780
rect 11186 3836 11250 3840
rect 11186 3780 11190 3836
rect 11190 3780 11246 3836
rect 11246 3780 11250 3836
rect 11186 3776 11250 3780
rect 6684 3768 6748 3772
rect 6684 3712 6698 3768
rect 6698 3712 6748 3768
rect 6684 3708 6748 3712
rect 3450 3292 3514 3296
rect 3450 3236 3454 3292
rect 3454 3236 3510 3292
rect 3510 3236 3514 3292
rect 3450 3232 3514 3236
rect 3530 3292 3594 3296
rect 3530 3236 3534 3292
rect 3534 3236 3590 3292
rect 3590 3236 3594 3292
rect 3530 3232 3594 3236
rect 3610 3292 3674 3296
rect 3610 3236 3614 3292
rect 3614 3236 3670 3292
rect 3670 3236 3674 3292
rect 3610 3232 3674 3236
rect 3690 3292 3754 3296
rect 3690 3236 3694 3292
rect 3694 3236 3750 3292
rect 3750 3236 3754 3292
rect 3690 3232 3754 3236
rect 8448 3292 8512 3296
rect 8448 3236 8452 3292
rect 8452 3236 8508 3292
rect 8508 3236 8512 3292
rect 8448 3232 8512 3236
rect 8528 3292 8592 3296
rect 8528 3236 8532 3292
rect 8532 3236 8588 3292
rect 8588 3236 8592 3292
rect 8528 3232 8592 3236
rect 8608 3292 8672 3296
rect 8608 3236 8612 3292
rect 8612 3236 8668 3292
rect 8668 3236 8672 3292
rect 8608 3232 8672 3236
rect 8688 3292 8752 3296
rect 8688 3236 8692 3292
rect 8692 3236 8748 3292
rect 8748 3236 8752 3292
rect 8688 3232 8752 3236
rect 13445 3292 13509 3296
rect 13445 3236 13449 3292
rect 13449 3236 13505 3292
rect 13505 3236 13509 3292
rect 13445 3232 13509 3236
rect 13525 3292 13589 3296
rect 13525 3236 13529 3292
rect 13529 3236 13585 3292
rect 13585 3236 13589 3292
rect 13525 3232 13589 3236
rect 13605 3292 13669 3296
rect 13605 3236 13609 3292
rect 13609 3236 13665 3292
rect 13665 3236 13669 3292
rect 13605 3232 13669 3236
rect 13685 3292 13749 3296
rect 13685 3236 13689 3292
rect 13689 3236 13745 3292
rect 13745 3236 13749 3292
rect 13685 3232 13749 3236
rect 5949 2748 6013 2752
rect 5949 2692 5953 2748
rect 5953 2692 6009 2748
rect 6009 2692 6013 2748
rect 5949 2688 6013 2692
rect 6029 2748 6093 2752
rect 6029 2692 6033 2748
rect 6033 2692 6089 2748
rect 6089 2692 6093 2748
rect 6029 2688 6093 2692
rect 6109 2748 6173 2752
rect 6109 2692 6113 2748
rect 6113 2692 6169 2748
rect 6169 2692 6173 2748
rect 6109 2688 6173 2692
rect 6189 2748 6253 2752
rect 6189 2692 6193 2748
rect 6193 2692 6249 2748
rect 6249 2692 6253 2748
rect 6189 2688 6253 2692
rect 10946 2748 11010 2752
rect 10946 2692 10950 2748
rect 10950 2692 11006 2748
rect 11006 2692 11010 2748
rect 10946 2688 11010 2692
rect 11026 2748 11090 2752
rect 11026 2692 11030 2748
rect 11030 2692 11086 2748
rect 11086 2692 11090 2748
rect 11026 2688 11090 2692
rect 11106 2748 11170 2752
rect 11106 2692 11110 2748
rect 11110 2692 11166 2748
rect 11166 2692 11170 2748
rect 11106 2688 11170 2692
rect 11186 2748 11250 2752
rect 11186 2692 11190 2748
rect 11190 2692 11246 2748
rect 11246 2692 11250 2748
rect 11186 2688 11250 2692
rect 12572 2680 12636 2684
rect 12572 2624 12622 2680
rect 12622 2624 12636 2680
rect 12572 2620 12636 2624
rect 4108 2544 4172 2548
rect 4108 2488 4122 2544
rect 4122 2488 4172 2544
rect 4108 2484 4172 2488
rect 11468 2484 11532 2548
rect 3450 2204 3514 2208
rect 3450 2148 3454 2204
rect 3454 2148 3510 2204
rect 3510 2148 3514 2204
rect 3450 2144 3514 2148
rect 3530 2204 3594 2208
rect 3530 2148 3534 2204
rect 3534 2148 3590 2204
rect 3590 2148 3594 2204
rect 3530 2144 3594 2148
rect 3610 2204 3674 2208
rect 3610 2148 3614 2204
rect 3614 2148 3670 2204
rect 3670 2148 3674 2204
rect 3610 2144 3674 2148
rect 3690 2204 3754 2208
rect 3690 2148 3694 2204
rect 3694 2148 3750 2204
rect 3750 2148 3754 2204
rect 3690 2144 3754 2148
rect 8448 2204 8512 2208
rect 8448 2148 8452 2204
rect 8452 2148 8508 2204
rect 8508 2148 8512 2204
rect 8448 2144 8512 2148
rect 8528 2204 8592 2208
rect 8528 2148 8532 2204
rect 8532 2148 8588 2204
rect 8588 2148 8592 2204
rect 8528 2144 8592 2148
rect 8608 2204 8672 2208
rect 8608 2148 8612 2204
rect 8612 2148 8668 2204
rect 8668 2148 8672 2204
rect 8608 2144 8672 2148
rect 8688 2204 8752 2208
rect 8688 2148 8692 2204
rect 8692 2148 8748 2204
rect 8748 2148 8752 2204
rect 8688 2144 8752 2148
rect 13445 2204 13509 2208
rect 13445 2148 13449 2204
rect 13449 2148 13505 2204
rect 13505 2148 13509 2204
rect 13445 2144 13509 2148
rect 13525 2204 13589 2208
rect 13525 2148 13529 2204
rect 13529 2148 13585 2204
rect 13585 2148 13589 2204
rect 13525 2144 13589 2148
rect 13605 2204 13669 2208
rect 13605 2148 13609 2204
rect 13609 2148 13665 2204
rect 13665 2148 13669 2204
rect 13605 2144 13669 2148
rect 13685 2204 13749 2208
rect 13685 2148 13689 2204
rect 13689 2148 13745 2204
rect 13745 2148 13749 2204
rect 13685 2144 13749 2148
<< metal4 >>
rect 3442 17440 3763 17456
rect 3442 17376 3450 17440
rect 3514 17376 3530 17440
rect 3594 17376 3610 17440
rect 3674 17376 3690 17440
rect 3754 17376 3763 17440
rect 3442 16352 3763 17376
rect 3442 16288 3450 16352
rect 3514 16288 3530 16352
rect 3594 16288 3610 16352
rect 3674 16288 3690 16352
rect 3754 16288 3763 16352
rect 3442 15264 3763 16288
rect 3442 15200 3450 15264
rect 3514 15200 3530 15264
rect 3594 15200 3610 15264
rect 3674 15200 3690 15264
rect 3754 15200 3763 15264
rect 3442 14176 3763 15200
rect 3442 14112 3450 14176
rect 3514 14112 3530 14176
rect 3594 14112 3610 14176
rect 3674 14112 3690 14176
rect 3754 14112 3763 14176
rect 3442 13088 3763 14112
rect 3442 13024 3450 13088
rect 3514 13024 3530 13088
rect 3594 13024 3610 13088
rect 3674 13024 3690 13088
rect 3754 13024 3763 13088
rect 3442 12000 3763 13024
rect 3442 11936 3450 12000
rect 3514 11936 3530 12000
rect 3594 11936 3610 12000
rect 3674 11936 3690 12000
rect 3754 11936 3763 12000
rect 3442 10912 3763 11936
rect 3442 10848 3450 10912
rect 3514 10848 3530 10912
rect 3594 10848 3610 10912
rect 3674 10848 3690 10912
rect 3754 10848 3763 10912
rect 3442 9824 3763 10848
rect 3442 9760 3450 9824
rect 3514 9760 3530 9824
rect 3594 9760 3610 9824
rect 3674 9760 3690 9824
rect 3754 9760 3763 9824
rect 3442 8736 3763 9760
rect 3442 8672 3450 8736
rect 3514 8672 3530 8736
rect 3594 8672 3610 8736
rect 3674 8672 3690 8736
rect 3754 8672 3763 8736
rect 3442 7648 3763 8672
rect 3442 7584 3450 7648
rect 3514 7584 3530 7648
rect 3594 7584 3610 7648
rect 3674 7584 3690 7648
rect 3754 7584 3763 7648
rect 3442 6560 3763 7584
rect 3442 6496 3450 6560
rect 3514 6496 3530 6560
rect 3594 6496 3610 6560
rect 3674 6496 3690 6560
rect 3754 6496 3763 6560
rect 3442 5472 3763 6496
rect 3442 5408 3450 5472
rect 3514 5408 3530 5472
rect 3594 5408 3610 5472
rect 3674 5408 3690 5472
rect 3754 5408 3763 5472
rect 3442 4384 3763 5408
rect 5941 16896 6261 17456
rect 5941 16832 5949 16896
rect 6013 16832 6029 16896
rect 6093 16832 6109 16896
rect 6173 16832 6189 16896
rect 6253 16832 6261 16896
rect 5941 15808 6261 16832
rect 5941 15744 5949 15808
rect 6013 15744 6029 15808
rect 6093 15744 6109 15808
rect 6173 15744 6189 15808
rect 6253 15744 6261 15808
rect 5941 14720 6261 15744
rect 5941 14656 5949 14720
rect 6013 14656 6029 14720
rect 6093 14656 6109 14720
rect 6173 14656 6189 14720
rect 6253 14656 6261 14720
rect 5941 13632 6261 14656
rect 5941 13568 5949 13632
rect 6013 13568 6029 13632
rect 6093 13568 6109 13632
rect 6173 13568 6189 13632
rect 6253 13568 6261 13632
rect 5941 12544 6261 13568
rect 5941 12480 5949 12544
rect 6013 12480 6029 12544
rect 6093 12480 6109 12544
rect 6173 12480 6189 12544
rect 6253 12480 6261 12544
rect 5941 11456 6261 12480
rect 5941 11392 5949 11456
rect 6013 11392 6029 11456
rect 6093 11392 6109 11456
rect 6173 11392 6189 11456
rect 6253 11392 6261 11456
rect 5941 10368 6261 11392
rect 5941 10304 5949 10368
rect 6013 10304 6029 10368
rect 6093 10304 6109 10368
rect 6173 10304 6189 10368
rect 6253 10304 6261 10368
rect 5941 9280 6261 10304
rect 5941 9216 5949 9280
rect 6013 9216 6029 9280
rect 6093 9216 6109 9280
rect 6173 9216 6189 9280
rect 6253 9216 6261 9280
rect 5941 8192 6261 9216
rect 5941 8128 5949 8192
rect 6013 8128 6029 8192
rect 6093 8128 6109 8192
rect 6173 8128 6189 8192
rect 6253 8128 6261 8192
rect 5941 7104 6261 8128
rect 5941 7040 5949 7104
rect 6013 7040 6029 7104
rect 6093 7040 6109 7104
rect 6173 7040 6189 7104
rect 6253 7040 6261 7104
rect 5941 6016 6261 7040
rect 8440 17440 8760 17456
rect 8440 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8760 17440
rect 8440 16352 8760 17376
rect 8440 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8760 16352
rect 8440 15264 8760 16288
rect 8440 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8760 15264
rect 8440 14176 8760 15200
rect 8440 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8760 14176
rect 8440 13088 8760 14112
rect 8440 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8760 13088
rect 8440 12000 8760 13024
rect 8440 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8760 12000
rect 8440 10912 8760 11936
rect 8440 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8760 10912
rect 8440 9824 8760 10848
rect 8440 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8760 9824
rect 8440 8736 8760 9760
rect 10938 16896 11259 17456
rect 10938 16832 10946 16896
rect 11010 16832 11026 16896
rect 11090 16832 11106 16896
rect 11170 16832 11186 16896
rect 11250 16832 11259 16896
rect 10938 15808 11259 16832
rect 13437 17440 13757 17456
rect 13437 17376 13445 17440
rect 13509 17376 13525 17440
rect 13589 17376 13605 17440
rect 13669 17376 13685 17440
rect 13749 17376 13757 17440
rect 13437 16352 13757 17376
rect 13437 16288 13445 16352
rect 13509 16288 13525 16352
rect 13589 16288 13605 16352
rect 13669 16288 13685 16352
rect 13749 16288 13757 16352
rect 12755 16148 12821 16149
rect 12755 16084 12756 16148
rect 12820 16084 12821 16148
rect 12755 16083 12821 16084
rect 10938 15744 10946 15808
rect 11010 15744 11026 15808
rect 11090 15744 11106 15808
rect 11170 15744 11186 15808
rect 11250 15744 11259 15808
rect 10938 14720 11259 15744
rect 10938 14656 10946 14720
rect 11010 14656 11026 14720
rect 11090 14656 11106 14720
rect 11170 14656 11186 14720
rect 11250 14656 11259 14720
rect 10938 13632 11259 14656
rect 10938 13568 10946 13632
rect 11010 13568 11026 13632
rect 11090 13568 11106 13632
rect 11170 13568 11186 13632
rect 11250 13568 11259 13632
rect 10938 12544 11259 13568
rect 12758 13021 12818 16083
rect 13437 15264 13757 16288
rect 13437 15200 13445 15264
rect 13509 15200 13525 15264
rect 13589 15200 13605 15264
rect 13669 15200 13685 15264
rect 13749 15200 13757 15264
rect 13437 14176 13757 15200
rect 13437 14112 13445 14176
rect 13509 14112 13525 14176
rect 13589 14112 13605 14176
rect 13669 14112 13685 14176
rect 13749 14112 13757 14176
rect 13437 13088 13757 14112
rect 13437 13024 13445 13088
rect 13509 13024 13525 13088
rect 13589 13024 13605 13088
rect 13669 13024 13685 13088
rect 13749 13024 13757 13088
rect 12755 13020 12821 13021
rect 12755 12956 12756 13020
rect 12820 12956 12821 13020
rect 12755 12955 12821 12956
rect 10938 12480 10946 12544
rect 11010 12480 11026 12544
rect 11090 12480 11106 12544
rect 11170 12480 11186 12544
rect 11250 12480 11259 12544
rect 10938 11456 11259 12480
rect 10938 11392 10946 11456
rect 11010 11392 11026 11456
rect 11090 11392 11106 11456
rect 11170 11392 11186 11456
rect 11250 11392 11259 11456
rect 10938 10368 11259 11392
rect 10938 10304 10946 10368
rect 11010 10304 11026 10368
rect 11090 10304 11106 10368
rect 11170 10304 11186 10368
rect 11250 10304 11259 10368
rect 10938 9280 11259 10304
rect 10938 9216 10946 9280
rect 11010 9216 11026 9280
rect 11090 9216 11106 9280
rect 11170 9216 11186 9280
rect 11250 9216 11259 9280
rect 8891 8940 8957 8941
rect 8891 8876 8892 8940
rect 8956 8876 8957 8940
rect 8891 8875 8957 8876
rect 8440 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8760 8736
rect 8440 7648 8760 8672
rect 8440 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8760 7648
rect 6683 6628 6749 6629
rect 6683 6564 6684 6628
rect 6748 6564 6749 6628
rect 6683 6563 6749 6564
rect 5941 5952 5949 6016
rect 6013 5952 6029 6016
rect 6093 5952 6109 6016
rect 6173 5952 6189 6016
rect 6253 5952 6261 6016
rect 5941 4928 6261 5952
rect 5941 4864 5949 4928
rect 6013 4864 6029 4928
rect 6093 4864 6109 4928
rect 6173 4864 6189 4928
rect 6253 4864 6261 4928
rect 4107 4860 4173 4861
rect 4107 4796 4108 4860
rect 4172 4796 4173 4860
rect 4107 4795 4173 4796
rect 3442 4320 3450 4384
rect 3514 4320 3530 4384
rect 3594 4320 3610 4384
rect 3674 4320 3690 4384
rect 3754 4320 3763 4384
rect 3442 3296 3763 4320
rect 3442 3232 3450 3296
rect 3514 3232 3530 3296
rect 3594 3232 3610 3296
rect 3674 3232 3690 3296
rect 3754 3232 3763 3296
rect 3442 2208 3763 3232
rect 4110 2549 4170 4795
rect 5941 3840 6261 4864
rect 5941 3776 5949 3840
rect 6013 3776 6029 3840
rect 6093 3776 6109 3840
rect 6173 3776 6189 3840
rect 6253 3776 6261 3840
rect 5941 2752 6261 3776
rect 6686 3773 6746 6563
rect 8440 6560 8760 7584
rect 8440 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8760 6560
rect 8440 5472 8760 6496
rect 8894 5541 8954 8875
rect 10938 8192 11259 9216
rect 10938 8128 10946 8192
rect 11010 8128 11026 8192
rect 11090 8128 11106 8192
rect 11170 8128 11186 8192
rect 11250 8128 11259 8192
rect 10938 7104 11259 8128
rect 10938 7040 10946 7104
rect 11010 7040 11026 7104
rect 11090 7040 11106 7104
rect 11170 7040 11186 7104
rect 11250 7040 11259 7104
rect 10938 6016 11259 7040
rect 10938 5952 10946 6016
rect 11010 5952 11026 6016
rect 11090 5952 11106 6016
rect 11170 5952 11186 6016
rect 11250 5952 11259 6016
rect 8891 5540 8957 5541
rect 8891 5476 8892 5540
rect 8956 5476 8957 5540
rect 8891 5475 8957 5476
rect 8440 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8760 5472
rect 8440 4384 8760 5408
rect 8440 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8760 4384
rect 6683 3772 6749 3773
rect 6683 3708 6684 3772
rect 6748 3708 6749 3772
rect 6683 3707 6749 3708
rect 5941 2688 5949 2752
rect 6013 2688 6029 2752
rect 6093 2688 6109 2752
rect 6173 2688 6189 2752
rect 6253 2688 6261 2752
rect 4107 2548 4173 2549
rect 4107 2484 4108 2548
rect 4172 2484 4173 2548
rect 4107 2483 4173 2484
rect 3442 2144 3450 2208
rect 3514 2144 3530 2208
rect 3594 2144 3610 2208
rect 3674 2144 3690 2208
rect 3754 2144 3763 2208
rect 3442 2128 3763 2144
rect 5941 2128 6261 2688
rect 8440 3296 8760 4320
rect 8440 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8760 3296
rect 8440 2208 8760 3232
rect 8440 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8760 2208
rect 8440 2128 8760 2144
rect 10938 4928 11259 5952
rect 13437 12000 13757 13024
rect 13437 11936 13445 12000
rect 13509 11936 13525 12000
rect 13589 11936 13605 12000
rect 13669 11936 13685 12000
rect 13749 11936 13757 12000
rect 13437 10912 13757 11936
rect 13437 10848 13445 10912
rect 13509 10848 13525 10912
rect 13589 10848 13605 10912
rect 13669 10848 13685 10912
rect 13749 10848 13757 10912
rect 13437 9824 13757 10848
rect 13437 9760 13445 9824
rect 13509 9760 13525 9824
rect 13589 9760 13605 9824
rect 13669 9760 13685 9824
rect 13749 9760 13757 9824
rect 13437 8736 13757 9760
rect 13437 8672 13445 8736
rect 13509 8672 13525 8736
rect 13589 8672 13605 8736
rect 13669 8672 13685 8736
rect 13749 8672 13757 8736
rect 13437 7648 13757 8672
rect 13437 7584 13445 7648
rect 13509 7584 13525 7648
rect 13589 7584 13605 7648
rect 13669 7584 13685 7648
rect 13749 7584 13757 7648
rect 13437 6560 13757 7584
rect 13437 6496 13445 6560
rect 13509 6496 13525 6560
rect 13589 6496 13605 6560
rect 13669 6496 13685 6560
rect 13749 6496 13757 6560
rect 13437 5472 13757 6496
rect 13437 5408 13445 5472
rect 13509 5408 13525 5472
rect 13589 5408 13605 5472
rect 13669 5408 13685 5472
rect 13749 5408 13757 5472
rect 11467 5404 11533 5405
rect 11467 5340 11468 5404
rect 11532 5340 11533 5404
rect 11467 5339 11533 5340
rect 10938 4864 10946 4928
rect 11010 4864 11026 4928
rect 11090 4864 11106 4928
rect 11170 4864 11186 4928
rect 11250 4864 11259 4928
rect 10938 3840 11259 4864
rect 10938 3776 10946 3840
rect 11010 3776 11026 3840
rect 11090 3776 11106 3840
rect 11170 3776 11186 3840
rect 11250 3776 11259 3840
rect 10938 2752 11259 3776
rect 10938 2688 10946 2752
rect 11010 2688 11026 2752
rect 11090 2688 11106 2752
rect 11170 2688 11186 2752
rect 11250 2688 11259 2752
rect 10938 2128 11259 2688
rect 11470 2549 11530 5339
rect 13437 4384 13757 5408
rect 13437 4320 13445 4384
rect 13509 4320 13525 4384
rect 13589 4320 13605 4384
rect 13669 4320 13685 4384
rect 13749 4320 13757 4384
rect 12571 4316 12637 4317
rect 12571 4252 12572 4316
rect 12636 4252 12637 4316
rect 12571 4251 12637 4252
rect 12574 2685 12634 4251
rect 13437 3296 13757 4320
rect 13437 3232 13445 3296
rect 13509 3232 13525 3296
rect 13589 3232 13605 3296
rect 13669 3232 13685 3296
rect 13749 3232 13757 3296
rect 12571 2684 12637 2685
rect 12571 2620 12572 2684
rect 12636 2620 12637 2684
rect 12571 2619 12637 2620
rect 11467 2548 11533 2549
rect 11467 2484 11468 2548
rect 11532 2484 11533 2548
rect 11467 2483 11533 2484
rect 13437 2208 13757 3232
rect 13437 2144 13445 2208
rect 13509 2144 13525 2208
rect 13589 2144 13605 2208
rect 13669 2144 13685 2208
rect 13749 2144 13757 2208
rect 13437 2128 13757 2144
use sky130_fd_sc_hd__clkbuf_2  output58 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 2116 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output57
timestamp 1624635492
transform -1 0 1748 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output46
timestamp 1624635492
transform -1 0 1748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1624635492
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _34_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1748 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output61
timestamp 1624635492
transform -1 0 3220 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output60
timestamp 1624635492
transform -1 0 2852 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output59
timestamp 1624635492
transform -1 0 2484 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2024 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _36_
timestamp 1624635492
transform 1 0 3496 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp 1624635492
transform 1 0 3864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_2_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 4416 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_3_
timestamp 1624635492
transform 1 0 4508 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_1_
timestamp 1624635492
transform -1 0 4416 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output47
timestamp 1624635492
transform -1 0 4508 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output62
timestamp 1624635492
transform -1 0 3588 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 5520 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_1_
timestamp 1624635492
transform 1 0 5520 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_0_
timestamp 1624635492
transform 1 0 5520 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _31_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5244 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_58 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 6440 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1624635492
transform 1 0 6348 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output48
timestamp 1624635492
transform -1 0 6900 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1624635492
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1624635492
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 8004 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _44_
timestamp 1624635492
transform 1 0 8004 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 9752 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_4  input3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input14
timestamp 1624635492
transform -1 0 8556 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output49
timestamp 1624635492
transform -1 0 7268 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output50
timestamp 1624635492
transform -1 0 7636 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output51
timestamp 1624635492
transform -1 0 8004 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 11224 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1624635492
transform 1 0 10028 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1624635492
transform 1 0 9200 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1624635492
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_1_
timestamp 1624635492
transform -1 0 12880 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_2_
timestamp 1624635492
transform 1 0 12052 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1624635492
transform 1 0 10856 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1624635492
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1624635492
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1624635492
transform 1 0 11684 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1624635492
transform -1 0 12052 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115
timestamp 1624635492
transform 1 0 11684 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 12880 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_0_
timestamp 1624635492
transform 1 0 12880 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1624635492
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1624635492
transform -1 0 14076 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1624635492
transform -1 0 14444 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1624635492
transform -1 0 14720 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_S_FTB01 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 14996 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624635492
transform -1 0 16008 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624635492
transform -1 0 16008 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 14536 0 -1 2720
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  output107 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1624635492
transform -1 0 14904 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1624635492
transform -1 0 15732 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_150
timestamp 1624635492
transform 1 0 14904 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 2116 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624635492
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output88
timestamp 1624635492
transform -1 0 1748 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output104
timestamp 1624635492
transform -1 0 2116 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 5796 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1624635492
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output63
timestamp 1624635492
transform -1 0 4232 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_34
timestamp 1624635492
transform 1 0 4232 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp 1624635492
transform 1 0 5796 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l1_in_0_
timestamp 1624635492
transform 1 0 6440 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output52
timestamp 1624635492
transform 1 0 6072 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _46_
timestamp 1624635492
transform 1 0 7268 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 7544 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _47_
timestamp 1624635492
transform 1 0 9108 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1624635492
transform 1 0 9384 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1624635492
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input15
timestamp 1624635492
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_0_
timestamp 1624635492
transform -1 0 13340 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1624635492
transform 1 0 10856 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1624635492
transform -1 0 12052 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1624635492
transform -1 0 12420 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_105
timestamp 1624635492
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_123
timestamp 1624635492
transform 1 0 12420 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1624635492
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1624635492
transform -1 0 14812 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1624635492
transform -1 0 13708 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1624635492
transform -1 0 14076 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1624635492
transform -1 0 14260 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_144
timestamp 1624635492
transform 1 0 14352 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624635492
transform -1 0 16008 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1624635492
transform -1 0 15180 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1624635492
transform -1 0 15640 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_153
timestamp 1624635492
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_158
timestamp 1624635492
transform 1 0 15640 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1624635492
transform 1 0 1748 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _37_
timestamp 1624635492
transform 1 0 2024 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1624635492
transform -1 0 2668 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624635492
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output64
timestamp 1624635492
transform 1 0 2668 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output89
timestamp 1624635492
transform -1 0 1748 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_13
timestamp 1624635492
transform 1 0 2300 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 4508 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  output65
timestamp 1624635492
transform -1 0 4876 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 4876 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 6440 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_0_
timestamp 1624635492
transform 1 0 5060 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1624635492
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output55
timestamp 1624635492
transform 1 0 5980 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_52
timestamp 1624635492
transform 1 0 5888 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_0_
timestamp 1624635492
transform 1 0 7912 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output54
timestamp 1624635492
transform -1 0 9108 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1624635492
transform 1 0 10120 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1624635492
transform -1 0 10120 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1624635492
transform -1 0 9292 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1624635492
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _45_
timestamp 1624635492
transform 1 0 11684 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_1_
timestamp 1624635492
transform -1 0 12788 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1624635492
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1624635492
transform -1 0 11316 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_0_
timestamp 1624635492
transform -1 0 13616 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_1_
timestamp 1624635492
transform 1 0 13616 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1624635492
transform -1 0 14628 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624635492
transform -1 0 16008 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1624635492
transform -1 0 15732 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1624635492
transform -1 0 15364 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output45
timestamp 1624635492
transform 1 0 14628 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 1472 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 1748 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_0_
timestamp 1624635492
transform 1 0 2024 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_1_
timestamp 1624635492
transform 1 0 2852 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624635492
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1624635492
transform 1 0 1380 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1624635492
transform 1 0 4692 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l4_in_0_
timestamp 1624635492
transform 1 0 3864 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1624635492
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_28
timestamp 1624635492
transform 1 0 3680 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _43_
timestamp 1624635492
transform 1 0 4968 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1624635492
transform -1 0 6072 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1624635492
transform 1 0 6164 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1624635492
transform -1 0 6808 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1624635492
transform -1 0 5796 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1624635492
transform 1 0 5244 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output53
timestamp 1624635492
transform -1 0 7176 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_54
timestamp 1624635492
transform 1 0 6072 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_58
timestamp 1624635492
transform 1 0 6440 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_0_
timestamp 1624635492
transform 1 0 8188 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_1_
timestamp 1624635492
transform 1 0 7360 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 11776 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1624635492
transform 1 0 9476 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1624635492
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output56
timestamp 1624635492
transform -1 0 9476 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 11776 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_2_
timestamp 1624635492
transform 1 0 14352 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_3_
timestamp 1624635492
transform -1 0 14260 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1624635492
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1624635492
transform -1 0 13432 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624635492
transform -1 0 16008 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1624635492
transform -1 0 15732 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1624635492
transform -1 0 15364 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_0_
timestamp 1624635492
transform -1 0 2576 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l4_in_0_
timestamp 1624635492
transform 1 0 2576 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1624635492
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output90
timestamp 1624635492
transform -1 0 1748 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1624635492
transform 1 0 3404 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 3864 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 3680 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_1_
timestamp 1624635492
transform 1 0 6440 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l4_in_0_
timestamp 1624635492
transform 1 0 5520 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1624635492
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1624635492
transform -1 0 5520 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 9752 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_0_
timestamp 1624635492
transform 1 0 7268 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 8096 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1624635492
transform 1 0 9752 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1624635492
transform 1 0 10028 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 11960 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1624635492
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 11132 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1624635492
transform -1 0 11316 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1624635492
transform -1 0 11868 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1624635492
transform -1 0 11500 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_113
timestamp 1624635492
transform 1 0 11500 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_117
timestamp 1624635492
transform 1 0 11868 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 13432 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1624635492
transform 1 0 14904 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 15456 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1624635492
transform -1 0 16008 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1624635492
transform -1 0 15640 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_158
timestamp 1624635492
transform 1 0 15640 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_10
timestamp 1624635492
transform 1 0 2024 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1624635492
transform 1 0 1380 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1624635492
transform -1 0 1564 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1624635492
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1624635492
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 1748 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 1472 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_0_
timestamp 1624635492
transform -1 0 2944 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_1_
timestamp 1624635492
transform 1 0 2944 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 3036 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1624635492
transform 1 0 3404 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1624635492
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 3588 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1624635492
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_1_
timestamp 1624635492
transform 1 0 3772 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_2_
timestamp 1624635492
transform 1 0 3864 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_7_38
timestamp 1624635492
transform 1 0 4600 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 4692 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_2_
timestamp 1624635492
transform 1 0 4692 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1624635492
transform -1 0 5244 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 6716 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_3_
timestamp 1624635492
transform 1 0 5520 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1624635492
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 6440 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 6716 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1624635492
transform -1 0 6900 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_60
timestamp 1624635492
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1624635492
transform 1 0 8556 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 8372 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_2_
timestamp 1624635492
transform 1 0 6900 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_3_
timestamp 1624635492
transform 1 0 7728 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 8372 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1624635492
transform 1 0 8556 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 8740 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1624635492
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 9108 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1624635492
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_85
timestamp 1624635492
transform 1 0 8924 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 9660 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 9292 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1624635492
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 9568 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_93
timestamp 1624635492
transform 1 0 9660 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1624635492
transform -1 0 10764 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_1_
timestamp 1624635492
transform 1 0 10580 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l1_in_0_
timestamp 1624635492
transform -1 0 10580 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9752 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 11316 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 11500 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1624635492
transform -1 0 11316 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 10948 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 10764 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1624635492
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_115
timestamp 1624635492
transform 1 0 11684 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_121
timestamp 1624635492
transform 1 0 12236 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 12052 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 11684 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 12328 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1624635492
transform -1 0 12052 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_3_
timestamp 1624635492
transform -1 0 12604 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1624635492
transform 1 0 12604 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 12512 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_126
timestamp 1624635492
transform 1 0 12696 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__A0
timestamp 1624635492
transform -1 0 13524 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A1
timestamp 1624635492
transform -1 0 13340 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 12972 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 12788 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l4_in_0_
timestamp 1624635492
transform -1 0 13800 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_7_135 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 13524 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_142
timestamp 1624635492
transform 1 0 14168 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 14260 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1624635492
transform -1 0 14168 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1624635492
transform -1 0 13984 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1624635492
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_145
timestamp 1624635492
transform 1 0 14444 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_146
timestamp 1624635492
transform 1 0 14536 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_S_FTB01_A
timestamp 1624635492
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1624635492
transform -1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1624635492
transform -1 0 15548 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1624635492
transform -1 0 15180 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1624635492
transform -1 0 15364 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output108
timestamp 1624635492
transform 1 0 15364 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_157 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 15548 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1624635492
transform -1 0 16008 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1624635492
transform -1 0 16008 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 1840 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1624635492
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output91
timestamp 1624635492
transform -1 0 1748 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7
timestamp 1624635492
transform 1 0 1748 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_26
timestamp 1624635492
transform 1 0 3496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1624635492
transform 1 0 3312 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1624635492
transform -1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1624635492
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_32
timestamp 1624635492
transform 1 0 4048 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 3864 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1624635492
transform 1 0 4140 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 4324 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 4508 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 4692 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_41
timestamp 1624635492
transform 1 0 4876 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_1_
timestamp 1624635492
transform 1 0 5520 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 6348 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 6624 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1624635492
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 5336 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1624635492
transform -1 0 5336 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 4968 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1624635492
transform -1 0 7544 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 7544 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_66
timestamp 1624635492
transform 1 0 7176 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9108 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_0_
timestamp 1624635492
transform 1 0 10580 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1624635492
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 11592 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 11408 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_1_
timestamp 1624635492
transform 1 0 13064 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1624635492
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_139 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 13892 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_144 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 14352 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1624635492
transform -1 0 16008 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_156
timestamp 1624635492
transform 1 0 15456 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 2944 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 1748 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1624635492
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output92
timestamp 1624635492
transform -1 0 1748 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1624635492
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A1
timestamp 1624635492
transform -1 0 2944 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output104_A
timestamp 1624635492
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_10
timestamp 1624635492
transform 1 0 2024 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_15
timestamp 1624635492
transform 1 0 2484 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_2_
timestamp 1624635492
transform 1 0 4416 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_0_
timestamp 1624635492
transform 1 0 5520 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1624635492
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 6440 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 5244 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1624635492
transform 1 0 6624 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1624635492
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_47
timestamp 1624635492
transform 1 0 5428 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 6992 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l4_in_0_
timestamp 1624635492
transform 1 0 8464 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9660 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1624635492
transform 1 0 12604 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_2_
timestamp 1624635492
transform -1 0 12604 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1624635492
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 11316 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 1624635492
transform 1 0 11500 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_115
timestamp 1624635492
transform 1 0 11684 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 12880 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_130
timestamp 1624635492
transform 1 0 13064 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_142
timestamp 1624635492
transform 1 0 14168 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1624635492
transform -1 0 16008 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_154
timestamp 1624635492
transform 1 0 15272 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_158
timestamp 1624635492
transform 1 0 15640 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 1748 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1624635492
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output93
timestamp 1624635492
transform -1 0 1748 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_10
timestamp 1624635492
transform 1 0 2024 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_1_
timestamp 1624635492
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1624635492
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 5152 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1624635492
transform 1 0 3864 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A1
timestamp 1624635492
transform -1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1624635492
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_22
timestamp 1624635492
transform 1 0 3128 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 6808 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_0_
timestamp 1624635492
transform -1 0 7820 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_1_
timestamp 1624635492
transform -1 0 9016 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 7820 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_76
timestamp 1624635492
transform 1 0 8096 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_3_
timestamp 1624635492
transform 1 0 9108 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_0_
timestamp 1624635492
transform -1 0 10948 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1624635492
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 9936 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l4_in_0_
timestamp 1624635492
transform 1 0 10948 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_2_
timestamp 1624635492
transform -1 0 12604 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_0_
timestamp 1624635492
transform -1 0 13432 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1624635492
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 13432 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 13616 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_138
timestamp 1624635492
transform 1 0 13800 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_142
timestamp 1624635492
transform 1 0 14168 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_144
timestamp 1624635492
transform 1 0 14352 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1624635492
transform -1 0 16008 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_156
timestamp 1624635492
transform 1 0 15456 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 2484 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 1564 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1624635492
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1624635492
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1840 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_14
timestamp 1624635492
transform 1 0 2392 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_0_
timestamp 1624635492
transform 1 0 3956 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 4876 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_40
timestamp 1624635492
transform 1 0 4784 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1624635492
transform 1 0 5888 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 6440 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_0_
timestamp 1624635492
transform 1 0 5060 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1624635492
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_1_
timestamp 1624635492
transform 1 0 8464 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 7912 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1624635492
transform -1 0 9568 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 9936 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 9936 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_92
timestamp 1624635492
transform 1 0 9568 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_1_
timestamp 1624635492
transform -1 0 12880 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1624635492
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 11868 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_112
timestamp 1624635492
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 12880 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_11_144
timestamp 1624635492
transform 1 0 14352 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1624635492
transform -1 0 16008 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_156
timestamp 1624635492
transform 1 0 15456 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l4_in_0_
timestamp 1624635492
transform 1 0 2944 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1624635492
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output94
timestamp 1624635492
transform -1 0 1748 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_7
timestamp 1624635492
transform 1 0 1748 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_19
timestamp 1624635492
transform 1 0 2852 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 3864 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1624635492
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 5336 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_0_
timestamp 1624635492
transform -1 0 7636 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_0_
timestamp 1624635492
transform -1 0 8648 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 7636 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 8648 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_2_
timestamp 1624635492
transform 1 0 9108 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_0_
timestamp 1624635492
transform 1 0 9936 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1624635492
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 10764 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_0_
timestamp 1624635492
transform -1 0 13340 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 12328 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_121
timestamp 1624635492
transform 1 0 12236 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1624635492
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 13340 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_135
timestamp 1624635492
transform 1 0 13524 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_144
timestamp 1624635492
transform 1 0 14352 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1624635492
transform -1 0 16008 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_156
timestamp 1624635492
transform 1 0 15456 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 1748 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1624635492
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1624635492
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output95
timestamp 1624635492
transform -1 0 1748 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1624635492
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1624635492
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_10
timestamp 1624635492
transform 1 0 2024 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_2_
timestamp 1624635492
transform 1 0 4508 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_1_
timestamp 1624635492
transform 1 0 3680 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_0_
timestamp 1624635492
transform 1 0 3864 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1624635492
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 4692 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_27
timestamp 1624635492
transform 1 0 3588 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_22
timestamp 1624635492
transform 1 0 3128 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_28
timestamp 1624635492
transform 1 0 3680 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1624635492
transform -1 0 5520 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 5796 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 7912 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_3_
timestamp 1624635492
transform 1 0 5336 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1624635492
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_43
timestamp 1624635492
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_48
timestamp 1624635492
transform 1 0 5520 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1624635492
transform 1 0 8740 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_2_
timestamp 1624635492
transform 1 0 7912 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 9844 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_13_74
timestamp 1624635492
transform 1 0 7912 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_67
timestamp 1624635492
transform 1 0 7268 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_73
timestamp 1624635492
transform 1 0 7820 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 11500 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_1_
timestamp 1624635492
transform 1 0 9936 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_0_
timestamp 1624635492
transform -1 0 10028 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1624635492
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_95
timestamp 1624635492
transform 1 0 9844 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_87
timestamp 1624635492
transform 1 0 9108 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 12972 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_1_
timestamp 1624635492
transform -1 0 12972 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1624635492
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 10764 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 10948 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_111
timestamp 1624635492
transform 1 0 11316 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_115
timestamp 1624635492
transform 1 0 11684 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_119
timestamp 1624635492
transform 1 0 12052 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_2_
timestamp 1624635492
transform -1 0 14168 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_3_
timestamp 1624635492
transform 1 0 14352 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_0_
timestamp 1624635492
transform 1 0 12972 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_1_
timestamp 1624635492
transform 1 0 13800 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1624635492
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 12972 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_131
timestamp 1624635492
transform 1 0 13156 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_142
timestamp 1624635492
transform 1 0 14168 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1624635492
transform -1 0 16008 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1624635492
transform -1 0 16008 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output86
timestamp 1624635492
transform 1 0 15364 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A1
timestamp 1624635492
transform -1 0 15364 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_147
timestamp 1624635492
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 1472 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_0_
timestamp 1624635492
transform 1 0 2852 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_0_
timestamp 1624635492
transform 1 0 2024 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1624635492
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1624635492
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_7
timestamp 1624635492
transform 1 0 1748 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 5428 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_30
timestamp 1624635492
transform 1 0 3864 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_2_
timestamp 1624635492
transform 1 0 5428 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1624635492
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 6440 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_56
timestamp 1624635492
transform 1 0 6256 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_60
timestamp 1624635492
transform 1 0 6624 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 9200 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_1_
timestamp 1624635492
transform -1 0 7728 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9844 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_2_
timestamp 1624635492
transform 1 0 10672 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_92
timestamp 1624635492
transform 1 0 9568 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l4_in_0_
timestamp 1624635492
transform 1 0 11684 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1624635492
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 12512 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1624635492
transform 1 0 11500 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1624635492
transform -1 0 14536 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 12788 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_126
timestamp 1624635492
transform 1 0 12696 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1624635492
transform -1 0 16008 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 14536 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_148
timestamp 1624635492
transform 1 0 14720 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_156
timestamp 1624635492
transform 1 0 15456 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_1_
timestamp 1624635492
transform 1 0 2852 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l4_in_0_
timestamp 1624635492
transform 1 0 1840 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1624635492
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output96
timestamp 1624635492
transform -1 0 1748 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1624635492
transform 1 0 1748 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_17
timestamp 1624635492
transform 1 0 2668 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 5336 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1624635492
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_28
timestamp 1624635492
transform 1 0 3680 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_1_
timestamp 1624635492
transform 1 0 6716 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_3_
timestamp 1624635492
transform 1 0 5336 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 6164 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_57
timestamp 1624635492
transform 1 0 6348 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_3_
timestamp 1624635492
transform 1 0 7912 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 8740 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_72
timestamp 1624635492
transform 1 0 7728 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_1_
timestamp 1624635492
transform -1 0 10212 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1624635492
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 10212 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1624635492
transform 1 0 8924 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_87
timestamp 1624635492
transform 1 0 9108 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_101
timestamp 1624635492
transform 1 0 10396 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 13064 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_16_113
timestamp 1624635492
transform 1 0 11500 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1624635492
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_130
timestamp 1624635492
transform 1 0 13064 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_142
timestamp 1624635492
transform 1 0 14168 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_144
timestamp 1624635492
transform 1 0 14352 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1624635492
transform -1 0 16008 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_156
timestamp 1624635492
transform 1 0 15456 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 2852 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1624635492
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_19
timestamp 1624635492
transform 1 0 2852 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l4_in_0_
timestamp 1624635492
transform 1 0 4692 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_1_
timestamp 1624635492
transform 1 0 3864 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 3680 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_25
timestamp 1624635492
transform 1 0 3404 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 6440 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1624635492
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 5520 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_51
timestamp 1624635492
transform 1 0 5796 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1624635492
transform 1 0 8740 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l4_in_0_
timestamp 1624635492
transform 1 0 7912 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9936 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 9752 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 9568 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_86
timestamp 1624635492
transform 1 0 9016 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_1_
timestamp 1624635492
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1624635492
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 11960 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A1
timestamp 1624635492
transform -1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 12328 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_124
timestamp 1624635492
transform 1 0 12512 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_136
timestamp 1624635492
transform 1 0 13616 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1624635492
transform -1 0 16008 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_148
timestamp 1624635492
transform 1 0 14720 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_156
timestamp 1624635492
transform 1 0 15456 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 2024 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 1748 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1624635492
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output97
timestamp 1624635492
transform -1 0 1748 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_0_
timestamp 1624635492
transform -1 0 5336 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1624635492
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 3496 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 3864 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_28
timestamp 1624635492
transform 1 0 3680 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_32
timestamp 1624635492
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_36
timestamp 1624635492
transform 1 0 4416 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_1_
timestamp 1624635492
transform 1 0 5336 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_3_
timestamp 1624635492
transform -1 0 7268 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 6164 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_57
timestamp 1624635492
transform 1 0 6348 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 7268 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 9016 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9108 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1624635492
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 10580 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 11224 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 10856 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_105
timestamp 1624635492
transform 1 0 10764 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 14076 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1624635492
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1624635492
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_126
timestamp 1624635492
transform 1 0 12696 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1624635492
transform 1 0 14076 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_144
timestamp 1624635492
transform 1 0 14352 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1624635492
transform -1 0 16008 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_156
timestamp 1624635492
transform 1 0 15456 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_7
timestamp 1624635492
transform 1 0 1748 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 1624635492
transform 1 0 1380 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output98
timestamp 1624635492
transform -1 0 1748 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1624635492
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1624635492
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 1748 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 1472 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_15
timestamp 1624635492
transform 1 0 2484 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_14
timestamp 1624635492
transform 1 0 2392 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_10
timestamp 1624635492
transform 1 0 2024 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_0_
timestamp 1624635492
transform 1 0 2668 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l1_in_0_
timestamp 1624635492
transform -1 0 3312 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 3312 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1624635492
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 3496 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 3956 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_40
timestamp 1624635492
transform 1 0 4784 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_28
timestamp 1624635492
transform 1 0 3680 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_30
timestamp 1624635492
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_33
timestamp 1624635492
transform 1 0 4140 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_41
timestamp 1624635492
transform 1 0 4876 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 6256 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_0_
timestamp 1624635492
transform 1 0 5428 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_1_
timestamp 1624635492
transform 1 0 6440 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_2_
timestamp 1624635492
transform 1 0 5520 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1624635492
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 5336 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 5060 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_45
timestamp 1624635492
transform 1 0 5244 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_2_
timestamp 1624635492
transform 1 0 7268 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 8096 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 7728 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 8648 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 7912 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_83
timestamp 1624635492
transform 1 0 8740 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_76
timestamp 1624635492
transform 1 0 8096 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1624635492
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_87
timestamp 1624635492
transform 1 0 9108 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 9752 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1624635492
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_0_
timestamp 1624635492
transform 1 0 9568 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_19_103
timestamp 1624635492
transform 1 0 10580 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9752 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_2_
timestamp 1624635492
transform -1 0 11500 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 11868 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_1_
timestamp 1624635492
transform 1 0 11684 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_2_
timestamp 1624635492
transform 1 0 12512 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_3_
timestamp 1624635492
transform 1 0 12144 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1624635492
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 11868 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 1624635492
transform 1 0 11500 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_119
timestamp 1624635492
transform 1 0 12052 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 13340 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1624635492
transform -1 0 13156 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 13524 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 13340 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1624635492
transform 1 0 13340 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 14076 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A1
timestamp 1624635492
transform -1 0 13892 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__A0
timestamp 1624635492
transform -1 0 14536 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 14168 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__A1
timestamp 1624635492
transform -1 0 14260 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 14352 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1624635492
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_146
timestamp 1624635492
transform 1 0 14536 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 14536 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 14720 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_N_FTB01_A
timestamp 1624635492
transform -1 0 14996 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_N_FTB01
timestamp 1624635492
transform 1 0 14996 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 14904 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_153
timestamp 1624635492
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1624635492
transform -1 0 15732 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1624635492
transform -1 0 15456 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1624635492
transform 1 0 15456 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1624635492
transform -1 0 16008 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1624635492
transform -1 0 16008 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_1_
timestamp 1624635492
transform 1 0 2944 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_0_
timestamp 1624635492
transform 1 0 2116 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 1748 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1624635492
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output99
timestamp 1624635492
transform -1 0 1748 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_10
timestamp 1624635492
transform 1 0 2024 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1624635492
transform -1 0 5152 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_2_
timestamp 1624635492
transform 1 0 4048 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_31
timestamp 1624635492
transform 1 0 3956 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_0_
timestamp 1624635492
transform 1 0 5336 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1624635492
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 6440 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 5152 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 6624 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_55
timestamp 1624635492
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_62
timestamp 1624635492
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 8464 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 8464 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 11408 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_1_
timestamp 1624635492
transform 1 0 11684 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_0_
timestamp 1624635492
transform -1 0 13432 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1624635492
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1624635492
transform -1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_124
timestamp 1624635492
transform 1 0 12512 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_1_
timestamp 1624635492
transform 1 0 13432 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1624635492
transform -1 0 14444 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_145
timestamp 1624635492
transform 1 0 14444 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 15732 0 1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1624635492
transform -1 0 16008 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1624635492
transform 1 0 1564 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 3404 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1624635492
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1624635492
transform -1 0 1564 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_8
timestamp 1624635492
transform 1 0 1840 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 3864 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1624635492
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_25
timestamp 1624635492
transform 1 0 3404 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_3_
timestamp 1624635492
transform 1 0 5336 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_0_
timestamp 1624635492
transform 1 0 6808 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 6440 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 6624 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 6440 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_0_
timestamp 1624635492
transform 1 0 7636 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l4_in_0_
timestamp 1624635492
transform 1 0 9200 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1624635492
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 10948 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1624635492
transform -1 0 10580 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 10212 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1624635492
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 10028 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_87
timestamp 1624635492
transform 1 0 9108 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_103
timestamp 1624635492
transform 1 0 10580 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 10948 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1624635492
transform -1 0 12788 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 12788 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1624635492
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1624635492
transform -1 0 14536 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1624635492
transform 1 0 14536 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1624635492
transform -1 0 16008 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1624635492
transform -1 0 15732 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output87
timestamp 1624635492
transform 1 0 14996 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1624635492
transform -1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1624635492
transform -1 0 2024 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l4_in_0_
timestamp 1624635492
transform 1 0 2116 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1624635492
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output100
timestamp 1624635492
transform -1 0 1748 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1624635492
transform -1 0 3128 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_10
timestamp 1624635492
transform 1 0 2024 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4416 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_1_
timestamp 1624635492
transform 1 0 3312 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1624635492
transform 1 0 3128 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_33
timestamp 1624635492
transform 1 0 4140 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_1_
timestamp 1624635492
transform 1 0 6716 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1624635492
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1624635492
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_52
timestamp 1624635492
transform 1 0 5888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_58
timestamp 1624635492
transform 1 0 6440 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_2_
timestamp 1624635492
transform 1 0 7728 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_3_
timestamp 1624635492
transform 1 0 8556 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 7544 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 9936 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1624635492
transform -1 0 9936 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1624635492
transform 1 0 9384 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 9568 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_2_
timestamp 1624635492
transform -1 0 12972 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1624635492
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1624635492
transform -1 0 12052 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1624635492
transform -1 0 11592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_119
timestamp 1624635492
transform 1 0 12052 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_0_
timestamp 1624635492
transform 1 0 12972 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_3_
timestamp 1624635492
transform -1 0 14904 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1624635492
transform -1 0 14076 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_138
timestamp 1624635492
transform 1 0 13800 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_1_
timestamp 1624635492
transform 1 0 14904 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1624635492
transform -1 0 16008 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 1748 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2024 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2300 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1624635492
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1624635492
transform 1 0 2576 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1624635492
transform 1 0 2852 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output101
timestamp 1624635492
transform -1 0 1748 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 6256 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1624635492
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1624635492
transform -1 0 3312 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1624635492
transform -1 0 3496 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1624635492
transform 1 0 3496 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1624635492
transform 1 0 4600 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_28
timestamp 1624635492
transform 1 0 3680 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_30
timestamp 1624635492
transform 1 0 3864 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_0_
timestamp 1624635492
transform -1 0 7268 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1624635492
transform 1 0 6256 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1624635492
transform -1 0 8556 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_1_
timestamp 1624635492
transform 1 0 7268 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1624635492
transform 1 0 8096 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1624635492
transform 1 0 8556 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1624635492
transform 1 0 8740 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_0_
timestamp 1624635492
transform -1 0 10028 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_1_
timestamp 1624635492
transform 1 0 10304 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1624635492
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1624635492
transform -1 0 10304 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_85
timestamp 1624635492
transform 1 0 8924 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_87
timestamp 1624635492
transform 1 0 9108 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_97
timestamp 1624635492
transform 1 0 10028 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l4_in_0_
timestamp 1624635492
transform 1 0 11132 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_1_
timestamp 1624635492
transform -1 0 12972 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1624635492
transform -1 0 12144 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_2_
timestamp 1624635492
transform -1 0 15180 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_0_
timestamp 1624635492
transform 1 0 12972 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1624635492
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1624635492
transform -1 0 14168 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_142
timestamp 1624635492
transform 1 0 14168 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1624635492
transform -1 0 16008 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1624635492
transform -1 0 15640 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_153
timestamp 1624635492
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_158
timestamp 1624635492
transform 1 0 15640 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1624635492
transform -1 0 2484 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1624635492
transform -1 0 2760 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1624635492
transform 1 0 2852 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp 1624635492
transform 1 0 1748 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1624635492
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output105
timestamp 1624635492
transform -1 0 1748 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1624635492
transform -1 0 2208 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_18
timestamp 1624635492
transform 1 0 2760 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1624635492
transform 1 0 3128 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1624635492
transform -1 0 3680 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 1624635492
transform -1 0 3956 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 1624635492
transform 1 0 4692 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1624635492
transform -1 0 4140 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1624635492
transform -1 0 4324 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1624635492
transform -1 0 4508 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1624635492
transform -1 0 4692 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1624635492
transform -1 0 5704 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1624635492
transform 1 0 5980 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1624635492
transform -1 0 5980 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l4_in_0_
timestamp 1624635492
transform 1 0 6440 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1624635492
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1624635492
transform -1 0 5152 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1624635492
transform -1 0 5428 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_44
timestamp 1624635492
transform 1 0 5152 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_56
timestamp 1624635492
transform 1 0 6256 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1624635492
transform 1 0 7268 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1624635492
transform 1 0 7544 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1624635492
transform 1 0 7820 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp 1624635492
transform -1 0 8556 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l1_in_0_
timestamp 1624635492
transform -1 0 9476 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1624635492
transform -1 0 8280 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_81
timestamp 1624635492
transform 1 0 8556 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1624635492
transform -1 0 9936 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_0_
timestamp 1624635492
transform -1 0 10764 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1624635492
transform -1 0 9660 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 12144 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_1_
timestamp 1624635492
transform -1 0 11592 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1624635492
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1624635492
transform -1 0 12052 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_119
timestamp 1624635492
transform 1 0 12052 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 13800 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1624635492
transform -1 0 13800 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1624635492
transform -1 0 16008 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1624635492
transform -1 0 15640 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_158
timestamp 1624635492
transform 1 0 15640 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output102
timestamp 1624635492
transform -1 0 1748 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output66
timestamp 1624635492
transform -1 0 1748 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1624635492
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1624635492
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output103
timestamp 1624635492
transform -1 0 2116 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output77
timestamp 1624635492
transform -1 0 2116 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1624635492
transform 1 0 2392 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output78
timestamp 1624635492
transform -1 0 2484 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1624635492
transform 1 0 2116 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output81
timestamp 1624635492
transform -1 0 2944 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output80
timestamp 1624635492
transform -1 0 3220 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output79
timestamp 1624635492
transform -1 0 2852 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_20
timestamp 1624635492
transform 1 0 2944 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_23
timestamp 1624635492
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output83
timestamp 1624635492
transform -1 0 3772 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output82
timestamp 1624635492
transform -1 0 3404 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output75
timestamp 1624635492
transform 1 0 3404 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output84
timestamp 1624635492
transform -1 0 4232 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output74
timestamp 1624635492
transform 1 0 3864 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1624635492
transform 1 0 3772 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1624635492
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output85
timestamp 1624635492
transform -1 0 4600 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output73
timestamp 1624635492
transform 1 0 4232 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output67
timestamp 1624635492
transform -1 0 4968 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1624635492
transform 1 0 4600 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1624635492
transform -1 0 5060 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_51
timestamp 1624635492
transform 1 0 5796 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_42
timestamp 1624635492
transform 1 0 4968 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output70
timestamp 1624635492
transform -1 0 6256 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output69
timestamp 1624635492
transform -1 0 5796 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output68
timestamp 1624635492
transform -1 0 5428 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1624635492
transform 1 0 5060 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1624635492
transform -1 0 6440 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output71
timestamp 1624635492
transform -1 0 6900 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1624635492
transform 1 0 6440 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 6808 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 5336 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1624635492
transform 1 0 8740 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input23
timestamp 1624635492
transform -1 0 9108 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 1624635492
transform -1 0 8556 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1624635492
transform -1 0 8188 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1624635492
transform -1 0 7820 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output72
timestamp 1624635492
transform -1 0 7268 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output76
timestamp 1624635492
transform -1 0 8740 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1624635492
transform -1 0 7452 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_78
timestamp 1624635492
transform 1 0 8280 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9108 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 9384 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1624635492
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1624635492
transform 1 0 9108 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input36
timestamp 1624635492
transform 1 0 10580 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1624635492
transform -1 0 9384 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_2_
timestamp 1624635492
transform 1 0 11040 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_3_
timestamp 1624635492
transform 1 0 11868 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l4_in_0_
timestamp 1624635492
transform 1 0 12328 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1624635492
transform 1 0 11776 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1624635492
transform -1 0 12328 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1624635492
transform -1 0 11776 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input35
timestamp 1624635492
transform 1 0 10856 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_107
timestamp 1624635492
transform 1 0 10948 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_117
timestamp 1624635492
transform 1 0 11868 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 14168 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1624635492
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1624635492
transform 1 0 14444 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1624635492
transform -1 0 13524 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1624635492
transform -1 0 13892 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1624635492
transform -1 0 14260 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1624635492
transform -1 0 14720 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1624635492
transform -1 0 14444 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_142
timestamp 1624635492
transform 1 0 14168 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_2  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 14904 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 14720 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1624635492
transform -1 0 16008 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1624635492
transform -1 0 16008 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1624635492
transform -1 0 14904 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output106
timestamp 1624635492
transform 1 0 15456 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1624635492
transform -1 0 15732 0 1 16864
box -38 -48 222 592
<< labels >>
rlabel metal2 s 202 19200 258 20000 6 IO_ISOL_N
port 0 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 ccff_head
port 1 nsew signal input
rlabel metal3 s 16400 1912 17200 2032 6 ccff_tail
port 2 nsew signal tristate
rlabel metal2 s 8574 0 8630 800 6 chany_bottom_in[0]
port 3 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 chany_bottom_in[10]
port 4 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 chany_bottom_in[11]
port 5 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 chany_bottom_in[12]
port 6 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 chany_bottom_in[13]
port 7 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 chany_bottom_in[14]
port 8 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 chany_bottom_in[15]
port 9 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 chany_bottom_in[16]
port 10 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 chany_bottom_in[17]
port 11 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 chany_bottom_in[18]
port 12 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 chany_bottom_in[19]
port 13 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 chany_bottom_in[1]
port 14 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 chany_bottom_in[2]
port 15 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 chany_bottom_in[3]
port 16 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 chany_bottom_in[4]
port 17 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 chany_bottom_in[5]
port 18 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 chany_bottom_in[6]
port 19 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 chany_bottom_in[7]
port 20 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 chany_bottom_in[8]
port 21 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 chany_bottom_in[9]
port 22 nsew signal input
rlabel metal2 s 202 0 258 800 6 chany_bottom_out[0]
port 23 nsew signal tristate
rlabel metal2 s 4342 0 4398 800 6 chany_bottom_out[10]
port 24 nsew signal tristate
rlabel metal2 s 4802 0 4858 800 6 chany_bottom_out[11]
port 25 nsew signal tristate
rlabel metal2 s 5170 0 5226 800 6 chany_bottom_out[12]
port 26 nsew signal tristate
rlabel metal2 s 5630 0 5686 800 6 chany_bottom_out[13]
port 27 nsew signal tristate
rlabel metal2 s 5998 0 6054 800 6 chany_bottom_out[14]
port 28 nsew signal tristate
rlabel metal2 s 6458 0 6514 800 6 chany_bottom_out[15]
port 29 nsew signal tristate
rlabel metal2 s 6826 0 6882 800 6 chany_bottom_out[16]
port 30 nsew signal tristate
rlabel metal2 s 7286 0 7342 800 6 chany_bottom_out[17]
port 31 nsew signal tristate
rlabel metal2 s 7746 0 7802 800 6 chany_bottom_out[18]
port 32 nsew signal tristate
rlabel metal2 s 8114 0 8170 800 6 chany_bottom_out[19]
port 33 nsew signal tristate
rlabel metal2 s 570 0 626 800 6 chany_bottom_out[1]
port 34 nsew signal tristate
rlabel metal2 s 1030 0 1086 800 6 chany_bottom_out[2]
port 35 nsew signal tristate
rlabel metal2 s 1398 0 1454 800 6 chany_bottom_out[3]
port 36 nsew signal tristate
rlabel metal2 s 1858 0 1914 800 6 chany_bottom_out[4]
port 37 nsew signal tristate
rlabel metal2 s 2226 0 2282 800 6 chany_bottom_out[5]
port 38 nsew signal tristate
rlabel metal2 s 2686 0 2742 800 6 chany_bottom_out[6]
port 39 nsew signal tristate
rlabel metal2 s 3054 0 3110 800 6 chany_bottom_out[7]
port 40 nsew signal tristate
rlabel metal2 s 3514 0 3570 800 6 chany_bottom_out[8]
port 41 nsew signal tristate
rlabel metal2 s 3974 0 4030 800 6 chany_bottom_out[9]
port 42 nsew signal tristate
rlabel metal2 s 8758 19200 8814 20000 6 chany_top_in[0]
port 43 nsew signal input
rlabel metal2 s 12898 19200 12954 20000 6 chany_top_in[10]
port 44 nsew signal input
rlabel metal2 s 13266 19200 13322 20000 6 chany_top_in[11]
port 45 nsew signal input
rlabel metal2 s 13634 19200 13690 20000 6 chany_top_in[12]
port 46 nsew signal input
rlabel metal2 s 14094 19200 14150 20000 6 chany_top_in[13]
port 47 nsew signal input
rlabel metal2 s 14462 19200 14518 20000 6 chany_top_in[14]
port 48 nsew signal input
rlabel metal2 s 14922 19200 14978 20000 6 chany_top_in[15]
port 49 nsew signal input
rlabel metal2 s 15290 19200 15346 20000 6 chany_top_in[16]
port 50 nsew signal input
rlabel metal2 s 15750 19200 15806 20000 6 chany_top_in[17]
port 51 nsew signal input
rlabel metal2 s 16118 19200 16174 20000 6 chany_top_in[18]
port 52 nsew signal input
rlabel metal2 s 16578 19200 16634 20000 6 chany_top_in[19]
port 53 nsew signal input
rlabel metal2 s 9126 19200 9182 20000 6 chany_top_in[1]
port 54 nsew signal input
rlabel metal2 s 9586 19200 9642 20000 6 chany_top_in[2]
port 55 nsew signal input
rlabel metal2 s 9954 19200 10010 20000 6 chany_top_in[3]
port 56 nsew signal input
rlabel metal2 s 10414 19200 10470 20000 6 chany_top_in[4]
port 57 nsew signal input
rlabel metal2 s 10782 19200 10838 20000 6 chany_top_in[5]
port 58 nsew signal input
rlabel metal2 s 11242 19200 11298 20000 6 chany_top_in[6]
port 59 nsew signal input
rlabel metal2 s 11610 19200 11666 20000 6 chany_top_in[7]
port 60 nsew signal input
rlabel metal2 s 12070 19200 12126 20000 6 chany_top_in[8]
port 61 nsew signal input
rlabel metal2 s 12438 19200 12494 20000 6 chany_top_in[9]
port 62 nsew signal input
rlabel metal2 s 570 19200 626 20000 6 chany_top_out[0]
port 63 nsew signal tristate
rlabel metal2 s 4618 19200 4674 20000 6 chany_top_out[10]
port 64 nsew signal tristate
rlabel metal2 s 5078 19200 5134 20000 6 chany_top_out[11]
port 65 nsew signal tristate
rlabel metal2 s 5446 19200 5502 20000 6 chany_top_out[12]
port 66 nsew signal tristate
rlabel metal2 s 5906 19200 5962 20000 6 chany_top_out[13]
port 67 nsew signal tristate
rlabel metal2 s 6274 19200 6330 20000 6 chany_top_out[14]
port 68 nsew signal tristate
rlabel metal2 s 6734 19200 6790 20000 6 chany_top_out[15]
port 69 nsew signal tristate
rlabel metal2 s 7102 19200 7158 20000 6 chany_top_out[16]
port 70 nsew signal tristate
rlabel metal2 s 7562 19200 7618 20000 6 chany_top_out[17]
port 71 nsew signal tristate
rlabel metal2 s 7930 19200 7986 20000 6 chany_top_out[18]
port 72 nsew signal tristate
rlabel metal2 s 8390 19200 8446 20000 6 chany_top_out[19]
port 73 nsew signal tristate
rlabel metal2 s 938 19200 994 20000 6 chany_top_out[1]
port 74 nsew signal tristate
rlabel metal2 s 1398 19200 1454 20000 6 chany_top_out[2]
port 75 nsew signal tristate
rlabel metal2 s 1766 19200 1822 20000 6 chany_top_out[3]
port 76 nsew signal tristate
rlabel metal2 s 2226 19200 2282 20000 6 chany_top_out[4]
port 77 nsew signal tristate
rlabel metal2 s 2594 19200 2650 20000 6 chany_top_out[5]
port 78 nsew signal tristate
rlabel metal2 s 3054 19200 3110 20000 6 chany_top_out[6]
port 79 nsew signal tristate
rlabel metal2 s 3422 19200 3478 20000 6 chany_top_out[7]
port 80 nsew signal tristate
rlabel metal2 s 3882 19200 3938 20000 6 chany_top_out[8]
port 81 nsew signal tristate
rlabel metal2 s 4250 19200 4306 20000 6 chany_top_out[9]
port 82 nsew signal tristate
rlabel metal3 s 16400 9800 17200 9920 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 83 nsew signal tristate
rlabel metal3 s 16400 13880 17200 14000 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 84 nsew signal input
rlabel metal3 s 16400 17824 17200 17944 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 85 nsew signal tristate
rlabel metal3 s 0 3272 800 3392 6 left_grid_pin_16_
port 86 nsew signal tristate
rlabel metal3 s 0 4224 800 4344 6 left_grid_pin_17_
port 87 nsew signal tristate
rlabel metal3 s 0 5176 800 5296 6 left_grid_pin_18_
port 88 nsew signal tristate
rlabel metal3 s 0 6128 800 6248 6 left_grid_pin_19_
port 89 nsew signal tristate
rlabel metal3 s 0 7080 800 7200 6 left_grid_pin_20_
port 90 nsew signal tristate
rlabel metal3 s 0 8032 800 8152 6 left_grid_pin_21_
port 91 nsew signal tristate
rlabel metal3 s 0 8984 800 9104 6 left_grid_pin_22_
port 92 nsew signal tristate
rlabel metal3 s 0 9936 800 10056 6 left_grid_pin_23_
port 93 nsew signal tristate
rlabel metal3 s 0 10888 800 11008 6 left_grid_pin_24_
port 94 nsew signal tristate
rlabel metal3 s 0 11840 800 11960 6 left_grid_pin_25_
port 95 nsew signal tristate
rlabel metal3 s 0 12792 800 12912 6 left_grid_pin_26_
port 96 nsew signal tristate
rlabel metal3 s 0 13744 800 13864 6 left_grid_pin_27_
port 97 nsew signal tristate
rlabel metal3 s 0 14696 800 14816 6 left_grid_pin_28_
port 98 nsew signal tristate
rlabel metal3 s 0 15648 800 15768 6 left_grid_pin_29_
port 99 nsew signal tristate
rlabel metal3 s 0 16600 800 16720 6 left_grid_pin_30_
port 100 nsew signal tristate
rlabel metal3 s 0 17552 800 17672 6 left_grid_pin_31_
port 101 nsew signal tristate
rlabel metal3 s 0 18504 800 18624 6 left_width_0_height_0__pin_0_
port 102 nsew signal input
rlabel metal3 s 0 416 800 536 6 left_width_0_height_0__pin_1_lower
port 103 nsew signal tristate
rlabel metal3 s 0 19456 800 19576 6 left_width_0_height_0__pin_1_upper
port 104 nsew signal tristate
rlabel metal2 s 16946 19200 17002 20000 6 prog_clk_0_N_out
port 105 nsew signal tristate
rlabel metal2 s 16946 0 17002 800 6 prog_clk_0_S_out
port 106 nsew signal tristate
rlabel metal3 s 0 2320 800 2440 6 prog_clk_0_W_in
port 107 nsew signal input
rlabel metal3 s 16400 5856 17200 5976 6 right_grid_pin_0_
port 108 nsew signal tristate
rlabel metal4 s 13437 2128 13757 17456 6 VPWR
port 109 nsew power bidirectional
rlabel metal4 s 8440 2128 8760 17456 6 VPWR
port 110 nsew power bidirectional
rlabel metal4 s 3443 2128 3763 17456 6 VPWR
port 111 nsew power bidirectional
rlabel metal4 s 10939 2128 11259 17456 6 VGND
port 112 nsew ground bidirectional
rlabel metal4 s 5941 2128 6261 17456 6 VGND
port 113 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 17200 20000
<< end >>
