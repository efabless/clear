magic
tech sky130A
magscale 1 2
timestamp 1680199036
<< viali >>
rect 13829 54281 13863 54315
rect 18981 54281 19015 54315
rect 2237 54145 2271 54179
rect 4813 54145 4847 54179
rect 7389 54145 7423 54179
rect 9597 54145 9631 54179
rect 12173 54145 12207 54179
rect 14473 54145 14507 54179
rect 15117 54145 15151 54179
rect 15393 54145 15427 54179
rect 17049 54145 17083 54179
rect 17325 54145 17359 54179
rect 17877 54145 17911 54179
rect 18153 54145 18187 54179
rect 19441 54145 19475 54179
rect 20729 54145 20763 54179
rect 21281 54145 21315 54179
rect 22017 54145 22051 54179
rect 22569 54145 22603 54179
rect 23213 54145 23247 54179
rect 23765 54145 23799 54179
rect 24593 54145 24627 54179
rect 25145 54145 25179 54179
rect 2513 54077 2547 54111
rect 5181 54077 5215 54111
rect 7849 54077 7883 54111
rect 9873 54077 9907 54111
rect 12633 54077 12667 54111
rect 19717 54077 19751 54111
rect 14933 54009 14967 54043
rect 17693 54009 17727 54043
rect 20913 54009 20947 54043
rect 24225 54009 24259 54043
rect 14289 53941 14323 53975
rect 16865 53941 16899 53975
rect 22201 53941 22235 53975
rect 23397 53941 23431 53975
rect 24777 53941 24811 53975
rect 25421 53941 25455 53975
rect 24501 53737 24535 53771
rect 24777 53737 24811 53771
rect 2053 53601 2087 53635
rect 4445 53601 4479 53635
rect 7113 53601 7147 53635
rect 11253 53601 11287 53635
rect 1777 53533 1811 53567
rect 4169 53533 4203 53567
rect 6837 53533 6871 53567
rect 10793 53533 10827 53567
rect 23121 53533 23155 53567
rect 23765 53533 23799 53567
rect 25053 53533 25087 53567
rect 23213 53397 23247 53431
rect 23949 53397 23983 53431
rect 25237 53397 25271 53431
rect 5181 53193 5215 53227
rect 23397 53193 23431 53227
rect 5365 53057 5399 53091
rect 24317 53057 24351 53091
rect 25053 53057 25087 53091
rect 25237 52921 25271 52955
rect 24501 52853 24535 52887
rect 6561 52649 6595 52683
rect 6745 52445 6779 52479
rect 24593 52445 24627 52479
rect 25329 52445 25363 52479
rect 24961 52377 24995 52411
rect 24869 51969 24903 52003
rect 25329 51969 25363 52003
rect 25145 51765 25179 51799
rect 8309 51561 8343 51595
rect 9229 51493 9263 51527
rect 7849 51357 7883 51391
rect 8493 51357 8527 51391
rect 9413 51357 9447 51391
rect 7665 51289 7699 51323
rect 24593 51289 24627 51323
rect 24961 51289 24995 51323
rect 25329 51289 25363 51323
rect 24593 50881 24627 50915
rect 24961 50881 24995 50915
rect 25053 50677 25087 50711
rect 7849 50473 7883 50507
rect 9597 50473 9631 50507
rect 8033 50405 8067 50439
rect 7573 50269 7607 50303
rect 9505 50269 9539 50303
rect 25513 50133 25547 50167
rect 24501 49793 24535 49827
rect 24777 49725 24811 49759
rect 10701 49317 10735 49351
rect 11713 49317 11747 49351
rect 10517 49113 10551 49147
rect 11529 49113 11563 49147
rect 24777 49113 24811 49147
rect 25145 49113 25179 49147
rect 25237 49045 25271 49079
rect 8401 48841 8435 48875
rect 6653 48637 6687 48671
rect 6929 48637 6963 48671
rect 8769 48501 8803 48535
rect 25421 48501 25455 48535
rect 10368 48093 10402 48127
rect 25145 48093 25179 48127
rect 25329 48025 25363 48059
rect 10471 47957 10505 47991
rect 9873 47753 9907 47787
rect 9413 47617 9447 47651
rect 24869 47617 24903 47651
rect 25329 47617 25363 47651
rect 9505 47413 9539 47447
rect 25145 47413 25179 47447
rect 11656 47005 11690 47039
rect 11759 46937 11793 46971
rect 25421 46869 25455 46903
rect 10793 46665 10827 46699
rect 14105 46597 14139 46631
rect 10333 46529 10367 46563
rect 12576 46529 12610 46563
rect 13921 46529 13955 46563
rect 25329 46529 25363 46563
rect 15761 46461 15795 46495
rect 10425 46325 10459 46359
rect 12679 46325 12713 46359
rect 25145 46325 25179 46359
rect 8493 46121 8527 46155
rect 8125 45985 8159 46019
rect 14841 45985 14875 46019
rect 15025 45985 15059 46019
rect 16497 45985 16531 46019
rect 7941 45917 7975 45951
rect 13312 45917 13346 45951
rect 24869 45917 24903 45951
rect 25329 45917 25363 45951
rect 13415 45781 13449 45815
rect 25145 45781 25179 45815
rect 12909 45509 12943 45543
rect 12725 45441 12759 45475
rect 14565 45373 14599 45407
rect 25421 45237 25455 45271
rect 10885 45033 10919 45067
rect 9137 44897 9171 44931
rect 15669 44897 15703 44931
rect 25329 44829 25363 44863
rect 9413 44761 9447 44795
rect 15853 44761 15887 44795
rect 17509 44761 17543 44795
rect 11253 44693 11287 44727
rect 25145 44693 25179 44727
rect 9597 44489 9631 44523
rect 9137 44353 9171 44387
rect 10609 44353 10643 44387
rect 24777 44353 24811 44387
rect 25145 44353 25179 44387
rect 8953 44285 8987 44319
rect 25329 44217 25363 44251
rect 10701 44149 10735 44183
rect 11069 44149 11103 44183
rect 20624 43945 20658 43979
rect 22385 43809 22419 43843
rect 20361 43741 20395 43775
rect 22109 43605 22143 43639
rect 25513 43605 25547 43639
rect 25145 43333 25179 43367
rect 25329 43129 25363 43163
rect 9781 42721 9815 42755
rect 10241 42721 10275 42755
rect 9597 42653 9631 42687
rect 24777 42585 24811 42619
rect 25145 42585 25179 42619
rect 25329 42585 25363 42619
rect 11161 42313 11195 42347
rect 9413 42109 9447 42143
rect 9689 42109 9723 42143
rect 11529 41973 11563 42007
rect 25421 41973 25455 42007
rect 10885 41769 10919 41803
rect 10425 41633 10459 41667
rect 10241 41565 10275 41599
rect 25145 41565 25179 41599
rect 25329 41497 25363 41531
rect 24869 41089 24903 41123
rect 25329 41089 25363 41123
rect 25145 40885 25179 40919
rect 25513 40341 25547 40375
rect 25145 40137 25179 40171
rect 25329 40001 25363 40035
rect 24869 39389 24903 39423
rect 25329 39389 25363 39423
rect 25145 39253 25179 39287
rect 25421 38709 25455 38743
rect 25329 38301 25363 38335
rect 25145 38165 25179 38199
rect 8677 37961 8711 37995
rect 8861 37825 8895 37859
rect 24777 37825 24811 37859
rect 25145 37825 25179 37859
rect 25329 37689 25363 37723
rect 25513 37077 25547 37111
rect 25145 36805 25179 36839
rect 25329 36601 25363 36635
rect 24869 36125 24903 36159
rect 25329 36125 25363 36159
rect 25145 35989 25179 36023
rect 11161 35785 11195 35819
rect 11529 35785 11563 35819
rect 22477 35785 22511 35819
rect 21189 35717 21223 35751
rect 21097 35649 21131 35683
rect 22385 35649 22419 35683
rect 9413 35581 9447 35615
rect 9689 35581 9723 35615
rect 21281 35581 21315 35615
rect 22569 35581 22603 35615
rect 20729 35513 20763 35547
rect 20361 35445 20395 35479
rect 22017 35445 22051 35479
rect 25421 35445 25455 35479
rect 23305 35105 23339 35139
rect 23213 35037 23247 35071
rect 25329 35037 25363 35071
rect 22477 34969 22511 35003
rect 23121 34969 23155 35003
rect 21833 34901 21867 34935
rect 22753 34901 22787 34935
rect 25145 34901 25179 34935
rect 25145 34697 25179 34731
rect 24869 34561 24903 34595
rect 25329 34561 25363 34595
rect 21373 34357 21407 34391
rect 9137 34153 9171 34187
rect 15393 34017 15427 34051
rect 21649 34017 21683 34051
rect 9321 33949 9355 33983
rect 19441 33949 19475 33983
rect 23673 33949 23707 33983
rect 24869 33949 24903 33983
rect 25329 33949 25363 33983
rect 14657 33881 14691 33915
rect 15853 33881 15887 33915
rect 19717 33881 19751 33915
rect 21925 33881 21959 33915
rect 21189 33813 21223 33847
rect 23397 33813 23431 33847
rect 25145 33813 25179 33847
rect 19809 33541 19843 33575
rect 24133 33541 24167 33575
rect 24317 33541 24351 33575
rect 19533 33473 19567 33507
rect 22017 33473 22051 33507
rect 24869 33473 24903 33507
rect 25329 33473 25363 33507
rect 21281 33405 21315 33439
rect 22293 33405 22327 33439
rect 23765 33405 23799 33439
rect 21557 33269 21591 33303
rect 24593 33269 24627 33303
rect 25145 33269 25179 33303
rect 16589 33065 16623 33099
rect 24041 33065 24075 33099
rect 16865 32997 16899 33031
rect 16037 32929 16071 32963
rect 16129 32929 16163 32963
rect 22293 32929 22327 32963
rect 22569 32929 22603 32963
rect 25145 32929 25179 32963
rect 20637 32861 20671 32895
rect 24961 32861 24995 32895
rect 25053 32861 25087 32895
rect 15945 32793 15979 32827
rect 19901 32793 19935 32827
rect 15577 32725 15611 32759
rect 19625 32725 19659 32759
rect 24593 32725 24627 32759
rect 16773 32521 16807 32555
rect 21097 32521 21131 32555
rect 25237 32521 25271 32555
rect 15393 32453 15427 32487
rect 22845 32453 22879 32487
rect 22109 32385 22143 32419
rect 23489 32385 23523 32419
rect 16129 32317 16163 32351
rect 19073 32317 19107 32351
rect 19349 32317 19383 32351
rect 23765 32317 23799 32351
rect 20821 32181 20855 32215
rect 21649 32181 21683 32215
rect 17036 31977 17070 32011
rect 22661 31977 22695 32011
rect 15577 31909 15611 31943
rect 23029 31909 23063 31943
rect 25145 31909 25179 31943
rect 16129 31841 16163 31875
rect 18521 31841 18555 31875
rect 19717 31841 19751 31875
rect 22109 31841 22143 31875
rect 22201 31841 22235 31875
rect 23581 31841 23615 31875
rect 16773 31773 16807 31807
rect 19441 31773 19475 31807
rect 23489 31773 23523 31807
rect 24869 31773 24903 31807
rect 25329 31773 25363 31807
rect 15945 31705 15979 31739
rect 18797 31705 18831 31739
rect 23397 31705 23431 31739
rect 16037 31637 16071 31671
rect 21189 31637 21223 31671
rect 21649 31637 21683 31671
rect 22017 31637 22051 31671
rect 24685 31637 24719 31671
rect 16497 31433 16531 31467
rect 19165 31433 19199 31467
rect 21281 31433 21315 31467
rect 15485 31365 15519 31399
rect 17693 31365 17727 31399
rect 19809 31365 19843 31399
rect 20453 31365 20487 31399
rect 22753 31365 22787 31399
rect 17417 31297 17451 31331
rect 19441 31297 19475 31331
rect 20545 31297 20579 31331
rect 22477 31297 22511 31331
rect 25329 31297 25363 31331
rect 13369 31229 13403 31263
rect 13645 31229 13679 31263
rect 16681 31229 16715 31263
rect 20637 31229 20671 31263
rect 21557 31229 21591 31263
rect 20085 31161 20119 31195
rect 24225 31161 24259 31195
rect 15117 31093 15151 31127
rect 24593 31093 24627 31127
rect 25145 31093 25179 31127
rect 9137 30889 9171 30923
rect 15577 30889 15611 30923
rect 15761 30889 15795 30923
rect 18521 30889 18555 30923
rect 22477 30889 22511 30923
rect 25513 30889 25547 30923
rect 16773 30753 16807 30787
rect 20729 30753 20763 30787
rect 9321 30685 9355 30719
rect 14381 30685 14415 30719
rect 15117 30617 15151 30651
rect 17049 30617 17083 30651
rect 21005 30617 21039 30651
rect 18797 30549 18831 30583
rect 20085 30549 20119 30583
rect 22845 30549 22879 30583
rect 24593 30549 24627 30583
rect 20269 30345 20303 30379
rect 14105 30277 14139 30311
rect 20361 30277 20395 30311
rect 22477 30277 22511 30311
rect 9137 30209 9171 30243
rect 11805 30209 11839 30243
rect 15853 30209 15887 30243
rect 16957 30209 16991 30243
rect 21281 30209 21315 30243
rect 22385 30209 22419 30243
rect 12081 30141 12115 30175
rect 14841 30141 14875 30175
rect 15945 30141 15979 30175
rect 16037 30141 16071 30175
rect 16773 30141 16807 30175
rect 20545 30141 20579 30175
rect 22661 30141 22695 30175
rect 23305 30141 23339 30175
rect 23581 30141 23615 30175
rect 25053 30141 25087 30175
rect 8953 30073 8987 30107
rect 25329 30073 25363 30107
rect 13553 30005 13587 30039
rect 15485 30005 15519 30039
rect 18889 30005 18923 30039
rect 19901 30005 19935 30039
rect 22017 30005 22051 30039
rect 16497 29801 16531 29835
rect 18797 29801 18831 29835
rect 12909 29733 12943 29767
rect 20177 29733 20211 29767
rect 25145 29733 25179 29767
rect 11161 29665 11195 29699
rect 15853 29665 15887 29699
rect 17049 29665 17083 29699
rect 20729 29665 20763 29699
rect 15669 29597 15703 29631
rect 23397 29597 23431 29631
rect 24041 29597 24075 29631
rect 25329 29597 25363 29631
rect 11437 29529 11471 29563
rect 13185 29529 13219 29563
rect 13645 29529 13679 29563
rect 15577 29529 15611 29563
rect 17325 29529 17359 29563
rect 20637 29529 20671 29563
rect 22937 29529 22971 29563
rect 15209 29461 15243 29495
rect 16313 29461 16347 29495
rect 19441 29461 19475 29495
rect 20545 29461 20579 29495
rect 23213 29461 23247 29495
rect 23857 29461 23891 29495
rect 24501 29461 24535 29495
rect 9505 29257 9539 29291
rect 12541 29257 12575 29291
rect 12633 29257 12667 29291
rect 15117 29257 15151 29291
rect 16037 29257 16071 29291
rect 17877 29257 17911 29291
rect 19165 29257 19199 29291
rect 19257 29257 19291 29291
rect 19993 29257 20027 29291
rect 23949 29257 23983 29291
rect 25421 29257 25455 29291
rect 9873 29189 9907 29223
rect 15945 29189 15979 29223
rect 24041 29189 24075 29223
rect 9965 29121 9999 29155
rect 13369 29121 13403 29155
rect 17233 29121 17267 29155
rect 22201 29121 22235 29155
rect 10057 29053 10091 29087
rect 12725 29053 12759 29087
rect 16129 29053 16163 29087
rect 17325 29053 17359 29087
rect 17417 29053 17451 29087
rect 19441 29053 19475 29087
rect 23029 29053 23063 29087
rect 24225 29053 24259 29087
rect 24777 29053 24811 29087
rect 12173 28985 12207 29019
rect 15577 28985 15611 29019
rect 16865 28985 16899 29019
rect 18061 28985 18095 29019
rect 18797 28985 18831 29019
rect 21833 28985 21867 29019
rect 23581 28985 23615 29019
rect 13632 28917 13666 28951
rect 25237 28917 25271 28951
rect 10885 28713 10919 28747
rect 13553 28713 13587 28747
rect 15945 28713 15979 28747
rect 18889 28713 18923 28747
rect 22845 28713 22879 28747
rect 9137 28577 9171 28611
rect 11437 28577 11471 28611
rect 13185 28577 13219 28611
rect 15301 28577 15335 28611
rect 15393 28577 15427 28611
rect 17417 28577 17451 28611
rect 20085 28577 20119 28611
rect 23305 28577 23339 28611
rect 23397 28577 23431 28611
rect 25145 28577 25179 28611
rect 17141 28509 17175 28543
rect 20637 28509 20671 28543
rect 23857 28509 23891 28543
rect 24961 28509 24995 28543
rect 9413 28441 9447 28475
rect 11713 28441 11747 28475
rect 15209 28441 15243 28475
rect 20913 28441 20947 28475
rect 25053 28441 25087 28475
rect 14841 28373 14875 28407
rect 16037 28373 16071 28407
rect 16221 28373 16255 28407
rect 19441 28373 19475 28407
rect 19809 28373 19843 28407
rect 19901 28373 19935 28407
rect 22385 28373 22419 28407
rect 23213 28373 23247 28407
rect 24041 28373 24075 28407
rect 24593 28373 24627 28407
rect 18981 28169 19015 28203
rect 19717 28169 19751 28203
rect 21557 28169 21591 28203
rect 22477 28169 22511 28203
rect 11069 28101 11103 28135
rect 13737 28101 13771 28135
rect 15577 28101 15611 28135
rect 16405 28101 16439 28135
rect 17233 28101 17267 28135
rect 21097 28101 21131 28135
rect 22385 28101 22419 28135
rect 15669 28033 15703 28067
rect 17325 28033 17359 28067
rect 20361 28033 20395 28067
rect 23213 28033 23247 28067
rect 11713 27965 11747 27999
rect 11989 27965 12023 27999
rect 15761 27965 15795 27999
rect 17417 27965 17451 27999
rect 18061 27965 18095 27999
rect 18613 27965 18647 27999
rect 22569 27965 22603 27999
rect 23489 27965 23523 27999
rect 25237 27965 25271 27999
rect 19349 27897 19383 27931
rect 13461 27829 13495 27863
rect 15209 27829 15243 27863
rect 16313 27829 16347 27863
rect 16865 27829 16899 27863
rect 18705 27829 18739 27863
rect 22017 27829 22051 27863
rect 24961 27829 24995 27863
rect 25421 27829 25455 27863
rect 20164 27625 20198 27659
rect 23857 27625 23891 27659
rect 12633 27557 12667 27591
rect 10517 27489 10551 27523
rect 10793 27489 10827 27523
rect 12265 27489 12299 27523
rect 13553 27489 13587 27523
rect 15761 27489 15795 27523
rect 18061 27489 18095 27523
rect 19901 27489 19935 27523
rect 22109 27489 22143 27523
rect 24133 27489 24167 27523
rect 25053 27489 25087 27523
rect 25145 27489 25179 27523
rect 13461 27421 13495 27455
rect 15669 27421 15703 27455
rect 16405 27421 16439 27455
rect 17877 27421 17911 27455
rect 24961 27421 24995 27455
rect 13369 27353 13403 27387
rect 15577 27353 15611 27387
rect 22385 27353 22419 27387
rect 13001 27285 13035 27319
rect 15209 27285 15243 27319
rect 16221 27285 16255 27319
rect 17509 27285 17543 27319
rect 17969 27285 18003 27319
rect 21649 27285 21683 27319
rect 24593 27285 24627 27319
rect 11069 27081 11103 27115
rect 11621 27081 11655 27115
rect 15669 27081 15703 27115
rect 22845 27081 22879 27115
rect 25329 27081 25363 27115
rect 9597 27013 9631 27047
rect 13369 27013 13403 27047
rect 15761 27013 15795 27047
rect 13093 26945 13127 26979
rect 17969 26945 18003 26979
rect 22753 26945 22787 26979
rect 9321 26877 9355 26911
rect 15853 26877 15887 26911
rect 18245 26877 18279 26911
rect 23029 26877 23063 26911
rect 23581 26877 23615 26911
rect 23857 26877 23891 26911
rect 14841 26741 14875 26775
rect 15301 26741 15335 26775
rect 19717 26741 19751 26775
rect 20085 26741 20119 26775
rect 21833 26741 21867 26775
rect 22385 26741 22419 26775
rect 10885 26537 10919 26571
rect 15301 26537 15335 26571
rect 16957 26537 16991 26571
rect 21189 26537 21223 26571
rect 23857 26537 23891 26571
rect 11253 26469 11287 26503
rect 15669 26469 15703 26503
rect 17233 26469 17267 26503
rect 22661 26469 22695 26503
rect 24593 26469 24627 26503
rect 9413 26401 9447 26435
rect 14749 26401 14783 26435
rect 14841 26401 14875 26435
rect 16221 26401 16255 26435
rect 16773 26401 16807 26435
rect 19441 26401 19475 26435
rect 19717 26401 19751 26435
rect 23213 26401 23247 26435
rect 25237 26401 25271 26435
rect 9137 26333 9171 26367
rect 14657 26333 14691 26367
rect 23121 26333 23155 26367
rect 24041 26333 24075 26367
rect 24961 26333 24995 26367
rect 16037 26265 16071 26299
rect 16129 26265 16163 26299
rect 17141 26265 17175 26299
rect 21465 26265 21499 26299
rect 22385 26265 22419 26299
rect 23029 26265 23063 26299
rect 25053 26265 25087 26299
rect 14289 26197 14323 26231
rect 18245 26197 18279 26231
rect 12633 25993 12667 26027
rect 14841 25993 14875 26027
rect 15301 25993 15335 26027
rect 17785 25993 17819 26027
rect 18153 25993 18187 26027
rect 22477 25993 22511 26027
rect 18245 25925 18279 25959
rect 22385 25925 22419 25959
rect 12541 25857 12575 25891
rect 13921 25857 13955 25891
rect 15209 25857 15243 25891
rect 16037 25857 16071 25891
rect 17049 25857 17083 25891
rect 17417 25857 17451 25891
rect 23489 25857 23523 25891
rect 23949 25857 23983 25891
rect 12725 25789 12759 25823
rect 14013 25789 14047 25823
rect 14105 25789 14139 25823
rect 15393 25789 15427 25823
rect 18429 25789 18463 25823
rect 22569 25789 22603 25823
rect 25145 25789 25179 25823
rect 12173 25721 12207 25755
rect 13553 25721 13587 25755
rect 22017 25721 22051 25755
rect 16865 25653 16899 25687
rect 19073 25653 19107 25687
rect 21557 25653 21591 25687
rect 23305 25653 23339 25687
rect 14289 25449 14323 25483
rect 15393 25449 15427 25483
rect 18153 25449 18187 25483
rect 19257 25449 19291 25483
rect 20821 25449 20855 25483
rect 21557 25449 21591 25483
rect 24501 25449 24535 25483
rect 13001 25381 13035 25415
rect 16957 25381 16991 25415
rect 24593 25381 24627 25415
rect 10885 25313 10919 25347
rect 11161 25313 11195 25347
rect 14841 25313 14875 25347
rect 16313 25313 16347 25347
rect 17141 25245 17175 25279
rect 17785 25245 17819 25279
rect 18337 25245 18371 25279
rect 21005 25245 21039 25279
rect 21741 25245 21775 25279
rect 22661 25245 22695 25279
rect 25329 25245 25363 25279
rect 14657 25177 14691 25211
rect 16129 25177 16163 25211
rect 19809 25177 19843 25211
rect 23857 25177 23891 25211
rect 24869 25177 24903 25211
rect 12633 25109 12667 25143
rect 14749 25109 14783 25143
rect 15761 25109 15795 25143
rect 16221 25109 16255 25143
rect 17601 25109 17635 25143
rect 18705 25109 18739 25143
rect 19901 25109 19935 25143
rect 20361 25109 20395 25143
rect 25145 25109 25179 25143
rect 17233 24905 17267 24939
rect 19073 24905 19107 24939
rect 12081 24837 12115 24871
rect 18521 24837 18555 24871
rect 22477 24837 22511 24871
rect 12173 24769 12207 24803
rect 13001 24769 13035 24803
rect 15393 24769 15427 24803
rect 17325 24769 17359 24803
rect 18429 24769 18463 24803
rect 19349 24769 19383 24803
rect 19717 24769 19751 24803
rect 22569 24769 22603 24803
rect 9413 24701 9447 24735
rect 9689 24701 9723 24735
rect 12357 24701 12391 24735
rect 13277 24701 13311 24735
rect 14749 24701 14783 24735
rect 17417 24701 17451 24735
rect 18613 24701 18647 24735
rect 19993 24701 20027 24735
rect 21465 24701 21499 24735
rect 22661 24701 22695 24735
rect 23581 24701 23615 24735
rect 23857 24701 23891 24735
rect 25329 24701 25363 24735
rect 11161 24565 11195 24599
rect 11713 24565 11747 24599
rect 15025 24565 15059 24599
rect 16865 24565 16899 24599
rect 18061 24565 18095 24599
rect 22109 24565 22143 24599
rect 21189 24361 21223 24395
rect 25329 24361 25363 24395
rect 14197 24293 14231 24327
rect 25145 24293 25179 24327
rect 11989 24225 12023 24259
rect 18797 24225 18831 24259
rect 19441 24225 19475 24259
rect 21925 24225 21959 24259
rect 24593 24225 24627 24259
rect 9137 24157 9171 24191
rect 11253 24157 11287 24191
rect 11437 24157 11471 24191
rect 17693 24157 17727 24191
rect 18521 24157 18555 24191
rect 9413 24089 9447 24123
rect 12265 24089 12299 24123
rect 15945 24089 15979 24123
rect 19717 24089 19751 24123
rect 22201 24089 22235 24123
rect 10885 24021 10919 24055
rect 13737 24021 13771 24055
rect 18153 24021 18187 24055
rect 18613 24021 18647 24055
rect 21557 24021 21591 24055
rect 23673 24021 23707 24055
rect 23949 24021 23983 24055
rect 25421 24021 25455 24055
rect 9781 23817 9815 23851
rect 10425 23817 10459 23851
rect 10793 23817 10827 23851
rect 14473 23817 14507 23851
rect 14933 23817 14967 23851
rect 17233 23817 17267 23851
rect 18889 23817 18923 23851
rect 24961 23817 24995 23851
rect 25513 23817 25547 23851
rect 13645 23749 13679 23783
rect 13737 23749 13771 23783
rect 8033 23681 8067 23715
rect 14841 23681 14875 23715
rect 17325 23681 17359 23715
rect 18245 23681 18279 23715
rect 19625 23681 19659 23715
rect 20821 23681 20855 23715
rect 22385 23681 22419 23715
rect 8309 23613 8343 23647
rect 10885 23613 10919 23647
rect 10977 23613 11011 23647
rect 13829 23613 13863 23647
rect 15025 23613 15059 23647
rect 15669 23613 15703 23647
rect 17417 23613 17451 23647
rect 18797 23613 18831 23647
rect 19717 23613 19751 23647
rect 19901 23613 19935 23647
rect 20913 23613 20947 23647
rect 21005 23613 21039 23647
rect 23213 23613 23247 23647
rect 23489 23613 23523 23647
rect 18061 23545 18095 23579
rect 10149 23477 10183 23511
rect 13277 23477 13311 23511
rect 16865 23477 16899 23511
rect 18521 23477 18555 23511
rect 19257 23477 19291 23511
rect 20453 23477 20487 23511
rect 21557 23477 21591 23511
rect 22201 23477 22235 23511
rect 25237 23477 25271 23511
rect 9137 23273 9171 23307
rect 14381 23273 14415 23307
rect 15853 23273 15887 23307
rect 14749 23205 14783 23239
rect 17877 23205 17911 23239
rect 18981 23205 19015 23239
rect 9689 23137 9723 23171
rect 11713 23137 11747 23171
rect 11805 23137 11839 23171
rect 13553 23137 13587 23171
rect 15301 23137 15335 23171
rect 18521 23137 18555 23171
rect 19993 23137 20027 23171
rect 20177 23137 20211 23171
rect 20729 23137 20763 23171
rect 25053 23137 25087 23171
rect 25237 23137 25271 23171
rect 13369 23069 13403 23103
rect 15117 23069 15151 23103
rect 18245 23069 18279 23103
rect 19901 23069 19935 23103
rect 21833 23069 21867 23103
rect 22845 23069 22879 23103
rect 24961 23069 24995 23103
rect 9505 23001 9539 23035
rect 11621 23001 11655 23035
rect 13461 23001 13495 23035
rect 14197 23001 14231 23035
rect 15209 23001 15243 23035
rect 23857 23001 23891 23035
rect 9597 22933 9631 22967
rect 11253 22933 11287 22967
rect 13001 22933 13035 22967
rect 18337 22933 18371 22967
rect 19533 22933 19567 22967
rect 21649 22933 21683 22967
rect 24593 22933 24627 22967
rect 10149 22729 10183 22763
rect 14473 22729 14507 22763
rect 16865 22729 16899 22763
rect 18705 22729 18739 22763
rect 19717 22729 19751 22763
rect 21189 22729 21223 22763
rect 18889 22661 18923 22695
rect 8125 22593 8159 22627
rect 12357 22593 12391 22627
rect 17049 22593 17083 22627
rect 21097 22593 21131 22627
rect 22109 22593 22143 22627
rect 23949 22593 23983 22627
rect 8401 22525 8435 22559
rect 12633 22525 12667 22559
rect 21281 22525 21315 22559
rect 23305 22525 23339 22559
rect 24777 22525 24811 22559
rect 9873 22389 9907 22423
rect 14105 22389 14139 22423
rect 20453 22389 20487 22423
rect 20729 22389 20763 22423
rect 21820 22185 21854 22219
rect 23765 22185 23799 22219
rect 11989 22117 12023 22151
rect 8953 22049 8987 22083
rect 11345 22049 11379 22083
rect 12449 22049 12483 22083
rect 12541 22049 12575 22083
rect 15301 22049 15335 22083
rect 15485 22049 15519 22083
rect 20177 22049 20211 22083
rect 20361 22049 20395 22083
rect 21557 22049 21591 22083
rect 23305 22049 23339 22083
rect 25053 22049 25087 22083
rect 25237 22049 25271 22083
rect 16129 21981 16163 22015
rect 23949 21981 23983 22015
rect 11161 21913 11195 21947
rect 16405 21913 16439 21947
rect 18153 21913 18187 21947
rect 24961 21913 24995 21947
rect 10333 21845 10367 21879
rect 10701 21845 10735 21879
rect 11069 21845 11103 21879
rect 12357 21845 12391 21879
rect 14841 21845 14875 21879
rect 15209 21845 15243 21879
rect 17877 21845 17911 21879
rect 19717 21845 19751 21879
rect 20085 21845 20119 21879
rect 20913 21845 20947 21879
rect 24593 21845 24627 21879
rect 9229 21641 9263 21675
rect 10425 21641 10459 21675
rect 11713 21641 11747 21675
rect 15761 21641 15795 21675
rect 21189 21641 21223 21675
rect 21373 21641 21407 21675
rect 22477 21641 22511 21675
rect 25053 21641 25087 21675
rect 13369 21573 13403 21607
rect 9597 21505 9631 21539
rect 10793 21505 10827 21539
rect 15669 21505 15703 21539
rect 18889 21505 18923 21539
rect 19901 21505 19935 21539
rect 20729 21505 20763 21539
rect 22385 21505 22419 21539
rect 23305 21505 23339 21539
rect 6929 21437 6963 21471
rect 7205 21437 7239 21471
rect 9689 21437 9723 21471
rect 9781 21437 9815 21471
rect 10885 21437 10919 21471
rect 10977 21437 11011 21471
rect 13093 21437 13127 21471
rect 19993 21437 20027 21471
rect 20177 21437 20211 21471
rect 22661 21437 22695 21471
rect 23581 21437 23615 21471
rect 15117 21369 15151 21403
rect 18705 21369 18739 21403
rect 8677 21301 8711 21335
rect 14841 21301 14875 21335
rect 19165 21301 19199 21335
rect 19533 21301 19567 21335
rect 21557 21301 21591 21335
rect 22017 21301 22051 21335
rect 25329 21301 25363 21335
rect 21465 21097 21499 21131
rect 12449 21029 12483 21063
rect 19441 21029 19475 21063
rect 20821 21029 20855 21063
rect 9965 20961 9999 20995
rect 15209 20961 15243 20995
rect 19993 20961 20027 20995
rect 22017 20961 22051 20995
rect 23857 20961 23891 20995
rect 25053 20961 25087 20995
rect 25145 20961 25179 20995
rect 10701 20893 10735 20927
rect 19809 20893 19843 20927
rect 20453 20893 20487 20927
rect 21005 20893 21039 20927
rect 22661 20893 22695 20927
rect 10977 20825 11011 20859
rect 15485 20825 15519 20859
rect 19901 20825 19935 20859
rect 21281 20825 21315 20859
rect 9045 20757 9079 20791
rect 12817 20757 12851 20791
rect 14657 20757 14691 20791
rect 16957 20757 16991 20791
rect 17325 20757 17359 20791
rect 18705 20757 18739 20791
rect 24593 20757 24627 20791
rect 24961 20757 24995 20791
rect 10425 20553 10459 20587
rect 10793 20553 10827 20587
rect 15393 20553 15427 20587
rect 15485 20553 15519 20587
rect 20913 20553 20947 20587
rect 21465 20553 21499 20587
rect 25329 20553 25363 20587
rect 8033 20485 8067 20519
rect 10057 20485 10091 20519
rect 17141 20485 17175 20519
rect 20821 20485 20855 20519
rect 16865 20417 16899 20451
rect 19257 20417 19291 20451
rect 19901 20417 19935 20451
rect 22201 20417 22235 20451
rect 22937 20417 22971 20451
rect 7757 20349 7791 20383
rect 9781 20349 9815 20383
rect 10885 20349 10919 20383
rect 10977 20349 11011 20383
rect 12725 20349 12759 20383
rect 13001 20349 13035 20383
rect 15577 20349 15611 20383
rect 18613 20349 18647 20383
rect 21097 20349 21131 20383
rect 23581 20349 23615 20383
rect 23857 20349 23891 20383
rect 22017 20281 22051 20315
rect 14473 20213 14507 20247
rect 15025 20213 15059 20247
rect 19073 20213 19107 20247
rect 19717 20213 19751 20247
rect 20453 20213 20487 20247
rect 22753 20213 22787 20247
rect 8493 20009 8527 20043
rect 11345 20009 11379 20043
rect 16037 20009 16071 20043
rect 16497 20009 16531 20043
rect 23857 20009 23891 20043
rect 11989 19873 12023 19907
rect 14565 19873 14599 19907
rect 16957 19873 16991 19907
rect 17969 19873 18003 19907
rect 18061 19873 18095 19907
rect 19901 19873 19935 19907
rect 22109 19873 22143 19907
rect 24409 19873 24443 19907
rect 9137 19805 9171 19839
rect 14289 19805 14323 19839
rect 16681 19805 16715 19839
rect 17877 19805 17911 19839
rect 18889 19805 18923 19839
rect 9413 19737 9447 19771
rect 11805 19737 11839 19771
rect 20177 19737 20211 19771
rect 22385 19737 22419 19771
rect 10885 19669 10919 19703
rect 11713 19669 11747 19703
rect 17509 19669 17543 19703
rect 18705 19669 18739 19703
rect 21649 19669 21683 19703
rect 24133 19669 24167 19703
rect 25421 19669 25455 19703
rect 8769 19465 8803 19499
rect 10977 19465 11011 19499
rect 11713 19465 11747 19499
rect 15945 19465 15979 19499
rect 16865 19465 16899 19499
rect 17325 19465 17359 19499
rect 18981 19465 19015 19499
rect 20085 19465 20119 19499
rect 20453 19465 20487 19499
rect 20545 19465 20579 19499
rect 22201 19465 22235 19499
rect 22661 19465 22695 19499
rect 25145 19465 25179 19499
rect 25421 19465 25455 19499
rect 9137 19397 9171 19431
rect 23673 19397 23707 19431
rect 15209 19329 15243 19363
rect 16129 19329 16163 19363
rect 17233 19329 17267 19363
rect 19165 19329 19199 19363
rect 21281 19329 21315 19363
rect 22569 19329 22603 19363
rect 23397 19329 23431 19363
rect 6561 19261 6595 19295
rect 6837 19261 6871 19295
rect 9229 19261 9263 19295
rect 9321 19261 9355 19295
rect 12541 19261 12575 19295
rect 12817 19261 12851 19295
rect 17417 19261 17451 19295
rect 20729 19261 20763 19295
rect 22845 19261 22879 19295
rect 15025 19193 15059 19227
rect 8309 19125 8343 19159
rect 11253 19125 11287 19159
rect 14289 19125 14323 19159
rect 14657 19125 14691 19159
rect 21833 19125 21867 19159
rect 8677 18921 8711 18955
rect 10057 18921 10091 18955
rect 11529 18921 11563 18955
rect 12725 18853 12759 18887
rect 6929 18785 6963 18819
rect 10609 18785 10643 18819
rect 12081 18785 12115 18819
rect 13277 18785 13311 18819
rect 17509 18785 17543 18819
rect 23857 18785 23891 18819
rect 6653 18717 6687 18751
rect 11989 18717 12023 18751
rect 13185 18717 13219 18751
rect 17233 18717 17267 18751
rect 17877 18717 17911 18751
rect 21465 18717 21499 18751
rect 22201 18717 22235 18751
rect 22753 18717 22787 18751
rect 24685 18717 24719 18751
rect 13829 18649 13863 18683
rect 24869 18649 24903 18683
rect 8401 18581 8435 18615
rect 9689 18581 9723 18615
rect 10425 18581 10459 18615
rect 10517 18581 10551 18615
rect 11897 18581 11931 18615
rect 13093 18581 13127 18615
rect 14289 18581 14323 18615
rect 16865 18581 16899 18615
rect 17325 18581 17359 18615
rect 18061 18581 18095 18615
rect 21281 18581 21315 18615
rect 22017 18581 22051 18615
rect 10425 18377 10459 18411
rect 13829 18377 13863 18411
rect 14197 18377 14231 18411
rect 14933 18377 14967 18411
rect 8033 18309 8067 18343
rect 11069 18309 11103 18343
rect 12449 18309 12483 18343
rect 17141 18309 17175 18343
rect 23305 18309 23339 18343
rect 10333 18241 10367 18275
rect 16313 18241 16347 18275
rect 16865 18241 16899 18275
rect 21281 18241 21315 18275
rect 22109 18241 22143 18275
rect 23949 18241 23983 18275
rect 7757 18173 7791 18207
rect 10517 18173 10551 18207
rect 13185 18173 13219 18207
rect 14289 18173 14323 18207
rect 14473 18173 14507 18207
rect 24685 18173 24719 18207
rect 9965 18105 9999 18139
rect 9505 18037 9539 18071
rect 16129 18037 16163 18071
rect 18613 18037 18647 18071
rect 18981 18037 19015 18071
rect 21097 18037 21131 18071
rect 7849 17833 7883 17867
rect 12265 17833 12299 17867
rect 18153 17833 18187 17867
rect 19349 17765 19383 17799
rect 20821 17765 20855 17799
rect 8401 17697 8435 17731
rect 10057 17697 10091 17731
rect 11805 17697 11839 17731
rect 12909 17697 12943 17731
rect 17417 17697 17451 17731
rect 17509 17697 17543 17731
rect 18705 17697 18739 17731
rect 23857 17697 23891 17731
rect 25053 17697 25087 17731
rect 25145 17697 25179 17731
rect 9781 17629 9815 17663
rect 12633 17629 12667 17663
rect 17325 17629 17359 17663
rect 19993 17629 20027 17663
rect 21005 17629 21039 17663
rect 22017 17629 22051 17663
rect 22845 17629 22879 17663
rect 8217 17561 8251 17595
rect 18521 17561 18555 17595
rect 18613 17561 18647 17595
rect 19441 17561 19475 17595
rect 22201 17561 22235 17595
rect 7205 17493 7239 17527
rect 8309 17493 8343 17527
rect 9137 17493 9171 17527
rect 12725 17493 12759 17527
rect 13461 17493 13495 17527
rect 15761 17493 15795 17527
rect 16405 17493 16439 17527
rect 16957 17493 16991 17527
rect 19809 17493 19843 17527
rect 24593 17493 24627 17527
rect 24961 17493 24995 17527
rect 8033 17289 8067 17323
rect 9045 17289 9079 17323
rect 9413 17289 9447 17323
rect 11621 17289 11655 17323
rect 13185 17289 13219 17323
rect 17417 17289 17451 17323
rect 20361 17289 20395 17323
rect 22753 17289 22787 17323
rect 10241 17221 10275 17255
rect 11897 17221 11931 17255
rect 16957 17221 16991 17255
rect 17969 17221 18003 17255
rect 18889 17221 18923 17255
rect 20729 17221 20763 17255
rect 10977 17153 11011 17187
rect 13277 17153 13311 17187
rect 14565 17153 14599 17187
rect 18153 17153 18187 17187
rect 21281 17153 21315 17187
rect 22661 17153 22695 17187
rect 23489 17153 23523 17187
rect 8125 17085 8159 17119
rect 8217 17085 8251 17119
rect 9505 17085 9539 17119
rect 9597 17085 9631 17119
rect 13461 17085 13495 17119
rect 14841 17085 14875 17119
rect 18613 17085 18647 17119
rect 22937 17085 22971 17119
rect 23765 17085 23799 17119
rect 12817 17017 12851 17051
rect 17141 17017 17175 17051
rect 7665 16949 7699 16983
rect 16313 16949 16347 16983
rect 22293 16949 22327 16983
rect 25237 16949 25271 16983
rect 13921 16745 13955 16779
rect 14289 16745 14323 16779
rect 24593 16745 24627 16779
rect 10793 16609 10827 16643
rect 11805 16609 11839 16643
rect 12081 16609 12115 16643
rect 15117 16609 15151 16643
rect 16221 16609 16255 16643
rect 16313 16609 16347 16643
rect 17969 16609 18003 16643
rect 19349 16609 19383 16643
rect 20269 16609 20303 16643
rect 16129 16541 16163 16575
rect 16957 16541 16991 16575
rect 17233 16541 17267 16575
rect 18889 16541 18923 16575
rect 19809 16541 19843 16575
rect 22661 16541 22695 16575
rect 23857 16541 23891 16575
rect 24777 16541 24811 16575
rect 10609 16473 10643 16507
rect 14933 16473 14967 16507
rect 20545 16473 20579 16507
rect 9873 16405 9907 16439
rect 10241 16405 10275 16439
rect 10701 16405 10735 16439
rect 13553 16405 13587 16439
rect 14565 16405 14599 16439
rect 15025 16405 15059 16439
rect 15761 16405 15795 16439
rect 18705 16405 18739 16439
rect 19625 16405 19659 16439
rect 22017 16405 22051 16439
rect 22385 16405 22419 16439
rect 25421 16405 25455 16439
rect 8309 16201 8343 16235
rect 8677 16201 8711 16235
rect 12173 16201 12207 16235
rect 12541 16201 12575 16235
rect 14565 16201 14599 16235
rect 15761 16201 15795 16235
rect 16865 16201 16899 16235
rect 24133 16201 24167 16235
rect 13737 16133 13771 16167
rect 17233 16133 17267 16167
rect 20085 16133 20119 16167
rect 6561 16065 6595 16099
rect 12633 16065 12667 16099
rect 14933 16065 14967 16099
rect 15025 16065 15059 16099
rect 18061 16065 18095 16099
rect 18705 16065 18739 16099
rect 19257 16065 19291 16099
rect 21097 16065 21131 16099
rect 22017 16065 22051 16099
rect 24777 16065 24811 16099
rect 6837 15997 6871 16031
rect 12725 15997 12759 16031
rect 13829 15997 13863 16031
rect 13921 15997 13955 16031
rect 15117 15997 15151 16031
rect 21189 15997 21223 16031
rect 21373 15997 21407 16031
rect 22293 15997 22327 16031
rect 24501 15997 24535 16031
rect 16313 15929 16347 15963
rect 13369 15861 13403 15895
rect 17325 15861 17359 15895
rect 17877 15861 17911 15895
rect 18521 15861 18555 15895
rect 20729 15861 20763 15895
rect 23765 15861 23799 15895
rect 9137 15657 9171 15691
rect 10241 15657 10275 15691
rect 11621 15657 11655 15691
rect 18153 15657 18187 15691
rect 18521 15657 18555 15691
rect 24041 15657 24075 15691
rect 25145 15657 25179 15691
rect 9689 15521 9723 15555
rect 12173 15521 12207 15555
rect 16405 15521 16439 15555
rect 16681 15521 16715 15555
rect 19441 15521 19475 15555
rect 22293 15521 22327 15555
rect 22569 15521 22603 15555
rect 24593 15521 24627 15555
rect 21833 15453 21867 15487
rect 9597 15385 9631 15419
rect 11989 15385 12023 15419
rect 19717 15385 19751 15419
rect 9505 15317 9539 15351
rect 12081 15317 12115 15351
rect 14289 15317 14323 15351
rect 15761 15317 15795 15351
rect 21189 15317 21223 15351
rect 21649 15317 21683 15351
rect 10149 15113 10183 15147
rect 12081 15113 12115 15147
rect 14105 15113 14139 15147
rect 15577 15113 15611 15147
rect 15945 15113 15979 15147
rect 20085 15113 20119 15147
rect 10609 15045 10643 15079
rect 18705 15045 18739 15079
rect 21281 15045 21315 15079
rect 23305 15045 23339 15079
rect 10517 14977 10551 15011
rect 19993 14977 20027 15011
rect 21005 14977 21039 15011
rect 22109 14977 22143 15011
rect 24133 14977 24167 15011
rect 7665 14909 7699 14943
rect 7941 14909 7975 14943
rect 9689 14909 9723 14943
rect 10701 14909 10735 14943
rect 14197 14909 14231 14943
rect 14381 14909 14415 14943
rect 16037 14909 16071 14943
rect 16221 14909 16255 14943
rect 20269 14909 20303 14943
rect 24777 14909 24811 14943
rect 13737 14841 13771 14875
rect 18889 14841 18923 14875
rect 19625 14841 19659 14875
rect 20821 14773 20855 14807
rect 8217 14569 8251 14603
rect 8585 14569 8619 14603
rect 12449 14569 12483 14603
rect 21465 14569 21499 14603
rect 9597 14501 9631 14535
rect 16497 14501 16531 14535
rect 6469 14433 6503 14467
rect 10241 14433 10275 14467
rect 13093 14433 13127 14467
rect 14841 14433 14875 14467
rect 17049 14433 17083 14467
rect 21925 14433 21959 14467
rect 22109 14433 22143 14467
rect 23857 14433 23891 14467
rect 9965 14365 9999 14399
rect 14657 14365 14691 14399
rect 15393 14365 15427 14399
rect 20453 14365 20487 14399
rect 22845 14365 22879 14399
rect 25053 14365 25087 14399
rect 6745 14297 6779 14331
rect 11989 14297 12023 14331
rect 16865 14297 16899 14331
rect 17693 14297 17727 14331
rect 12817 14229 12851 14263
rect 12909 14229 12943 14263
rect 13553 14229 13587 14263
rect 14289 14229 14323 14263
rect 14749 14229 14783 14263
rect 16957 14229 16991 14263
rect 20269 14229 20303 14263
rect 21833 14229 21867 14263
rect 24869 14229 24903 14263
rect 12173 14025 12207 14059
rect 13001 14025 13035 14059
rect 15577 14025 15611 14059
rect 15945 14025 15979 14059
rect 18613 14025 18647 14059
rect 19073 14025 19107 14059
rect 20177 14025 20211 14059
rect 25053 14025 25087 14059
rect 8033 13957 8067 13991
rect 9781 13957 9815 13991
rect 10241 13957 10275 13991
rect 18889 13957 18923 13991
rect 19533 13957 19567 13991
rect 7757 13889 7791 13923
rect 10977 13889 11011 13923
rect 20361 13889 20395 13923
rect 21097 13889 21131 13923
rect 22201 13889 22235 13923
rect 25237 13889 25271 13923
rect 11713 13821 11747 13855
rect 13093 13821 13127 13855
rect 13277 13821 13311 13855
rect 13829 13821 13863 13855
rect 16865 13821 16899 13855
rect 19717 13821 19751 13855
rect 22845 13821 22879 13855
rect 24593 13821 24627 13855
rect 20913 13753 20947 13787
rect 22017 13753 22051 13787
rect 12633 13685 12667 13719
rect 14092 13685 14126 13719
rect 17128 13685 17162 13719
rect 23102 13685 23136 13719
rect 8309 13481 8343 13515
rect 8677 13481 8711 13515
rect 9229 13481 9263 13515
rect 10688 13481 10722 13515
rect 14749 13481 14783 13515
rect 17417 13481 17451 13515
rect 24593 13481 24627 13515
rect 21603 13413 21637 13447
rect 25053 13413 25087 13447
rect 6561 13345 6595 13379
rect 6837 13345 6871 13379
rect 9781 13345 9815 13379
rect 10425 13345 10459 13379
rect 13461 13345 13495 13379
rect 15761 13345 15795 13379
rect 18061 13345 18095 13379
rect 23857 13345 23891 13379
rect 15669 13277 15703 13311
rect 19441 13277 19475 13311
rect 20637 13277 20671 13311
rect 21373 13277 21407 13311
rect 22845 13277 22879 13311
rect 24777 13277 24811 13311
rect 9597 13209 9631 13243
rect 12633 13209 12667 13243
rect 15577 13209 15611 13243
rect 17877 13209 17911 13243
rect 18613 13209 18647 13243
rect 18797 13209 18831 13243
rect 20269 13209 20303 13243
rect 9689 13141 9723 13175
rect 12173 13141 12207 13175
rect 13921 13141 13955 13175
rect 15209 13141 15243 13175
rect 16313 13141 16347 13175
rect 6653 12937 6687 12971
rect 9045 12937 9079 12971
rect 9413 12937 9447 12971
rect 10425 12937 10459 12971
rect 10793 12937 10827 12971
rect 12265 12937 12299 12971
rect 15025 12937 15059 12971
rect 15485 12937 15519 12971
rect 16129 12937 16163 12971
rect 17325 12937 17359 12971
rect 19257 12937 19291 12971
rect 21097 12937 21131 12971
rect 21189 12937 21223 12971
rect 22477 12937 22511 12971
rect 22753 12937 22787 12971
rect 25145 12937 25179 12971
rect 13001 12869 13035 12903
rect 14289 12869 14323 12903
rect 15393 12869 15427 12903
rect 23397 12869 23431 12903
rect 7021 12801 7055 12835
rect 8217 12801 8251 12835
rect 9505 12801 9539 12835
rect 10885 12801 10919 12835
rect 13093 12801 13127 12835
rect 14197 12801 14231 12835
rect 17233 12801 17267 12835
rect 18245 12801 18279 12835
rect 19165 12801 19199 12835
rect 20177 12801 20211 12835
rect 22201 12801 22235 12835
rect 7113 12733 7147 12767
rect 7205 12733 7239 12767
rect 8309 12733 8343 12767
rect 8401 12733 8435 12767
rect 9689 12733 9723 12767
rect 10977 12733 11011 12767
rect 13277 12733 13311 12767
rect 14381 12733 14415 12767
rect 15577 12733 15611 12767
rect 17509 12733 17543 12767
rect 19441 12733 19475 12767
rect 21373 12733 21407 12767
rect 23121 12733 23155 12767
rect 7849 12665 7883 12699
rect 19993 12665 20027 12699
rect 12633 12597 12667 12631
rect 13829 12597 13863 12631
rect 16865 12597 16899 12631
rect 18061 12597 18095 12631
rect 18797 12597 18831 12631
rect 20729 12597 20763 12631
rect 22017 12597 22051 12631
rect 24869 12597 24903 12631
rect 10241 12393 10275 12427
rect 11437 12393 11471 12427
rect 12633 12393 12667 12427
rect 16313 12393 16347 12427
rect 20085 12393 20119 12427
rect 22201 12393 22235 12427
rect 24593 12393 24627 12427
rect 14289 12325 14323 12359
rect 7389 12257 7423 12291
rect 8217 12257 8251 12291
rect 10793 12257 10827 12291
rect 11989 12257 12023 12291
rect 13277 12257 13311 12291
rect 14749 12257 14783 12291
rect 14933 12257 14967 12291
rect 18705 12257 18739 12291
rect 20453 12257 20487 12291
rect 20729 12257 20763 12291
rect 11805 12189 11839 12223
rect 13093 12189 13127 12223
rect 17325 12189 17359 12223
rect 19533 12189 19567 12223
rect 22845 12189 22879 12223
rect 24777 12189 24811 12223
rect 10701 12121 10735 12155
rect 18061 12121 18095 12155
rect 23857 12121 23891 12155
rect 10609 12053 10643 12087
rect 11897 12053 11931 12087
rect 13001 12053 13035 12087
rect 14657 12053 14691 12087
rect 16681 12053 16715 12087
rect 19625 12053 19659 12087
rect 9045 11849 9079 11883
rect 9873 11849 9907 11883
rect 11897 11849 11931 11883
rect 13093 11849 13127 11883
rect 14289 11849 14323 11883
rect 17325 11849 17359 11883
rect 18061 11849 18095 11883
rect 18429 11849 18463 11883
rect 9505 11781 9539 11815
rect 10241 11781 10275 11815
rect 10333 11781 10367 11815
rect 12265 11781 12299 11815
rect 20085 11781 20119 11815
rect 21373 11781 21407 11815
rect 23305 11781 23339 11815
rect 9321 11713 9355 11747
rect 13461 11713 13495 11747
rect 14657 11713 14691 11747
rect 17233 11713 17267 11747
rect 19349 11713 19383 11747
rect 21189 11713 21223 11747
rect 22293 11713 22327 11747
rect 24133 11713 24167 11747
rect 7297 11645 7331 11679
rect 7573 11645 7607 11679
rect 10425 11645 10459 11679
rect 12357 11645 12391 11679
rect 12449 11645 12483 11679
rect 13553 11645 13587 11679
rect 13737 11645 13771 11679
rect 14749 11645 14783 11679
rect 14933 11645 14967 11679
rect 17417 11645 17451 11679
rect 18521 11645 18555 11679
rect 18705 11645 18739 11679
rect 20729 11645 20763 11679
rect 24777 11645 24811 11679
rect 16865 11577 16899 11611
rect 19441 11509 19475 11543
rect 20177 11509 20211 11543
rect 12633 11305 12667 11339
rect 19625 11305 19659 11339
rect 25053 11305 25087 11339
rect 11437 11237 11471 11271
rect 13645 11237 13679 11271
rect 16681 11237 16715 11271
rect 17049 11237 17083 11271
rect 18153 11237 18187 11271
rect 21557 11237 21591 11271
rect 9413 11169 9447 11203
rect 11897 11169 11931 11203
rect 11989 11169 12023 11203
rect 13277 11169 13311 11203
rect 14933 11169 14967 11203
rect 18613 11169 18647 11203
rect 18797 11169 18831 11203
rect 20269 11169 20303 11203
rect 9137 11101 9171 11135
rect 13001 11101 13035 11135
rect 19257 11101 19291 11135
rect 19993 11101 20027 11135
rect 20913 11101 20947 11135
rect 21741 11101 21775 11135
rect 22845 11101 22879 11135
rect 25237 11101 25271 11135
rect 13093 11033 13127 11067
rect 15209 11033 15243 11067
rect 18521 11033 18555 11067
rect 23857 11033 23891 11067
rect 10885 10965 10919 10999
rect 11805 10965 11839 10999
rect 14289 10965 14323 10999
rect 20085 10965 20119 10999
rect 21005 10965 21039 10999
rect 22109 10965 22143 10999
rect 9965 10761 9999 10795
rect 12725 10761 12759 10795
rect 20729 10761 20763 10795
rect 8493 10693 8527 10727
rect 10333 10693 10367 10727
rect 10977 10693 11011 10727
rect 12817 10693 12851 10727
rect 17601 10693 17635 10727
rect 21189 10693 21223 10727
rect 23397 10693 23431 10727
rect 14197 10625 14231 10659
rect 14289 10625 14323 10659
rect 15945 10625 15979 10659
rect 17049 10625 17083 10659
rect 18429 10625 18463 10659
rect 19073 10625 19107 10659
rect 19901 10625 19935 10659
rect 21097 10625 21131 10659
rect 22201 10625 22235 10659
rect 23121 10625 23155 10659
rect 8217 10557 8251 10591
rect 11713 10557 11747 10591
rect 12909 10557 12943 10591
rect 14473 10557 14507 10591
rect 16037 10557 16071 10591
rect 16221 10557 16255 10591
rect 19993 10557 20027 10591
rect 20177 10557 20211 10591
rect 21281 10557 21315 10591
rect 22569 10557 22603 10591
rect 25145 10557 25179 10591
rect 13829 10489 13863 10523
rect 15577 10489 15611 10523
rect 18245 10489 18279 10523
rect 12357 10421 12391 10455
rect 16865 10421 16899 10455
rect 17693 10421 17727 10455
rect 18889 10421 18923 10455
rect 19533 10421 19567 10455
rect 22017 10421 22051 10455
rect 24869 10421 24903 10455
rect 11069 10217 11103 10251
rect 11621 10217 11655 10251
rect 12817 10217 12851 10251
rect 14565 10217 14599 10251
rect 24593 10217 24627 10251
rect 17969 10149 18003 10183
rect 20177 10149 20211 10183
rect 22293 10149 22327 10183
rect 9321 10081 9355 10115
rect 12173 10081 12207 10115
rect 13461 10081 13495 10115
rect 15117 10081 15151 10115
rect 18613 10081 18647 10115
rect 19717 10081 19751 10115
rect 20821 10081 20855 10115
rect 23305 10081 23339 10115
rect 23397 10081 23431 10115
rect 13185 10013 13219 10047
rect 20545 10013 20579 10047
rect 24777 10013 24811 10047
rect 9597 9945 9631 9979
rect 11989 9945 12023 9979
rect 14933 9945 14967 9979
rect 16865 9945 16899 9979
rect 19533 9945 19567 9979
rect 12081 9877 12115 9911
rect 13277 9877 13311 9911
rect 13921 9877 13955 9911
rect 15025 9877 15059 9911
rect 16129 9877 16163 9911
rect 16957 9877 16991 9911
rect 18337 9877 18371 9911
rect 18429 9877 18463 9911
rect 18981 9877 19015 9911
rect 22845 9877 22879 9911
rect 23213 9877 23247 9911
rect 22017 9673 22051 9707
rect 24409 9673 24443 9707
rect 11253 9605 11287 9639
rect 14381 9605 14415 9639
rect 15485 9605 15519 9639
rect 11713 9537 11747 9571
rect 14289 9537 14323 9571
rect 20085 9537 20119 9571
rect 21281 9537 21315 9571
rect 25053 9537 25087 9571
rect 11989 9469 12023 9503
rect 13461 9469 13495 9503
rect 14565 9469 14599 9503
rect 15577 9469 15611 9503
rect 15761 9469 15795 9503
rect 17325 9469 17359 9503
rect 17601 9469 17635 9503
rect 22661 9469 22695 9503
rect 22937 9469 22971 9503
rect 13921 9401 13955 9435
rect 15117 9401 15151 9435
rect 25329 9401 25363 9435
rect 19073 9333 19107 9367
rect 19441 9333 19475 9367
rect 24869 9333 24903 9367
rect 11161 9129 11195 9163
rect 14289 9129 14323 9163
rect 24593 9129 24627 9163
rect 13001 9061 13035 9095
rect 15945 9061 15979 9095
rect 9137 8993 9171 9027
rect 13553 8993 13587 9027
rect 14933 8993 14967 9027
rect 16497 8993 16531 9027
rect 17693 8993 17727 9027
rect 19625 8993 19659 9027
rect 14657 8925 14691 8959
rect 16313 8925 16347 8959
rect 22017 8925 22051 8959
rect 22661 8925 22695 8959
rect 24777 8925 24811 8959
rect 9413 8857 9447 8891
rect 13369 8857 13403 8891
rect 18705 8857 18739 8891
rect 18889 8857 18923 8891
rect 19901 8857 19935 8891
rect 23857 8857 23891 8891
rect 10885 8789 10919 8823
rect 13461 8789 13495 8823
rect 14749 8789 14783 8823
rect 16405 8789 16439 8823
rect 17141 8789 17175 8823
rect 17509 8789 17543 8823
rect 17601 8789 17635 8823
rect 21373 8789 21407 8823
rect 21833 8789 21867 8823
rect 22385 8789 22419 8823
rect 17325 8585 17359 8619
rect 13921 8517 13955 8551
rect 15117 8449 15151 8483
rect 17233 8449 17267 8483
rect 17877 8449 17911 8483
rect 18245 8449 18279 8483
rect 20085 8449 20119 8483
rect 22293 8449 22327 8483
rect 23949 8449 23983 8483
rect 11713 8381 11747 8415
rect 13185 8381 13219 8415
rect 14841 8381 14875 8415
rect 16129 8381 16163 8415
rect 17417 8381 17451 8415
rect 19441 8381 19475 8415
rect 21281 8381 21315 8415
rect 22569 8381 22603 8415
rect 24777 8381 24811 8415
rect 14105 8313 14139 8347
rect 16865 8313 16899 8347
rect 11069 8041 11103 8075
rect 13001 8041 13035 8075
rect 15853 8041 15887 8075
rect 24777 8041 24811 8075
rect 19993 7973 20027 8007
rect 11621 7905 11655 7939
rect 13645 7905 13679 7939
rect 14841 7905 14875 7939
rect 16497 7905 16531 7939
rect 18705 7905 18739 7939
rect 22385 7905 22419 7939
rect 11437 7837 11471 7871
rect 13369 7837 13403 7871
rect 14657 7837 14691 7871
rect 16313 7837 16347 7871
rect 17693 7837 17727 7871
rect 19625 7837 19659 7871
rect 20453 7837 20487 7871
rect 22109 7837 22143 7871
rect 11529 7769 11563 7803
rect 13461 7769 13495 7803
rect 14749 7769 14783 7803
rect 21465 7769 21499 7803
rect 24685 7769 24719 7803
rect 12357 7701 12391 7735
rect 14289 7701 14323 7735
rect 16221 7701 16255 7735
rect 19441 7701 19475 7735
rect 23857 7701 23891 7735
rect 24225 7701 24259 7735
rect 12265 7497 12299 7531
rect 12633 7497 12667 7531
rect 15485 7497 15519 7531
rect 17785 7497 17819 7531
rect 16313 7429 16347 7463
rect 21097 7429 21131 7463
rect 25145 7429 25179 7463
rect 9045 7361 9079 7395
rect 16129 7361 16163 7395
rect 17693 7361 17727 7395
rect 18521 7361 18555 7395
rect 22293 7361 22327 7395
rect 23949 7361 23983 7395
rect 9321 7293 9355 7327
rect 12725 7293 12759 7327
rect 12817 7293 12851 7327
rect 13737 7293 13771 7327
rect 14013 7293 14047 7327
rect 17877 7293 17911 7327
rect 18797 7293 18831 7327
rect 21189 7293 21223 7327
rect 21281 7293 21315 7327
rect 23305 7293 23339 7327
rect 10793 7157 10827 7191
rect 11161 7157 11195 7191
rect 16681 7157 16715 7191
rect 17049 7157 17083 7191
rect 17325 7157 17359 7191
rect 20269 7157 20303 7191
rect 20729 7157 20763 7191
rect 15025 6885 15059 6919
rect 10793 6817 10827 6851
rect 12541 6817 12575 6851
rect 12909 6817 12943 6851
rect 15577 6817 15611 6851
rect 18889 6817 18923 6851
rect 20085 6817 20119 6851
rect 25145 6817 25179 6851
rect 13737 6749 13771 6783
rect 14565 6749 14599 6783
rect 17141 6749 17175 6783
rect 19809 6749 19843 6783
rect 20453 6749 20487 6783
rect 20913 6749 20947 6783
rect 22661 6749 22695 6783
rect 23857 6749 23891 6783
rect 11069 6681 11103 6715
rect 15393 6681 15427 6715
rect 15485 6681 15519 6715
rect 16497 6681 16531 6715
rect 16681 6681 16715 6715
rect 17417 6681 17451 6715
rect 22017 6681 22051 6715
rect 25053 6681 25087 6715
rect 13553 6613 13587 6647
rect 14381 6613 14415 6647
rect 16129 6613 16163 6647
rect 19441 6613 19475 6647
rect 19901 6613 19935 6647
rect 24593 6613 24627 6647
rect 24961 6613 24995 6647
rect 10425 6409 10459 6443
rect 11713 6409 11747 6443
rect 13829 6409 13863 6443
rect 24869 6409 24903 6443
rect 12725 6341 12759 6375
rect 24225 6341 24259 6375
rect 10793 6273 10827 6307
rect 12081 6273 12115 6307
rect 12173 6273 12207 6307
rect 13737 6273 13771 6307
rect 14381 6273 14415 6307
rect 15117 6273 15151 6307
rect 17601 6273 17635 6307
rect 18245 6273 18279 6307
rect 20269 6273 20303 6307
rect 22017 6273 22051 6307
rect 25053 6273 25087 6307
rect 10885 6205 10919 6239
rect 10977 6205 11011 6239
rect 12357 6205 12391 6239
rect 12909 6205 12943 6239
rect 13921 6205 13955 6239
rect 16129 6205 16163 6239
rect 16865 6205 16899 6239
rect 19441 6205 19475 6239
rect 21281 6205 21315 6239
rect 22293 6205 22327 6239
rect 23765 6205 23799 6239
rect 13369 6069 13403 6103
rect 17693 6069 17727 6103
rect 25329 6069 25363 6103
rect 11805 5865 11839 5899
rect 14749 5865 14783 5899
rect 16208 5865 16242 5899
rect 17693 5865 17727 5899
rect 23857 5865 23891 5899
rect 18153 5797 18187 5831
rect 24869 5797 24903 5831
rect 10333 5729 10367 5763
rect 15209 5729 15243 5763
rect 15301 5729 15335 5763
rect 18705 5729 18739 5763
rect 19901 5729 19935 5763
rect 21741 5729 21775 5763
rect 10057 5661 10091 5695
rect 12081 5661 12115 5695
rect 13737 5661 13771 5695
rect 14473 5661 14507 5695
rect 15945 5661 15979 5695
rect 18613 5661 18647 5695
rect 19625 5661 19659 5695
rect 21281 5661 21315 5695
rect 23213 5661 23247 5695
rect 24041 5661 24075 5695
rect 24685 5661 24719 5695
rect 23397 5593 23431 5627
rect 13553 5525 13587 5559
rect 15117 5525 15151 5559
rect 18521 5525 18555 5559
rect 20545 5321 20579 5355
rect 21557 5321 21591 5355
rect 13461 5253 13495 5287
rect 22937 5253 22971 5287
rect 15761 5185 15795 5219
rect 17141 5185 17175 5219
rect 18797 5185 18831 5219
rect 21097 5185 21131 5219
rect 22109 5185 22143 5219
rect 23857 5185 23891 5219
rect 13185 5117 13219 5151
rect 15485 5117 15519 5151
rect 18153 5117 18187 5151
rect 19073 5117 19107 5151
rect 24317 5117 24351 5151
rect 21281 5049 21315 5083
rect 14933 4981 14967 5015
rect 16865 4777 16899 4811
rect 21281 4777 21315 4811
rect 24777 4777 24811 4811
rect 12265 4709 12299 4743
rect 14473 4709 14507 4743
rect 5089 4641 5123 4675
rect 13185 4641 13219 4675
rect 15117 4641 15151 4675
rect 17877 4641 17911 4675
rect 19533 4641 19567 4675
rect 19809 4641 19843 4675
rect 22201 4641 22235 4675
rect 7389 4573 7423 4607
rect 12449 4573 12483 4607
rect 12909 4573 12943 4607
rect 14657 4573 14691 4607
rect 17601 4573 17635 4607
rect 21925 4573 21959 4607
rect 23673 4573 23707 4607
rect 24685 4573 24719 4607
rect 5365 4505 5399 4539
rect 7113 4505 7147 4539
rect 15393 4505 15427 4539
rect 1501 4437 1535 4471
rect 11253 4437 11287 4471
rect 14197 4437 14231 4471
rect 23765 4437 23799 4471
rect 24225 4437 24259 4471
rect 11161 4233 11195 4267
rect 16129 4233 16163 4267
rect 21557 4233 21591 4267
rect 14197 4165 14231 4199
rect 22937 4165 22971 4199
rect 1777 4097 1811 4131
rect 2421 4097 2455 4131
rect 2697 4097 2731 4131
rect 4353 4097 4387 4131
rect 4629 4097 4663 4131
rect 9505 4097 9539 4131
rect 9781 4097 9815 4131
rect 10885 4097 10919 4131
rect 10977 4097 11011 4131
rect 12265 4097 12299 4131
rect 13921 4097 13955 4131
rect 17049 4097 17083 4131
rect 18797 4097 18831 4131
rect 20913 4097 20947 4131
rect 21005 4097 21039 4131
rect 22017 4097 22051 4131
rect 23857 4097 23891 4131
rect 13277 4029 13311 4063
rect 17325 4029 17359 4063
rect 19165 4029 19199 4063
rect 21189 4029 21223 4063
rect 24317 4029 24351 4063
rect 1593 3961 1627 3995
rect 2237 3961 2271 3995
rect 4169 3961 4203 3995
rect 9321 3961 9355 3995
rect 15669 3961 15703 3995
rect 2881 3893 2915 3927
rect 10609 3893 10643 3927
rect 11621 3893 11655 3927
rect 11805 3893 11839 3927
rect 20545 3893 20579 3927
rect 2881 3689 2915 3723
rect 4261 3689 4295 3723
rect 8401 3689 8435 3723
rect 17969 3689 18003 3723
rect 18797 3689 18831 3723
rect 23121 3689 23155 3723
rect 6377 3621 6411 3655
rect 7113 3621 7147 3655
rect 24961 3621 24995 3655
rect 1593 3553 1627 3587
rect 5181 3553 5215 3587
rect 11069 3553 11103 3587
rect 12817 3553 12851 3587
rect 14749 3553 14783 3587
rect 16589 3553 16623 3587
rect 19901 3553 19935 3587
rect 21741 3553 21775 3587
rect 23857 3553 23891 3587
rect 1869 3485 1903 3519
rect 3065 3485 3099 3519
rect 3525 3485 3559 3519
rect 4445 3485 4479 3519
rect 4905 3485 4939 3519
rect 6101 3485 6135 3519
rect 6561 3485 6595 3519
rect 7297 3485 7331 3519
rect 7757 3485 7791 3519
rect 8585 3485 8619 3519
rect 8953 3485 8987 3519
rect 9413 3485 9447 3519
rect 9873 3485 9907 3519
rect 10609 3485 10643 3519
rect 11345 3485 11379 3519
rect 12449 3485 12483 3519
rect 14473 3485 14507 3519
rect 16313 3485 16347 3519
rect 18153 3485 18187 3519
rect 19441 3485 19475 3519
rect 21281 3485 21315 3519
rect 23305 3485 23339 3519
rect 25145 3485 25179 3519
rect 18705 3417 18739 3451
rect 3433 3349 3467 3383
rect 7573 3349 7607 3383
rect 9689 3349 9723 3383
rect 10425 3349 10459 3383
rect 4537 3145 4571 3179
rect 4813 3145 4847 3179
rect 6561 3145 6595 3179
rect 10977 3145 11011 3179
rect 20637 3145 20671 3179
rect 21281 3145 21315 3179
rect 22753 3145 22787 3179
rect 24869 3145 24903 3179
rect 9413 3077 9447 3111
rect 22109 3077 22143 3111
rect 2145 3009 2179 3043
rect 3433 3009 3467 3043
rect 3709 3009 3743 3043
rect 5457 3009 5491 3043
rect 6745 3009 6779 3043
rect 7389 3009 7423 3043
rect 8125 3009 8159 3043
rect 9229 3009 9263 3043
rect 9873 3009 9907 3043
rect 10517 3009 10551 3043
rect 11161 3009 11195 3043
rect 11713 3009 11747 3043
rect 11989 3009 12023 3043
rect 13185 3009 13219 3043
rect 14841 3009 14875 3043
rect 17049 3009 17083 3043
rect 18889 3009 18923 3043
rect 20821 3009 20855 3043
rect 23581 3009 23615 3043
rect 2421 2941 2455 2975
rect 5181 2941 5215 2975
rect 7849 2941 7883 2975
rect 13645 2941 13679 2975
rect 15301 2941 15335 2975
rect 17325 2941 17359 2975
rect 19165 2941 19199 2975
rect 22293 2941 22327 2975
rect 9689 2873 9723 2907
rect 7205 2805 7239 2839
rect 9045 2805 9079 2839
rect 10333 2805 10367 2839
rect 4537 2601 4571 2635
rect 18705 2601 18739 2635
rect 21281 2601 21315 2635
rect 25421 2601 25455 2635
rect 24593 2533 24627 2567
rect 2881 2465 2915 2499
rect 5457 2465 5491 2499
rect 14105 2465 14139 2499
rect 14933 2465 14967 2499
rect 17325 2465 17359 2499
rect 22477 2465 22511 2499
rect 2605 2397 2639 2431
rect 3985 2397 4019 2431
rect 4721 2397 4755 2431
rect 5181 2397 5215 2431
rect 6561 2397 6595 2431
rect 7297 2397 7331 2431
rect 8033 2397 8067 2431
rect 8585 2397 8619 2431
rect 9321 2397 9355 2431
rect 9873 2397 9907 2431
rect 11897 2397 11931 2431
rect 12541 2397 12575 2431
rect 14657 2397 14691 2431
rect 16129 2397 16163 2431
rect 16865 2397 16899 2431
rect 18889 2397 18923 2431
rect 19625 2397 19659 2431
rect 20361 2397 20395 2431
rect 21465 2397 21499 2431
rect 22017 2397 22051 2431
rect 24041 2397 24075 2431
rect 24777 2397 24811 2431
rect 4261 2329 4295 2363
rect 7941 2329 7975 2363
rect 10977 2329 11011 2363
rect 13277 2329 13311 2363
rect 16313 2329 16347 2363
rect 3801 2261 3835 2295
rect 6377 2261 6411 2295
rect 6745 2261 6779 2295
rect 7113 2261 7147 2295
rect 7757 2261 7791 2295
rect 8401 2261 8435 2295
rect 9137 2261 9171 2295
rect 11713 2261 11747 2295
rect 23857 2261 23891 2295
<< metal1 >>
rect 1104 54426 25852 54448
rect 1104 54374 7950 54426
rect 8002 54374 8014 54426
rect 8066 54374 8078 54426
rect 8130 54374 8142 54426
rect 8194 54374 8206 54426
rect 8258 54374 17950 54426
rect 18002 54374 18014 54426
rect 18066 54374 18078 54426
rect 18130 54374 18142 54426
rect 18194 54374 18206 54426
rect 18258 54374 25852 54426
rect 1104 54352 25852 54374
rect 13814 54272 13820 54324
rect 13872 54272 13878 54324
rect 18966 54272 18972 54324
rect 19024 54272 19030 54324
rect 2225 54179 2283 54185
rect 2225 54145 2237 54179
rect 2271 54176 2283 54179
rect 4062 54176 4068 54188
rect 2271 54148 4068 54176
rect 2271 54145 2283 54148
rect 2225 54139 2283 54145
rect 4062 54136 4068 54148
rect 4120 54136 4126 54188
rect 4798 54136 4804 54188
rect 4856 54136 4862 54188
rect 7374 54136 7380 54188
rect 7432 54136 7438 54188
rect 9582 54136 9588 54188
rect 9640 54136 9646 54188
rect 11698 54136 11704 54188
rect 11756 54176 11762 54188
rect 12161 54179 12219 54185
rect 12161 54176 12173 54179
rect 11756 54148 12173 54176
rect 11756 54136 11762 54148
rect 12161 54145 12173 54148
rect 12207 54145 12219 54179
rect 13832 54176 13860 54272
rect 14568 54216 18276 54244
rect 14461 54179 14519 54185
rect 14461 54176 14473 54179
rect 13832 54148 14473 54176
rect 12161 54139 12219 54145
rect 14461 54145 14473 54148
rect 14507 54145 14519 54179
rect 14461 54139 14519 54145
rect 2406 54068 2412 54120
rect 2464 54108 2470 54120
rect 2501 54111 2559 54117
rect 2501 54108 2513 54111
rect 2464 54080 2513 54108
rect 2464 54068 2470 54080
rect 2501 54077 2513 54080
rect 2547 54077 2559 54111
rect 2501 54071 2559 54077
rect 5166 54068 5172 54120
rect 5224 54068 5230 54120
rect 7834 54068 7840 54120
rect 7892 54068 7898 54120
rect 9306 54068 9312 54120
rect 9364 54108 9370 54120
rect 9861 54111 9919 54117
rect 9861 54108 9873 54111
rect 9364 54080 9873 54108
rect 9364 54068 9370 54080
rect 9861 54077 9873 54080
rect 9907 54077 9919 54111
rect 9861 54071 9919 54077
rect 12342 54068 12348 54120
rect 12400 54108 12406 54120
rect 12621 54111 12679 54117
rect 12621 54108 12633 54111
rect 12400 54080 12633 54108
rect 12400 54068 12406 54080
rect 12621 54077 12633 54080
rect 12667 54077 12679 54111
rect 14568 54108 14596 54216
rect 14826 54136 14832 54188
rect 14884 54176 14890 54188
rect 15105 54179 15163 54185
rect 15105 54176 15117 54179
rect 14884 54148 15117 54176
rect 14884 54136 14890 54148
rect 15105 54145 15117 54148
rect 15151 54176 15163 54179
rect 15381 54179 15439 54185
rect 15381 54176 15393 54179
rect 15151 54148 15393 54176
rect 15151 54145 15163 54148
rect 15105 54139 15163 54145
rect 15381 54145 15393 54148
rect 15427 54145 15439 54179
rect 15381 54139 15439 54145
rect 16574 54136 16580 54188
rect 16632 54176 16638 54188
rect 17037 54179 17095 54185
rect 17037 54176 17049 54179
rect 16632 54148 17049 54176
rect 16632 54136 16638 54148
rect 17037 54145 17049 54148
rect 17083 54176 17095 54179
rect 17313 54179 17371 54185
rect 17313 54176 17325 54179
rect 17083 54148 17325 54176
rect 17083 54145 17095 54148
rect 17037 54139 17095 54145
rect 17313 54145 17325 54148
rect 17359 54145 17371 54179
rect 17313 54139 17371 54145
rect 17586 54136 17592 54188
rect 17644 54176 17650 54188
rect 17865 54179 17923 54185
rect 17865 54176 17877 54179
rect 17644 54148 17877 54176
rect 17644 54136 17650 54148
rect 17865 54145 17877 54148
rect 17911 54176 17923 54179
rect 18141 54179 18199 54185
rect 18141 54176 18153 54179
rect 17911 54148 18153 54176
rect 17911 54145 17923 54148
rect 17865 54139 17923 54145
rect 18141 54145 18153 54148
rect 18187 54145 18199 54179
rect 18141 54139 18199 54145
rect 12621 54071 12679 54077
rect 12728 54080 14596 54108
rect 8294 54000 8300 54052
rect 8352 54040 8358 54052
rect 12728 54040 12756 54080
rect 16666 54068 16672 54120
rect 16724 54108 16730 54120
rect 18248 54108 18276 54216
rect 18984 54176 19012 54272
rect 19429 54179 19487 54185
rect 19429 54176 19441 54179
rect 18984 54148 19441 54176
rect 19429 54145 19441 54148
rect 19475 54145 19487 54179
rect 19429 54139 19487 54145
rect 20714 54136 20720 54188
rect 20772 54176 20778 54188
rect 21269 54179 21327 54185
rect 21269 54176 21281 54179
rect 20772 54148 21281 54176
rect 20772 54136 20778 54148
rect 21269 54145 21281 54148
rect 21315 54145 21327 54179
rect 21269 54139 21327 54145
rect 21726 54136 21732 54188
rect 21784 54176 21790 54188
rect 22005 54179 22063 54185
rect 22005 54176 22017 54179
rect 21784 54148 22017 54176
rect 21784 54136 21790 54148
rect 22005 54145 22017 54148
rect 22051 54176 22063 54179
rect 22557 54179 22615 54185
rect 22557 54176 22569 54179
rect 22051 54148 22569 54176
rect 22051 54145 22063 54148
rect 22005 54139 22063 54145
rect 22557 54145 22569 54148
rect 22603 54145 22615 54179
rect 22557 54139 22615 54145
rect 23106 54136 23112 54188
rect 23164 54176 23170 54188
rect 23201 54179 23259 54185
rect 23201 54176 23213 54179
rect 23164 54148 23213 54176
rect 23164 54136 23170 54148
rect 23201 54145 23213 54148
rect 23247 54176 23259 54179
rect 23753 54179 23811 54185
rect 23753 54176 23765 54179
rect 23247 54148 23765 54176
rect 23247 54145 23259 54148
rect 23201 54139 23259 54145
rect 23753 54145 23765 54148
rect 23799 54145 23811 54179
rect 23753 54139 23811 54145
rect 24486 54136 24492 54188
rect 24544 54176 24550 54188
rect 24581 54179 24639 54185
rect 24581 54176 24593 54179
rect 24544 54148 24593 54176
rect 24544 54136 24550 54148
rect 24581 54145 24593 54148
rect 24627 54176 24639 54179
rect 25133 54179 25191 54185
rect 25133 54176 25145 54179
rect 24627 54148 25145 54176
rect 24627 54145 24639 54148
rect 24581 54139 24639 54145
rect 25133 54145 25145 54148
rect 25179 54145 25191 54179
rect 25133 54139 25191 54145
rect 19705 54111 19763 54117
rect 19705 54108 19717 54111
rect 16724 54080 17816 54108
rect 18248 54080 19717 54108
rect 16724 54068 16730 54080
rect 8352 54012 12756 54040
rect 8352 54000 8358 54012
rect 13906 54000 13912 54052
rect 13964 54040 13970 54052
rect 14921 54043 14979 54049
rect 14921 54040 14933 54043
rect 13964 54012 14933 54040
rect 13964 54000 13970 54012
rect 14921 54009 14933 54012
rect 14967 54009 14979 54043
rect 14921 54003 14979 54009
rect 16114 54000 16120 54052
rect 16172 54040 16178 54052
rect 17681 54043 17739 54049
rect 17681 54040 17693 54043
rect 16172 54012 17693 54040
rect 16172 54000 16178 54012
rect 17681 54009 17693 54012
rect 17727 54009 17739 54043
rect 17788 54040 17816 54080
rect 19705 54077 19717 54080
rect 19751 54077 19763 54111
rect 19705 54071 19763 54077
rect 20901 54043 20959 54049
rect 20901 54040 20913 54043
rect 17788 54012 20913 54040
rect 17681 54003 17739 54009
rect 20901 54009 20913 54012
rect 20947 54009 20959 54043
rect 20901 54003 20959 54009
rect 24213 54043 24271 54049
rect 24213 54009 24225 54043
rect 24259 54040 24271 54043
rect 25038 54040 25044 54052
rect 24259 54012 25044 54040
rect 24259 54009 24271 54012
rect 24213 54003 24271 54009
rect 25038 54000 25044 54012
rect 25096 54000 25102 54052
rect 12710 53932 12716 53984
rect 12768 53972 12774 53984
rect 14277 53975 14335 53981
rect 14277 53972 14289 53975
rect 12768 53944 14289 53972
rect 12768 53932 12774 53944
rect 14277 53941 14289 53944
rect 14323 53941 14335 53975
rect 14277 53935 14335 53941
rect 15654 53932 15660 53984
rect 15712 53972 15718 53984
rect 16853 53975 16911 53981
rect 16853 53972 16865 53975
rect 15712 53944 16865 53972
rect 15712 53932 15718 53944
rect 16853 53941 16865 53944
rect 16899 53941 16911 53975
rect 16853 53935 16911 53941
rect 22186 53932 22192 53984
rect 22244 53932 22250 53984
rect 22646 53932 22652 53984
rect 22704 53972 22710 53984
rect 23385 53975 23443 53981
rect 23385 53972 23397 53975
rect 22704 53944 23397 53972
rect 22704 53932 22710 53944
rect 23385 53941 23397 53944
rect 23431 53941 23443 53975
rect 23385 53935 23443 53941
rect 24670 53932 24676 53984
rect 24728 53972 24734 53984
rect 24765 53975 24823 53981
rect 24765 53972 24777 53975
rect 24728 53944 24777 53972
rect 24728 53932 24734 53944
rect 24765 53941 24777 53944
rect 24811 53941 24823 53975
rect 24765 53935 24823 53941
rect 25130 53932 25136 53984
rect 25188 53972 25194 53984
rect 25409 53975 25467 53981
rect 25409 53972 25421 53975
rect 25188 53944 25421 53972
rect 25188 53932 25194 53944
rect 25409 53941 25421 53944
rect 25455 53941 25467 53975
rect 25409 53935 25467 53941
rect 1104 53882 25852 53904
rect 1104 53830 2950 53882
rect 3002 53830 3014 53882
rect 3066 53830 3078 53882
rect 3130 53830 3142 53882
rect 3194 53830 3206 53882
rect 3258 53830 12950 53882
rect 13002 53830 13014 53882
rect 13066 53830 13078 53882
rect 13130 53830 13142 53882
rect 13194 53830 13206 53882
rect 13258 53830 22950 53882
rect 23002 53830 23014 53882
rect 23066 53830 23078 53882
rect 23130 53830 23142 53882
rect 23194 53830 23206 53882
rect 23258 53830 25852 53882
rect 1104 53808 25852 53830
rect 24489 53771 24547 53777
rect 24489 53737 24501 53771
rect 24535 53768 24547 53771
rect 24578 53768 24584 53780
rect 24535 53740 24584 53768
rect 24535 53737 24547 53740
rect 24489 53731 24547 53737
rect 10686 53660 10692 53712
rect 10744 53660 10750 53712
rect 1026 53592 1032 53644
rect 1084 53632 1090 53644
rect 2041 53635 2099 53641
rect 2041 53632 2053 53635
rect 1084 53604 2053 53632
rect 1084 53592 1090 53604
rect 2041 53601 2053 53604
rect 2087 53601 2099 53635
rect 2041 53595 2099 53601
rect 3786 53592 3792 53644
rect 3844 53632 3850 53644
rect 4433 53635 4491 53641
rect 4433 53632 4445 53635
rect 3844 53604 4445 53632
rect 3844 53592 3850 53604
rect 4433 53601 4445 53604
rect 4479 53601 4491 53635
rect 4433 53595 4491 53601
rect 6546 53592 6552 53644
rect 6604 53632 6610 53644
rect 7101 53635 7159 53641
rect 7101 53632 7113 53635
rect 6604 53604 7113 53632
rect 6604 53592 6610 53604
rect 7101 53601 7113 53604
rect 7147 53601 7159 53635
rect 10704 53632 10732 53660
rect 11241 53635 11299 53641
rect 11241 53632 11253 53635
rect 10704 53604 11253 53632
rect 7101 53595 7159 53601
rect 11241 53601 11253 53604
rect 11287 53601 11299 53635
rect 11241 53595 11299 53601
rect 1765 53567 1823 53573
rect 1765 53533 1777 53567
rect 1811 53533 1823 53567
rect 1765 53527 1823 53533
rect 1780 53496 1808 53527
rect 4154 53524 4160 53576
rect 4212 53524 4218 53576
rect 6825 53567 6883 53573
rect 6825 53533 6837 53567
rect 6871 53564 6883 53567
rect 7834 53564 7840 53576
rect 6871 53536 7840 53564
rect 6871 53533 6883 53536
rect 6825 53527 6883 53533
rect 7834 53524 7840 53536
rect 7892 53524 7898 53576
rect 10686 53524 10692 53576
rect 10744 53564 10750 53576
rect 10781 53567 10839 53573
rect 10781 53564 10793 53567
rect 10744 53536 10793 53564
rect 10744 53524 10750 53536
rect 10781 53533 10793 53536
rect 10827 53533 10839 53567
rect 10781 53527 10839 53533
rect 23109 53567 23167 53573
rect 23109 53533 23121 53567
rect 23155 53564 23167 53567
rect 23382 53564 23388 53576
rect 23155 53536 23388 53564
rect 23155 53533 23167 53536
rect 23109 53527 23167 53533
rect 23382 53524 23388 53536
rect 23440 53524 23446 53576
rect 23753 53567 23811 53573
rect 23753 53533 23765 53567
rect 23799 53564 23811 53567
rect 24504 53564 24532 53731
rect 24578 53728 24584 53740
rect 24636 53728 24642 53780
rect 24762 53728 24768 53780
rect 24820 53728 24826 53780
rect 23799 53536 24532 53564
rect 23799 53533 23811 53536
rect 23753 53527 23811 53533
rect 25038 53524 25044 53576
rect 25096 53524 25102 53576
rect 5534 53496 5540 53508
rect 1780 53468 5540 53496
rect 5534 53456 5540 53468
rect 5592 53456 5598 53508
rect 22830 53388 22836 53440
rect 22888 53428 22894 53440
rect 23201 53431 23259 53437
rect 23201 53428 23213 53431
rect 22888 53400 23213 53428
rect 22888 53388 22894 53400
rect 23201 53397 23213 53400
rect 23247 53397 23259 53431
rect 23201 53391 23259 53397
rect 23934 53388 23940 53440
rect 23992 53388 23998 53440
rect 25225 53431 25283 53437
rect 25225 53397 25237 53431
rect 25271 53428 25283 53431
rect 26510 53428 26516 53440
rect 25271 53400 26516 53428
rect 25271 53397 25283 53400
rect 25225 53391 25283 53397
rect 26510 53388 26516 53400
rect 26568 53388 26574 53440
rect 1104 53338 25852 53360
rect 1104 53286 7950 53338
rect 8002 53286 8014 53338
rect 8066 53286 8078 53338
rect 8130 53286 8142 53338
rect 8194 53286 8206 53338
rect 8258 53286 17950 53338
rect 18002 53286 18014 53338
rect 18066 53286 18078 53338
rect 18130 53286 18142 53338
rect 18194 53286 18206 53338
rect 18258 53286 25852 53338
rect 1104 53264 25852 53286
rect 4062 53184 4068 53236
rect 4120 53224 4126 53236
rect 5169 53227 5227 53233
rect 5169 53224 5181 53227
rect 4120 53196 5181 53224
rect 4120 53184 4126 53196
rect 5169 53193 5181 53196
rect 5215 53193 5227 53227
rect 5169 53187 5227 53193
rect 23382 53184 23388 53236
rect 23440 53184 23446 53236
rect 5353 53091 5411 53097
rect 5353 53057 5365 53091
rect 5399 53088 5411 53091
rect 7742 53088 7748 53100
rect 5399 53060 7748 53088
rect 5399 53057 5411 53060
rect 5353 53051 5411 53057
rect 7742 53048 7748 53060
rect 7800 53048 7806 53100
rect 24305 53091 24363 53097
rect 24305 53057 24317 53091
rect 24351 53088 24363 53091
rect 24762 53088 24768 53100
rect 24351 53060 24768 53088
rect 24351 53057 24363 53060
rect 24305 53051 24363 53057
rect 24762 53048 24768 53060
rect 24820 53048 24826 53100
rect 25038 53048 25044 53100
rect 25096 53048 25102 53100
rect 15562 52912 15568 52964
rect 15620 52952 15626 52964
rect 25225 52955 25283 52961
rect 25225 52952 25237 52955
rect 15620 52924 25237 52952
rect 15620 52912 15626 52924
rect 25225 52921 25237 52924
rect 25271 52921 25283 52955
rect 25225 52915 25283 52921
rect 24486 52844 24492 52896
rect 24544 52844 24550 52896
rect 1104 52794 25852 52816
rect 1104 52742 2950 52794
rect 3002 52742 3014 52794
rect 3066 52742 3078 52794
rect 3130 52742 3142 52794
rect 3194 52742 3206 52794
rect 3258 52742 12950 52794
rect 13002 52742 13014 52794
rect 13066 52742 13078 52794
rect 13130 52742 13142 52794
rect 13194 52742 13206 52794
rect 13258 52742 22950 52794
rect 23002 52742 23014 52794
rect 23066 52742 23078 52794
rect 23130 52742 23142 52794
rect 23194 52742 23206 52794
rect 23258 52742 25852 52794
rect 1104 52720 25852 52742
rect 4154 52640 4160 52692
rect 4212 52680 4218 52692
rect 6549 52683 6607 52689
rect 6549 52680 6561 52683
rect 4212 52652 6561 52680
rect 4212 52640 4218 52652
rect 6549 52649 6561 52652
rect 6595 52649 6607 52683
rect 6549 52643 6607 52649
rect 16390 52640 16396 52692
rect 16448 52680 16454 52692
rect 24486 52680 24492 52692
rect 16448 52652 24492 52680
rect 16448 52640 16454 52652
rect 24486 52640 24492 52652
rect 24544 52640 24550 52692
rect 6733 52479 6791 52485
rect 6733 52445 6745 52479
rect 6779 52476 6791 52479
rect 9398 52476 9404 52488
rect 6779 52448 9404 52476
rect 6779 52445 6791 52448
rect 6733 52439 6791 52445
rect 9398 52436 9404 52448
rect 9456 52436 9462 52488
rect 24581 52479 24639 52485
rect 24581 52445 24593 52479
rect 24627 52476 24639 52479
rect 25317 52479 25375 52485
rect 24627 52448 24992 52476
rect 24627 52445 24639 52448
rect 24581 52439 24639 52445
rect 24964 52420 24992 52448
rect 25317 52445 25329 52479
rect 25363 52476 25375 52479
rect 26786 52476 26792 52488
rect 25363 52448 26792 52476
rect 25363 52445 25375 52448
rect 25317 52439 25375 52445
rect 26786 52436 26792 52448
rect 26844 52436 26850 52488
rect 24946 52368 24952 52420
rect 25004 52368 25010 52420
rect 1104 52250 25852 52272
rect 1104 52198 7950 52250
rect 8002 52198 8014 52250
rect 8066 52198 8078 52250
rect 8130 52198 8142 52250
rect 8194 52198 8206 52250
rect 8258 52198 17950 52250
rect 18002 52198 18014 52250
rect 18066 52198 18078 52250
rect 18130 52198 18142 52250
rect 18194 52198 18206 52250
rect 18258 52198 25852 52250
rect 1104 52176 25852 52198
rect 24857 52003 24915 52009
rect 24857 51969 24869 52003
rect 24903 52000 24915 52003
rect 25317 52003 25375 52009
rect 25317 52000 25329 52003
rect 24903 51972 25329 52000
rect 24903 51969 24915 51972
rect 24857 51963 24915 51969
rect 25317 51969 25329 51972
rect 25363 52000 25375 52003
rect 25866 52000 25872 52012
rect 25363 51972 25872 52000
rect 25363 51969 25375 51972
rect 25317 51963 25375 51969
rect 25866 51960 25872 51972
rect 25924 51960 25930 52012
rect 24854 51756 24860 51808
rect 24912 51796 24918 51808
rect 25133 51799 25191 51805
rect 25133 51796 25145 51799
rect 24912 51768 25145 51796
rect 24912 51756 24918 51768
rect 25133 51765 25145 51768
rect 25179 51765 25191 51799
rect 25133 51759 25191 51765
rect 1104 51706 25852 51728
rect 1104 51654 2950 51706
rect 3002 51654 3014 51706
rect 3066 51654 3078 51706
rect 3130 51654 3142 51706
rect 3194 51654 3206 51706
rect 3258 51654 12950 51706
rect 13002 51654 13014 51706
rect 13066 51654 13078 51706
rect 13130 51654 13142 51706
rect 13194 51654 13206 51706
rect 13258 51654 22950 51706
rect 23002 51654 23014 51706
rect 23066 51654 23078 51706
rect 23130 51654 23142 51706
rect 23194 51654 23206 51706
rect 23258 51654 25852 51706
rect 1104 51632 25852 51654
rect 7374 51552 7380 51604
rect 7432 51592 7438 51604
rect 8297 51595 8355 51601
rect 8297 51592 8309 51595
rect 7432 51564 8309 51592
rect 7432 51552 7438 51564
rect 8297 51561 8309 51564
rect 8343 51561 8355 51595
rect 8297 51555 8355 51561
rect 7834 51484 7840 51536
rect 7892 51524 7898 51536
rect 9217 51527 9275 51533
rect 9217 51524 9229 51527
rect 7892 51496 9229 51524
rect 7892 51484 7898 51496
rect 9217 51493 9229 51496
rect 9263 51493 9275 51527
rect 9217 51487 9275 51493
rect 4798 51348 4804 51400
rect 4856 51388 4862 51400
rect 7837 51391 7895 51397
rect 7837 51388 7849 51391
rect 4856 51360 7849 51388
rect 4856 51348 4862 51360
rect 7837 51357 7849 51360
rect 7883 51357 7895 51391
rect 7837 51351 7895 51357
rect 8478 51348 8484 51400
rect 8536 51348 8542 51400
rect 9401 51391 9459 51397
rect 9401 51357 9413 51391
rect 9447 51388 9459 51391
rect 10502 51388 10508 51400
rect 9447 51360 10508 51388
rect 9447 51357 9459 51360
rect 9401 51351 9459 51357
rect 10502 51348 10508 51360
rect 10560 51348 10566 51400
rect 7653 51323 7711 51329
rect 7653 51289 7665 51323
rect 7699 51320 7711 51323
rect 10778 51320 10784 51332
rect 7699 51292 10784 51320
rect 7699 51289 7711 51292
rect 7653 51283 7711 51289
rect 10778 51280 10784 51292
rect 10836 51280 10842 51332
rect 24581 51323 24639 51329
rect 24581 51289 24593 51323
rect 24627 51320 24639 51323
rect 24946 51320 24952 51332
rect 24627 51292 24952 51320
rect 24627 51289 24639 51292
rect 24581 51283 24639 51289
rect 24946 51280 24952 51292
rect 25004 51280 25010 51332
rect 25317 51323 25375 51329
rect 25317 51289 25329 51323
rect 25363 51320 25375 51323
rect 26878 51320 26884 51332
rect 25363 51292 26884 51320
rect 25363 51289 25375 51292
rect 25317 51283 25375 51289
rect 26878 51280 26884 51292
rect 26936 51280 26942 51332
rect 1104 51162 25852 51184
rect 1104 51110 7950 51162
rect 8002 51110 8014 51162
rect 8066 51110 8078 51162
rect 8130 51110 8142 51162
rect 8194 51110 8206 51162
rect 8258 51110 17950 51162
rect 18002 51110 18014 51162
rect 18066 51110 18078 51162
rect 18130 51110 18142 51162
rect 18194 51110 18206 51162
rect 18258 51110 25852 51162
rect 1104 51088 25852 51110
rect 24581 50915 24639 50921
rect 24581 50881 24593 50915
rect 24627 50912 24639 50915
rect 24946 50912 24952 50924
rect 24627 50884 24952 50912
rect 24627 50881 24639 50884
rect 24581 50875 24639 50881
rect 24946 50872 24952 50884
rect 25004 50872 25010 50924
rect 25038 50668 25044 50720
rect 25096 50668 25102 50720
rect 1104 50618 25852 50640
rect 1104 50566 2950 50618
rect 3002 50566 3014 50618
rect 3066 50566 3078 50618
rect 3130 50566 3142 50618
rect 3194 50566 3206 50618
rect 3258 50566 12950 50618
rect 13002 50566 13014 50618
rect 13066 50566 13078 50618
rect 13130 50566 13142 50618
rect 13194 50566 13206 50618
rect 13258 50566 22950 50618
rect 23002 50566 23014 50618
rect 23066 50566 23078 50618
rect 23130 50566 23142 50618
rect 23194 50566 23206 50618
rect 23258 50566 25852 50618
rect 1104 50544 25852 50566
rect 5534 50464 5540 50516
rect 5592 50504 5598 50516
rect 7837 50507 7895 50513
rect 7837 50504 7849 50507
rect 5592 50476 7849 50504
rect 5592 50464 5598 50476
rect 7837 50473 7849 50476
rect 7883 50504 7895 50507
rect 8386 50504 8392 50516
rect 7883 50476 8392 50504
rect 7883 50473 7895 50476
rect 7837 50467 7895 50473
rect 8386 50464 8392 50476
rect 8444 50464 8450 50516
rect 9582 50464 9588 50516
rect 9640 50464 9646 50516
rect 16022 50464 16028 50516
rect 16080 50504 16086 50516
rect 25038 50504 25044 50516
rect 16080 50476 25044 50504
rect 16080 50464 16086 50476
rect 25038 50464 25044 50476
rect 25096 50464 25102 50516
rect 7742 50396 7748 50448
rect 7800 50436 7806 50448
rect 8021 50439 8079 50445
rect 8021 50436 8033 50439
rect 7800 50408 8033 50436
rect 7800 50396 7806 50408
rect 8021 50405 8033 50408
rect 8067 50405 8079 50439
rect 8021 50399 8079 50405
rect 7561 50303 7619 50309
rect 7561 50269 7573 50303
rect 7607 50300 7619 50303
rect 8294 50300 8300 50312
rect 7607 50272 8300 50300
rect 7607 50269 7619 50272
rect 7561 50263 7619 50269
rect 8294 50260 8300 50272
rect 8352 50260 8358 50312
rect 9493 50303 9551 50309
rect 9493 50269 9505 50303
rect 9539 50300 9551 50303
rect 9582 50300 9588 50312
rect 9539 50272 9588 50300
rect 9539 50269 9551 50272
rect 9493 50263 9551 50269
rect 9582 50260 9588 50272
rect 9640 50260 9646 50312
rect 25498 50124 25504 50176
rect 25556 50124 25562 50176
rect 1104 50074 25852 50096
rect 1104 50022 7950 50074
rect 8002 50022 8014 50074
rect 8066 50022 8078 50074
rect 8130 50022 8142 50074
rect 8194 50022 8206 50074
rect 8258 50022 17950 50074
rect 18002 50022 18014 50074
rect 18066 50022 18078 50074
rect 18130 50022 18142 50074
rect 18194 50022 18206 50074
rect 18258 50022 25852 50074
rect 1104 50000 25852 50022
rect 24489 49827 24547 49833
rect 24489 49793 24501 49827
rect 24535 49824 24547 49827
rect 25498 49824 25504 49836
rect 24535 49796 25504 49824
rect 24535 49793 24547 49796
rect 24489 49787 24547 49793
rect 25498 49784 25504 49796
rect 25556 49784 25562 49836
rect 23658 49716 23664 49768
rect 23716 49756 23722 49768
rect 24765 49759 24823 49765
rect 24765 49756 24777 49759
rect 23716 49728 24777 49756
rect 23716 49716 23722 49728
rect 24765 49725 24777 49728
rect 24811 49725 24823 49759
rect 24765 49719 24823 49725
rect 1104 49530 25852 49552
rect 1104 49478 2950 49530
rect 3002 49478 3014 49530
rect 3066 49478 3078 49530
rect 3130 49478 3142 49530
rect 3194 49478 3206 49530
rect 3258 49478 12950 49530
rect 13002 49478 13014 49530
rect 13066 49478 13078 49530
rect 13130 49478 13142 49530
rect 13194 49478 13206 49530
rect 13258 49478 22950 49530
rect 23002 49478 23014 49530
rect 23066 49478 23078 49530
rect 23130 49478 23142 49530
rect 23194 49478 23206 49530
rect 23258 49478 25852 49530
rect 1104 49456 25852 49478
rect 10686 49308 10692 49360
rect 10744 49308 10750 49360
rect 11698 49308 11704 49360
rect 11756 49308 11762 49360
rect 10226 49104 10232 49156
rect 10284 49144 10290 49156
rect 10505 49147 10563 49153
rect 10505 49144 10517 49147
rect 10284 49116 10517 49144
rect 10284 49104 10290 49116
rect 10505 49113 10517 49116
rect 10551 49113 10563 49147
rect 10505 49107 10563 49113
rect 10870 49104 10876 49156
rect 10928 49144 10934 49156
rect 11517 49147 11575 49153
rect 11517 49144 11529 49147
rect 10928 49116 11529 49144
rect 10928 49104 10934 49116
rect 11517 49113 11529 49116
rect 11563 49113 11575 49147
rect 11517 49107 11575 49113
rect 24765 49147 24823 49153
rect 24765 49113 24777 49147
rect 24811 49144 24823 49147
rect 25130 49144 25136 49156
rect 24811 49116 25136 49144
rect 24811 49113 24823 49116
rect 24765 49107 24823 49113
rect 25130 49104 25136 49116
rect 25188 49104 25194 49156
rect 25222 49036 25228 49088
rect 25280 49036 25286 49088
rect 1104 48986 25852 49008
rect 1104 48934 7950 48986
rect 8002 48934 8014 48986
rect 8066 48934 8078 48986
rect 8130 48934 8142 48986
rect 8194 48934 8206 48986
rect 8258 48934 17950 48986
rect 18002 48934 18014 48986
rect 18066 48934 18078 48986
rect 18130 48934 18142 48986
rect 18194 48934 18206 48986
rect 18258 48934 25852 48986
rect 1104 48912 25852 48934
rect 8386 48832 8392 48884
rect 8444 48832 8450 48884
rect 8050 48708 9628 48736
rect 6641 48671 6699 48677
rect 6641 48637 6653 48671
rect 6687 48637 6699 48671
rect 6641 48631 6699 48637
rect 6917 48671 6975 48677
rect 6917 48637 6929 48671
rect 6963 48668 6975 48671
rect 9490 48668 9496 48680
rect 6963 48640 9496 48668
rect 6963 48637 6975 48640
rect 6917 48631 6975 48637
rect 6656 48532 6684 48631
rect 9490 48628 9496 48640
rect 9548 48628 9554 48680
rect 9122 48600 9128 48612
rect 8036 48572 9128 48600
rect 8036 48532 8064 48572
rect 9122 48560 9128 48572
rect 9180 48560 9186 48612
rect 6656 48504 8064 48532
rect 8757 48535 8815 48541
rect 8757 48501 8769 48535
rect 8803 48532 8815 48535
rect 9600 48532 9628 48708
rect 9950 48532 9956 48544
rect 8803 48504 9956 48532
rect 8803 48501 8815 48504
rect 8757 48495 8815 48501
rect 9950 48492 9956 48504
rect 10008 48492 10014 48544
rect 25130 48492 25136 48544
rect 25188 48532 25194 48544
rect 25409 48535 25467 48541
rect 25409 48532 25421 48535
rect 25188 48504 25421 48532
rect 25188 48492 25194 48504
rect 25409 48501 25421 48504
rect 25455 48501 25467 48535
rect 25409 48495 25467 48501
rect 1104 48442 25852 48464
rect 1104 48390 2950 48442
rect 3002 48390 3014 48442
rect 3066 48390 3078 48442
rect 3130 48390 3142 48442
rect 3194 48390 3206 48442
rect 3258 48390 12950 48442
rect 13002 48390 13014 48442
rect 13066 48390 13078 48442
rect 13130 48390 13142 48442
rect 13194 48390 13206 48442
rect 13258 48390 22950 48442
rect 23002 48390 23014 48442
rect 23066 48390 23078 48442
rect 23130 48390 23142 48442
rect 23194 48390 23206 48442
rect 23258 48390 25852 48442
rect 1104 48368 25852 48390
rect 7742 48084 7748 48136
rect 7800 48124 7806 48136
rect 10356 48127 10414 48133
rect 10356 48124 10368 48127
rect 7800 48096 10368 48124
rect 7800 48084 7806 48096
rect 10356 48093 10368 48096
rect 10402 48093 10414 48127
rect 10356 48087 10414 48093
rect 25130 48084 25136 48136
rect 25188 48084 25194 48136
rect 25317 48059 25375 48065
rect 25317 48025 25329 48059
rect 25363 48056 25375 48059
rect 26326 48056 26332 48068
rect 25363 48028 26332 48056
rect 25363 48025 25375 48028
rect 25317 48019 25375 48025
rect 26326 48016 26332 48028
rect 26384 48016 26390 48068
rect 10459 47991 10517 47997
rect 10459 47957 10471 47991
rect 10505 47988 10517 47991
rect 12618 47988 12624 48000
rect 10505 47960 12624 47988
rect 10505 47957 10517 47960
rect 10459 47951 10517 47957
rect 12618 47948 12624 47960
rect 12676 47948 12682 48000
rect 1104 47898 25852 47920
rect 1104 47846 7950 47898
rect 8002 47846 8014 47898
rect 8066 47846 8078 47898
rect 8130 47846 8142 47898
rect 8194 47846 8206 47898
rect 8258 47846 17950 47898
rect 18002 47846 18014 47898
rect 18066 47846 18078 47898
rect 18130 47846 18142 47898
rect 18194 47846 18206 47898
rect 18258 47846 25852 47898
rect 1104 47824 25852 47846
rect 9214 47744 9220 47796
rect 9272 47784 9278 47796
rect 9398 47784 9404 47796
rect 9272 47756 9404 47784
rect 9272 47744 9278 47756
rect 9398 47744 9404 47756
rect 9456 47784 9462 47796
rect 9861 47787 9919 47793
rect 9861 47784 9873 47787
rect 9456 47756 9873 47784
rect 9456 47744 9462 47756
rect 9861 47753 9873 47756
rect 9907 47753 9919 47787
rect 9861 47747 9919 47753
rect 8294 47608 8300 47660
rect 8352 47648 8358 47660
rect 9401 47651 9459 47657
rect 9401 47648 9413 47651
rect 8352 47620 9413 47648
rect 8352 47608 8358 47620
rect 9401 47617 9413 47620
rect 9447 47648 9459 47651
rect 10318 47648 10324 47660
rect 9447 47620 10324 47648
rect 9447 47617 9459 47620
rect 9401 47611 9459 47617
rect 10318 47608 10324 47620
rect 10376 47608 10382 47660
rect 24857 47651 24915 47657
rect 24857 47617 24869 47651
rect 24903 47648 24915 47651
rect 25314 47648 25320 47660
rect 24903 47620 25320 47648
rect 24903 47617 24915 47620
rect 24857 47611 24915 47617
rect 25314 47608 25320 47620
rect 25372 47608 25378 47660
rect 9490 47404 9496 47456
rect 9548 47404 9554 47456
rect 25133 47447 25191 47453
rect 25133 47413 25145 47447
rect 25179 47444 25191 47447
rect 26418 47444 26424 47456
rect 25179 47416 26424 47444
rect 25179 47413 25191 47416
rect 25133 47407 25191 47413
rect 26418 47404 26424 47416
rect 26476 47404 26482 47456
rect 1104 47354 25852 47376
rect 1104 47302 2950 47354
rect 3002 47302 3014 47354
rect 3066 47302 3078 47354
rect 3130 47302 3142 47354
rect 3194 47302 3206 47354
rect 3258 47302 12950 47354
rect 13002 47302 13014 47354
rect 13066 47302 13078 47354
rect 13130 47302 13142 47354
rect 13194 47302 13206 47354
rect 13258 47302 22950 47354
rect 23002 47302 23014 47354
rect 23066 47302 23078 47354
rect 23130 47302 23142 47354
rect 23194 47302 23206 47354
rect 23258 47302 25852 47354
rect 1104 47280 25852 47302
rect 9214 46996 9220 47048
rect 9272 47036 9278 47048
rect 11644 47039 11702 47045
rect 11644 47036 11656 47039
rect 9272 47008 11656 47036
rect 9272 46996 9278 47008
rect 11644 47005 11656 47008
rect 11690 47005 11702 47039
rect 11644 46999 11702 47005
rect 11747 46971 11805 46977
rect 11747 46937 11759 46971
rect 11793 46968 11805 46971
rect 13722 46968 13728 46980
rect 11793 46940 13728 46968
rect 11793 46937 11805 46940
rect 11747 46931 11805 46937
rect 13722 46928 13728 46940
rect 13780 46928 13786 46980
rect 25314 46860 25320 46912
rect 25372 46900 25378 46912
rect 25409 46903 25467 46909
rect 25409 46900 25421 46903
rect 25372 46872 25421 46900
rect 25372 46860 25378 46872
rect 25409 46869 25421 46872
rect 25455 46869 25467 46903
rect 25409 46863 25467 46869
rect 1104 46810 25852 46832
rect 1104 46758 7950 46810
rect 8002 46758 8014 46810
rect 8066 46758 8078 46810
rect 8130 46758 8142 46810
rect 8194 46758 8206 46810
rect 8258 46758 17950 46810
rect 18002 46758 18014 46810
rect 18066 46758 18078 46810
rect 18130 46758 18142 46810
rect 18194 46758 18206 46810
rect 18258 46758 25852 46810
rect 1104 46736 25852 46758
rect 9766 46656 9772 46708
rect 9824 46696 9830 46708
rect 10778 46696 10784 46708
rect 9824 46668 10784 46696
rect 9824 46656 9830 46668
rect 10778 46656 10784 46668
rect 10836 46656 10842 46708
rect 10318 46520 10324 46572
rect 10376 46520 10382 46572
rect 10796 46560 10824 46656
rect 13722 46588 13728 46640
rect 13780 46628 13786 46640
rect 14093 46631 14151 46637
rect 14093 46628 14105 46631
rect 13780 46600 14105 46628
rect 13780 46588 13786 46600
rect 14093 46597 14105 46600
rect 14139 46597 14151 46631
rect 14093 46591 14151 46597
rect 12564 46563 12622 46569
rect 12564 46560 12576 46563
rect 10796 46532 12576 46560
rect 12564 46529 12576 46532
rect 12610 46529 12622 46563
rect 12564 46523 12622 46529
rect 13906 46520 13912 46572
rect 13964 46520 13970 46572
rect 25314 46520 25320 46572
rect 25372 46520 25378 46572
rect 15746 46452 15752 46504
rect 15804 46452 15810 46504
rect 10410 46316 10416 46368
rect 10468 46316 10474 46368
rect 12667 46359 12725 46365
rect 12667 46325 12679 46359
rect 12713 46356 12725 46359
rect 15010 46356 15016 46368
rect 12713 46328 15016 46356
rect 12713 46325 12725 46328
rect 12667 46319 12725 46325
rect 15010 46316 15016 46328
rect 15068 46316 15074 46368
rect 25133 46359 25191 46365
rect 25133 46325 25145 46359
rect 25179 46356 25191 46359
rect 25406 46356 25412 46368
rect 25179 46328 25412 46356
rect 25179 46325 25191 46328
rect 25133 46319 25191 46325
rect 25406 46316 25412 46328
rect 25464 46316 25470 46368
rect 1104 46266 25852 46288
rect 1104 46214 2950 46266
rect 3002 46214 3014 46266
rect 3066 46214 3078 46266
rect 3130 46214 3142 46266
rect 3194 46214 3206 46266
rect 3258 46214 12950 46266
rect 13002 46214 13014 46266
rect 13066 46214 13078 46266
rect 13130 46214 13142 46266
rect 13194 46214 13206 46266
rect 13258 46214 22950 46266
rect 23002 46214 23014 46266
rect 23066 46214 23078 46266
rect 23130 46214 23142 46266
rect 23194 46214 23206 46266
rect 23258 46214 25852 46266
rect 1104 46192 25852 46214
rect 8478 46112 8484 46164
rect 8536 46112 8542 46164
rect 15654 46084 15660 46096
rect 14844 46056 15660 46084
rect 7742 45976 7748 46028
rect 7800 46016 7806 46028
rect 14844 46025 14872 46056
rect 15654 46044 15660 46056
rect 15712 46044 15718 46096
rect 8113 46019 8171 46025
rect 8113 46016 8125 46019
rect 7800 45988 8125 46016
rect 7800 45976 7806 45988
rect 8113 45985 8125 45988
rect 8159 45985 8171 46019
rect 8113 45979 8171 45985
rect 14829 46019 14887 46025
rect 14829 45985 14841 46019
rect 14875 45985 14887 46019
rect 14829 45979 14887 45985
rect 15010 45976 15016 46028
rect 15068 45976 15074 46028
rect 16482 45976 16488 46028
rect 16540 45976 16546 46028
rect 7834 45908 7840 45960
rect 7892 45948 7898 45960
rect 7929 45951 7987 45957
rect 7929 45948 7941 45951
rect 7892 45920 7941 45948
rect 7892 45908 7898 45920
rect 7929 45917 7941 45920
rect 7975 45917 7987 45951
rect 7929 45911 7987 45917
rect 12526 45908 12532 45960
rect 12584 45948 12590 45960
rect 13300 45951 13358 45957
rect 13300 45948 13312 45951
rect 12584 45920 13312 45948
rect 12584 45908 12590 45920
rect 13300 45917 13312 45920
rect 13346 45917 13358 45951
rect 13300 45911 13358 45917
rect 24857 45951 24915 45957
rect 24857 45917 24869 45951
rect 24903 45948 24915 45951
rect 25314 45948 25320 45960
rect 24903 45920 25320 45948
rect 24903 45917 24915 45920
rect 24857 45911 24915 45917
rect 25314 45908 25320 45920
rect 25372 45908 25378 45960
rect 13403 45815 13461 45821
rect 13403 45781 13415 45815
rect 13449 45812 13461 45815
rect 15102 45812 15108 45824
rect 13449 45784 15108 45812
rect 13449 45781 13461 45784
rect 13403 45775 13461 45781
rect 15102 45772 15108 45784
rect 15160 45772 15166 45824
rect 24854 45772 24860 45824
rect 24912 45812 24918 45824
rect 25133 45815 25191 45821
rect 25133 45812 25145 45815
rect 24912 45784 25145 45812
rect 24912 45772 24918 45784
rect 25133 45781 25145 45784
rect 25179 45781 25191 45815
rect 25133 45775 25191 45781
rect 1104 45722 25852 45744
rect 1104 45670 7950 45722
rect 8002 45670 8014 45722
rect 8066 45670 8078 45722
rect 8130 45670 8142 45722
rect 8194 45670 8206 45722
rect 8258 45670 17950 45722
rect 18002 45670 18014 45722
rect 18066 45670 18078 45722
rect 18130 45670 18142 45722
rect 18194 45670 18206 45722
rect 18258 45670 25852 45722
rect 1104 45648 25852 45670
rect 10502 45500 10508 45552
rect 10560 45540 10566 45552
rect 12526 45540 12532 45552
rect 10560 45512 12532 45540
rect 10560 45500 10566 45512
rect 12526 45500 12532 45512
rect 12584 45500 12590 45552
rect 12618 45500 12624 45552
rect 12676 45540 12682 45552
rect 12897 45543 12955 45549
rect 12897 45540 12909 45543
rect 12676 45512 12909 45540
rect 12676 45500 12682 45512
rect 12897 45509 12909 45512
rect 12943 45509 12955 45543
rect 12897 45503 12955 45509
rect 12710 45432 12716 45484
rect 12768 45432 12774 45484
rect 14550 45364 14556 45416
rect 14608 45364 14614 45416
rect 25314 45228 25320 45280
rect 25372 45268 25378 45280
rect 25409 45271 25467 45277
rect 25409 45268 25421 45271
rect 25372 45240 25421 45268
rect 25372 45228 25378 45240
rect 25409 45237 25421 45240
rect 25455 45237 25467 45271
rect 25409 45231 25467 45237
rect 1104 45178 25852 45200
rect 1104 45126 2950 45178
rect 3002 45126 3014 45178
rect 3066 45126 3078 45178
rect 3130 45126 3142 45178
rect 3194 45126 3206 45178
rect 3258 45126 12950 45178
rect 13002 45126 13014 45178
rect 13066 45126 13078 45178
rect 13130 45126 13142 45178
rect 13194 45126 13206 45178
rect 13258 45126 22950 45178
rect 23002 45126 23014 45178
rect 23066 45126 23078 45178
rect 23130 45126 23142 45178
rect 23194 45126 23206 45178
rect 23258 45126 25852 45178
rect 1104 45104 25852 45126
rect 9398 45024 9404 45076
rect 9456 45064 9462 45076
rect 10873 45067 10931 45073
rect 10873 45064 10885 45067
rect 9456 45036 10885 45064
rect 9456 45024 9462 45036
rect 10873 45033 10885 45036
rect 10919 45033 10931 45067
rect 10873 45027 10931 45033
rect 9122 44888 9128 44940
rect 9180 44928 9186 44940
rect 9398 44928 9404 44940
rect 9180 44900 9404 44928
rect 9180 44888 9186 44900
rect 9398 44888 9404 44900
rect 9456 44888 9462 44940
rect 9950 44888 9956 44940
rect 10008 44928 10014 44940
rect 15657 44931 15715 44937
rect 10008 44900 10640 44928
rect 10008 44888 10014 44900
rect 9401 44795 9459 44801
rect 9401 44761 9413 44795
rect 9447 44792 9459 44795
rect 9674 44792 9680 44804
rect 9447 44764 9680 44792
rect 9447 44761 9459 44764
rect 9401 44755 9459 44761
rect 9674 44752 9680 44764
rect 9732 44752 9738 44804
rect 10612 44792 10640 44900
rect 15657 44897 15669 44931
rect 15703 44928 15715 44931
rect 16114 44928 16120 44940
rect 15703 44900 16120 44928
rect 15703 44897 15715 44900
rect 15657 44891 15715 44897
rect 16114 44888 16120 44900
rect 16172 44888 16178 44940
rect 25314 44820 25320 44872
rect 25372 44820 25378 44872
rect 10612 44778 11284 44792
rect 10626 44764 11284 44778
rect 9692 44724 9720 44752
rect 10410 44724 10416 44736
rect 9692 44696 10416 44724
rect 10410 44684 10416 44696
rect 10468 44684 10474 44736
rect 11256 44733 11284 44764
rect 15102 44752 15108 44804
rect 15160 44792 15166 44804
rect 15841 44795 15899 44801
rect 15841 44792 15853 44795
rect 15160 44764 15853 44792
rect 15160 44752 15166 44764
rect 15841 44761 15853 44764
rect 15887 44761 15899 44795
rect 15841 44755 15899 44761
rect 17497 44795 17555 44801
rect 17497 44761 17509 44795
rect 17543 44792 17555 44795
rect 19978 44792 19984 44804
rect 17543 44764 19984 44792
rect 17543 44761 17555 44764
rect 17497 44755 17555 44761
rect 19978 44752 19984 44764
rect 20036 44752 20042 44804
rect 11241 44727 11299 44733
rect 11241 44693 11253 44727
rect 11287 44724 11299 44727
rect 11514 44724 11520 44736
rect 11287 44696 11520 44724
rect 11287 44693 11299 44696
rect 11241 44687 11299 44693
rect 11514 44684 11520 44696
rect 11572 44684 11578 44736
rect 25038 44684 25044 44736
rect 25096 44724 25102 44736
rect 25133 44727 25191 44733
rect 25133 44724 25145 44727
rect 25096 44696 25145 44724
rect 25096 44684 25102 44696
rect 25133 44693 25145 44696
rect 25179 44693 25191 44727
rect 25133 44687 25191 44693
rect 1104 44634 25852 44656
rect 1104 44582 7950 44634
rect 8002 44582 8014 44634
rect 8066 44582 8078 44634
rect 8130 44582 8142 44634
rect 8194 44582 8206 44634
rect 8258 44582 17950 44634
rect 18002 44582 18014 44634
rect 18066 44582 18078 44634
rect 18130 44582 18142 44634
rect 18194 44582 18206 44634
rect 18258 44582 25852 44634
rect 1104 44560 25852 44582
rect 9582 44480 9588 44532
rect 9640 44480 9646 44532
rect 9125 44387 9183 44393
rect 9125 44353 9137 44387
rect 9171 44384 9183 44387
rect 9214 44384 9220 44396
rect 9171 44356 9220 44384
rect 9171 44353 9183 44356
rect 9125 44347 9183 44353
rect 9214 44344 9220 44356
rect 9272 44344 9278 44396
rect 10318 44344 10324 44396
rect 10376 44384 10382 44396
rect 10597 44387 10655 44393
rect 10597 44384 10609 44387
rect 10376 44356 10609 44384
rect 10376 44344 10382 44356
rect 10597 44353 10609 44356
rect 10643 44353 10655 44387
rect 10597 44347 10655 44353
rect 24762 44344 24768 44396
rect 24820 44384 24826 44396
rect 25133 44387 25191 44393
rect 25133 44384 25145 44387
rect 24820 44356 25145 44384
rect 24820 44344 24826 44356
rect 25133 44353 25145 44356
rect 25179 44353 25191 44387
rect 25133 44347 25191 44353
rect 8941 44319 8999 44325
rect 8941 44285 8953 44319
rect 8987 44316 8999 44319
rect 9030 44316 9036 44328
rect 8987 44288 9036 44316
rect 8987 44285 8999 44288
rect 8941 44279 8999 44285
rect 9030 44276 9036 44288
rect 9088 44276 9094 44328
rect 10502 44208 10508 44260
rect 10560 44248 10566 44260
rect 25317 44251 25375 44257
rect 10560 44220 11008 44248
rect 10560 44208 10566 44220
rect 10980 44192 11008 44220
rect 25317 44217 25329 44251
rect 25363 44248 25375 44251
rect 25866 44248 25872 44260
rect 25363 44220 25872 44248
rect 25363 44217 25375 44220
rect 25317 44211 25375 44217
rect 25866 44208 25872 44220
rect 25924 44208 25930 44260
rect 10686 44140 10692 44192
rect 10744 44140 10750 44192
rect 10962 44140 10968 44192
rect 11020 44180 11026 44192
rect 11057 44183 11115 44189
rect 11057 44180 11069 44183
rect 11020 44152 11069 44180
rect 11020 44140 11026 44152
rect 11057 44149 11069 44152
rect 11103 44149 11115 44183
rect 11057 44143 11115 44149
rect 1104 44090 25852 44112
rect 1104 44038 2950 44090
rect 3002 44038 3014 44090
rect 3066 44038 3078 44090
rect 3130 44038 3142 44090
rect 3194 44038 3206 44090
rect 3258 44038 12950 44090
rect 13002 44038 13014 44090
rect 13066 44038 13078 44090
rect 13130 44038 13142 44090
rect 13194 44038 13206 44090
rect 13258 44038 22950 44090
rect 23002 44038 23014 44090
rect 23066 44038 23078 44090
rect 23130 44038 23142 44090
rect 23194 44038 23206 44090
rect 23258 44038 25852 44090
rect 1104 44016 25852 44038
rect 20612 43979 20670 43985
rect 20612 43945 20624 43979
rect 20658 43976 20670 43979
rect 24946 43976 24952 43988
rect 20658 43948 24952 43976
rect 20658 43945 20670 43948
rect 20612 43939 20670 43945
rect 24946 43936 24952 43948
rect 25004 43936 25010 43988
rect 21082 43800 21088 43852
rect 21140 43840 21146 43852
rect 22373 43843 22431 43849
rect 22373 43840 22385 43843
rect 21140 43812 22385 43840
rect 21140 43800 21146 43812
rect 22373 43809 22385 43812
rect 22419 43809 22431 43843
rect 22373 43803 22431 43809
rect 19518 43732 19524 43784
rect 19576 43772 19582 43784
rect 20349 43775 20407 43781
rect 20349 43772 20361 43775
rect 19576 43744 20361 43772
rect 19576 43732 19582 43744
rect 20349 43741 20361 43744
rect 20395 43741 20407 43775
rect 20349 43735 20407 43741
rect 21082 43664 21088 43716
rect 21140 43664 21146 43716
rect 22094 43596 22100 43648
rect 22152 43596 22158 43648
rect 25498 43596 25504 43648
rect 25556 43596 25562 43648
rect 1104 43546 25852 43568
rect 1104 43494 7950 43546
rect 8002 43494 8014 43546
rect 8066 43494 8078 43546
rect 8130 43494 8142 43546
rect 8194 43494 8206 43546
rect 8258 43494 17950 43546
rect 18002 43494 18014 43546
rect 18066 43494 18078 43546
rect 18130 43494 18142 43546
rect 18194 43494 18206 43546
rect 18258 43494 25852 43546
rect 1104 43472 25852 43494
rect 25133 43367 25191 43373
rect 25133 43333 25145 43367
rect 25179 43364 25191 43367
rect 25498 43364 25504 43376
rect 25179 43336 25504 43364
rect 25179 43333 25191 43336
rect 25133 43327 25191 43333
rect 25498 43324 25504 43336
rect 25556 43324 25562 43376
rect 25317 43163 25375 43169
rect 25317 43129 25329 43163
rect 25363 43160 25375 43163
rect 25958 43160 25964 43172
rect 25363 43132 25964 43160
rect 25363 43129 25375 43132
rect 25317 43123 25375 43129
rect 25958 43120 25964 43132
rect 26016 43120 26022 43172
rect 1104 43002 25852 43024
rect 1104 42950 2950 43002
rect 3002 42950 3014 43002
rect 3066 42950 3078 43002
rect 3130 42950 3142 43002
rect 3194 42950 3206 43002
rect 3258 42950 12950 43002
rect 13002 42950 13014 43002
rect 13066 42950 13078 43002
rect 13130 42950 13142 43002
rect 13194 42950 13206 43002
rect 13258 42950 22950 43002
rect 23002 42950 23014 43002
rect 23066 42950 23078 43002
rect 23130 42950 23142 43002
rect 23194 42950 23206 43002
rect 23258 42950 25852 43002
rect 1104 42928 25852 42950
rect 9766 42712 9772 42764
rect 9824 42712 9830 42764
rect 10226 42712 10232 42764
rect 10284 42712 10290 42764
rect 8938 42644 8944 42696
rect 8996 42684 9002 42696
rect 9585 42687 9643 42693
rect 9585 42684 9597 42687
rect 8996 42656 9597 42684
rect 8996 42644 9002 42656
rect 9585 42653 9597 42656
rect 9631 42653 9643 42687
rect 9585 42647 9643 42653
rect 24765 42619 24823 42625
rect 24765 42585 24777 42619
rect 24811 42616 24823 42619
rect 25130 42616 25136 42628
rect 24811 42588 25136 42616
rect 24811 42585 24823 42588
rect 24765 42579 24823 42585
rect 25130 42576 25136 42588
rect 25188 42576 25194 42628
rect 25317 42619 25375 42625
rect 25317 42585 25329 42619
rect 25363 42616 25375 42619
rect 25682 42616 25688 42628
rect 25363 42588 25688 42616
rect 25363 42585 25375 42588
rect 25317 42579 25375 42585
rect 25682 42576 25688 42588
rect 25740 42576 25746 42628
rect 1104 42458 25852 42480
rect 1104 42406 7950 42458
rect 8002 42406 8014 42458
rect 8066 42406 8078 42458
rect 8130 42406 8142 42458
rect 8194 42406 8206 42458
rect 8258 42406 17950 42458
rect 18002 42406 18014 42458
rect 18066 42406 18078 42458
rect 18130 42406 18142 42458
rect 18194 42406 18206 42458
rect 18258 42406 25852 42458
rect 1104 42384 25852 42406
rect 9674 42304 9680 42356
rect 9732 42344 9738 42356
rect 11149 42347 11207 42353
rect 11149 42344 11161 42347
rect 9732 42316 11161 42344
rect 9732 42304 9738 42316
rect 11149 42313 11161 42316
rect 11195 42313 11207 42347
rect 11149 42307 11207 42313
rect 11514 42276 11520 42288
rect 10902 42248 11520 42276
rect 11514 42236 11520 42248
rect 11572 42236 11578 42288
rect 9398 42100 9404 42152
rect 9456 42100 9462 42152
rect 9677 42143 9735 42149
rect 9677 42109 9689 42143
rect 9723 42140 9735 42143
rect 9766 42140 9772 42152
rect 9723 42112 9772 42140
rect 9723 42109 9735 42112
rect 9677 42103 9735 42109
rect 9766 42100 9772 42112
rect 9824 42140 9830 42152
rect 10686 42140 10692 42152
rect 9824 42112 10692 42140
rect 9824 42100 9830 42112
rect 10686 42100 10692 42112
rect 10744 42100 10750 42152
rect 11514 41964 11520 42016
rect 11572 41964 11578 42016
rect 25130 41964 25136 42016
rect 25188 42004 25194 42016
rect 25409 42007 25467 42013
rect 25409 42004 25421 42007
rect 25188 41976 25421 42004
rect 25188 41964 25194 41976
rect 25409 41973 25421 41976
rect 25455 41973 25467 42007
rect 25409 41967 25467 41973
rect 1104 41914 25852 41936
rect 1104 41862 2950 41914
rect 3002 41862 3014 41914
rect 3066 41862 3078 41914
rect 3130 41862 3142 41914
rect 3194 41862 3206 41914
rect 3258 41862 12950 41914
rect 13002 41862 13014 41914
rect 13066 41862 13078 41914
rect 13130 41862 13142 41914
rect 13194 41862 13206 41914
rect 13258 41862 22950 41914
rect 23002 41862 23014 41914
rect 23066 41862 23078 41914
rect 23130 41862 23142 41914
rect 23194 41862 23206 41914
rect 23258 41862 25852 41914
rect 1104 41840 25852 41862
rect 10870 41760 10876 41812
rect 10928 41760 10934 41812
rect 10413 41667 10471 41673
rect 10413 41633 10425 41667
rect 10459 41664 10471 41667
rect 10962 41664 10968 41676
rect 10459 41636 10968 41664
rect 10459 41633 10471 41636
rect 10413 41627 10471 41633
rect 10962 41624 10968 41636
rect 11020 41624 11026 41676
rect 9214 41556 9220 41608
rect 9272 41596 9278 41608
rect 10229 41599 10287 41605
rect 10229 41596 10241 41599
rect 9272 41568 10241 41596
rect 9272 41556 9278 41568
rect 10229 41565 10241 41568
rect 10275 41565 10287 41599
rect 10229 41559 10287 41565
rect 25130 41556 25136 41608
rect 25188 41556 25194 41608
rect 25317 41531 25375 41537
rect 25317 41497 25329 41531
rect 25363 41528 25375 41531
rect 26142 41528 26148 41540
rect 25363 41500 26148 41528
rect 25363 41497 25375 41500
rect 25317 41491 25375 41497
rect 26142 41488 26148 41500
rect 26200 41488 26206 41540
rect 1104 41370 25852 41392
rect 1104 41318 7950 41370
rect 8002 41318 8014 41370
rect 8066 41318 8078 41370
rect 8130 41318 8142 41370
rect 8194 41318 8206 41370
rect 8258 41318 17950 41370
rect 18002 41318 18014 41370
rect 18066 41318 18078 41370
rect 18130 41318 18142 41370
rect 18194 41318 18206 41370
rect 18258 41318 25852 41370
rect 1104 41296 25852 41318
rect 24857 41123 24915 41129
rect 24857 41089 24869 41123
rect 24903 41120 24915 41123
rect 25314 41120 25320 41132
rect 24903 41092 25320 41120
rect 24903 41089 24915 41092
rect 24857 41083 24915 41089
rect 25314 41080 25320 41092
rect 25372 41080 25378 41132
rect 25133 40919 25191 40925
rect 25133 40885 25145 40919
rect 25179 40916 25191 40919
rect 25590 40916 25596 40928
rect 25179 40888 25596 40916
rect 25179 40885 25191 40888
rect 25133 40879 25191 40885
rect 25590 40876 25596 40888
rect 25648 40876 25654 40928
rect 1104 40826 25852 40848
rect 1104 40774 2950 40826
rect 3002 40774 3014 40826
rect 3066 40774 3078 40826
rect 3130 40774 3142 40826
rect 3194 40774 3206 40826
rect 3258 40774 12950 40826
rect 13002 40774 13014 40826
rect 13066 40774 13078 40826
rect 13130 40774 13142 40826
rect 13194 40774 13206 40826
rect 13258 40774 22950 40826
rect 23002 40774 23014 40826
rect 23066 40774 23078 40826
rect 23130 40774 23142 40826
rect 23194 40774 23206 40826
rect 23258 40774 25852 40826
rect 1104 40752 25852 40774
rect 25498 40332 25504 40384
rect 25556 40332 25562 40384
rect 1104 40282 25852 40304
rect 1104 40230 7950 40282
rect 8002 40230 8014 40282
rect 8066 40230 8078 40282
rect 8130 40230 8142 40282
rect 8194 40230 8206 40282
rect 8258 40230 17950 40282
rect 18002 40230 18014 40282
rect 18066 40230 18078 40282
rect 18130 40230 18142 40282
rect 18194 40230 18206 40282
rect 18258 40230 25852 40282
rect 1104 40208 25852 40230
rect 23382 40128 23388 40180
rect 23440 40168 23446 40180
rect 25133 40171 25191 40177
rect 25133 40168 25145 40171
rect 23440 40140 25145 40168
rect 23440 40128 23446 40140
rect 25133 40137 25145 40140
rect 25179 40137 25191 40171
rect 25133 40131 25191 40137
rect 25498 40100 25504 40112
rect 25332 40072 25504 40100
rect 25332 40041 25360 40072
rect 25498 40060 25504 40072
rect 25556 40060 25562 40112
rect 25317 40035 25375 40041
rect 25317 40001 25329 40035
rect 25363 40001 25375 40035
rect 25317 39995 25375 40001
rect 1104 39738 25852 39760
rect 1104 39686 2950 39738
rect 3002 39686 3014 39738
rect 3066 39686 3078 39738
rect 3130 39686 3142 39738
rect 3194 39686 3206 39738
rect 3258 39686 12950 39738
rect 13002 39686 13014 39738
rect 13066 39686 13078 39738
rect 13130 39686 13142 39738
rect 13194 39686 13206 39738
rect 13258 39686 22950 39738
rect 23002 39686 23014 39738
rect 23066 39686 23078 39738
rect 23130 39686 23142 39738
rect 23194 39686 23206 39738
rect 23258 39686 25852 39738
rect 1104 39664 25852 39686
rect 24857 39423 24915 39429
rect 24857 39389 24869 39423
rect 24903 39420 24915 39423
rect 25314 39420 25320 39432
rect 24903 39392 25320 39420
rect 24903 39389 24915 39392
rect 24857 39383 24915 39389
rect 25314 39380 25320 39392
rect 25372 39380 25378 39432
rect 22066 39324 25176 39352
rect 21910 39244 21916 39296
rect 21968 39284 21974 39296
rect 22066 39284 22094 39324
rect 25148 39293 25176 39324
rect 21968 39256 22094 39284
rect 25133 39287 25191 39293
rect 21968 39244 21974 39256
rect 25133 39253 25145 39287
rect 25179 39253 25191 39287
rect 25133 39247 25191 39253
rect 1104 39194 25852 39216
rect 1104 39142 7950 39194
rect 8002 39142 8014 39194
rect 8066 39142 8078 39194
rect 8130 39142 8142 39194
rect 8194 39142 8206 39194
rect 8258 39142 17950 39194
rect 18002 39142 18014 39194
rect 18066 39142 18078 39194
rect 18130 39142 18142 39194
rect 18194 39142 18206 39194
rect 18258 39142 25852 39194
rect 1104 39120 25852 39142
rect 25314 38700 25320 38752
rect 25372 38740 25378 38752
rect 25409 38743 25467 38749
rect 25409 38740 25421 38743
rect 25372 38712 25421 38740
rect 25372 38700 25378 38712
rect 25409 38709 25421 38712
rect 25455 38709 25467 38743
rect 25409 38703 25467 38709
rect 1104 38650 25852 38672
rect 1104 38598 2950 38650
rect 3002 38598 3014 38650
rect 3066 38598 3078 38650
rect 3130 38598 3142 38650
rect 3194 38598 3206 38650
rect 3258 38598 12950 38650
rect 13002 38598 13014 38650
rect 13066 38598 13078 38650
rect 13130 38598 13142 38650
rect 13194 38598 13206 38650
rect 13258 38598 22950 38650
rect 23002 38598 23014 38650
rect 23066 38598 23078 38650
rect 23130 38598 23142 38650
rect 23194 38598 23206 38650
rect 23258 38598 25852 38650
rect 1104 38576 25852 38598
rect 25314 38292 25320 38344
rect 25372 38292 25378 38344
rect 25038 38156 25044 38208
rect 25096 38196 25102 38208
rect 25133 38199 25191 38205
rect 25133 38196 25145 38199
rect 25096 38168 25145 38196
rect 25096 38156 25102 38168
rect 25133 38165 25145 38168
rect 25179 38165 25191 38199
rect 25133 38159 25191 38165
rect 1104 38106 25852 38128
rect 1104 38054 7950 38106
rect 8002 38054 8014 38106
rect 8066 38054 8078 38106
rect 8130 38054 8142 38106
rect 8194 38054 8206 38106
rect 8258 38054 17950 38106
rect 18002 38054 18014 38106
rect 18066 38054 18078 38106
rect 18130 38054 18142 38106
rect 18194 38054 18206 38106
rect 18258 38054 25852 38106
rect 1104 38032 25852 38054
rect 7834 37952 7840 38004
rect 7892 37992 7898 38004
rect 8665 37995 8723 38001
rect 8665 37992 8677 37995
rect 7892 37964 8677 37992
rect 7892 37952 7898 37964
rect 8665 37961 8677 37964
rect 8711 37961 8723 37995
rect 8665 37955 8723 37961
rect 8846 37816 8852 37868
rect 8904 37816 8910 37868
rect 24765 37859 24823 37865
rect 24765 37825 24777 37859
rect 24811 37856 24823 37859
rect 25130 37856 25136 37868
rect 24811 37828 25136 37856
rect 24811 37825 24823 37828
rect 24765 37819 24823 37825
rect 25130 37816 25136 37828
rect 25188 37816 25194 37868
rect 25317 37723 25375 37729
rect 25317 37689 25329 37723
rect 25363 37720 25375 37723
rect 26050 37720 26056 37732
rect 25363 37692 26056 37720
rect 25363 37689 25375 37692
rect 25317 37683 25375 37689
rect 26050 37680 26056 37692
rect 26108 37680 26114 37732
rect 1104 37562 25852 37584
rect 1104 37510 2950 37562
rect 3002 37510 3014 37562
rect 3066 37510 3078 37562
rect 3130 37510 3142 37562
rect 3194 37510 3206 37562
rect 3258 37510 12950 37562
rect 13002 37510 13014 37562
rect 13066 37510 13078 37562
rect 13130 37510 13142 37562
rect 13194 37510 13206 37562
rect 13258 37510 22950 37562
rect 23002 37510 23014 37562
rect 23066 37510 23078 37562
rect 23130 37510 23142 37562
rect 23194 37510 23206 37562
rect 23258 37510 25852 37562
rect 1104 37488 25852 37510
rect 25498 37068 25504 37120
rect 25556 37068 25562 37120
rect 1104 37018 25852 37040
rect 1104 36966 7950 37018
rect 8002 36966 8014 37018
rect 8066 36966 8078 37018
rect 8130 36966 8142 37018
rect 8194 36966 8206 37018
rect 8258 36966 17950 37018
rect 18002 36966 18014 37018
rect 18066 36966 18078 37018
rect 18130 36966 18142 37018
rect 18194 36966 18206 37018
rect 18258 36966 25852 37018
rect 1104 36944 25852 36966
rect 25133 36839 25191 36845
rect 25133 36805 25145 36839
rect 25179 36836 25191 36839
rect 25498 36836 25504 36848
rect 25179 36808 25504 36836
rect 25179 36805 25191 36808
rect 25133 36799 25191 36805
rect 25498 36796 25504 36808
rect 25556 36796 25562 36848
rect 25317 36635 25375 36641
rect 25317 36601 25329 36635
rect 25363 36632 25375 36635
rect 26694 36632 26700 36644
rect 25363 36604 26700 36632
rect 25363 36601 25375 36604
rect 25317 36595 25375 36601
rect 26694 36592 26700 36604
rect 26752 36592 26758 36644
rect 1104 36474 25852 36496
rect 1104 36422 2950 36474
rect 3002 36422 3014 36474
rect 3066 36422 3078 36474
rect 3130 36422 3142 36474
rect 3194 36422 3206 36474
rect 3258 36422 12950 36474
rect 13002 36422 13014 36474
rect 13066 36422 13078 36474
rect 13130 36422 13142 36474
rect 13194 36422 13206 36474
rect 13258 36422 22950 36474
rect 23002 36422 23014 36474
rect 23066 36422 23078 36474
rect 23130 36422 23142 36474
rect 23194 36422 23206 36474
rect 23258 36422 25852 36474
rect 1104 36400 25852 36422
rect 24857 36159 24915 36165
rect 24857 36125 24869 36159
rect 24903 36156 24915 36159
rect 25314 36156 25320 36168
rect 24903 36128 25320 36156
rect 24903 36125 24915 36128
rect 24857 36119 24915 36125
rect 25314 36116 25320 36128
rect 25372 36116 25378 36168
rect 25133 36023 25191 36029
rect 25133 35989 25145 36023
rect 25179 36020 25191 36023
rect 26602 36020 26608 36032
rect 25179 35992 26608 36020
rect 25179 35989 25191 35992
rect 25133 35983 25191 35989
rect 26602 35980 26608 35992
rect 26660 35980 26666 36032
rect 1104 35930 25852 35952
rect 1104 35878 7950 35930
rect 8002 35878 8014 35930
rect 8066 35878 8078 35930
rect 8130 35878 8142 35930
rect 8194 35878 8206 35930
rect 8258 35878 17950 35930
rect 18002 35878 18014 35930
rect 18066 35878 18078 35930
rect 18130 35878 18142 35930
rect 18194 35878 18206 35930
rect 18258 35878 25852 35930
rect 1104 35856 25852 35878
rect 9766 35776 9772 35828
rect 9824 35816 9830 35828
rect 11149 35819 11207 35825
rect 11149 35816 11161 35819
rect 9824 35788 11161 35816
rect 9824 35776 9830 35788
rect 11149 35785 11161 35788
rect 11195 35785 11207 35819
rect 11149 35779 11207 35785
rect 11514 35776 11520 35828
rect 11572 35776 11578 35828
rect 22465 35819 22523 35825
rect 22465 35785 22477 35819
rect 22511 35816 22523 35819
rect 24854 35816 24860 35828
rect 22511 35788 24860 35816
rect 22511 35785 22523 35788
rect 22465 35779 22523 35785
rect 24854 35776 24860 35788
rect 24912 35776 24918 35828
rect 11532 35748 11560 35776
rect 12710 35748 12716 35760
rect 10902 35720 12716 35748
rect 12710 35708 12716 35720
rect 12768 35708 12774 35760
rect 21177 35751 21235 35757
rect 21177 35717 21189 35751
rect 21223 35748 21235 35751
rect 25406 35748 25412 35760
rect 21223 35720 25412 35748
rect 21223 35717 21235 35720
rect 21177 35711 21235 35717
rect 25406 35708 25412 35720
rect 25464 35708 25470 35760
rect 21085 35683 21143 35689
rect 21085 35649 21097 35683
rect 21131 35649 21143 35683
rect 21085 35643 21143 35649
rect 9398 35572 9404 35624
rect 9456 35572 9462 35624
rect 9674 35572 9680 35624
rect 9732 35572 9738 35624
rect 19334 35504 19340 35556
rect 19392 35544 19398 35556
rect 20717 35547 20775 35553
rect 20717 35544 20729 35547
rect 19392 35516 20729 35544
rect 19392 35504 19398 35516
rect 20717 35513 20729 35516
rect 20763 35513 20775 35547
rect 20717 35507 20775 35513
rect 21100 35544 21128 35643
rect 21818 35640 21824 35692
rect 21876 35680 21882 35692
rect 22373 35683 22431 35689
rect 22373 35680 22385 35683
rect 21876 35652 22385 35680
rect 21876 35640 21882 35652
rect 22373 35649 22385 35652
rect 22419 35649 22431 35683
rect 22373 35643 22431 35649
rect 21266 35572 21272 35624
rect 21324 35572 21330 35624
rect 22462 35572 22468 35624
rect 22520 35612 22526 35624
rect 22557 35615 22615 35621
rect 22557 35612 22569 35615
rect 22520 35584 22569 35612
rect 22520 35572 22526 35584
rect 22557 35581 22569 35584
rect 22603 35581 22615 35615
rect 22557 35575 22615 35581
rect 22370 35544 22376 35556
rect 21100 35516 22376 35544
rect 15746 35436 15752 35488
rect 15804 35476 15810 35488
rect 20349 35479 20407 35485
rect 20349 35476 20361 35479
rect 15804 35448 20361 35476
rect 15804 35436 15810 35448
rect 20349 35445 20361 35448
rect 20395 35476 20407 35479
rect 21100 35476 21128 35516
rect 22370 35504 22376 35516
rect 22428 35504 22434 35556
rect 20395 35448 21128 35476
rect 20395 35445 20407 35448
rect 20349 35439 20407 35445
rect 22002 35436 22008 35488
rect 22060 35436 22066 35488
rect 25314 35436 25320 35488
rect 25372 35476 25378 35488
rect 25409 35479 25467 35485
rect 25409 35476 25421 35479
rect 25372 35448 25421 35476
rect 25372 35436 25378 35448
rect 25409 35445 25421 35448
rect 25455 35445 25467 35479
rect 25409 35439 25467 35445
rect 1104 35386 25852 35408
rect 1104 35334 2950 35386
rect 3002 35334 3014 35386
rect 3066 35334 3078 35386
rect 3130 35334 3142 35386
rect 3194 35334 3206 35386
rect 3258 35334 12950 35386
rect 13002 35334 13014 35386
rect 13066 35334 13078 35386
rect 13130 35334 13142 35386
rect 13194 35334 13206 35386
rect 13258 35334 22950 35386
rect 23002 35334 23014 35386
rect 23066 35334 23078 35386
rect 23130 35334 23142 35386
rect 23194 35334 23206 35386
rect 23258 35334 25852 35386
rect 1104 35312 25852 35334
rect 23290 35096 23296 35148
rect 23348 35096 23354 35148
rect 23201 35071 23259 35077
rect 23201 35037 23213 35071
rect 23247 35068 23259 35071
rect 24946 35068 24952 35080
rect 23247 35040 24952 35068
rect 23247 35037 23259 35040
rect 23201 35031 23259 35037
rect 24946 35028 24952 35040
rect 25004 35028 25010 35080
rect 25314 35028 25320 35080
rect 25372 35028 25378 35080
rect 19978 34960 19984 35012
rect 20036 35000 20042 35012
rect 20622 35000 20628 35012
rect 20036 34972 20628 35000
rect 20036 34960 20042 34972
rect 20622 34960 20628 34972
rect 20680 35000 20686 35012
rect 22465 35003 22523 35009
rect 22465 35000 22477 35003
rect 20680 34972 22477 35000
rect 20680 34960 20686 34972
rect 22465 34969 22477 34972
rect 22511 35000 22523 35003
rect 23109 35003 23167 35009
rect 23109 35000 23121 35003
rect 22511 34972 23121 35000
rect 22511 34969 22523 34972
rect 22465 34963 22523 34969
rect 23109 34969 23121 34972
rect 23155 34969 23167 35003
rect 23109 34963 23167 34969
rect 16482 34892 16488 34944
rect 16540 34932 16546 34944
rect 21818 34932 21824 34944
rect 16540 34904 21824 34932
rect 16540 34892 16546 34904
rect 21818 34892 21824 34904
rect 21876 34892 21882 34944
rect 22554 34892 22560 34944
rect 22612 34932 22618 34944
rect 22741 34935 22799 34941
rect 22741 34932 22753 34935
rect 22612 34904 22753 34932
rect 22612 34892 22618 34904
rect 22741 34901 22753 34904
rect 22787 34901 22799 34935
rect 22741 34895 22799 34901
rect 25133 34935 25191 34941
rect 25133 34901 25145 34935
rect 25179 34932 25191 34935
rect 25774 34932 25780 34944
rect 25179 34904 25780 34932
rect 25179 34901 25191 34904
rect 25133 34895 25191 34901
rect 25774 34892 25780 34904
rect 25832 34892 25838 34944
rect 1104 34842 25852 34864
rect 1104 34790 7950 34842
rect 8002 34790 8014 34842
rect 8066 34790 8078 34842
rect 8130 34790 8142 34842
rect 8194 34790 8206 34842
rect 8258 34790 17950 34842
rect 18002 34790 18014 34842
rect 18066 34790 18078 34842
rect 18130 34790 18142 34842
rect 18194 34790 18206 34842
rect 18258 34790 25852 34842
rect 1104 34768 25852 34790
rect 20714 34688 20720 34740
rect 20772 34728 20778 34740
rect 25133 34731 25191 34737
rect 25133 34728 25145 34731
rect 20772 34700 25145 34728
rect 20772 34688 20778 34700
rect 25133 34697 25145 34700
rect 25179 34697 25191 34731
rect 25133 34691 25191 34697
rect 24857 34595 24915 34601
rect 24857 34561 24869 34595
rect 24903 34592 24915 34595
rect 25314 34592 25320 34604
rect 24903 34564 25320 34592
rect 24903 34561 24915 34564
rect 24857 34555 24915 34561
rect 25314 34552 25320 34564
rect 25372 34552 25378 34604
rect 20438 34416 20444 34468
rect 20496 34456 20502 34468
rect 23934 34456 23940 34468
rect 20496 34428 23940 34456
rect 20496 34416 20502 34428
rect 23934 34416 23940 34428
rect 23992 34416 23998 34468
rect 21082 34348 21088 34400
rect 21140 34388 21146 34400
rect 21358 34388 21364 34400
rect 21140 34360 21364 34388
rect 21140 34348 21146 34360
rect 21358 34348 21364 34360
rect 21416 34348 21422 34400
rect 1104 34298 25852 34320
rect 1104 34246 2950 34298
rect 3002 34246 3014 34298
rect 3066 34246 3078 34298
rect 3130 34246 3142 34298
rect 3194 34246 3206 34298
rect 3258 34246 12950 34298
rect 13002 34246 13014 34298
rect 13066 34246 13078 34298
rect 13130 34246 13142 34298
rect 13194 34246 13206 34298
rect 13258 34246 22950 34298
rect 23002 34246 23014 34298
rect 23066 34246 23078 34298
rect 23130 34246 23142 34298
rect 23194 34246 23206 34298
rect 23258 34246 25852 34298
rect 1104 34224 25852 34246
rect 9030 34144 9036 34196
rect 9088 34184 9094 34196
rect 9125 34187 9183 34193
rect 9125 34184 9137 34187
rect 9088 34156 9137 34184
rect 9088 34144 9094 34156
rect 9125 34153 9137 34156
rect 9171 34153 9183 34187
rect 9125 34147 9183 34153
rect 21358 34144 21364 34196
rect 21416 34184 21422 34196
rect 21416 34156 22968 34184
rect 21416 34144 21422 34156
rect 9398 34008 9404 34060
rect 9456 34048 9462 34060
rect 15381 34051 15439 34057
rect 15381 34048 15393 34051
rect 9456 34020 15393 34048
rect 9456 34008 9462 34020
rect 15381 34017 15393 34020
rect 15427 34017 15439 34051
rect 15381 34011 15439 34017
rect 19702 34008 19708 34060
rect 19760 34048 19766 34060
rect 21637 34051 21695 34057
rect 21637 34048 21649 34051
rect 19760 34020 21649 34048
rect 19760 34008 19766 34020
rect 21637 34017 21649 34020
rect 21683 34048 21695 34051
rect 22278 34048 22284 34060
rect 21683 34020 22284 34048
rect 21683 34017 21695 34020
rect 21637 34011 21695 34017
rect 22278 34008 22284 34020
rect 22336 34008 22342 34060
rect 9306 33940 9312 33992
rect 9364 33940 9370 33992
rect 19426 33940 19432 33992
rect 19484 33940 19490 33992
rect 22940 33980 22968 34156
rect 23566 33980 23572 33992
rect 22940 33952 23572 33980
rect 23566 33940 23572 33952
rect 23624 33980 23630 33992
rect 23661 33983 23719 33989
rect 23661 33980 23673 33983
rect 23624 33952 23673 33980
rect 23624 33940 23630 33952
rect 23661 33949 23673 33952
rect 23707 33949 23719 33983
rect 23661 33943 23719 33949
rect 24857 33983 24915 33989
rect 24857 33949 24869 33983
rect 24903 33980 24915 33983
rect 25314 33980 25320 33992
rect 24903 33952 25320 33980
rect 24903 33949 24915 33952
rect 24857 33943 24915 33949
rect 25314 33940 25320 33952
rect 25372 33940 25378 33992
rect 14645 33915 14703 33921
rect 14645 33881 14657 33915
rect 14691 33912 14703 33915
rect 15378 33912 15384 33924
rect 14691 33884 15384 33912
rect 14691 33881 14703 33884
rect 14645 33875 14703 33881
rect 15378 33872 15384 33884
rect 15436 33912 15442 33924
rect 15841 33915 15899 33921
rect 15841 33912 15853 33915
rect 15436 33884 15853 33912
rect 15436 33872 15442 33884
rect 15841 33881 15853 33884
rect 15887 33881 15899 33915
rect 15841 33875 15899 33881
rect 19705 33915 19763 33921
rect 19705 33881 19717 33915
rect 19751 33912 19763 33915
rect 19794 33912 19800 33924
rect 19751 33884 19800 33912
rect 19751 33881 19763 33884
rect 19705 33875 19763 33881
rect 19794 33872 19800 33884
rect 19852 33872 19858 33924
rect 21913 33915 21971 33921
rect 20930 33884 21312 33912
rect 21284 33856 21312 33884
rect 21913 33881 21925 33915
rect 21959 33912 21971 33915
rect 21959 33884 22094 33912
rect 21959 33881 21971 33884
rect 21913 33875 21971 33881
rect 21174 33804 21180 33856
rect 21232 33804 21238 33856
rect 21266 33804 21272 33856
rect 21324 33804 21330 33856
rect 22066 33844 22094 33884
rect 22922 33844 22928 33856
rect 22066 33816 22928 33844
rect 22922 33804 22928 33816
rect 22980 33804 22986 33856
rect 23198 33804 23204 33856
rect 23256 33844 23262 33856
rect 23385 33847 23443 33853
rect 23385 33844 23397 33847
rect 23256 33816 23397 33844
rect 23256 33804 23262 33816
rect 23385 33813 23397 33816
rect 23431 33813 23443 33847
rect 23385 33807 23443 33813
rect 25133 33847 25191 33853
rect 25133 33813 25145 33847
rect 25179 33844 25191 33847
rect 26234 33844 26240 33856
rect 25179 33816 26240 33844
rect 25179 33813 25191 33816
rect 25133 33807 25191 33813
rect 26234 33804 26240 33816
rect 26292 33804 26298 33856
rect 1104 33754 25852 33776
rect 1104 33702 7950 33754
rect 8002 33702 8014 33754
rect 8066 33702 8078 33754
rect 8130 33702 8142 33754
rect 8194 33702 8206 33754
rect 8258 33702 17950 33754
rect 18002 33702 18014 33754
rect 18066 33702 18078 33754
rect 18130 33702 18142 33754
rect 18194 33702 18206 33754
rect 18258 33702 25852 33754
rect 1104 33680 25852 33702
rect 22462 33640 22468 33652
rect 19812 33612 22468 33640
rect 19812 33581 19840 33612
rect 22462 33600 22468 33612
rect 22520 33640 22526 33652
rect 23198 33640 23204 33652
rect 22520 33612 23204 33640
rect 22520 33600 22526 33612
rect 23198 33600 23204 33612
rect 23256 33600 23262 33652
rect 19797 33575 19855 33581
rect 19797 33541 19809 33575
rect 19843 33541 19855 33575
rect 21266 33572 21272 33584
rect 21022 33544 21272 33572
rect 19797 33535 19855 33541
rect 21266 33532 21272 33544
rect 21324 33532 21330 33584
rect 22278 33572 22284 33584
rect 22020 33544 22284 33572
rect 19518 33464 19524 33516
rect 19576 33464 19582 33516
rect 22020 33513 22048 33544
rect 22278 33532 22284 33544
rect 22336 33532 22342 33584
rect 23566 33572 23572 33584
rect 23506 33544 23572 33572
rect 23566 33532 23572 33544
rect 23624 33572 23630 33584
rect 24121 33575 24179 33581
rect 24121 33572 24133 33575
rect 23624 33544 24133 33572
rect 23624 33532 23630 33544
rect 24121 33541 24133 33544
rect 24167 33572 24179 33575
rect 24305 33575 24363 33581
rect 24305 33572 24317 33575
rect 24167 33544 24317 33572
rect 24167 33541 24179 33544
rect 24121 33535 24179 33541
rect 24305 33541 24317 33544
rect 24351 33541 24363 33575
rect 24305 33535 24363 33541
rect 22005 33507 22063 33513
rect 22005 33473 22017 33507
rect 22051 33473 22063 33507
rect 22005 33467 22063 33473
rect 24857 33507 24915 33513
rect 24857 33473 24869 33507
rect 24903 33504 24915 33507
rect 25317 33507 25375 33513
rect 25317 33504 25329 33507
rect 24903 33476 25329 33504
rect 24903 33473 24915 33476
rect 24857 33467 24915 33473
rect 25317 33473 25329 33476
rect 25363 33504 25375 33507
rect 25498 33504 25504 33516
rect 25363 33476 25504 33504
rect 25363 33473 25375 33476
rect 25317 33467 25375 33473
rect 25498 33464 25504 33476
rect 25556 33464 25562 33516
rect 19794 33396 19800 33448
rect 19852 33436 19858 33448
rect 20530 33436 20536 33448
rect 19852 33408 20536 33436
rect 19852 33396 19858 33408
rect 20530 33396 20536 33408
rect 20588 33436 20594 33448
rect 21269 33439 21327 33445
rect 21269 33436 21281 33439
rect 20588 33408 21281 33436
rect 20588 33396 20594 33408
rect 21269 33405 21281 33408
rect 21315 33405 21327 33439
rect 21269 33399 21327 33405
rect 22281 33439 22339 33445
rect 22281 33405 22293 33439
rect 22327 33436 22339 33439
rect 22370 33436 22376 33448
rect 22327 33408 22376 33436
rect 22327 33405 22339 33408
rect 22281 33399 22339 33405
rect 22370 33396 22376 33408
rect 22428 33396 22434 33448
rect 22738 33396 22744 33448
rect 22796 33436 22802 33448
rect 22922 33436 22928 33448
rect 22796 33408 22928 33436
rect 22796 33396 22802 33408
rect 22922 33396 22928 33408
rect 22980 33436 22986 33448
rect 23753 33439 23811 33445
rect 23753 33436 23765 33439
rect 22980 33408 23765 33436
rect 22980 33396 22986 33408
rect 23753 33405 23765 33408
rect 23799 33405 23811 33439
rect 23753 33399 23811 33405
rect 21266 33260 21272 33312
rect 21324 33300 21330 33312
rect 21545 33303 21603 33309
rect 21545 33300 21557 33303
rect 21324 33272 21557 33300
rect 21324 33260 21330 33272
rect 21545 33269 21557 33272
rect 21591 33269 21603 33303
rect 21545 33263 21603 33269
rect 24578 33260 24584 33312
rect 24636 33260 24642 33312
rect 25133 33303 25191 33309
rect 25133 33269 25145 33303
rect 25179 33300 25191 33303
rect 25406 33300 25412 33312
rect 25179 33272 25412 33300
rect 25179 33269 25191 33272
rect 25133 33263 25191 33269
rect 25406 33260 25412 33272
rect 25464 33260 25470 33312
rect 1104 33210 25852 33232
rect 1104 33158 2950 33210
rect 3002 33158 3014 33210
rect 3066 33158 3078 33210
rect 3130 33158 3142 33210
rect 3194 33158 3206 33210
rect 3258 33158 12950 33210
rect 13002 33158 13014 33210
rect 13066 33158 13078 33210
rect 13130 33158 13142 33210
rect 13194 33158 13206 33210
rect 13258 33158 22950 33210
rect 23002 33158 23014 33210
rect 23066 33158 23078 33210
rect 23130 33158 23142 33210
rect 23194 33158 23206 33210
rect 23258 33158 25852 33210
rect 1104 33136 25852 33158
rect 16574 33096 16580 33108
rect 16040 33068 16580 33096
rect 16040 32969 16068 33068
rect 16574 33056 16580 33068
rect 16632 33096 16638 33108
rect 17310 33096 17316 33108
rect 16632 33068 17316 33096
rect 16632 33056 16638 33068
rect 17310 33056 17316 33068
rect 17368 33056 17374 33108
rect 22370 33056 22376 33108
rect 22428 33096 22434 33108
rect 23290 33096 23296 33108
rect 22428 33068 23296 33096
rect 22428 33056 22434 33068
rect 23290 33056 23296 33068
rect 23348 33096 23354 33108
rect 24029 33099 24087 33105
rect 24029 33096 24041 33099
rect 23348 33068 24041 33096
rect 23348 33056 23354 33068
rect 24029 33065 24041 33068
rect 24075 33065 24087 33099
rect 24029 33059 24087 33065
rect 16850 32988 16856 33040
rect 16908 33028 16914 33040
rect 17126 33028 17132 33040
rect 16908 33000 17132 33028
rect 16908 32988 16914 33000
rect 17126 32988 17132 33000
rect 17184 33028 17190 33040
rect 17184 33000 22232 33028
rect 17184 32988 17190 33000
rect 16025 32963 16083 32969
rect 16025 32929 16037 32963
rect 16071 32929 16083 32963
rect 16025 32923 16083 32929
rect 16114 32920 16120 32972
rect 16172 32960 16178 32972
rect 22094 32960 22100 32972
rect 16172 32932 22100 32960
rect 16172 32920 16178 32932
rect 22094 32920 22100 32932
rect 22152 32920 22158 32972
rect 19426 32852 19432 32904
rect 19484 32892 19490 32904
rect 20625 32895 20683 32901
rect 20625 32892 20637 32895
rect 19484 32864 20637 32892
rect 19484 32852 19490 32864
rect 20625 32861 20637 32864
rect 20671 32861 20683 32895
rect 20625 32855 20683 32861
rect 15933 32827 15991 32833
rect 15933 32793 15945 32827
rect 15979 32824 15991 32827
rect 19889 32827 19947 32833
rect 15979 32796 16574 32824
rect 15979 32793 15991 32796
rect 15933 32787 15991 32793
rect 12618 32716 12624 32768
rect 12676 32756 12682 32768
rect 15565 32759 15623 32765
rect 15565 32756 15577 32759
rect 12676 32728 15577 32756
rect 12676 32716 12682 32728
rect 15565 32725 15577 32728
rect 15611 32725 15623 32759
rect 16546 32756 16574 32796
rect 19889 32793 19901 32827
rect 19935 32824 19947 32827
rect 22204 32824 22232 33000
rect 24946 32988 24952 33040
rect 25004 33028 25010 33040
rect 25004 33000 25176 33028
rect 25004 32988 25010 33000
rect 22278 32920 22284 32972
rect 22336 32920 22342 32972
rect 25148 32969 25176 33000
rect 22557 32963 22615 32969
rect 22557 32929 22569 32963
rect 22603 32960 22615 32963
rect 25133 32963 25191 32969
rect 22603 32932 24256 32960
rect 22603 32929 22615 32932
rect 22557 32923 22615 32929
rect 19935 32796 19969 32824
rect 22204 32796 22968 32824
rect 19935 32793 19947 32796
rect 19889 32787 19947 32793
rect 16850 32756 16856 32768
rect 16546 32728 16856 32756
rect 15565 32719 15623 32725
rect 16850 32716 16856 32728
rect 16908 32716 16914 32768
rect 19610 32716 19616 32768
rect 19668 32756 19674 32768
rect 19904 32756 19932 32787
rect 21818 32756 21824 32768
rect 19668 32728 21824 32756
rect 19668 32716 19674 32728
rect 21818 32716 21824 32728
rect 21876 32716 21882 32768
rect 22370 32716 22376 32768
rect 22428 32756 22434 32768
rect 22830 32756 22836 32768
rect 22428 32728 22836 32756
rect 22428 32716 22434 32728
rect 22830 32716 22836 32728
rect 22888 32716 22894 32768
rect 22940 32756 22968 32796
rect 23566 32784 23572 32836
rect 23624 32784 23630 32836
rect 24228 32824 24256 32932
rect 25133 32929 25145 32963
rect 25179 32929 25191 32963
rect 25133 32923 25191 32929
rect 24578 32852 24584 32904
rect 24636 32892 24642 32904
rect 24762 32892 24768 32904
rect 24636 32864 24768 32892
rect 24636 32852 24642 32864
rect 24762 32852 24768 32864
rect 24820 32892 24826 32904
rect 24949 32895 25007 32901
rect 24949 32892 24961 32895
rect 24820 32864 24961 32892
rect 24820 32852 24826 32864
rect 24949 32861 24961 32864
rect 24995 32861 25007 32895
rect 24949 32855 25007 32861
rect 25041 32895 25099 32901
rect 25041 32861 25053 32895
rect 25087 32892 25099 32895
rect 25590 32892 25596 32904
rect 25087 32864 25596 32892
rect 25087 32861 25099 32864
rect 25041 32855 25099 32861
rect 25590 32852 25596 32864
rect 25648 32852 25654 32904
rect 24228 32796 25084 32824
rect 25056 32768 25084 32796
rect 24486 32756 24492 32768
rect 22940 32728 24492 32756
rect 24486 32716 24492 32728
rect 24544 32716 24550 32768
rect 24578 32716 24584 32768
rect 24636 32716 24642 32768
rect 25038 32716 25044 32768
rect 25096 32716 25102 32768
rect 1104 32666 25852 32688
rect 1104 32614 7950 32666
rect 8002 32614 8014 32666
rect 8066 32614 8078 32666
rect 8130 32614 8142 32666
rect 8194 32614 8206 32666
rect 8258 32614 17950 32666
rect 18002 32614 18014 32666
rect 18066 32614 18078 32666
rect 18130 32614 18142 32666
rect 18194 32614 18206 32666
rect 18258 32614 25852 32666
rect 1104 32592 25852 32614
rect 16761 32555 16819 32561
rect 16761 32552 16773 32555
rect 16546 32524 16773 32552
rect 15378 32444 15384 32496
rect 15436 32484 15442 32496
rect 16546 32484 16574 32524
rect 16761 32521 16773 32524
rect 16807 32552 16819 32555
rect 19610 32552 19616 32564
rect 16807 32524 19616 32552
rect 16807 32521 16819 32524
rect 16761 32515 16819 32521
rect 19610 32512 19616 32524
rect 19668 32512 19674 32564
rect 21085 32555 21143 32561
rect 21085 32552 21097 32555
rect 19720 32524 21097 32552
rect 15436 32456 16574 32484
rect 19720 32484 19748 32524
rect 21085 32521 21097 32524
rect 21131 32552 21143 32555
rect 21266 32552 21272 32564
rect 21131 32524 21272 32552
rect 21131 32521 21143 32524
rect 21085 32515 21143 32521
rect 21266 32512 21272 32524
rect 21324 32512 21330 32564
rect 23566 32512 23572 32564
rect 23624 32512 23630 32564
rect 25038 32512 25044 32564
rect 25096 32552 25102 32564
rect 25225 32555 25283 32561
rect 25225 32552 25237 32555
rect 25096 32524 25237 32552
rect 25096 32512 25102 32524
rect 25225 32521 25237 32524
rect 25271 32521 25283 32555
rect 25225 32515 25283 32521
rect 19794 32484 19800 32496
rect 19720 32456 19800 32484
rect 15436 32444 15442 32456
rect 19794 32444 19800 32456
rect 19852 32444 19858 32496
rect 22278 32444 22284 32496
rect 22336 32484 22342 32496
rect 22833 32487 22891 32493
rect 22833 32484 22845 32487
rect 22336 32456 22845 32484
rect 22336 32444 22342 32456
rect 22833 32453 22845 32456
rect 22879 32484 22891 32487
rect 23584 32484 23612 32512
rect 22879 32456 23520 32484
rect 23584 32456 24242 32484
rect 22879 32453 22891 32456
rect 22833 32447 22891 32453
rect 21818 32376 21824 32428
rect 21876 32416 21882 32428
rect 23492 32425 23520 32456
rect 25498 32444 25504 32496
rect 25556 32484 25562 32496
rect 25774 32484 25780 32496
rect 25556 32456 25780 32484
rect 25556 32444 25562 32456
rect 25774 32444 25780 32456
rect 25832 32444 25838 32496
rect 22097 32419 22155 32425
rect 22097 32416 22109 32419
rect 21876 32388 22109 32416
rect 21876 32376 21882 32388
rect 22097 32385 22109 32388
rect 22143 32385 22155 32419
rect 22097 32379 22155 32385
rect 23477 32419 23535 32425
rect 23477 32385 23489 32419
rect 23523 32385 23535 32419
rect 23477 32379 23535 32385
rect 13354 32308 13360 32360
rect 13412 32348 13418 32360
rect 16117 32351 16175 32357
rect 16117 32348 16129 32351
rect 13412 32320 16129 32348
rect 13412 32308 13418 32320
rect 16117 32317 16129 32320
rect 16163 32348 16175 32351
rect 16758 32348 16764 32360
rect 16163 32320 16764 32348
rect 16163 32317 16175 32320
rect 16117 32311 16175 32317
rect 16758 32308 16764 32320
rect 16816 32308 16822 32360
rect 19061 32351 19119 32357
rect 19061 32317 19073 32351
rect 19107 32317 19119 32351
rect 19061 32311 19119 32317
rect 19337 32351 19395 32357
rect 19337 32317 19349 32351
rect 19383 32348 19395 32351
rect 21174 32348 21180 32360
rect 19383 32320 21180 32348
rect 19383 32317 19395 32320
rect 19337 32311 19395 32317
rect 19076 32212 19104 32311
rect 21174 32308 21180 32320
rect 21232 32308 21238 32360
rect 23753 32351 23811 32357
rect 23753 32317 23765 32351
rect 23799 32348 23811 32351
rect 24946 32348 24952 32360
rect 23799 32320 24952 32348
rect 23799 32317 23811 32320
rect 23753 32311 23811 32317
rect 24946 32308 24952 32320
rect 25004 32308 25010 32360
rect 24854 32240 24860 32292
rect 24912 32280 24918 32292
rect 25038 32280 25044 32292
rect 24912 32252 25044 32280
rect 24912 32240 24918 32252
rect 25038 32240 25044 32252
rect 25096 32240 25102 32292
rect 19426 32212 19432 32224
rect 19076 32184 19432 32212
rect 19426 32172 19432 32184
rect 19484 32172 19490 32224
rect 20809 32215 20867 32221
rect 20809 32181 20821 32215
rect 20855 32212 20867 32215
rect 20898 32212 20904 32224
rect 20855 32184 20904 32212
rect 20855 32181 20867 32184
rect 20809 32175 20867 32181
rect 20898 32172 20904 32184
rect 20956 32172 20962 32224
rect 21637 32215 21695 32221
rect 21637 32181 21649 32215
rect 21683 32212 21695 32215
rect 21818 32212 21824 32224
rect 21683 32184 21824 32212
rect 21683 32181 21695 32184
rect 21637 32175 21695 32181
rect 21818 32172 21824 32184
rect 21876 32172 21882 32224
rect 22094 32172 22100 32224
rect 22152 32212 22158 32224
rect 26786 32212 26792 32224
rect 22152 32184 26792 32212
rect 22152 32172 22158 32184
rect 26786 32172 26792 32184
rect 26844 32172 26850 32224
rect 1104 32122 25852 32144
rect 1104 32070 2950 32122
rect 3002 32070 3014 32122
rect 3066 32070 3078 32122
rect 3130 32070 3142 32122
rect 3194 32070 3206 32122
rect 3258 32070 12950 32122
rect 13002 32070 13014 32122
rect 13066 32070 13078 32122
rect 13130 32070 13142 32122
rect 13194 32070 13206 32122
rect 13258 32070 22950 32122
rect 23002 32070 23014 32122
rect 23066 32070 23078 32122
rect 23130 32070 23142 32122
rect 23194 32070 23206 32122
rect 23258 32070 25852 32122
rect 1104 32048 25852 32070
rect 17024 32011 17082 32017
rect 17024 31977 17036 32011
rect 17070 32008 17082 32011
rect 18506 32008 18512 32020
rect 17070 31980 18512 32008
rect 17070 31977 17082 31980
rect 17024 31971 17082 31977
rect 18506 31968 18512 31980
rect 18564 31968 18570 32020
rect 22094 32008 22100 32020
rect 18616 31980 22100 32008
rect 12526 31900 12532 31952
rect 12584 31940 12590 31952
rect 15565 31943 15623 31949
rect 15565 31940 15577 31943
rect 12584 31912 15577 31940
rect 12584 31900 12590 31912
rect 15565 31909 15577 31912
rect 15611 31909 15623 31943
rect 15565 31903 15623 31909
rect 18046 31900 18052 31952
rect 18104 31940 18110 31952
rect 18616 31940 18644 31980
rect 22094 31968 22100 31980
rect 22152 31968 22158 32020
rect 22462 31968 22468 32020
rect 22520 32008 22526 32020
rect 22649 32011 22707 32017
rect 22649 32008 22661 32011
rect 22520 31980 22661 32008
rect 22520 31968 22526 31980
rect 22649 31977 22661 31980
rect 22695 32008 22707 32011
rect 23198 32008 23204 32020
rect 22695 31980 23204 32008
rect 22695 31977 22707 31980
rect 22649 31971 22707 31977
rect 23198 31968 23204 31980
rect 23256 31968 23262 32020
rect 18104 31912 18644 31940
rect 20732 31912 22232 31940
rect 18104 31900 18110 31912
rect 16114 31832 16120 31884
rect 16172 31832 16178 31884
rect 17678 31832 17684 31884
rect 17736 31872 17742 31884
rect 18509 31875 18567 31881
rect 18509 31872 18521 31875
rect 17736 31844 18521 31872
rect 17736 31832 17742 31844
rect 18509 31841 18521 31844
rect 18555 31841 18567 31875
rect 18509 31835 18567 31841
rect 19702 31832 19708 31884
rect 19760 31872 19766 31884
rect 20732 31872 20760 31912
rect 19760 31844 20760 31872
rect 19760 31832 19766 31844
rect 21910 31832 21916 31884
rect 21968 31872 21974 31884
rect 22204 31881 22232 31912
rect 22738 31900 22744 31952
rect 22796 31940 22802 31952
rect 23017 31943 23075 31949
rect 23017 31940 23029 31943
rect 22796 31912 23029 31940
rect 22796 31900 22802 31912
rect 23017 31909 23029 31912
rect 23063 31909 23075 31943
rect 23017 31903 23075 31909
rect 23382 31900 23388 31952
rect 23440 31940 23446 31952
rect 23440 31912 23704 31940
rect 23440 31900 23446 31912
rect 22097 31875 22155 31881
rect 22097 31872 22109 31875
rect 21968 31844 22109 31872
rect 21968 31832 21974 31844
rect 22097 31841 22109 31844
rect 22143 31841 22155 31875
rect 22097 31835 22155 31841
rect 22189 31875 22247 31881
rect 22189 31841 22201 31875
rect 22235 31841 22247 31875
rect 23569 31875 23627 31881
rect 23569 31872 23581 31875
rect 22189 31835 22247 31841
rect 23032 31844 23581 31872
rect 23032 31816 23060 31844
rect 23569 31841 23581 31844
rect 23615 31841 23627 31875
rect 23569 31835 23627 31841
rect 16758 31764 16764 31816
rect 16816 31764 16822 31816
rect 19426 31764 19432 31816
rect 19484 31764 19490 31816
rect 23014 31764 23020 31816
rect 23072 31764 23078 31816
rect 23477 31807 23535 31813
rect 23477 31773 23489 31807
rect 23523 31804 23535 31807
rect 23676 31804 23704 31912
rect 25038 31900 25044 31952
rect 25096 31940 25102 31952
rect 25133 31943 25191 31949
rect 25133 31940 25145 31943
rect 25096 31912 25145 31940
rect 25096 31900 25102 31912
rect 25133 31909 25145 31912
rect 25179 31909 25191 31943
rect 25133 31903 25191 31909
rect 23523 31776 23704 31804
rect 24857 31807 24915 31813
rect 23523 31773 23535 31776
rect 23477 31767 23535 31773
rect 24857 31773 24869 31807
rect 24903 31804 24915 31807
rect 25314 31804 25320 31816
rect 24903 31776 25320 31804
rect 24903 31773 24915 31776
rect 24857 31767 24915 31773
rect 25314 31764 25320 31776
rect 25372 31764 25378 31816
rect 15933 31739 15991 31745
rect 15933 31705 15945 31739
rect 15979 31736 15991 31739
rect 16666 31736 16672 31748
rect 15979 31708 16672 31736
rect 15979 31705 15991 31708
rect 15933 31699 15991 31705
rect 16666 31696 16672 31708
rect 16724 31696 16730 31748
rect 18785 31739 18843 31745
rect 18785 31736 18797 31739
rect 18262 31708 18797 31736
rect 18785 31705 18797 31708
rect 18831 31736 18843 31739
rect 19794 31736 19800 31748
rect 18831 31708 19800 31736
rect 18831 31705 18843 31708
rect 18785 31699 18843 31705
rect 19794 31696 19800 31708
rect 19852 31736 19858 31748
rect 19852 31708 20194 31736
rect 19852 31696 19858 31708
rect 23198 31696 23204 31748
rect 23256 31736 23262 31748
rect 23385 31739 23443 31745
rect 23385 31736 23397 31739
rect 23256 31708 23397 31736
rect 23256 31696 23262 31708
rect 23385 31705 23397 31708
rect 23431 31705 23443 31739
rect 23385 31699 23443 31705
rect 16025 31671 16083 31677
rect 16025 31637 16037 31671
rect 16071 31668 16083 31671
rect 16482 31668 16488 31680
rect 16071 31640 16488 31668
rect 16071 31637 16083 31640
rect 16025 31631 16083 31637
rect 16482 31628 16488 31640
rect 16540 31628 16546 31680
rect 20990 31628 20996 31680
rect 21048 31668 21054 31680
rect 21177 31671 21235 31677
rect 21177 31668 21189 31671
rect 21048 31640 21189 31668
rect 21048 31628 21054 31640
rect 21177 31637 21189 31640
rect 21223 31637 21235 31671
rect 21177 31631 21235 31637
rect 21634 31628 21640 31680
rect 21692 31628 21698 31680
rect 21726 31628 21732 31680
rect 21784 31668 21790 31680
rect 22002 31668 22008 31680
rect 21784 31640 22008 31668
rect 21784 31628 21790 31640
rect 22002 31628 22008 31640
rect 22060 31628 22066 31680
rect 22462 31628 22468 31680
rect 22520 31668 22526 31680
rect 22646 31668 22652 31680
rect 22520 31640 22652 31668
rect 22520 31628 22526 31640
rect 22646 31628 22652 31640
rect 22704 31628 22710 31680
rect 24670 31628 24676 31680
rect 24728 31628 24734 31680
rect 1104 31578 25852 31600
rect 1104 31526 7950 31578
rect 8002 31526 8014 31578
rect 8066 31526 8078 31578
rect 8130 31526 8142 31578
rect 8194 31526 8206 31578
rect 8258 31526 17950 31578
rect 18002 31526 18014 31578
rect 18066 31526 18078 31578
rect 18130 31526 18142 31578
rect 18194 31526 18206 31578
rect 18258 31526 25852 31578
rect 1104 31504 25852 31526
rect 16482 31424 16488 31476
rect 16540 31464 16546 31476
rect 17862 31464 17868 31476
rect 16540 31436 17868 31464
rect 16540 31424 16546 31436
rect 17862 31424 17868 31436
rect 17920 31424 17926 31476
rect 19153 31467 19211 31473
rect 19153 31433 19165 31467
rect 19199 31464 19211 31467
rect 19702 31464 19708 31476
rect 19199 31436 19708 31464
rect 19199 31433 19211 31436
rect 19153 31427 19211 31433
rect 19702 31424 19708 31436
rect 19760 31424 19766 31476
rect 21266 31424 21272 31476
rect 21324 31424 21330 31476
rect 23566 31424 23572 31476
rect 23624 31464 23630 31476
rect 23624 31436 24072 31464
rect 23624 31424 23630 31436
rect 14918 31396 14924 31408
rect 14858 31368 14924 31396
rect 14918 31356 14924 31368
rect 14976 31396 14982 31408
rect 15473 31399 15531 31405
rect 15473 31396 15485 31399
rect 14976 31368 15485 31396
rect 14976 31356 14982 31368
rect 15473 31365 15485 31368
rect 15519 31365 15531 31399
rect 15473 31359 15531 31365
rect 17681 31399 17739 31405
rect 17681 31365 17693 31399
rect 17727 31396 17739 31399
rect 17770 31396 17776 31408
rect 17727 31368 17776 31396
rect 17727 31365 17739 31368
rect 17681 31359 17739 31365
rect 17770 31356 17776 31368
rect 17828 31356 17834 31408
rect 19797 31399 19855 31405
rect 19797 31365 19809 31399
rect 19843 31396 19855 31399
rect 20441 31399 20499 31405
rect 20441 31396 20453 31399
rect 19843 31368 20453 31396
rect 19843 31365 19855 31368
rect 19797 31359 19855 31365
rect 20441 31365 20453 31368
rect 20487 31396 20499 31399
rect 20622 31396 20628 31408
rect 20487 31368 20628 31396
rect 20487 31365 20499 31368
rect 20441 31359 20499 31365
rect 20622 31356 20628 31368
rect 20680 31396 20686 31408
rect 21358 31396 21364 31408
rect 20680 31368 21364 31396
rect 20680 31356 20686 31368
rect 21358 31356 21364 31368
rect 21416 31356 21422 31408
rect 22646 31356 22652 31408
rect 22704 31396 22710 31408
rect 22741 31399 22799 31405
rect 22741 31396 22753 31399
rect 22704 31368 22753 31396
rect 22704 31356 22710 31368
rect 22741 31365 22753 31368
rect 22787 31396 22799 31399
rect 23014 31396 23020 31408
rect 22787 31368 23020 31396
rect 22787 31365 22799 31368
rect 22741 31359 22799 31365
rect 23014 31356 23020 31368
rect 23072 31356 23078 31408
rect 24044 31396 24072 31436
rect 24670 31396 24676 31408
rect 23966 31368 24676 31396
rect 24670 31356 24676 31368
rect 24728 31356 24734 31408
rect 16758 31288 16764 31340
rect 16816 31328 16822 31340
rect 17405 31331 17463 31337
rect 17405 31328 17417 31331
rect 16816 31300 17417 31328
rect 16816 31288 16822 31300
rect 17405 31297 17417 31300
rect 17451 31297 17463 31331
rect 19429 31331 19487 31337
rect 19429 31328 19441 31331
rect 18814 31300 19441 31328
rect 17405 31291 17463 31297
rect 19429 31297 19441 31300
rect 19475 31328 19487 31331
rect 19702 31328 19708 31340
rect 19475 31300 19708 31328
rect 19475 31297 19487 31300
rect 19429 31291 19487 31297
rect 19702 31288 19708 31300
rect 19760 31288 19766 31340
rect 20533 31331 20591 31337
rect 20533 31297 20545 31331
rect 20579 31328 20591 31331
rect 20579 31300 22232 31328
rect 20579 31297 20591 31300
rect 20533 31291 20591 31297
rect 13354 31220 13360 31272
rect 13412 31220 13418 31272
rect 13633 31263 13691 31269
rect 13633 31229 13645 31263
rect 13679 31260 13691 31263
rect 16114 31260 16120 31272
rect 13679 31232 16120 31260
rect 13679 31229 13691 31232
rect 13633 31223 13691 31229
rect 16114 31220 16120 31232
rect 16172 31220 16178 31272
rect 16666 31220 16672 31272
rect 16724 31260 16730 31272
rect 17218 31260 17224 31272
rect 16724 31232 17224 31260
rect 16724 31220 16730 31232
rect 17218 31220 17224 31232
rect 17276 31260 17282 31272
rect 20438 31260 20444 31272
rect 17276 31232 20444 31260
rect 17276 31220 17282 31232
rect 20438 31220 20444 31232
rect 20496 31220 20502 31272
rect 20622 31220 20628 31272
rect 20680 31220 20686 31272
rect 21545 31263 21603 31269
rect 21545 31229 21557 31263
rect 21591 31260 21603 31263
rect 22002 31260 22008 31272
rect 21591 31232 22008 31260
rect 21591 31229 21603 31232
rect 21545 31223 21603 31229
rect 22002 31220 22008 31232
rect 22060 31260 22066 31272
rect 22094 31260 22100 31272
rect 22060 31232 22100 31260
rect 22060 31220 22066 31232
rect 22094 31220 22100 31232
rect 22152 31220 22158 31272
rect 22204 31260 22232 31300
rect 22278 31288 22284 31340
rect 22336 31328 22342 31340
rect 22465 31331 22523 31337
rect 22465 31328 22477 31331
rect 22336 31300 22477 31328
rect 22336 31288 22342 31300
rect 22465 31297 22477 31300
rect 22511 31297 22523 31331
rect 22465 31291 22523 31297
rect 25317 31331 25375 31337
rect 25317 31297 25329 31331
rect 25363 31328 25375 31331
rect 25498 31328 25504 31340
rect 25363 31300 25504 31328
rect 25363 31297 25375 31300
rect 25317 31291 25375 31297
rect 25498 31288 25504 31300
rect 25556 31288 25562 31340
rect 25130 31260 25136 31272
rect 22204 31232 25136 31260
rect 25130 31220 25136 31232
rect 25188 31220 25194 31272
rect 20073 31195 20131 31201
rect 20073 31192 20085 31195
rect 18708 31164 20085 31192
rect 12342 31084 12348 31136
rect 12400 31124 12406 31136
rect 15105 31127 15163 31133
rect 15105 31124 15117 31127
rect 12400 31096 15117 31124
rect 12400 31084 12406 31096
rect 15105 31093 15117 31096
rect 15151 31093 15163 31127
rect 15105 31087 15163 31093
rect 17494 31084 17500 31136
rect 17552 31124 17558 31136
rect 18708 31124 18736 31164
rect 20073 31161 20085 31164
rect 20119 31161 20131 31195
rect 20073 31155 20131 31161
rect 23750 31152 23756 31204
rect 23808 31192 23814 31204
rect 24213 31195 24271 31201
rect 24213 31192 24225 31195
rect 23808 31164 24225 31192
rect 23808 31152 23814 31164
rect 24213 31161 24225 31164
rect 24259 31161 24271 31195
rect 24213 31155 24271 31161
rect 17552 31096 18736 31124
rect 17552 31084 17558 31096
rect 18782 31084 18788 31136
rect 18840 31124 18846 31136
rect 20622 31124 20628 31136
rect 18840 31096 20628 31124
rect 18840 31084 18846 31096
rect 20622 31084 20628 31096
rect 20680 31084 20686 31136
rect 24581 31127 24639 31133
rect 24581 31093 24593 31127
rect 24627 31124 24639 31127
rect 24670 31124 24676 31136
rect 24627 31096 24676 31124
rect 24627 31093 24639 31096
rect 24581 31087 24639 31093
rect 24670 31084 24676 31096
rect 24728 31084 24734 31136
rect 25130 31084 25136 31136
rect 25188 31084 25194 31136
rect 1104 31034 25852 31056
rect 1104 30982 2950 31034
rect 3002 30982 3014 31034
rect 3066 30982 3078 31034
rect 3130 30982 3142 31034
rect 3194 30982 3206 31034
rect 3258 30982 12950 31034
rect 13002 30982 13014 31034
rect 13066 30982 13078 31034
rect 13130 30982 13142 31034
rect 13194 30982 13206 31034
rect 13258 30982 22950 31034
rect 23002 30982 23014 31034
rect 23066 30982 23078 31034
rect 23130 30982 23142 31034
rect 23194 30982 23206 31034
rect 23258 30982 25852 31034
rect 1104 30960 25852 30982
rect 9125 30923 9183 30929
rect 9125 30889 9137 30923
rect 9171 30920 9183 30923
rect 9214 30920 9220 30932
rect 9171 30892 9220 30920
rect 9171 30889 9183 30892
rect 9125 30883 9183 30889
rect 9214 30880 9220 30892
rect 9272 30880 9278 30932
rect 15378 30880 15384 30932
rect 15436 30920 15442 30932
rect 15565 30923 15623 30929
rect 15565 30920 15577 30923
rect 15436 30892 15577 30920
rect 15436 30880 15442 30892
rect 15565 30889 15577 30892
rect 15611 30920 15623 30923
rect 15749 30923 15807 30929
rect 15749 30920 15761 30923
rect 15611 30892 15761 30920
rect 15611 30889 15623 30892
rect 15565 30883 15623 30889
rect 15749 30889 15761 30892
rect 15795 30889 15807 30923
rect 15749 30883 15807 30889
rect 18506 30880 18512 30932
rect 18564 30920 18570 30932
rect 18782 30920 18788 30932
rect 18564 30892 18788 30920
rect 18564 30880 18570 30892
rect 18782 30880 18788 30892
rect 18840 30880 18846 30932
rect 18874 30880 18880 30932
rect 18932 30920 18938 30932
rect 19702 30920 19708 30932
rect 18932 30892 19708 30920
rect 18932 30880 18938 30892
rect 19702 30880 19708 30892
rect 19760 30880 19766 30932
rect 22465 30923 22523 30929
rect 22465 30889 22477 30923
rect 22511 30920 22523 30923
rect 22646 30920 22652 30932
rect 22511 30892 22652 30920
rect 22511 30889 22523 30892
rect 22465 30883 22523 30889
rect 22646 30880 22652 30892
rect 22704 30880 22710 30932
rect 25498 30880 25504 30932
rect 25556 30880 25562 30932
rect 18064 30824 19334 30852
rect 16761 30787 16819 30793
rect 16761 30753 16773 30787
rect 16807 30784 16819 30787
rect 18064 30784 18092 30824
rect 16807 30756 18092 30784
rect 19306 30784 19334 30824
rect 19426 30784 19432 30796
rect 19306 30756 19432 30784
rect 16807 30753 16819 30756
rect 16761 30747 16819 30753
rect 19426 30744 19432 30756
rect 19484 30784 19490 30796
rect 20717 30787 20775 30793
rect 20717 30784 20729 30787
rect 19484 30756 20729 30784
rect 19484 30744 19490 30756
rect 20717 30753 20729 30756
rect 20763 30753 20775 30787
rect 20717 30747 20775 30753
rect 8754 30676 8760 30728
rect 8812 30716 8818 30728
rect 9309 30719 9367 30725
rect 9309 30716 9321 30719
rect 8812 30688 9321 30716
rect 8812 30676 8818 30688
rect 9309 30685 9321 30688
rect 9355 30685 9367 30719
rect 9309 30679 9367 30685
rect 14090 30676 14096 30728
rect 14148 30716 14154 30728
rect 14369 30719 14427 30725
rect 14369 30716 14381 30719
rect 14148 30688 14381 30716
rect 14148 30676 14154 30688
rect 14369 30685 14381 30688
rect 14415 30716 14427 30719
rect 15378 30716 15384 30728
rect 14415 30688 15384 30716
rect 14415 30685 14427 30688
rect 14369 30679 14427 30685
rect 15378 30676 15384 30688
rect 15436 30676 15442 30728
rect 15102 30608 15108 30660
rect 15160 30608 15166 30660
rect 17037 30651 17095 30657
rect 17037 30617 17049 30651
rect 17083 30617 17095 30651
rect 18262 30620 18828 30648
rect 17037 30611 17095 30617
rect 17052 30580 17080 30611
rect 18800 30592 18828 30620
rect 20990 30608 20996 30660
rect 21048 30608 21054 30660
rect 21266 30608 21272 30660
rect 21324 30648 21330 30660
rect 21324 30620 21482 30648
rect 21324 30608 21330 30620
rect 18690 30580 18696 30592
rect 17052 30552 18696 30580
rect 18690 30540 18696 30552
rect 18748 30540 18754 30592
rect 18782 30540 18788 30592
rect 18840 30540 18846 30592
rect 20070 30540 20076 30592
rect 20128 30540 20134 30592
rect 21376 30580 21404 30620
rect 22833 30583 22891 30589
rect 22833 30580 22845 30583
rect 21376 30552 22845 30580
rect 22833 30549 22845 30552
rect 22879 30549 22891 30583
rect 22833 30543 22891 30549
rect 22922 30540 22928 30592
rect 22980 30580 22986 30592
rect 24581 30583 24639 30589
rect 24581 30580 24593 30583
rect 22980 30552 24593 30580
rect 22980 30540 22986 30552
rect 24581 30549 24593 30552
rect 24627 30549 24639 30583
rect 24581 30543 24639 30549
rect 1104 30490 25852 30512
rect 1104 30438 7950 30490
rect 8002 30438 8014 30490
rect 8066 30438 8078 30490
rect 8130 30438 8142 30490
rect 8194 30438 8206 30490
rect 8258 30438 17950 30490
rect 18002 30438 18014 30490
rect 18066 30438 18078 30490
rect 18130 30438 18142 30490
rect 18194 30438 18206 30490
rect 18258 30438 25852 30490
rect 1104 30416 25852 30438
rect 13354 30376 13360 30388
rect 12406 30348 13360 30376
rect 12406 30308 12434 30348
rect 13354 30336 13360 30348
rect 13412 30336 13418 30388
rect 18248 30348 18460 30376
rect 11808 30280 12434 30308
rect 8478 30200 8484 30252
rect 8536 30240 8542 30252
rect 11808 30249 11836 30280
rect 12710 30268 12716 30320
rect 12768 30268 12774 30320
rect 14090 30268 14096 30320
rect 14148 30268 14154 30320
rect 14550 30268 14556 30320
rect 14608 30308 14614 30320
rect 18248 30308 18276 30348
rect 14608 30280 18276 30308
rect 18432 30308 18460 30348
rect 20070 30336 20076 30388
rect 20128 30376 20134 30388
rect 20257 30379 20315 30385
rect 20257 30376 20269 30379
rect 20128 30348 20269 30376
rect 20128 30336 20134 30348
rect 20257 30345 20269 30348
rect 20303 30345 20315 30379
rect 20257 30339 20315 30345
rect 22646 30336 22652 30388
rect 22704 30376 22710 30388
rect 23290 30376 23296 30388
rect 22704 30348 23296 30376
rect 22704 30336 22710 30348
rect 23290 30336 23296 30348
rect 23348 30336 23354 30388
rect 19978 30308 19984 30320
rect 18432 30280 19984 30308
rect 14608 30268 14614 30280
rect 19978 30268 19984 30280
rect 20036 30268 20042 30320
rect 20349 30311 20407 30317
rect 20349 30277 20361 30311
rect 20395 30308 20407 30311
rect 21910 30308 21916 30320
rect 20395 30280 21916 30308
rect 20395 30277 20407 30280
rect 20349 30271 20407 30277
rect 21910 30268 21916 30280
rect 21968 30268 21974 30320
rect 22465 30311 22523 30317
rect 22465 30277 22477 30311
rect 22511 30308 22523 30311
rect 22554 30308 22560 30320
rect 22511 30280 22560 30308
rect 22511 30277 22523 30280
rect 22465 30271 22523 30277
rect 22554 30268 22560 30280
rect 22612 30268 22618 30320
rect 9125 30243 9183 30249
rect 9125 30240 9137 30243
rect 8536 30212 9137 30240
rect 8536 30200 8542 30212
rect 9125 30209 9137 30212
rect 9171 30209 9183 30243
rect 9125 30203 9183 30209
rect 11793 30243 11851 30249
rect 11793 30209 11805 30243
rect 11839 30209 11851 30243
rect 11793 30203 11851 30209
rect 15841 30243 15899 30249
rect 15841 30209 15853 30243
rect 15887 30240 15899 30243
rect 16942 30240 16948 30252
rect 15887 30212 16948 30240
rect 15887 30209 15899 30212
rect 15841 30203 15899 30209
rect 16942 30200 16948 30212
rect 17000 30240 17006 30252
rect 21269 30243 21327 30249
rect 17000 30212 20668 30240
rect 17000 30200 17006 30212
rect 12066 30132 12072 30184
rect 12124 30132 12130 30184
rect 13354 30132 13360 30184
rect 13412 30172 13418 30184
rect 14829 30175 14887 30181
rect 14829 30172 14841 30175
rect 13412 30144 14841 30172
rect 13412 30132 13418 30144
rect 14829 30141 14841 30144
rect 14875 30141 14887 30175
rect 14829 30135 14887 30141
rect 15933 30175 15991 30181
rect 15933 30141 15945 30175
rect 15979 30141 15991 30175
rect 15933 30135 15991 30141
rect 8938 30064 8944 30116
rect 8996 30064 9002 30116
rect 15948 30104 15976 30135
rect 16022 30132 16028 30184
rect 16080 30132 16086 30184
rect 16758 30172 16764 30184
rect 16132 30144 16764 30172
rect 16132 30104 16160 30144
rect 16758 30132 16764 30144
rect 16816 30172 16822 30184
rect 20254 30172 20260 30184
rect 16816 30144 20260 30172
rect 16816 30132 16822 30144
rect 20254 30132 20260 30144
rect 20312 30132 20318 30184
rect 20530 30132 20536 30184
rect 20588 30132 20594 30184
rect 20640 30172 20668 30212
rect 21269 30209 21281 30243
rect 21315 30240 21327 30243
rect 22373 30243 22431 30249
rect 22373 30240 22385 30243
rect 21315 30212 22385 30240
rect 21315 30209 21327 30212
rect 21269 30203 21327 30209
rect 22373 30209 22385 30212
rect 22419 30209 22431 30243
rect 22373 30203 22431 30209
rect 24670 30200 24676 30252
rect 24728 30200 24734 30252
rect 22278 30172 22284 30184
rect 20640 30144 22284 30172
rect 22278 30132 22284 30144
rect 22336 30132 22342 30184
rect 22649 30175 22707 30181
rect 22649 30141 22661 30175
rect 22695 30172 22707 30175
rect 22830 30172 22836 30184
rect 22695 30144 22836 30172
rect 22695 30141 22707 30144
rect 22649 30135 22707 30141
rect 22830 30132 22836 30144
rect 22888 30132 22894 30184
rect 23290 30132 23296 30184
rect 23348 30132 23354 30184
rect 23569 30175 23627 30181
rect 23569 30141 23581 30175
rect 23615 30172 23627 30175
rect 23658 30172 23664 30184
rect 23615 30144 23664 30172
rect 23615 30141 23627 30144
rect 23569 30135 23627 30141
rect 23658 30132 23664 30144
rect 23716 30132 23722 30184
rect 15948 30076 16160 30104
rect 16482 30064 16488 30116
rect 16540 30104 16546 30116
rect 22462 30104 22468 30116
rect 16540 30076 22468 30104
rect 16540 30064 16546 30076
rect 22462 30064 22468 30076
rect 22520 30064 22526 30116
rect 24688 30104 24716 30200
rect 24946 30132 24952 30184
rect 25004 30172 25010 30184
rect 25041 30175 25099 30181
rect 25041 30172 25053 30175
rect 25004 30144 25053 30172
rect 25004 30132 25010 30144
rect 25041 30141 25053 30144
rect 25087 30141 25099 30175
rect 25041 30135 25099 30141
rect 25317 30107 25375 30113
rect 25317 30104 25329 30107
rect 24688 30076 25329 30104
rect 25317 30073 25329 30076
rect 25363 30073 25375 30107
rect 25317 30067 25375 30073
rect 11330 29996 11336 30048
rect 11388 30036 11394 30048
rect 13541 30039 13599 30045
rect 13541 30036 13553 30039
rect 11388 30008 13553 30036
rect 11388 29996 11394 30008
rect 13541 30005 13553 30008
rect 13587 30036 13599 30039
rect 13630 30036 13636 30048
rect 13587 30008 13636 30036
rect 13587 30005 13599 30008
rect 13541 29999 13599 30005
rect 13630 29996 13636 30008
rect 13688 29996 13694 30048
rect 15473 30039 15531 30045
rect 15473 30005 15485 30039
rect 15519 30036 15531 30039
rect 15930 30036 15936 30048
rect 15519 30008 15936 30036
rect 15519 30005 15531 30008
rect 15473 29999 15531 30005
rect 15930 29996 15936 30008
rect 15988 29996 15994 30048
rect 18782 29996 18788 30048
rect 18840 30036 18846 30048
rect 18877 30039 18935 30045
rect 18877 30036 18889 30039
rect 18840 30008 18889 30036
rect 18840 29996 18846 30008
rect 18877 30005 18889 30008
rect 18923 30005 18935 30039
rect 18877 29999 18935 30005
rect 19794 29996 19800 30048
rect 19852 30036 19858 30048
rect 19889 30039 19947 30045
rect 19889 30036 19901 30039
rect 19852 30008 19901 30036
rect 19852 29996 19858 30008
rect 19889 30005 19901 30008
rect 19935 30005 19947 30039
rect 19889 29999 19947 30005
rect 21910 29996 21916 30048
rect 21968 30036 21974 30048
rect 22005 30039 22063 30045
rect 22005 30036 22017 30039
rect 21968 30008 22017 30036
rect 21968 29996 21974 30008
rect 22005 30005 22017 30008
rect 22051 30005 22063 30039
rect 22005 29999 22063 30005
rect 1104 29946 25852 29968
rect 1104 29894 2950 29946
rect 3002 29894 3014 29946
rect 3066 29894 3078 29946
rect 3130 29894 3142 29946
rect 3194 29894 3206 29946
rect 3258 29894 12950 29946
rect 13002 29894 13014 29946
rect 13066 29894 13078 29946
rect 13130 29894 13142 29946
rect 13194 29894 13206 29946
rect 13258 29894 22950 29946
rect 23002 29894 23014 29946
rect 23066 29894 23078 29946
rect 23130 29894 23142 29946
rect 23194 29894 23206 29946
rect 23258 29894 25852 29946
rect 1104 29872 25852 29894
rect 12066 29792 12072 29844
rect 12124 29832 12130 29844
rect 12124 29804 12940 29832
rect 12124 29792 12130 29804
rect 12912 29773 12940 29804
rect 16482 29792 16488 29844
rect 16540 29792 16546 29844
rect 18690 29792 18696 29844
rect 18748 29832 18754 29844
rect 18785 29835 18843 29841
rect 18785 29832 18797 29835
rect 18748 29804 18797 29832
rect 18748 29792 18754 29804
rect 18785 29801 18797 29804
rect 18831 29801 18843 29835
rect 26510 29832 26516 29844
rect 18785 29795 18843 29801
rect 22066 29804 26516 29832
rect 12897 29767 12955 29773
rect 12897 29733 12909 29767
rect 12943 29764 12955 29767
rect 12943 29736 15884 29764
rect 12943 29733 12955 29736
rect 12897 29727 12955 29733
rect 11149 29699 11207 29705
rect 11149 29665 11161 29699
rect 11195 29696 11207 29699
rect 11422 29696 11428 29708
rect 11195 29668 11428 29696
rect 11195 29665 11207 29668
rect 11149 29659 11207 29665
rect 11422 29656 11428 29668
rect 11480 29696 11486 29708
rect 13354 29696 13360 29708
rect 11480 29668 13360 29696
rect 11480 29656 11486 29668
rect 13354 29656 13360 29668
rect 13412 29656 13418 29708
rect 15856 29705 15884 29736
rect 18414 29724 18420 29776
rect 18472 29764 18478 29776
rect 20165 29767 20223 29773
rect 20165 29764 20177 29767
rect 18472 29736 20177 29764
rect 18472 29724 18478 29736
rect 20165 29733 20177 29736
rect 20211 29733 20223 29767
rect 20165 29727 20223 29733
rect 20254 29724 20260 29776
rect 20312 29764 20318 29776
rect 22066 29764 22094 29804
rect 26510 29792 26516 29804
rect 26568 29792 26574 29844
rect 20312 29736 22094 29764
rect 20312 29724 20318 29736
rect 23198 29724 23204 29776
rect 23256 29764 23262 29776
rect 25133 29767 25191 29773
rect 25133 29764 25145 29767
rect 23256 29736 25145 29764
rect 23256 29724 23262 29736
rect 25133 29733 25145 29736
rect 25179 29733 25191 29767
rect 25133 29727 25191 29733
rect 15841 29699 15899 29705
rect 15841 29665 15853 29699
rect 15887 29696 15899 29699
rect 16022 29696 16028 29708
rect 15887 29668 16028 29696
rect 15887 29665 15899 29668
rect 15841 29659 15899 29665
rect 16022 29656 16028 29668
rect 16080 29656 16086 29708
rect 17037 29699 17095 29705
rect 17037 29665 17049 29699
rect 17083 29696 17095 29699
rect 19334 29696 19340 29708
rect 17083 29668 19340 29696
rect 17083 29665 17095 29668
rect 17037 29659 17095 29665
rect 19334 29656 19340 29668
rect 19392 29656 19398 29708
rect 20717 29699 20775 29705
rect 20717 29696 20729 29699
rect 19444 29668 20729 29696
rect 15657 29631 15715 29637
rect 15657 29597 15669 29631
rect 15703 29628 15715 29631
rect 16482 29628 16488 29640
rect 15703 29600 16488 29628
rect 15703 29597 15715 29600
rect 15657 29591 15715 29597
rect 16482 29588 16488 29600
rect 16540 29588 16546 29640
rect 18874 29588 18880 29640
rect 18932 29628 18938 29640
rect 19444 29628 19472 29668
rect 20717 29665 20729 29668
rect 20763 29665 20775 29699
rect 20717 29659 20775 29665
rect 18932 29600 19472 29628
rect 23385 29631 23443 29637
rect 18932 29588 18938 29600
rect 23385 29597 23397 29631
rect 23431 29597 23443 29631
rect 23385 29591 23443 29597
rect 24029 29631 24087 29637
rect 24029 29597 24041 29631
rect 24075 29628 24087 29631
rect 24486 29628 24492 29640
rect 24075 29600 24492 29628
rect 24075 29597 24087 29600
rect 24029 29591 24087 29597
rect 11054 29520 11060 29572
rect 11112 29560 11118 29572
rect 11425 29563 11483 29569
rect 11425 29560 11437 29563
rect 11112 29532 11437 29560
rect 11112 29520 11118 29532
rect 11425 29529 11437 29532
rect 11471 29529 11483 29563
rect 12710 29560 12716 29572
rect 12650 29532 12716 29560
rect 11425 29523 11483 29529
rect 12710 29520 12716 29532
rect 12768 29560 12774 29572
rect 13173 29563 13231 29569
rect 13173 29560 13185 29563
rect 12768 29532 13185 29560
rect 12768 29520 12774 29532
rect 13173 29529 13185 29532
rect 13219 29560 13231 29563
rect 13633 29563 13691 29569
rect 13633 29560 13645 29563
rect 13219 29532 13645 29560
rect 13219 29529 13231 29532
rect 13173 29523 13231 29529
rect 13633 29529 13645 29532
rect 13679 29560 13691 29563
rect 13722 29560 13728 29572
rect 13679 29532 13728 29560
rect 13679 29529 13691 29532
rect 13633 29523 13691 29529
rect 13722 29520 13728 29532
rect 13780 29520 13786 29572
rect 15562 29520 15568 29572
rect 15620 29560 15626 29572
rect 17313 29563 17371 29569
rect 15620 29532 16344 29560
rect 15620 29520 15626 29532
rect 16316 29504 16344 29532
rect 17313 29529 17325 29563
rect 17359 29529 17371 29563
rect 18782 29560 18788 29572
rect 18538 29532 18788 29560
rect 17313 29523 17371 29529
rect 15194 29452 15200 29504
rect 15252 29452 15258 29504
rect 16298 29452 16304 29504
rect 16356 29452 16362 29504
rect 17328 29492 17356 29523
rect 18782 29520 18788 29532
rect 18840 29520 18846 29572
rect 20625 29563 20683 29569
rect 20625 29529 20637 29563
rect 20671 29560 20683 29563
rect 20714 29560 20720 29572
rect 20671 29532 20720 29560
rect 20671 29529 20683 29532
rect 20625 29523 20683 29529
rect 20714 29520 20720 29532
rect 20772 29520 20778 29572
rect 22925 29563 22983 29569
rect 22925 29529 22937 29563
rect 22971 29560 22983 29563
rect 23400 29560 23428 29591
rect 24486 29588 24492 29600
rect 24544 29588 24550 29640
rect 25314 29588 25320 29640
rect 25372 29588 25378 29640
rect 24946 29560 24952 29572
rect 22971 29532 24952 29560
rect 22971 29529 22983 29532
rect 22925 29523 22983 29529
rect 24946 29520 24952 29532
rect 25004 29520 25010 29572
rect 18874 29492 18880 29504
rect 17328 29464 18880 29492
rect 18874 29452 18880 29464
rect 18932 29452 18938 29504
rect 19150 29452 19156 29504
rect 19208 29492 19214 29504
rect 19429 29495 19487 29501
rect 19429 29492 19441 29495
rect 19208 29464 19441 29492
rect 19208 29452 19214 29464
rect 19429 29461 19441 29464
rect 19475 29461 19487 29495
rect 19429 29455 19487 29461
rect 19978 29452 19984 29504
rect 20036 29492 20042 29504
rect 20533 29495 20591 29501
rect 20533 29492 20545 29495
rect 20036 29464 20545 29492
rect 20036 29452 20042 29464
rect 20533 29461 20545 29464
rect 20579 29461 20591 29495
rect 20533 29455 20591 29461
rect 22646 29452 22652 29504
rect 22704 29492 22710 29504
rect 23201 29495 23259 29501
rect 23201 29492 23213 29495
rect 22704 29464 23213 29492
rect 22704 29452 22710 29464
rect 23201 29461 23213 29464
rect 23247 29461 23259 29495
rect 23201 29455 23259 29461
rect 23845 29495 23903 29501
rect 23845 29461 23857 29495
rect 23891 29492 23903 29495
rect 24302 29492 24308 29504
rect 23891 29464 24308 29492
rect 23891 29461 23903 29464
rect 23845 29455 23903 29461
rect 24302 29452 24308 29464
rect 24360 29452 24366 29504
rect 24486 29452 24492 29504
rect 24544 29452 24550 29504
rect 1104 29402 25852 29424
rect 1104 29350 7950 29402
rect 8002 29350 8014 29402
rect 8066 29350 8078 29402
rect 8130 29350 8142 29402
rect 8194 29350 8206 29402
rect 8258 29350 17950 29402
rect 18002 29350 18014 29402
rect 18066 29350 18078 29402
rect 18130 29350 18142 29402
rect 18194 29350 18206 29402
rect 18258 29350 25852 29402
rect 1104 29328 25852 29350
rect 8846 29248 8852 29300
rect 8904 29288 8910 29300
rect 9493 29291 9551 29297
rect 9493 29288 9505 29291
rect 8904 29260 9505 29288
rect 8904 29248 8910 29260
rect 9493 29257 9505 29260
rect 9539 29257 9551 29291
rect 9493 29251 9551 29257
rect 12526 29248 12532 29300
rect 12584 29248 12590 29300
rect 12618 29248 12624 29300
rect 12676 29248 12682 29300
rect 13446 29248 13452 29300
rect 13504 29288 13510 29300
rect 15105 29291 15163 29297
rect 15105 29288 15117 29291
rect 13504 29260 15117 29288
rect 13504 29248 13510 29260
rect 15105 29257 15117 29260
rect 15151 29257 15163 29291
rect 15105 29251 15163 29257
rect 9861 29223 9919 29229
rect 9861 29189 9873 29223
rect 9907 29220 9919 29223
rect 10318 29220 10324 29232
rect 9907 29192 10324 29220
rect 9907 29189 9919 29192
rect 9861 29183 9919 29189
rect 10318 29180 10324 29192
rect 10376 29180 10382 29232
rect 14918 29220 14924 29232
rect 14858 29192 14924 29220
rect 14918 29180 14924 29192
rect 14976 29180 14982 29232
rect 15120 29220 15148 29251
rect 15194 29248 15200 29300
rect 15252 29288 15258 29300
rect 16025 29291 16083 29297
rect 16025 29288 16037 29291
rect 15252 29260 16037 29288
rect 15252 29248 15258 29260
rect 16025 29257 16037 29260
rect 16071 29257 16083 29291
rect 16025 29251 16083 29257
rect 16298 29248 16304 29300
rect 16356 29288 16362 29300
rect 16356 29260 17356 29288
rect 16356 29248 16362 29260
rect 15838 29220 15844 29232
rect 15120 29192 15844 29220
rect 15838 29180 15844 29192
rect 15896 29180 15902 29232
rect 15930 29180 15936 29232
rect 15988 29180 15994 29232
rect 17126 29180 17132 29232
rect 17184 29220 17190 29232
rect 17328 29220 17356 29260
rect 17402 29248 17408 29300
rect 17460 29288 17466 29300
rect 17865 29291 17923 29297
rect 17865 29288 17877 29291
rect 17460 29260 17877 29288
rect 17460 29248 17466 29260
rect 17865 29257 17877 29260
rect 17911 29257 17923 29291
rect 17865 29251 17923 29257
rect 19150 29248 19156 29300
rect 19208 29248 19214 29300
rect 19245 29291 19303 29297
rect 19245 29257 19257 29291
rect 19291 29288 19303 29291
rect 19426 29288 19432 29300
rect 19291 29260 19432 29288
rect 19291 29257 19303 29260
rect 19245 29251 19303 29257
rect 19426 29248 19432 29260
rect 19484 29248 19490 29300
rect 19978 29248 19984 29300
rect 20036 29288 20042 29300
rect 20162 29288 20168 29300
rect 20036 29260 20168 29288
rect 20036 29248 20042 29260
rect 20162 29248 20168 29260
rect 20220 29288 20226 29300
rect 23937 29291 23995 29297
rect 23937 29288 23949 29291
rect 20220 29260 23949 29288
rect 20220 29248 20226 29260
rect 23937 29257 23949 29260
rect 23983 29288 23995 29291
rect 24118 29288 24124 29300
rect 23983 29260 24124 29288
rect 23983 29257 23995 29260
rect 23937 29251 23995 29257
rect 24118 29248 24124 29260
rect 24176 29288 24182 29300
rect 24762 29288 24768 29300
rect 24176 29260 24768 29288
rect 24176 29248 24182 29260
rect 24762 29248 24768 29260
rect 24820 29248 24826 29300
rect 25314 29248 25320 29300
rect 25372 29288 25378 29300
rect 25409 29291 25467 29297
rect 25409 29288 25421 29291
rect 25372 29260 25421 29288
rect 25372 29248 25378 29260
rect 25409 29257 25421 29260
rect 25455 29257 25467 29291
rect 25409 29251 25467 29257
rect 24029 29223 24087 29229
rect 17184 29192 17264 29220
rect 17328 29192 23888 29220
rect 17184 29180 17190 29192
rect 9953 29155 10011 29161
rect 9953 29121 9965 29155
rect 9999 29152 10011 29155
rect 10226 29152 10232 29164
rect 9999 29124 10232 29152
rect 9999 29121 10011 29124
rect 9953 29115 10011 29121
rect 10226 29112 10232 29124
rect 10284 29112 10290 29164
rect 13354 29112 13360 29164
rect 13412 29112 13418 29164
rect 17236 29161 17264 29192
rect 17221 29155 17279 29161
rect 17221 29121 17233 29155
rect 17267 29152 17279 29155
rect 22189 29155 22247 29161
rect 22189 29152 22201 29155
rect 17267 29124 17540 29152
rect 17267 29121 17279 29124
rect 17221 29115 17279 29121
rect 9674 29044 9680 29096
rect 9732 29084 9738 29096
rect 10045 29087 10103 29093
rect 10045 29084 10057 29087
rect 9732 29056 10057 29084
rect 9732 29044 9738 29056
rect 10045 29053 10057 29056
rect 10091 29084 10103 29087
rect 10870 29084 10876 29096
rect 10091 29056 10876 29084
rect 10091 29053 10103 29056
rect 10045 29047 10103 29053
rect 10870 29044 10876 29056
rect 10928 29044 10934 29096
rect 11146 29044 11152 29096
rect 11204 29084 11210 29096
rect 12342 29084 12348 29096
rect 11204 29056 12348 29084
rect 11204 29044 11210 29056
rect 12342 29044 12348 29056
rect 12400 29084 12406 29096
rect 12713 29087 12771 29093
rect 12713 29084 12725 29087
rect 12400 29056 12725 29084
rect 12400 29044 12406 29056
rect 12713 29053 12725 29056
rect 12759 29053 12771 29087
rect 12713 29047 12771 29053
rect 13630 29044 13636 29096
rect 13688 29084 13694 29096
rect 16117 29087 16175 29093
rect 16117 29084 16129 29087
rect 13688 29056 16129 29084
rect 13688 29044 13694 29056
rect 16117 29053 16129 29056
rect 16163 29053 16175 29087
rect 16117 29047 16175 29053
rect 17310 29044 17316 29096
rect 17368 29044 17374 29096
rect 17402 29044 17408 29096
rect 17460 29044 17466 29096
rect 17512 29028 17540 29124
rect 22066 29124 22201 29152
rect 19429 29087 19487 29093
rect 19429 29053 19441 29087
rect 19475 29084 19487 29087
rect 20898 29084 20904 29096
rect 19475 29056 20904 29084
rect 19475 29053 19487 29056
rect 19429 29047 19487 29053
rect 20898 29044 20904 29056
rect 20956 29044 20962 29096
rect 12161 29019 12219 29025
rect 12161 28985 12173 29019
rect 12207 29016 12219 29019
rect 12250 29016 12256 29028
rect 12207 28988 12256 29016
rect 12207 28985 12219 28988
rect 12161 28979 12219 28985
rect 12250 28976 12256 28988
rect 12308 28976 12314 29028
rect 15565 29019 15623 29025
rect 15565 29016 15577 29019
rect 14660 28988 15577 29016
rect 13620 28951 13678 28957
rect 13620 28917 13632 28951
rect 13666 28948 13678 28951
rect 14090 28948 14096 28960
rect 13666 28920 14096 28948
rect 13666 28917 13678 28920
rect 13620 28911 13678 28917
rect 14090 28908 14096 28920
rect 14148 28908 14154 28960
rect 14182 28908 14188 28960
rect 14240 28948 14246 28960
rect 14660 28948 14688 28988
rect 15565 28985 15577 28988
rect 15611 28985 15623 29019
rect 15565 28979 15623 28985
rect 15746 28976 15752 29028
rect 15804 29016 15810 29028
rect 16853 29019 16911 29025
rect 16853 29016 16865 29019
rect 15804 28988 16865 29016
rect 15804 28976 15810 28988
rect 16853 28985 16865 28988
rect 16899 28985 16911 29019
rect 16853 28979 16911 28985
rect 17494 28976 17500 29028
rect 17552 29016 17558 29028
rect 18049 29019 18107 29025
rect 18049 29016 18061 29019
rect 17552 28988 18061 29016
rect 17552 28976 17558 28988
rect 18049 28985 18061 28988
rect 18095 28985 18107 29019
rect 18049 28979 18107 28985
rect 18785 29019 18843 29025
rect 18785 28985 18797 29019
rect 18831 29016 18843 29019
rect 19058 29016 19064 29028
rect 18831 28988 19064 29016
rect 18831 28985 18843 28988
rect 18785 28979 18843 28985
rect 19058 28976 19064 28988
rect 19116 28976 19122 29028
rect 21818 28976 21824 29028
rect 21876 29016 21882 29028
rect 22066 29016 22094 29124
rect 22189 29121 22201 29124
rect 22235 29121 22247 29155
rect 22189 29115 22247 29121
rect 23017 29087 23075 29093
rect 23017 29053 23029 29087
rect 23063 29084 23075 29087
rect 23382 29084 23388 29096
rect 23063 29056 23388 29084
rect 23063 29053 23075 29056
rect 23017 29047 23075 29053
rect 23382 29044 23388 29056
rect 23440 29044 23446 29096
rect 23860 29084 23888 29192
rect 24029 29189 24041 29223
rect 24075 29220 24087 29223
rect 26418 29220 26424 29232
rect 24075 29192 26424 29220
rect 24075 29189 24087 29192
rect 24029 29183 24087 29189
rect 26418 29180 26424 29192
rect 26476 29180 26482 29232
rect 26878 29152 26884 29164
rect 24044 29124 26884 29152
rect 24044 29084 24072 29124
rect 26878 29112 26884 29124
rect 26936 29112 26942 29164
rect 23860 29056 24072 29084
rect 24210 29044 24216 29096
rect 24268 29044 24274 29096
rect 24765 29087 24823 29093
rect 24765 29053 24777 29087
rect 24811 29084 24823 29087
rect 24946 29084 24952 29096
rect 24811 29056 24952 29084
rect 24811 29053 24823 29056
rect 24765 29047 24823 29053
rect 24946 29044 24952 29056
rect 25004 29044 25010 29096
rect 21876 28988 22094 29016
rect 23569 29019 23627 29025
rect 21876 28976 21882 28988
rect 23569 28985 23581 29019
rect 23615 29016 23627 29019
rect 24394 29016 24400 29028
rect 23615 28988 24400 29016
rect 23615 28985 23627 28988
rect 23569 28979 23627 28985
rect 24394 28976 24400 28988
rect 24452 28976 24458 29028
rect 14240 28920 14688 28948
rect 14240 28908 14246 28920
rect 22094 28908 22100 28960
rect 22152 28948 22158 28960
rect 22462 28948 22468 28960
rect 22152 28920 22468 28948
rect 22152 28908 22158 28920
rect 22462 28908 22468 28920
rect 22520 28908 22526 28960
rect 25222 28908 25228 28960
rect 25280 28908 25286 28960
rect 1104 28858 25852 28880
rect 1104 28806 2950 28858
rect 3002 28806 3014 28858
rect 3066 28806 3078 28858
rect 3130 28806 3142 28858
rect 3194 28806 3206 28858
rect 3258 28806 12950 28858
rect 13002 28806 13014 28858
rect 13066 28806 13078 28858
rect 13130 28806 13142 28858
rect 13194 28806 13206 28858
rect 13258 28806 22950 28858
rect 23002 28806 23014 28858
rect 23066 28806 23078 28858
rect 23130 28806 23142 28858
rect 23194 28806 23206 28858
rect 23258 28806 25852 28858
rect 1104 28784 25852 28806
rect 10870 28704 10876 28756
rect 10928 28704 10934 28756
rect 13541 28747 13599 28753
rect 13541 28713 13553 28747
rect 13587 28744 13599 28747
rect 13722 28744 13728 28756
rect 13587 28716 13728 28744
rect 13587 28713 13599 28716
rect 13541 28707 13599 28713
rect 13722 28704 13728 28716
rect 13780 28744 13786 28756
rect 15010 28744 15016 28756
rect 13780 28716 15016 28744
rect 13780 28704 13786 28716
rect 15010 28704 15016 28716
rect 15068 28744 15074 28756
rect 15933 28747 15991 28753
rect 15933 28744 15945 28747
rect 15068 28716 15945 28744
rect 15068 28704 15074 28716
rect 15933 28713 15945 28716
rect 15979 28744 15991 28747
rect 18782 28744 18788 28756
rect 15979 28716 18788 28744
rect 15979 28713 15991 28716
rect 15933 28707 15991 28713
rect 18782 28704 18788 28716
rect 18840 28704 18846 28756
rect 18874 28704 18880 28756
rect 18932 28704 18938 28756
rect 21082 28704 21088 28756
rect 21140 28744 21146 28756
rect 22833 28747 22891 28753
rect 22833 28744 22845 28747
rect 21140 28716 22845 28744
rect 21140 28704 21146 28716
rect 22833 28713 22845 28716
rect 22879 28713 22891 28747
rect 25498 28744 25504 28756
rect 22833 28707 22891 28713
rect 23216 28716 25504 28744
rect 16206 28676 16212 28688
rect 15304 28648 16212 28676
rect 9125 28611 9183 28617
rect 9125 28577 9137 28611
rect 9171 28608 9183 28611
rect 11422 28608 11428 28620
rect 9171 28580 11428 28608
rect 9171 28577 9183 28580
rect 9125 28571 9183 28577
rect 11422 28568 11428 28580
rect 11480 28568 11486 28620
rect 13173 28611 13231 28617
rect 13173 28577 13185 28611
rect 13219 28608 13231 28611
rect 14090 28608 14096 28620
rect 13219 28580 14096 28608
rect 13219 28577 13231 28580
rect 13173 28571 13231 28577
rect 14090 28568 14096 28580
rect 14148 28568 14154 28620
rect 15304 28617 15332 28648
rect 16206 28636 16212 28648
rect 16264 28636 16270 28688
rect 22554 28636 22560 28688
rect 22612 28676 22618 28688
rect 23216 28676 23244 28716
rect 25498 28704 25504 28716
rect 25556 28704 25562 28756
rect 25406 28676 25412 28688
rect 22612 28648 23244 28676
rect 23308 28648 25412 28676
rect 22612 28636 22618 28648
rect 15289 28611 15347 28617
rect 15289 28577 15301 28611
rect 15335 28577 15347 28611
rect 15289 28571 15347 28577
rect 15378 28568 15384 28620
rect 15436 28568 15442 28620
rect 17405 28611 17463 28617
rect 17405 28577 17417 28611
rect 17451 28608 17463 28611
rect 18966 28608 18972 28620
rect 17451 28580 18972 28608
rect 17451 28577 17463 28580
rect 17405 28571 17463 28577
rect 18966 28568 18972 28580
rect 19024 28568 19030 28620
rect 20073 28611 20131 28617
rect 20073 28577 20085 28611
rect 20119 28608 20131 28611
rect 20990 28608 20996 28620
rect 20119 28580 20996 28608
rect 20119 28577 20131 28580
rect 20073 28571 20131 28577
rect 20990 28568 20996 28580
rect 21048 28568 21054 28620
rect 21450 28568 21456 28620
rect 21508 28608 21514 28620
rect 23308 28617 23336 28648
rect 25406 28636 25412 28648
rect 25464 28636 25470 28688
rect 23293 28611 23351 28617
rect 21508 28580 21956 28608
rect 21508 28568 21514 28580
rect 15102 28500 15108 28552
rect 15160 28540 15166 28552
rect 17129 28543 17187 28549
rect 17129 28540 17141 28543
rect 15160 28512 17141 28540
rect 15160 28500 15166 28512
rect 17129 28509 17141 28512
rect 17175 28509 17187 28543
rect 17129 28503 17187 28509
rect 19334 28500 19340 28552
rect 19392 28540 19398 28552
rect 20622 28540 20628 28552
rect 19392 28512 20628 28540
rect 19392 28500 19398 28512
rect 20622 28500 20628 28512
rect 20680 28500 20686 28552
rect 21928 28540 21956 28580
rect 23293 28577 23305 28611
rect 23339 28577 23351 28611
rect 23293 28571 23351 28577
rect 23385 28611 23443 28617
rect 23385 28577 23397 28611
rect 23431 28608 23443 28611
rect 23566 28608 23572 28620
rect 23431 28580 23572 28608
rect 23431 28577 23443 28580
rect 23385 28571 23443 28577
rect 23566 28568 23572 28580
rect 23624 28568 23630 28620
rect 24854 28568 24860 28620
rect 24912 28608 24918 28620
rect 25133 28611 25191 28617
rect 25133 28608 25145 28611
rect 24912 28580 25145 28608
rect 24912 28568 24918 28580
rect 25133 28577 25145 28580
rect 25179 28577 25191 28611
rect 25133 28571 25191 28577
rect 23845 28543 23903 28549
rect 23845 28540 23857 28543
rect 21928 28512 23857 28540
rect 23845 28509 23857 28512
rect 23891 28540 23903 28543
rect 23934 28540 23940 28552
rect 23891 28512 23940 28540
rect 23891 28509 23903 28512
rect 23845 28503 23903 28509
rect 23934 28500 23940 28512
rect 23992 28500 23998 28552
rect 24578 28500 24584 28552
rect 24636 28500 24642 28552
rect 24946 28500 24952 28552
rect 25004 28500 25010 28552
rect 9401 28475 9459 28481
rect 9401 28441 9413 28475
rect 9447 28472 9459 28475
rect 9447 28444 9812 28472
rect 10626 28444 11284 28472
rect 9447 28441 9459 28444
rect 9401 28435 9459 28441
rect 9784 28416 9812 28444
rect 11256 28416 11284 28444
rect 11330 28432 11336 28484
rect 11388 28472 11394 28484
rect 11701 28475 11759 28481
rect 11701 28472 11713 28475
rect 11388 28444 11713 28472
rect 11388 28432 11394 28444
rect 11701 28441 11713 28444
rect 11747 28441 11759 28475
rect 13722 28472 13728 28484
rect 12926 28444 13728 28472
rect 11701 28435 11759 28441
rect 9766 28364 9772 28416
rect 9824 28364 9830 28416
rect 11238 28364 11244 28416
rect 11296 28404 11302 28416
rect 12618 28404 12624 28416
rect 11296 28376 12624 28404
rect 11296 28364 11302 28376
rect 12618 28364 12624 28376
rect 12676 28404 12682 28416
rect 13004 28404 13032 28444
rect 13722 28432 13728 28444
rect 13780 28432 13786 28484
rect 15197 28475 15255 28481
rect 15197 28441 15209 28475
rect 15243 28472 15255 28475
rect 18782 28472 18788 28484
rect 15243 28444 16068 28472
rect 18630 28444 18788 28472
rect 15243 28441 15255 28444
rect 15197 28435 15255 28441
rect 16040 28416 16068 28444
rect 18782 28432 18788 28444
rect 18840 28432 18846 28484
rect 20898 28432 20904 28484
rect 20956 28432 20962 28484
rect 21450 28432 21456 28484
rect 21508 28432 21514 28484
rect 24210 28472 24216 28484
rect 22388 28444 24216 28472
rect 12676 28376 13032 28404
rect 12676 28364 12682 28376
rect 14826 28364 14832 28416
rect 14884 28364 14890 28416
rect 16022 28364 16028 28416
rect 16080 28364 16086 28416
rect 16206 28364 16212 28416
rect 16264 28364 16270 28416
rect 19429 28407 19487 28413
rect 19429 28373 19441 28407
rect 19475 28404 19487 28407
rect 19518 28404 19524 28416
rect 19475 28376 19524 28404
rect 19475 28373 19487 28376
rect 19429 28367 19487 28373
rect 19518 28364 19524 28376
rect 19576 28364 19582 28416
rect 19702 28364 19708 28416
rect 19760 28404 19766 28416
rect 19797 28407 19855 28413
rect 19797 28404 19809 28407
rect 19760 28376 19809 28404
rect 19760 28364 19766 28376
rect 19797 28373 19809 28376
rect 19843 28373 19855 28407
rect 19797 28367 19855 28373
rect 19889 28407 19947 28413
rect 19889 28373 19901 28407
rect 19935 28404 19947 28407
rect 21634 28404 21640 28416
rect 19935 28376 21640 28404
rect 19935 28373 19947 28376
rect 19889 28367 19947 28373
rect 21634 28364 21640 28376
rect 21692 28364 21698 28416
rect 22388 28413 22416 28444
rect 24210 28432 24216 28444
rect 24268 28432 24274 28484
rect 24596 28472 24624 28500
rect 25041 28475 25099 28481
rect 25041 28472 25053 28475
rect 24596 28444 25053 28472
rect 25041 28441 25053 28444
rect 25087 28441 25099 28475
rect 25041 28435 25099 28441
rect 22373 28407 22431 28413
rect 22373 28373 22385 28407
rect 22419 28373 22431 28407
rect 22373 28367 22431 28373
rect 22462 28364 22468 28416
rect 22520 28404 22526 28416
rect 23201 28407 23259 28413
rect 23201 28404 23213 28407
rect 22520 28376 23213 28404
rect 22520 28364 22526 28376
rect 23201 28373 23213 28376
rect 23247 28404 23259 28407
rect 24029 28407 24087 28413
rect 24029 28404 24041 28407
rect 23247 28376 24041 28404
rect 23247 28373 23259 28376
rect 23201 28367 23259 28373
rect 24029 28373 24041 28376
rect 24075 28373 24087 28407
rect 24029 28367 24087 28373
rect 24486 28364 24492 28416
rect 24544 28404 24550 28416
rect 24581 28407 24639 28413
rect 24581 28404 24593 28407
rect 24544 28376 24593 28404
rect 24544 28364 24550 28376
rect 24581 28373 24593 28376
rect 24627 28373 24639 28407
rect 24581 28367 24639 28373
rect 1104 28314 25852 28336
rect 1104 28262 7950 28314
rect 8002 28262 8014 28314
rect 8066 28262 8078 28314
rect 8130 28262 8142 28314
rect 8194 28262 8206 28314
rect 8258 28262 17950 28314
rect 18002 28262 18014 28314
rect 18066 28262 18078 28314
rect 18130 28262 18142 28314
rect 18194 28262 18206 28314
rect 18258 28262 25852 28314
rect 1104 28240 25852 28262
rect 3418 28160 3424 28212
rect 3476 28200 3482 28212
rect 3476 28172 18736 28200
rect 3476 28160 3482 28172
rect 11057 28135 11115 28141
rect 11057 28101 11069 28135
rect 11103 28132 11115 28135
rect 11238 28132 11244 28144
rect 11103 28104 11244 28132
rect 11103 28101 11115 28104
rect 11057 28095 11115 28101
rect 11238 28092 11244 28104
rect 11296 28092 11302 28144
rect 13722 28132 13728 28144
rect 13202 28104 13728 28132
rect 13722 28092 13728 28104
rect 13780 28092 13786 28144
rect 15565 28135 15623 28141
rect 15565 28101 15577 28135
rect 15611 28132 15623 28135
rect 15930 28132 15936 28144
rect 15611 28104 15936 28132
rect 15611 28101 15623 28104
rect 15565 28095 15623 28101
rect 15930 28092 15936 28104
rect 15988 28132 15994 28144
rect 16390 28132 16396 28144
rect 15988 28104 16396 28132
rect 15988 28092 15994 28104
rect 16390 28092 16396 28104
rect 16448 28092 16454 28144
rect 17218 28092 17224 28144
rect 17276 28092 17282 28144
rect 18708 28132 18736 28172
rect 18782 28160 18788 28212
rect 18840 28200 18846 28212
rect 18969 28203 19027 28209
rect 18969 28200 18981 28203
rect 18840 28172 18981 28200
rect 18840 28160 18846 28172
rect 18969 28169 18981 28172
rect 19015 28169 19027 28203
rect 18969 28163 19027 28169
rect 19702 28160 19708 28212
rect 19760 28160 19766 28212
rect 21545 28203 21603 28209
rect 21545 28200 21557 28203
rect 19812 28172 21557 28200
rect 19812 28132 19840 28172
rect 21545 28169 21557 28172
rect 21591 28200 21603 28203
rect 22465 28203 22523 28209
rect 21591 28172 22094 28200
rect 21591 28169 21603 28172
rect 21545 28163 21603 28169
rect 18708 28104 19840 28132
rect 20622 28092 20628 28144
rect 20680 28132 20686 28144
rect 21085 28135 21143 28141
rect 21085 28132 21097 28135
rect 20680 28104 21097 28132
rect 20680 28092 20686 28104
rect 21085 28101 21097 28104
rect 21131 28101 21143 28135
rect 22066 28132 22094 28172
rect 22465 28169 22477 28203
rect 22511 28200 22523 28203
rect 26234 28200 26240 28212
rect 22511 28172 26240 28200
rect 22511 28169 22523 28172
rect 22465 28163 22523 28169
rect 26234 28160 26240 28172
rect 26292 28160 26298 28212
rect 22373 28135 22431 28141
rect 22373 28132 22385 28135
rect 22066 28104 22385 28132
rect 21085 28095 21143 28101
rect 22373 28101 22385 28104
rect 22419 28132 22431 28135
rect 22554 28132 22560 28144
rect 22419 28104 22560 28132
rect 22419 28101 22431 28104
rect 22373 28095 22431 28101
rect 22554 28092 22560 28104
rect 22612 28092 22618 28144
rect 23382 28132 23388 28144
rect 23216 28104 23388 28132
rect 15654 28024 15660 28076
rect 15712 28064 15718 28076
rect 16298 28064 16304 28076
rect 15712 28036 16304 28064
rect 15712 28024 15718 28036
rect 16298 28024 16304 28036
rect 16356 28024 16362 28076
rect 17313 28067 17371 28073
rect 17313 28033 17325 28067
rect 17359 28064 17371 28067
rect 17862 28064 17868 28076
rect 17359 28036 17868 28064
rect 17359 28033 17371 28036
rect 17313 28027 17371 28033
rect 17862 28024 17868 28036
rect 17920 28064 17926 28076
rect 20349 28067 20407 28073
rect 17920 28036 18644 28064
rect 17920 28024 17926 28036
rect 11698 27956 11704 28008
rect 11756 27956 11762 28008
rect 11974 27956 11980 28008
rect 12032 27956 12038 28008
rect 15749 27999 15807 28005
rect 15749 27965 15761 27999
rect 15795 27965 15807 27999
rect 15749 27959 15807 27965
rect 10778 27888 10784 27940
rect 10836 27928 10842 27940
rect 15378 27928 15384 27940
rect 10836 27900 11836 27928
rect 10836 27888 10842 27900
rect 11808 27860 11836 27900
rect 13464 27900 15384 27928
rect 13464 27869 13492 27900
rect 15378 27888 15384 27900
rect 15436 27928 15442 27940
rect 15764 27928 15792 27959
rect 17402 27956 17408 28008
rect 17460 27956 17466 28008
rect 17954 27956 17960 28008
rect 18012 27996 18018 28008
rect 18616 28005 18644 28036
rect 20349 28033 20361 28067
rect 20395 28064 20407 28067
rect 21818 28064 21824 28076
rect 20395 28036 21824 28064
rect 20395 28033 20407 28036
rect 20349 28027 20407 28033
rect 18049 27999 18107 28005
rect 18049 27996 18061 27999
rect 18012 27968 18061 27996
rect 18012 27956 18018 27968
rect 18049 27965 18061 27968
rect 18095 27965 18107 27999
rect 18049 27959 18107 27965
rect 18601 27999 18659 28005
rect 18601 27965 18613 27999
rect 18647 27996 18659 27999
rect 18782 27996 18788 28008
rect 18647 27968 18788 27996
rect 18647 27965 18659 27968
rect 18601 27959 18659 27965
rect 18782 27956 18788 27968
rect 18840 27956 18846 28008
rect 15436 27900 15792 27928
rect 15436 27888 15442 27900
rect 17678 27888 17684 27940
rect 17736 27928 17742 27940
rect 19337 27931 19395 27937
rect 19337 27928 19349 27931
rect 17736 27900 19349 27928
rect 17736 27888 17742 27900
rect 19337 27897 19349 27900
rect 19383 27928 19395 27931
rect 20364 27928 20392 28027
rect 21818 28024 21824 28036
rect 21876 28024 21882 28076
rect 23216 28073 23244 28104
rect 23382 28092 23388 28104
rect 23440 28092 23446 28144
rect 23934 28092 23940 28144
rect 23992 28092 23998 28144
rect 23201 28067 23259 28073
rect 23201 28033 23213 28067
rect 23247 28033 23259 28067
rect 23201 28027 23259 28033
rect 22554 27956 22560 28008
rect 22612 27956 22618 28008
rect 23474 27956 23480 28008
rect 23532 27956 23538 28008
rect 23934 27956 23940 28008
rect 23992 27996 23998 28008
rect 25222 27996 25228 28008
rect 23992 27968 25228 27996
rect 23992 27956 23998 27968
rect 25222 27956 25228 27968
rect 25280 27956 25286 28008
rect 19383 27900 20392 27928
rect 19383 27897 19395 27900
rect 19337 27891 19395 27897
rect 13449 27863 13507 27869
rect 13449 27860 13461 27863
rect 11808 27832 13461 27860
rect 13449 27829 13461 27832
rect 13495 27829 13507 27863
rect 13449 27823 13507 27829
rect 13814 27820 13820 27872
rect 13872 27860 13878 27872
rect 15197 27863 15255 27869
rect 15197 27860 15209 27863
rect 13872 27832 15209 27860
rect 13872 27820 13878 27832
rect 15197 27829 15209 27832
rect 15243 27829 15255 27863
rect 15197 27823 15255 27829
rect 16298 27820 16304 27872
rect 16356 27820 16362 27872
rect 16850 27820 16856 27872
rect 16908 27820 16914 27872
rect 17218 27820 17224 27872
rect 17276 27860 17282 27872
rect 18506 27860 18512 27872
rect 17276 27832 18512 27860
rect 17276 27820 17282 27832
rect 18506 27820 18512 27832
rect 18564 27860 18570 27872
rect 18693 27863 18751 27869
rect 18693 27860 18705 27863
rect 18564 27832 18705 27860
rect 18564 27820 18570 27832
rect 18693 27829 18705 27832
rect 18739 27829 18751 27863
rect 18693 27823 18751 27829
rect 20714 27820 20720 27872
rect 20772 27860 20778 27872
rect 22005 27863 22063 27869
rect 22005 27860 22017 27863
rect 20772 27832 22017 27860
rect 20772 27820 20778 27832
rect 22005 27829 22017 27832
rect 22051 27829 22063 27863
rect 22005 27823 22063 27829
rect 22370 27820 22376 27872
rect 22428 27860 22434 27872
rect 24949 27863 25007 27869
rect 24949 27860 24961 27863
rect 22428 27832 24961 27860
rect 22428 27820 22434 27832
rect 24949 27829 24961 27832
rect 24995 27829 25007 27863
rect 24949 27823 25007 27829
rect 25406 27820 25412 27872
rect 25464 27820 25470 27872
rect 1104 27770 25852 27792
rect 1104 27718 2950 27770
rect 3002 27718 3014 27770
rect 3066 27718 3078 27770
rect 3130 27718 3142 27770
rect 3194 27718 3206 27770
rect 3258 27718 12950 27770
rect 13002 27718 13014 27770
rect 13066 27718 13078 27770
rect 13130 27718 13142 27770
rect 13194 27718 13206 27770
rect 13258 27718 22950 27770
rect 23002 27718 23014 27770
rect 23066 27718 23078 27770
rect 23130 27718 23142 27770
rect 23194 27718 23206 27770
rect 23258 27718 25852 27770
rect 1104 27696 25852 27718
rect 11422 27656 11428 27668
rect 10612 27628 11428 27656
rect 10505 27523 10563 27529
rect 10505 27489 10517 27523
rect 10551 27520 10563 27523
rect 10612 27520 10640 27628
rect 11422 27616 11428 27628
rect 11480 27616 11486 27668
rect 11790 27616 11796 27668
rect 11848 27656 11854 27668
rect 15102 27656 15108 27668
rect 11848 27628 15108 27656
rect 11848 27616 11854 27628
rect 12434 27588 12440 27600
rect 11900 27560 12440 27588
rect 10551 27492 10640 27520
rect 10551 27489 10563 27492
rect 10505 27483 10563 27489
rect 10778 27480 10784 27532
rect 10836 27480 10842 27532
rect 11900 27438 11928 27560
rect 12434 27548 12440 27560
rect 12492 27588 12498 27600
rect 12618 27588 12624 27600
rect 12492 27560 12624 27588
rect 12492 27548 12498 27560
rect 12618 27548 12624 27560
rect 12676 27548 12682 27600
rect 13078 27548 13084 27600
rect 13136 27588 13142 27600
rect 13188 27588 13216 27628
rect 15102 27616 15108 27628
rect 15160 27616 15166 27668
rect 20152 27659 20210 27665
rect 20152 27625 20164 27659
rect 20198 27656 20210 27659
rect 23566 27656 23572 27668
rect 20198 27628 23572 27656
rect 20198 27625 20210 27628
rect 20152 27619 20210 27625
rect 23566 27616 23572 27628
rect 23624 27656 23630 27668
rect 23845 27659 23903 27665
rect 23845 27656 23857 27659
rect 23624 27628 23857 27656
rect 23624 27616 23630 27628
rect 23845 27625 23857 27628
rect 23891 27625 23903 27659
rect 23845 27619 23903 27625
rect 13136 27560 13216 27588
rect 13136 27548 13142 27560
rect 23474 27548 23480 27600
rect 23532 27588 23538 27600
rect 24762 27588 24768 27600
rect 23532 27560 24768 27588
rect 23532 27548 23538 27560
rect 24762 27548 24768 27560
rect 24820 27588 24826 27600
rect 24820 27560 25176 27588
rect 24820 27548 24826 27560
rect 12253 27523 12311 27529
rect 12253 27489 12265 27523
rect 12299 27520 12311 27523
rect 13541 27523 13599 27529
rect 13541 27520 13553 27523
rect 12299 27492 13553 27520
rect 12299 27489 12311 27492
rect 12253 27483 12311 27489
rect 13541 27489 13553 27492
rect 13587 27489 13599 27523
rect 13541 27483 13599 27489
rect 9582 27276 9588 27328
rect 9640 27316 9646 27328
rect 12268 27316 12296 27483
rect 15102 27480 15108 27532
rect 15160 27520 15166 27532
rect 15749 27523 15807 27529
rect 15749 27520 15761 27523
rect 15160 27492 15761 27520
rect 15160 27480 15166 27492
rect 15749 27489 15761 27492
rect 15795 27489 15807 27523
rect 15749 27483 15807 27489
rect 17770 27480 17776 27532
rect 17828 27520 17834 27532
rect 18049 27523 18107 27529
rect 18049 27520 18061 27523
rect 17828 27492 18061 27520
rect 17828 27480 17834 27492
rect 18049 27489 18061 27492
rect 18095 27489 18107 27523
rect 18049 27483 18107 27489
rect 19889 27523 19947 27529
rect 19889 27489 19901 27523
rect 19935 27520 19947 27523
rect 22097 27523 22155 27529
rect 22097 27520 22109 27523
rect 19935 27492 22109 27520
rect 19935 27489 19947 27492
rect 19889 27483 19947 27489
rect 22097 27489 22109 27492
rect 22143 27520 22155 27523
rect 23382 27520 23388 27532
rect 22143 27492 23388 27520
rect 22143 27489 22155 27492
rect 22097 27483 22155 27489
rect 23382 27480 23388 27492
rect 23440 27480 23446 27532
rect 24118 27480 24124 27532
rect 24176 27480 24182 27532
rect 25038 27480 25044 27532
rect 25096 27480 25102 27532
rect 25148 27529 25176 27560
rect 25133 27523 25191 27529
rect 25133 27489 25145 27523
rect 25179 27489 25191 27523
rect 25133 27483 25191 27489
rect 13449 27455 13507 27461
rect 13449 27421 13461 27455
rect 13495 27452 13507 27455
rect 14826 27452 14832 27464
rect 13495 27424 14832 27452
rect 13495 27421 13507 27424
rect 13449 27415 13507 27421
rect 14826 27412 14832 27424
rect 14884 27412 14890 27464
rect 15657 27455 15715 27461
rect 15657 27421 15669 27455
rect 15703 27452 15715 27455
rect 16206 27452 16212 27464
rect 15703 27424 16212 27452
rect 15703 27421 15715 27424
rect 15657 27415 15715 27421
rect 16206 27412 16212 27424
rect 16264 27452 16270 27464
rect 16393 27455 16451 27461
rect 16393 27452 16405 27455
rect 16264 27424 16405 27452
rect 16264 27412 16270 27424
rect 16393 27421 16405 27424
rect 16439 27421 16451 27455
rect 16393 27415 16451 27421
rect 17865 27455 17923 27461
rect 17865 27421 17877 27455
rect 17911 27452 17923 27455
rect 17954 27452 17960 27464
rect 17911 27424 17960 27452
rect 17911 27421 17923 27424
rect 17865 27415 17923 27421
rect 17954 27412 17960 27424
rect 18012 27412 18018 27464
rect 23934 27452 23940 27464
rect 23506 27424 23940 27452
rect 23934 27412 23940 27424
rect 23992 27412 23998 27464
rect 24949 27455 25007 27461
rect 24949 27421 24961 27455
rect 24995 27452 25007 27455
rect 25406 27452 25412 27464
rect 24995 27424 25412 27452
rect 24995 27421 25007 27424
rect 24949 27415 25007 27421
rect 25406 27412 25412 27424
rect 25464 27412 25470 27464
rect 13357 27387 13415 27393
rect 13357 27353 13369 27387
rect 13403 27384 13415 27387
rect 13814 27384 13820 27396
rect 13403 27356 13820 27384
rect 13403 27353 13415 27356
rect 13357 27347 13415 27353
rect 13814 27344 13820 27356
rect 13872 27344 13878 27396
rect 15565 27387 15623 27393
rect 15565 27353 15577 27387
rect 15611 27384 15623 27387
rect 21450 27384 21456 27396
rect 15611 27356 16068 27384
rect 21390 27356 21456 27384
rect 15611 27353 15623 27356
rect 15565 27347 15623 27353
rect 16040 27328 16068 27356
rect 21450 27344 21456 27356
rect 21508 27384 21514 27396
rect 21818 27384 21824 27396
rect 21508 27356 21824 27384
rect 21508 27344 21514 27356
rect 21818 27344 21824 27356
rect 21876 27344 21882 27396
rect 22370 27344 22376 27396
rect 22428 27344 22434 27396
rect 9640 27288 12296 27316
rect 9640 27276 9646 27288
rect 12618 27276 12624 27328
rect 12676 27316 12682 27328
rect 12989 27319 13047 27325
rect 12989 27316 13001 27319
rect 12676 27288 13001 27316
rect 12676 27276 12682 27288
rect 12989 27285 13001 27288
rect 13035 27285 13047 27319
rect 12989 27279 13047 27285
rect 13722 27276 13728 27328
rect 13780 27316 13786 27328
rect 15197 27319 15255 27325
rect 15197 27316 15209 27319
rect 13780 27288 15209 27316
rect 13780 27276 13786 27288
rect 15197 27285 15209 27288
rect 15243 27285 15255 27319
rect 15197 27279 15255 27285
rect 16022 27276 16028 27328
rect 16080 27316 16086 27328
rect 16209 27319 16267 27325
rect 16209 27316 16221 27319
rect 16080 27288 16221 27316
rect 16080 27276 16086 27288
rect 16209 27285 16221 27288
rect 16255 27285 16267 27319
rect 16209 27279 16267 27285
rect 16482 27276 16488 27328
rect 16540 27316 16546 27328
rect 17497 27319 17555 27325
rect 17497 27316 17509 27319
rect 16540 27288 17509 27316
rect 16540 27276 16546 27288
rect 17497 27285 17509 27288
rect 17543 27285 17555 27319
rect 17497 27279 17555 27285
rect 17586 27276 17592 27328
rect 17644 27316 17650 27328
rect 17957 27319 18015 27325
rect 17957 27316 17969 27319
rect 17644 27288 17969 27316
rect 17644 27276 17650 27288
rect 17957 27285 17969 27288
rect 18003 27285 18015 27319
rect 17957 27279 18015 27285
rect 21634 27276 21640 27328
rect 21692 27276 21698 27328
rect 24578 27276 24584 27328
rect 24636 27276 24642 27328
rect 24854 27276 24860 27328
rect 24912 27316 24918 27328
rect 25314 27316 25320 27328
rect 24912 27288 25320 27316
rect 24912 27276 24918 27288
rect 25314 27276 25320 27288
rect 25372 27276 25378 27328
rect 1104 27226 25852 27248
rect 1104 27174 7950 27226
rect 8002 27174 8014 27226
rect 8066 27174 8078 27226
rect 8130 27174 8142 27226
rect 8194 27174 8206 27226
rect 8258 27174 17950 27226
rect 18002 27174 18014 27226
rect 18066 27174 18078 27226
rect 18130 27174 18142 27226
rect 18194 27174 18206 27226
rect 18258 27174 25852 27226
rect 1104 27152 25852 27174
rect 11054 27072 11060 27124
rect 11112 27072 11118 27124
rect 11609 27115 11667 27121
rect 11609 27081 11621 27115
rect 11655 27112 11667 27115
rect 12434 27112 12440 27124
rect 11655 27084 12440 27112
rect 11655 27081 11667 27084
rect 11609 27075 11667 27081
rect 9582 27004 9588 27056
rect 9640 27004 9646 27056
rect 11238 27044 11244 27056
rect 10810 27016 11244 27044
rect 11238 27004 11244 27016
rect 11296 27044 11302 27056
rect 11624 27044 11652 27075
rect 12434 27072 12440 27084
rect 12492 27112 12498 27124
rect 13538 27112 13544 27124
rect 12492 27084 13544 27112
rect 12492 27072 12498 27084
rect 13538 27072 13544 27084
rect 13596 27112 13602 27124
rect 15657 27115 15715 27121
rect 13596 27084 13768 27112
rect 13596 27072 13602 27084
rect 11296 27016 11652 27044
rect 13357 27047 13415 27053
rect 11296 27004 11302 27016
rect 13357 27013 13369 27047
rect 13403 27044 13415 27047
rect 13446 27044 13452 27056
rect 13403 27016 13452 27044
rect 13403 27013 13415 27016
rect 13357 27007 13415 27013
rect 13446 27004 13452 27016
rect 13504 27004 13510 27056
rect 13740 27044 13768 27084
rect 15657 27081 15669 27115
rect 15703 27112 15715 27115
rect 16850 27112 16856 27124
rect 15703 27084 16856 27112
rect 15703 27081 15715 27084
rect 15657 27075 15715 27081
rect 16850 27072 16856 27084
rect 16908 27072 16914 27124
rect 19242 27112 19248 27124
rect 18064 27084 19248 27112
rect 13740 27016 13846 27044
rect 15746 27004 15752 27056
rect 15804 27004 15810 27056
rect 18064 27044 18092 27084
rect 19242 27072 19248 27084
rect 19300 27072 19306 27124
rect 22738 27072 22744 27124
rect 22796 27112 22802 27124
rect 22833 27115 22891 27121
rect 22833 27112 22845 27115
rect 22796 27084 22845 27112
rect 22796 27072 22802 27084
rect 22833 27081 22845 27084
rect 22879 27081 22891 27115
rect 23658 27112 23664 27124
rect 22833 27075 22891 27081
rect 23032 27084 23664 27112
rect 20070 27044 20076 27056
rect 17972 27016 18092 27044
rect 19458 27016 20076 27044
rect 12710 26936 12716 26988
rect 12768 26976 12774 26988
rect 13078 26976 13084 26988
rect 12768 26948 13084 26976
rect 12768 26936 12774 26948
rect 13078 26936 13084 26948
rect 13136 26936 13142 26988
rect 14734 26936 14740 26988
rect 14792 26976 14798 26988
rect 16758 26976 16764 26988
rect 14792 26948 16764 26976
rect 14792 26936 14798 26948
rect 16758 26936 16764 26948
rect 16816 26936 16822 26988
rect 17972 26985 18000 27016
rect 20070 27004 20076 27016
rect 20128 27004 20134 27056
rect 17957 26979 18015 26985
rect 17957 26945 17969 26979
rect 18003 26945 18015 26979
rect 17957 26939 18015 26945
rect 22741 26979 22799 26985
rect 22741 26945 22753 26979
rect 22787 26976 22799 26979
rect 22922 26976 22928 26988
rect 22787 26948 22928 26976
rect 22787 26945 22799 26948
rect 22741 26939 22799 26945
rect 22922 26936 22928 26948
rect 22980 26936 22986 26988
rect 9309 26911 9367 26917
rect 9309 26877 9321 26911
rect 9355 26877 9367 26911
rect 9309 26871 9367 26877
rect 15841 26911 15899 26917
rect 15841 26877 15853 26911
rect 15887 26877 15899 26911
rect 15841 26871 15899 26877
rect 18233 26911 18291 26917
rect 18233 26877 18245 26911
rect 18279 26908 18291 26911
rect 22094 26908 22100 26920
rect 18279 26880 22100 26908
rect 18279 26877 18291 26880
rect 18233 26871 18291 26877
rect 9324 26772 9352 26871
rect 15856 26840 15884 26871
rect 22094 26868 22100 26880
rect 22152 26908 22158 26920
rect 22554 26908 22560 26920
rect 22152 26880 22560 26908
rect 22152 26868 22158 26880
rect 22554 26868 22560 26880
rect 22612 26868 22618 26920
rect 23032 26917 23060 27084
rect 23658 27072 23664 27084
rect 23716 27072 23722 27124
rect 24762 27072 24768 27124
rect 24820 27112 24826 27124
rect 25317 27115 25375 27121
rect 25317 27112 25329 27115
rect 24820 27084 25329 27112
rect 24820 27072 24826 27084
rect 25317 27081 25329 27084
rect 25363 27081 25375 27115
rect 25317 27075 25375 27081
rect 23934 27004 23940 27056
rect 23992 27044 23998 27056
rect 23992 27016 24334 27044
rect 23992 27004 23998 27016
rect 25222 27004 25228 27056
rect 25280 27044 25286 27056
rect 25498 27044 25504 27056
rect 25280 27016 25504 27044
rect 25280 27004 25286 27016
rect 25498 27004 25504 27016
rect 25556 27004 25562 27056
rect 25774 26936 25780 26988
rect 25832 26976 25838 26988
rect 26050 26976 26056 26988
rect 25832 26948 26056 26976
rect 25832 26936 25838 26948
rect 26050 26936 26056 26948
rect 26108 26936 26114 26988
rect 23017 26911 23075 26917
rect 23017 26877 23029 26911
rect 23063 26877 23075 26911
rect 23017 26871 23075 26877
rect 23382 26868 23388 26920
rect 23440 26908 23446 26920
rect 23569 26911 23627 26917
rect 23569 26908 23581 26911
rect 23440 26880 23581 26908
rect 23440 26868 23446 26880
rect 23569 26877 23581 26880
rect 23615 26877 23627 26911
rect 23569 26871 23627 26877
rect 23845 26911 23903 26917
rect 23845 26877 23857 26911
rect 23891 26908 23903 26911
rect 25498 26908 25504 26920
rect 23891 26880 25504 26908
rect 23891 26877 23903 26880
rect 23845 26871 23903 26877
rect 25498 26868 25504 26880
rect 25556 26868 25562 26920
rect 14844 26812 15884 26840
rect 9674 26772 9680 26784
rect 9324 26744 9680 26772
rect 9674 26732 9680 26744
rect 9732 26732 9738 26784
rect 12066 26732 12072 26784
rect 12124 26772 12130 26784
rect 14844 26781 14872 26812
rect 22462 26800 22468 26852
rect 22520 26840 22526 26852
rect 22830 26840 22836 26852
rect 22520 26812 22836 26840
rect 22520 26800 22526 26812
rect 22830 26800 22836 26812
rect 22888 26800 22894 26852
rect 14829 26775 14887 26781
rect 14829 26772 14841 26775
rect 12124 26744 14841 26772
rect 12124 26732 12130 26744
rect 14829 26741 14841 26744
rect 14875 26741 14887 26775
rect 14829 26735 14887 26741
rect 14918 26732 14924 26784
rect 14976 26772 14982 26784
rect 15289 26775 15347 26781
rect 15289 26772 15301 26775
rect 14976 26744 15301 26772
rect 14976 26732 14982 26744
rect 15289 26741 15301 26744
rect 15335 26741 15347 26775
rect 15289 26735 15347 26741
rect 18966 26732 18972 26784
rect 19024 26772 19030 26784
rect 19705 26775 19763 26781
rect 19705 26772 19717 26775
rect 19024 26744 19717 26772
rect 19024 26732 19030 26744
rect 19705 26741 19717 26744
rect 19751 26741 19763 26775
rect 19705 26735 19763 26741
rect 20070 26732 20076 26784
rect 20128 26772 20134 26784
rect 21818 26772 21824 26784
rect 20128 26744 21824 26772
rect 20128 26732 20134 26744
rect 21818 26732 21824 26744
rect 21876 26732 21882 26784
rect 22186 26732 22192 26784
rect 22244 26772 22250 26784
rect 22373 26775 22431 26781
rect 22373 26772 22385 26775
rect 22244 26744 22385 26772
rect 22244 26732 22250 26744
rect 22373 26741 22385 26744
rect 22419 26741 22431 26775
rect 22373 26735 22431 26741
rect 1104 26682 25852 26704
rect 1104 26630 2950 26682
rect 3002 26630 3014 26682
rect 3066 26630 3078 26682
rect 3130 26630 3142 26682
rect 3194 26630 3206 26682
rect 3258 26630 12950 26682
rect 13002 26630 13014 26682
rect 13066 26630 13078 26682
rect 13130 26630 13142 26682
rect 13194 26630 13206 26682
rect 13258 26630 22950 26682
rect 23002 26630 23014 26682
rect 23066 26630 23078 26682
rect 23130 26630 23142 26682
rect 23194 26630 23206 26682
rect 23258 26630 25852 26682
rect 1104 26608 25852 26630
rect 10873 26571 10931 26577
rect 10873 26537 10885 26571
rect 10919 26568 10931 26571
rect 11974 26568 11980 26580
rect 10919 26540 11980 26568
rect 10919 26537 10931 26540
rect 10873 26531 10931 26537
rect 11974 26528 11980 26540
rect 12032 26568 12038 26580
rect 12342 26568 12348 26580
rect 12032 26540 12348 26568
rect 12032 26528 12038 26540
rect 12342 26528 12348 26540
rect 12400 26528 12406 26580
rect 13538 26528 13544 26580
rect 13596 26568 13602 26580
rect 15289 26571 15347 26577
rect 15289 26568 15301 26571
rect 13596 26540 15301 26568
rect 13596 26528 13602 26540
rect 15289 26537 15301 26540
rect 15335 26537 15347 26571
rect 15289 26531 15347 26537
rect 16942 26528 16948 26580
rect 17000 26528 17006 26580
rect 21177 26571 21235 26577
rect 21177 26537 21189 26571
rect 21223 26568 21235 26571
rect 22094 26568 22100 26580
rect 21223 26540 22100 26568
rect 21223 26537 21235 26540
rect 21177 26531 21235 26537
rect 22094 26528 22100 26540
rect 22152 26528 22158 26580
rect 23845 26571 23903 26577
rect 23845 26537 23857 26571
rect 23891 26568 23903 26571
rect 24946 26568 24952 26580
rect 23891 26540 24952 26568
rect 23891 26537 23903 26540
rect 23845 26531 23903 26537
rect 24946 26528 24952 26540
rect 25004 26528 25010 26580
rect 25222 26568 25228 26580
rect 25148 26540 25228 26568
rect 11238 26460 11244 26512
rect 11296 26460 11302 26512
rect 13630 26460 13636 26512
rect 13688 26500 13694 26512
rect 15657 26503 15715 26509
rect 15657 26500 15669 26503
rect 13688 26472 15669 26500
rect 13688 26460 13694 26472
rect 15657 26469 15669 26472
rect 15703 26469 15715 26503
rect 15657 26463 15715 26469
rect 15930 26460 15936 26512
rect 15988 26500 15994 26512
rect 17218 26500 17224 26512
rect 15988 26472 17224 26500
rect 15988 26460 15994 26472
rect 17218 26460 17224 26472
rect 17276 26460 17282 26512
rect 22462 26460 22468 26512
rect 22520 26500 22526 26512
rect 22649 26503 22707 26509
rect 22649 26500 22661 26503
rect 22520 26472 22661 26500
rect 22520 26460 22526 26472
rect 22649 26469 22661 26472
rect 22695 26469 22707 26503
rect 22649 26463 22707 26469
rect 24581 26503 24639 26509
rect 24581 26469 24593 26503
rect 24627 26500 24639 26503
rect 25038 26500 25044 26512
rect 24627 26472 25044 26500
rect 24627 26469 24639 26472
rect 24581 26463 24639 26469
rect 25038 26460 25044 26472
rect 25096 26460 25102 26512
rect 7742 26392 7748 26444
rect 7800 26432 7806 26444
rect 9401 26435 9459 26441
rect 9401 26432 9413 26435
rect 7800 26404 9413 26432
rect 7800 26392 7806 26404
rect 9401 26401 9413 26404
rect 9447 26432 9459 26435
rect 11146 26432 11152 26444
rect 9447 26404 11152 26432
rect 9447 26401 9459 26404
rect 9401 26395 9459 26401
rect 11146 26392 11152 26404
rect 11204 26392 11210 26444
rect 14458 26392 14464 26444
rect 14516 26432 14522 26444
rect 14734 26432 14740 26444
rect 14516 26404 14740 26432
rect 14516 26392 14522 26404
rect 14734 26392 14740 26404
rect 14792 26392 14798 26444
rect 14826 26392 14832 26444
rect 14884 26392 14890 26444
rect 15102 26392 15108 26444
rect 15160 26432 15166 26444
rect 16209 26435 16267 26441
rect 16209 26432 16221 26435
rect 15160 26404 16221 26432
rect 15160 26392 15166 26404
rect 16209 26401 16221 26404
rect 16255 26401 16267 26435
rect 16209 26395 16267 26401
rect 16758 26392 16764 26444
rect 16816 26392 16822 26444
rect 19426 26392 19432 26444
rect 19484 26392 19490 26444
rect 19705 26435 19763 26441
rect 19705 26401 19717 26435
rect 19751 26432 19763 26435
rect 20990 26432 20996 26444
rect 19751 26404 20996 26432
rect 19751 26401 19763 26404
rect 19705 26395 19763 26401
rect 20990 26392 20996 26404
rect 21048 26432 21054 26444
rect 21634 26432 21640 26444
rect 21048 26404 21640 26432
rect 21048 26392 21054 26404
rect 21634 26392 21640 26404
rect 21692 26392 21698 26444
rect 22370 26392 22376 26444
rect 22428 26432 22434 26444
rect 23201 26435 23259 26441
rect 23201 26432 23213 26435
rect 22428 26404 23213 26432
rect 22428 26392 22434 26404
rect 23201 26401 23213 26404
rect 23247 26401 23259 26435
rect 23201 26395 23259 26401
rect 9125 26367 9183 26373
rect 9125 26333 9137 26367
rect 9171 26333 9183 26367
rect 9125 26327 9183 26333
rect 9140 26296 9168 26327
rect 10962 26324 10968 26376
rect 11020 26364 11026 26376
rect 12710 26364 12716 26376
rect 11020 26336 12716 26364
rect 11020 26324 11026 26336
rect 12710 26324 12716 26336
rect 12768 26324 12774 26376
rect 14645 26367 14703 26373
rect 14645 26333 14657 26367
rect 14691 26333 14703 26367
rect 16942 26364 16948 26376
rect 14645 26327 14703 26333
rect 15856 26336 16948 26364
rect 9674 26296 9680 26308
rect 9140 26268 9680 26296
rect 9646 26256 9680 26268
rect 9732 26256 9738 26308
rect 11238 26296 11244 26308
rect 10626 26268 11244 26296
rect 11238 26256 11244 26268
rect 11296 26256 11302 26308
rect 11790 26256 11796 26308
rect 11848 26296 11854 26308
rect 14660 26296 14688 26327
rect 15856 26296 15884 26336
rect 16942 26324 16948 26336
rect 17000 26324 17006 26376
rect 23109 26367 23167 26373
rect 23109 26333 23121 26367
rect 23155 26364 23167 26367
rect 23290 26364 23296 26376
rect 23155 26336 23296 26364
rect 23155 26333 23167 26336
rect 23109 26327 23167 26333
rect 23290 26324 23296 26336
rect 23348 26324 23354 26376
rect 24026 26324 24032 26376
rect 24084 26324 24090 26376
rect 24949 26367 25007 26373
rect 24949 26333 24961 26367
rect 24995 26364 25007 26367
rect 25148 26364 25176 26540
rect 25222 26528 25228 26540
rect 25280 26528 25286 26580
rect 25590 26528 25596 26580
rect 25648 26568 25654 26580
rect 25866 26568 25872 26580
rect 25648 26540 25872 26568
rect 25648 26528 25654 26540
rect 25866 26528 25872 26540
rect 25924 26528 25930 26580
rect 25222 26392 25228 26444
rect 25280 26392 25286 26444
rect 25590 26364 25596 26376
rect 24995 26336 25596 26364
rect 24995 26333 25007 26336
rect 24949 26327 25007 26333
rect 25590 26324 25596 26336
rect 25648 26324 25654 26376
rect 11848 26268 14320 26296
rect 14660 26268 15884 26296
rect 11848 26256 11854 26268
rect 9646 26228 9674 26256
rect 10870 26228 10876 26240
rect 9646 26200 10876 26228
rect 10870 26188 10876 26200
rect 10928 26188 10934 26240
rect 14292 26237 14320 26268
rect 15930 26256 15936 26308
rect 15988 26296 15994 26308
rect 16025 26299 16083 26305
rect 16025 26296 16037 26299
rect 15988 26268 16037 26296
rect 15988 26256 15994 26268
rect 16025 26265 16037 26268
rect 16071 26265 16083 26299
rect 16025 26259 16083 26265
rect 16117 26299 16175 26305
rect 16117 26265 16129 26299
rect 16163 26296 16175 26299
rect 16298 26296 16304 26308
rect 16163 26268 16304 26296
rect 16163 26265 16175 26268
rect 16117 26259 16175 26265
rect 16298 26256 16304 26268
rect 16356 26296 16362 26308
rect 17129 26299 17187 26305
rect 17129 26296 17141 26299
rect 16356 26268 17141 26296
rect 16356 26256 16362 26268
rect 17129 26265 17141 26268
rect 17175 26296 17187 26299
rect 17402 26296 17408 26308
rect 17175 26268 17408 26296
rect 17175 26265 17187 26268
rect 17129 26259 17187 26265
rect 17402 26256 17408 26268
rect 17460 26256 17466 26308
rect 21082 26296 21088 26308
rect 20930 26268 21088 26296
rect 21082 26256 21088 26268
rect 21140 26296 21146 26308
rect 21453 26299 21511 26305
rect 21453 26296 21465 26299
rect 21140 26268 21465 26296
rect 21140 26256 21146 26268
rect 21453 26265 21465 26268
rect 21499 26296 21511 26299
rect 21818 26296 21824 26308
rect 21499 26268 21824 26296
rect 21499 26265 21511 26268
rect 21453 26259 21511 26265
rect 21818 26256 21824 26268
rect 21876 26256 21882 26308
rect 22373 26299 22431 26305
rect 22373 26265 22385 26299
rect 22419 26296 22431 26299
rect 22830 26296 22836 26308
rect 22419 26268 22836 26296
rect 22419 26265 22431 26268
rect 22373 26259 22431 26265
rect 22830 26256 22836 26268
rect 22888 26296 22894 26308
rect 23017 26299 23075 26305
rect 23017 26296 23029 26299
rect 22888 26268 23029 26296
rect 22888 26256 22894 26268
rect 23017 26265 23029 26268
rect 23063 26265 23075 26299
rect 23017 26259 23075 26265
rect 23474 26256 23480 26308
rect 23532 26296 23538 26308
rect 24578 26296 24584 26308
rect 23532 26268 24584 26296
rect 23532 26256 23538 26268
rect 24578 26256 24584 26268
rect 24636 26256 24642 26308
rect 25041 26299 25099 26305
rect 25041 26265 25053 26299
rect 25087 26296 25099 26299
rect 25130 26296 25136 26308
rect 25087 26268 25136 26296
rect 25087 26265 25099 26268
rect 25041 26259 25099 26265
rect 25130 26256 25136 26268
rect 25188 26256 25194 26308
rect 14277 26231 14335 26237
rect 14277 26197 14289 26231
rect 14323 26197 14335 26231
rect 14277 26191 14335 26197
rect 18233 26231 18291 26237
rect 18233 26197 18245 26231
rect 18279 26228 18291 26231
rect 18322 26228 18328 26240
rect 18279 26200 18328 26228
rect 18279 26197 18291 26200
rect 18233 26191 18291 26197
rect 18322 26188 18328 26200
rect 18380 26188 18386 26240
rect 1104 26138 25852 26160
rect 1104 26086 7950 26138
rect 8002 26086 8014 26138
rect 8066 26086 8078 26138
rect 8130 26086 8142 26138
rect 8194 26086 8206 26138
rect 8258 26086 17950 26138
rect 18002 26086 18014 26138
rect 18066 26086 18078 26138
rect 18130 26086 18142 26138
rect 18194 26086 18206 26138
rect 18258 26086 25852 26138
rect 1104 26064 25852 26086
rect 12618 25984 12624 26036
rect 12676 25984 12682 26036
rect 13814 25984 13820 26036
rect 13872 26024 13878 26036
rect 14829 26027 14887 26033
rect 14829 26024 14841 26027
rect 13872 25996 14841 26024
rect 13872 25984 13878 25996
rect 14829 25993 14841 25996
rect 14875 25993 14887 26027
rect 14829 25987 14887 25993
rect 15289 26027 15347 26033
rect 15289 25993 15301 26027
rect 15335 26024 15347 26027
rect 15335 25996 16160 26024
rect 15335 25993 15347 25996
rect 15289 25987 15347 25993
rect 9674 25916 9680 25968
rect 9732 25956 9738 25968
rect 9732 25928 14320 25956
rect 9732 25916 9738 25928
rect 12526 25848 12532 25900
rect 12584 25848 12590 25900
rect 13909 25891 13967 25897
rect 13909 25857 13921 25891
rect 13955 25888 13967 25891
rect 14182 25888 14188 25900
rect 13955 25860 14188 25888
rect 13955 25857 13967 25860
rect 13909 25851 13967 25857
rect 14182 25848 14188 25860
rect 14240 25848 14246 25900
rect 11054 25780 11060 25832
rect 11112 25820 11118 25832
rect 12713 25823 12771 25829
rect 11112 25792 12572 25820
rect 11112 25780 11118 25792
rect 12161 25755 12219 25761
rect 12161 25721 12173 25755
rect 12207 25752 12219 25755
rect 12544 25752 12572 25792
rect 12713 25789 12725 25823
rect 12759 25789 12771 25823
rect 12713 25783 12771 25789
rect 12728 25752 12756 25783
rect 13998 25780 14004 25832
rect 14056 25780 14062 25832
rect 14090 25780 14096 25832
rect 14148 25780 14154 25832
rect 14292 25820 14320 25928
rect 15197 25891 15255 25897
rect 15197 25857 15209 25891
rect 15243 25888 15255 25891
rect 16025 25891 16083 25897
rect 16025 25888 16037 25891
rect 15243 25860 16037 25888
rect 15243 25857 15255 25860
rect 15197 25851 15255 25857
rect 16025 25857 16037 25860
rect 16071 25857 16083 25891
rect 16025 25851 16083 25857
rect 15381 25823 15439 25829
rect 15381 25820 15393 25823
rect 14292 25792 15393 25820
rect 15381 25789 15393 25792
rect 15427 25789 15439 25823
rect 16132 25820 16160 25996
rect 16298 25984 16304 26036
rect 16356 26024 16362 26036
rect 17773 26027 17831 26033
rect 17773 26024 17785 26027
rect 16356 25996 17785 26024
rect 16356 25984 16362 25996
rect 17773 25993 17785 25996
rect 17819 25993 17831 26027
rect 17773 25987 17831 25993
rect 18141 26027 18199 26033
rect 18141 25993 18153 26027
rect 18187 26024 18199 26027
rect 18322 26024 18328 26036
rect 18187 25996 18328 26024
rect 18187 25993 18199 25996
rect 18141 25987 18199 25993
rect 18322 25984 18328 25996
rect 18380 25984 18386 26036
rect 19150 25984 19156 26036
rect 19208 26024 19214 26036
rect 22278 26024 22284 26036
rect 19208 25996 22284 26024
rect 19208 25984 19214 25996
rect 22278 25984 22284 25996
rect 22336 25984 22342 26036
rect 22465 26027 22523 26033
rect 22465 25993 22477 26027
rect 22511 26024 22523 26027
rect 22646 26024 22652 26036
rect 22511 25996 22652 26024
rect 22511 25993 22523 25996
rect 22465 25987 22523 25993
rect 22646 25984 22652 25996
rect 22704 25984 22710 26036
rect 25406 26024 25412 26036
rect 23400 25996 25412 26024
rect 18233 25959 18291 25965
rect 18233 25925 18245 25959
rect 18279 25956 18291 25959
rect 18414 25956 18420 25968
rect 18279 25928 18420 25956
rect 18279 25925 18291 25928
rect 18233 25919 18291 25925
rect 18414 25916 18420 25928
rect 18472 25916 18478 25968
rect 22373 25959 22431 25965
rect 22373 25956 22385 25959
rect 22066 25928 22385 25956
rect 16574 25848 16580 25900
rect 16632 25888 16638 25900
rect 17037 25891 17095 25897
rect 17037 25888 17049 25891
rect 16632 25860 17049 25888
rect 16632 25848 16638 25860
rect 17037 25857 17049 25860
rect 17083 25857 17095 25891
rect 17037 25851 17095 25857
rect 17405 25891 17463 25897
rect 17405 25857 17417 25891
rect 17451 25888 17463 25891
rect 17586 25888 17592 25900
rect 17451 25860 17592 25888
rect 17451 25857 17463 25860
rect 17405 25851 17463 25857
rect 17420 25820 17448 25851
rect 17586 25848 17592 25860
rect 17644 25888 17650 25900
rect 17644 25860 18828 25888
rect 17644 25848 17650 25860
rect 16132 25792 17448 25820
rect 18417 25823 18475 25829
rect 15381 25783 15439 25789
rect 18417 25789 18429 25823
rect 18463 25820 18475 25823
rect 18690 25820 18696 25832
rect 18463 25792 18696 25820
rect 18463 25789 18475 25792
rect 18417 25783 18475 25789
rect 18690 25780 18696 25792
rect 18748 25780 18754 25832
rect 18800 25820 18828 25860
rect 21450 25848 21456 25900
rect 21508 25888 21514 25900
rect 22066 25888 22094 25928
rect 22373 25925 22385 25928
rect 22419 25956 22431 25959
rect 23400 25956 23428 25996
rect 25406 25984 25412 25996
rect 25464 25984 25470 26036
rect 24854 25956 24860 25968
rect 22419 25928 23428 25956
rect 23492 25928 24860 25956
rect 22419 25925 22431 25928
rect 22373 25919 22431 25925
rect 23492 25897 23520 25928
rect 24854 25916 24860 25928
rect 24912 25916 24918 25968
rect 21508 25860 22094 25888
rect 23477 25891 23535 25897
rect 21508 25848 21514 25860
rect 23477 25857 23489 25891
rect 23523 25857 23535 25891
rect 23477 25851 23535 25857
rect 23934 25848 23940 25900
rect 23992 25848 23998 25900
rect 18800 25792 22508 25820
rect 12207 25724 12434 25752
rect 12544 25724 12756 25752
rect 13541 25755 13599 25761
rect 12207 25721 12219 25724
rect 12161 25715 12219 25721
rect 12406 25684 12434 25724
rect 13541 25721 13553 25755
rect 13587 25752 13599 25755
rect 17586 25752 17592 25764
rect 13587 25724 17592 25752
rect 13587 25721 13599 25724
rect 13541 25715 13599 25721
rect 17586 25712 17592 25724
rect 17644 25712 17650 25764
rect 19978 25712 19984 25764
rect 20036 25752 20042 25764
rect 22005 25755 22063 25761
rect 22005 25752 22017 25755
rect 20036 25724 22017 25752
rect 20036 25712 20042 25724
rect 22005 25721 22017 25724
rect 22051 25721 22063 25755
rect 22480 25752 22508 25792
rect 22554 25780 22560 25832
rect 22612 25780 22618 25832
rect 25130 25780 25136 25832
rect 25188 25780 25194 25832
rect 24762 25752 24768 25764
rect 22480 25724 24768 25752
rect 22005 25715 22063 25721
rect 24762 25712 24768 25724
rect 24820 25712 24826 25764
rect 16574 25684 16580 25696
rect 12406 25656 16580 25684
rect 16574 25644 16580 25656
rect 16632 25644 16638 25696
rect 16850 25644 16856 25696
rect 16908 25644 16914 25696
rect 18598 25644 18604 25696
rect 18656 25684 18662 25696
rect 19061 25687 19119 25693
rect 19061 25684 19073 25687
rect 18656 25656 19073 25684
rect 18656 25644 18662 25656
rect 19061 25653 19073 25656
rect 19107 25684 19119 25687
rect 19150 25684 19156 25696
rect 19107 25656 19156 25684
rect 19107 25653 19119 25656
rect 19061 25647 19119 25653
rect 19150 25644 19156 25656
rect 19208 25644 19214 25696
rect 21450 25644 21456 25696
rect 21508 25684 21514 25696
rect 21545 25687 21603 25693
rect 21545 25684 21557 25687
rect 21508 25656 21557 25684
rect 21508 25644 21514 25656
rect 21545 25653 21557 25656
rect 21591 25653 21603 25687
rect 21545 25647 21603 25653
rect 23290 25644 23296 25696
rect 23348 25644 23354 25696
rect 1104 25594 25852 25616
rect 1104 25542 2950 25594
rect 3002 25542 3014 25594
rect 3066 25542 3078 25594
rect 3130 25542 3142 25594
rect 3194 25542 3206 25594
rect 3258 25542 12950 25594
rect 13002 25542 13014 25594
rect 13066 25542 13078 25594
rect 13130 25542 13142 25594
rect 13194 25542 13206 25594
rect 13258 25542 22950 25594
rect 23002 25542 23014 25594
rect 23066 25542 23078 25594
rect 23130 25542 23142 25594
rect 23194 25542 23206 25594
rect 23258 25542 25852 25594
rect 1104 25520 25852 25542
rect 11698 25440 11704 25492
rect 11756 25480 11762 25492
rect 14277 25483 14335 25489
rect 14277 25480 14289 25483
rect 11756 25452 14289 25480
rect 11756 25440 11762 25452
rect 14277 25449 14289 25452
rect 14323 25449 14335 25483
rect 14277 25443 14335 25449
rect 15381 25483 15439 25489
rect 15381 25449 15393 25483
rect 15427 25480 15439 25483
rect 15562 25480 15568 25492
rect 15427 25452 15568 25480
rect 15427 25449 15439 25452
rect 15381 25443 15439 25449
rect 15562 25440 15568 25452
rect 15620 25440 15626 25492
rect 18141 25483 18199 25489
rect 18141 25480 18153 25483
rect 16592 25452 18153 25480
rect 12986 25372 12992 25424
rect 13044 25412 13050 25424
rect 13538 25412 13544 25424
rect 13044 25384 13544 25412
rect 13044 25372 13050 25384
rect 13538 25372 13544 25384
rect 13596 25372 13602 25424
rect 15102 25412 15108 25424
rect 14752 25384 15108 25412
rect 14752 25356 14780 25384
rect 15102 25372 15108 25384
rect 15160 25372 15166 25424
rect 10870 25304 10876 25356
rect 10928 25304 10934 25356
rect 11149 25347 11207 25353
rect 11149 25313 11161 25347
rect 11195 25344 11207 25347
rect 14734 25344 14740 25356
rect 11195 25316 14740 25344
rect 11195 25313 11207 25316
rect 11149 25307 11207 25313
rect 14734 25304 14740 25316
rect 14792 25304 14798 25356
rect 14826 25304 14832 25356
rect 14884 25304 14890 25356
rect 16301 25347 16359 25353
rect 16301 25344 16313 25347
rect 14936 25316 16313 25344
rect 13354 25236 13360 25288
rect 13412 25276 13418 25288
rect 14936 25276 14964 25316
rect 16301 25313 16313 25316
rect 16347 25313 16359 25347
rect 16301 25307 16359 25313
rect 13412 25248 14964 25276
rect 13412 25236 13418 25248
rect 12986 25208 12992 25220
rect 12374 25180 12992 25208
rect 12986 25168 12992 25180
rect 13044 25168 13050 25220
rect 14645 25211 14703 25217
rect 14645 25177 14657 25211
rect 14691 25208 14703 25211
rect 15562 25208 15568 25220
rect 14691 25180 15568 25208
rect 14691 25177 14703 25180
rect 14645 25171 14703 25177
rect 15562 25168 15568 25180
rect 15620 25168 15626 25220
rect 16117 25211 16175 25217
rect 16117 25177 16129 25211
rect 16163 25208 16175 25211
rect 16592 25208 16620 25452
rect 18141 25449 18153 25452
rect 18187 25480 18199 25483
rect 18506 25480 18512 25492
rect 18187 25452 18512 25480
rect 18187 25449 18199 25452
rect 18141 25443 18199 25449
rect 18506 25440 18512 25452
rect 18564 25480 18570 25492
rect 19245 25483 19303 25489
rect 19245 25480 19257 25483
rect 18564 25452 19257 25480
rect 18564 25440 18570 25452
rect 19245 25449 19257 25452
rect 19291 25480 19303 25483
rect 20070 25480 20076 25492
rect 19291 25452 20076 25480
rect 19291 25449 19303 25452
rect 19245 25443 19303 25449
rect 20070 25440 20076 25452
rect 20128 25440 20134 25492
rect 20809 25483 20867 25489
rect 20809 25449 20821 25483
rect 20855 25480 20867 25483
rect 21545 25483 21603 25489
rect 20855 25452 21496 25480
rect 20855 25449 20867 25452
rect 20809 25443 20867 25449
rect 16945 25415 17003 25421
rect 16945 25381 16957 25415
rect 16991 25412 17003 25415
rect 21468 25412 21496 25452
rect 21545 25449 21557 25483
rect 21591 25480 21603 25483
rect 23934 25480 23940 25492
rect 21591 25452 23940 25480
rect 21591 25449 21603 25452
rect 21545 25443 21603 25449
rect 23934 25440 23940 25452
rect 23992 25440 23998 25492
rect 24489 25483 24547 25489
rect 24489 25449 24501 25483
rect 24535 25480 24547 25483
rect 24854 25480 24860 25492
rect 24535 25452 24860 25480
rect 24535 25449 24547 25452
rect 24489 25443 24547 25449
rect 24854 25440 24860 25452
rect 24912 25440 24918 25492
rect 16991 25384 21404 25412
rect 21468 25384 22094 25412
rect 16991 25381 17003 25384
rect 16945 25375 17003 25381
rect 16850 25304 16856 25356
rect 16908 25344 16914 25356
rect 21376 25344 21404 25384
rect 16908 25316 21036 25344
rect 21376 25316 21772 25344
rect 16908 25304 16914 25316
rect 17126 25236 17132 25288
rect 17184 25236 17190 25288
rect 17586 25236 17592 25288
rect 17644 25276 17650 25288
rect 17773 25279 17831 25285
rect 17773 25276 17785 25279
rect 17644 25248 17785 25276
rect 17644 25236 17650 25248
rect 17773 25245 17785 25248
rect 17819 25245 17831 25279
rect 17773 25239 17831 25245
rect 18325 25279 18383 25285
rect 18325 25245 18337 25279
rect 18371 25276 18383 25279
rect 18598 25276 18604 25288
rect 18371 25248 18604 25276
rect 18371 25245 18383 25248
rect 18325 25239 18383 25245
rect 18598 25236 18604 25248
rect 18656 25236 18662 25288
rect 21008 25285 21036 25316
rect 21744 25285 21772 25316
rect 20993 25279 21051 25285
rect 20993 25245 21005 25279
rect 21039 25245 21051 25279
rect 20993 25239 21051 25245
rect 21729 25279 21787 25285
rect 21729 25245 21741 25279
rect 21775 25245 21787 25279
rect 22066 25276 22094 25384
rect 24026 25372 24032 25424
rect 24084 25412 24090 25424
rect 24581 25415 24639 25421
rect 24581 25412 24593 25415
rect 24084 25384 24593 25412
rect 24084 25372 24090 25384
rect 24581 25381 24593 25384
rect 24627 25381 24639 25415
rect 24581 25375 24639 25381
rect 22649 25279 22707 25285
rect 22649 25276 22661 25279
rect 22066 25248 22661 25276
rect 21729 25239 21787 25245
rect 22649 25245 22661 25248
rect 22695 25245 22707 25279
rect 22649 25239 22707 25245
rect 25314 25236 25320 25288
rect 25372 25236 25378 25288
rect 19150 25208 19156 25220
rect 16163 25180 16620 25208
rect 17604 25180 19156 25208
rect 16163 25177 16175 25180
rect 16117 25171 16175 25177
rect 12618 25100 12624 25152
rect 12676 25100 12682 25152
rect 14737 25143 14795 25149
rect 14737 25109 14749 25143
rect 14783 25140 14795 25143
rect 15378 25140 15384 25152
rect 14783 25112 15384 25140
rect 14783 25109 14795 25112
rect 14737 25103 14795 25109
rect 15378 25100 15384 25112
rect 15436 25100 15442 25152
rect 15746 25100 15752 25152
rect 15804 25100 15810 25152
rect 16206 25100 16212 25152
rect 16264 25100 16270 25152
rect 17604 25149 17632 25180
rect 19150 25168 19156 25180
rect 19208 25168 19214 25220
rect 19797 25211 19855 25217
rect 19797 25177 19809 25211
rect 19843 25208 19855 25211
rect 19843 25180 20392 25208
rect 19843 25177 19855 25180
rect 19797 25171 19855 25177
rect 17589 25143 17647 25149
rect 17589 25109 17601 25143
rect 17635 25109 17647 25143
rect 17589 25103 17647 25109
rect 18506 25100 18512 25152
rect 18564 25140 18570 25152
rect 18693 25143 18751 25149
rect 18693 25140 18705 25143
rect 18564 25112 18705 25140
rect 18564 25100 18570 25112
rect 18693 25109 18705 25112
rect 18739 25109 18751 25143
rect 18693 25103 18751 25109
rect 19886 25100 19892 25152
rect 19944 25100 19950 25152
rect 20364 25149 20392 25180
rect 23842 25168 23848 25220
rect 23900 25168 23906 25220
rect 24857 25211 24915 25217
rect 24857 25177 24869 25211
rect 24903 25208 24915 25211
rect 25406 25208 25412 25220
rect 24903 25180 25412 25208
rect 24903 25177 24915 25180
rect 24857 25171 24915 25177
rect 25406 25168 25412 25180
rect 25464 25168 25470 25220
rect 20349 25143 20407 25149
rect 20349 25109 20361 25143
rect 20395 25140 20407 25143
rect 23750 25140 23756 25152
rect 20395 25112 23756 25140
rect 20395 25109 20407 25112
rect 20349 25103 20407 25109
rect 23750 25100 23756 25112
rect 23808 25100 23814 25152
rect 25130 25100 25136 25152
rect 25188 25100 25194 25152
rect 1104 25050 25852 25072
rect 1104 24998 7950 25050
rect 8002 24998 8014 25050
rect 8066 24998 8078 25050
rect 8130 24998 8142 25050
rect 8194 24998 8206 25050
rect 8258 24998 17950 25050
rect 18002 24998 18014 25050
rect 18066 24998 18078 25050
rect 18130 24998 18142 25050
rect 18194 24998 18206 25050
rect 18258 24998 25852 25050
rect 1104 24976 25852 24998
rect 17126 24936 17132 24948
rect 15212 24908 17132 24936
rect 10134 24828 10140 24880
rect 10192 24828 10198 24880
rect 11238 24828 11244 24880
rect 11296 24868 11302 24880
rect 12069 24871 12127 24877
rect 12069 24868 12081 24871
rect 11296 24840 12081 24868
rect 11296 24828 11302 24840
rect 12069 24837 12081 24840
rect 12115 24837 12127 24871
rect 12069 24831 12127 24837
rect 13538 24828 13544 24880
rect 13596 24868 13602 24880
rect 13596 24840 13754 24868
rect 13596 24828 13602 24840
rect 12161 24803 12219 24809
rect 12161 24769 12173 24803
rect 12207 24800 12219 24803
rect 12250 24800 12256 24812
rect 12207 24772 12256 24800
rect 12207 24769 12219 24772
rect 12161 24763 12219 24769
rect 12250 24760 12256 24772
rect 12308 24760 12314 24812
rect 12710 24760 12716 24812
rect 12768 24800 12774 24812
rect 12989 24803 13047 24809
rect 12989 24800 13001 24803
rect 12768 24772 13001 24800
rect 12768 24760 12774 24772
rect 12989 24769 13001 24772
rect 13035 24769 13047 24803
rect 15212 24800 15240 24908
rect 17126 24896 17132 24908
rect 17184 24896 17190 24948
rect 17218 24896 17224 24948
rect 17276 24936 17282 24948
rect 18322 24936 18328 24948
rect 17276 24908 18328 24936
rect 17276 24896 17282 24908
rect 18322 24896 18328 24908
rect 18380 24936 18386 24948
rect 19061 24939 19119 24945
rect 19061 24936 19073 24939
rect 18380 24908 19073 24936
rect 18380 24896 18386 24908
rect 19061 24905 19073 24908
rect 19107 24905 19119 24939
rect 19061 24899 19119 24905
rect 16206 24828 16212 24880
rect 16264 24868 16270 24880
rect 18509 24871 18567 24877
rect 18509 24868 18521 24871
rect 16264 24840 18521 24868
rect 16264 24828 16270 24840
rect 18509 24837 18521 24840
rect 18555 24868 18567 24871
rect 18598 24868 18604 24880
rect 18555 24840 18604 24868
rect 18555 24837 18567 24840
rect 18509 24831 18567 24837
rect 18598 24828 18604 24840
rect 18656 24828 18662 24880
rect 22465 24871 22523 24877
rect 22465 24837 22477 24871
rect 22511 24868 22523 24871
rect 24118 24868 24124 24880
rect 22511 24840 24124 24868
rect 22511 24837 22523 24840
rect 22465 24831 22523 24837
rect 24118 24828 24124 24840
rect 24176 24828 24182 24880
rect 25406 24868 25412 24880
rect 25070 24840 25412 24868
rect 25406 24828 25412 24840
rect 25464 24828 25470 24880
rect 12989 24763 13047 24769
rect 14568 24772 15240 24800
rect 9401 24735 9459 24741
rect 9401 24701 9413 24735
rect 9447 24701 9459 24735
rect 9401 24695 9459 24701
rect 9677 24735 9735 24741
rect 9677 24701 9689 24735
rect 9723 24732 9735 24735
rect 11146 24732 11152 24744
rect 9723 24704 11152 24732
rect 9723 24701 9735 24704
rect 9677 24695 9735 24701
rect 9416 24596 9444 24695
rect 11146 24692 11152 24704
rect 11204 24692 11210 24744
rect 12342 24692 12348 24744
rect 12400 24692 12406 24744
rect 13265 24735 13323 24741
rect 13265 24701 13277 24735
rect 13311 24732 13323 24735
rect 13906 24732 13912 24744
rect 13311 24704 13912 24732
rect 13311 24701 13323 24704
rect 13265 24695 13323 24701
rect 13906 24692 13912 24704
rect 13964 24692 13970 24744
rect 10870 24624 10876 24676
rect 10928 24664 10934 24676
rect 10928 24636 11192 24664
rect 10928 24624 10934 24636
rect 11054 24596 11060 24608
rect 9416 24568 11060 24596
rect 11054 24556 11060 24568
rect 11112 24556 11118 24608
rect 11164 24605 11192 24636
rect 11149 24599 11207 24605
rect 11149 24565 11161 24599
rect 11195 24565 11207 24599
rect 11149 24559 11207 24565
rect 11701 24599 11759 24605
rect 11701 24565 11713 24599
rect 11747 24596 11759 24599
rect 14568 24596 14596 24772
rect 15378 24760 15384 24812
rect 15436 24800 15442 24812
rect 16390 24800 16396 24812
rect 15436 24772 16396 24800
rect 15436 24760 15442 24772
rect 16390 24760 16396 24772
rect 16448 24800 16454 24812
rect 17313 24803 17371 24809
rect 17313 24800 17325 24803
rect 16448 24772 17325 24800
rect 16448 24760 16454 24772
rect 17313 24769 17325 24772
rect 17359 24800 17371 24803
rect 17359 24772 17908 24800
rect 17359 24769 17371 24772
rect 17313 24763 17371 24769
rect 14734 24692 14740 24744
rect 14792 24692 14798 24744
rect 15010 24692 15016 24744
rect 15068 24732 15074 24744
rect 17405 24735 17463 24741
rect 17405 24732 17417 24735
rect 15068 24704 17417 24732
rect 15068 24692 15074 24704
rect 17405 24701 17417 24704
rect 17451 24701 17463 24735
rect 17880 24732 17908 24772
rect 18414 24760 18420 24812
rect 18472 24760 18478 24812
rect 18690 24800 18696 24812
rect 18524 24772 18696 24800
rect 18524 24732 18552 24772
rect 18690 24760 18696 24772
rect 18748 24800 18754 24812
rect 19337 24803 19395 24809
rect 19337 24800 19349 24803
rect 18748 24772 19349 24800
rect 18748 24760 18754 24772
rect 19337 24769 19349 24772
rect 19383 24769 19395 24803
rect 19337 24763 19395 24769
rect 19426 24760 19432 24812
rect 19484 24800 19490 24812
rect 19705 24803 19763 24809
rect 19705 24800 19717 24803
rect 19484 24772 19717 24800
rect 19484 24760 19490 24772
rect 19705 24769 19717 24772
rect 19751 24769 19763 24803
rect 19705 24763 19763 24769
rect 21082 24760 21088 24812
rect 21140 24760 21146 24812
rect 22557 24803 22615 24809
rect 22557 24769 22569 24803
rect 22603 24800 22615 24803
rect 23474 24800 23480 24812
rect 22603 24772 23480 24800
rect 22603 24769 22615 24772
rect 22557 24763 22615 24769
rect 23474 24760 23480 24772
rect 23532 24760 23538 24812
rect 17880 24704 18552 24732
rect 18601 24735 18659 24741
rect 17405 24695 17463 24701
rect 18601 24701 18613 24735
rect 18647 24701 18659 24735
rect 18601 24695 18659 24701
rect 19981 24735 20039 24741
rect 19981 24701 19993 24735
rect 20027 24732 20039 24735
rect 20438 24732 20444 24744
rect 20027 24704 20444 24732
rect 20027 24701 20039 24704
rect 19981 24695 20039 24701
rect 17034 24624 17040 24676
rect 17092 24664 17098 24676
rect 18616 24664 18644 24695
rect 20438 24692 20444 24704
rect 20496 24692 20502 24744
rect 21453 24735 21511 24741
rect 21453 24701 21465 24735
rect 21499 24732 21511 24735
rect 22370 24732 22376 24744
rect 21499 24704 22376 24732
rect 21499 24701 21511 24704
rect 21453 24695 21511 24701
rect 22370 24692 22376 24704
rect 22428 24692 22434 24744
rect 22646 24692 22652 24744
rect 22704 24692 22710 24744
rect 23569 24735 23627 24741
rect 23569 24701 23581 24735
rect 23615 24701 23627 24735
rect 23569 24695 23627 24701
rect 23845 24735 23903 24741
rect 23845 24701 23857 24735
rect 23891 24732 23903 24735
rect 25222 24732 25228 24744
rect 23891 24704 25228 24732
rect 23891 24701 23903 24704
rect 23845 24695 23903 24701
rect 17092 24636 18644 24664
rect 17092 24624 17098 24636
rect 22186 24624 22192 24676
rect 22244 24664 22250 24676
rect 23382 24664 23388 24676
rect 22244 24636 23388 24664
rect 22244 24624 22250 24636
rect 23382 24624 23388 24636
rect 23440 24664 23446 24676
rect 23584 24664 23612 24695
rect 25222 24692 25228 24704
rect 25280 24692 25286 24744
rect 25317 24735 25375 24741
rect 25317 24701 25329 24735
rect 25363 24732 25375 24735
rect 25498 24732 25504 24744
rect 25363 24704 25504 24732
rect 25363 24701 25375 24704
rect 25317 24695 25375 24701
rect 25498 24692 25504 24704
rect 25556 24692 25562 24744
rect 23440 24636 23612 24664
rect 23440 24624 23446 24636
rect 11747 24568 14596 24596
rect 11747 24565 11759 24568
rect 11701 24559 11759 24565
rect 14734 24556 14740 24608
rect 14792 24596 14798 24608
rect 15013 24599 15071 24605
rect 15013 24596 15025 24599
rect 14792 24568 15025 24596
rect 14792 24556 14798 24568
rect 15013 24565 15025 24568
rect 15059 24565 15071 24599
rect 15013 24559 15071 24565
rect 15470 24556 15476 24608
rect 15528 24596 15534 24608
rect 16853 24599 16911 24605
rect 16853 24596 16865 24599
rect 15528 24568 16865 24596
rect 15528 24556 15534 24568
rect 16853 24565 16865 24568
rect 16899 24565 16911 24599
rect 16853 24559 16911 24565
rect 17862 24556 17868 24608
rect 17920 24596 17926 24608
rect 18049 24599 18107 24605
rect 18049 24596 18061 24599
rect 17920 24568 18061 24596
rect 17920 24556 17926 24568
rect 18049 24565 18061 24568
rect 18095 24565 18107 24599
rect 18049 24559 18107 24565
rect 22097 24599 22155 24605
rect 22097 24565 22109 24599
rect 22143 24596 22155 24599
rect 22370 24596 22376 24608
rect 22143 24568 22376 24596
rect 22143 24565 22155 24568
rect 22097 24559 22155 24565
rect 22370 24556 22376 24568
rect 22428 24556 22434 24608
rect 1104 24506 25852 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 25852 24506
rect 1104 24432 25852 24454
rect 10870 24352 10876 24404
rect 10928 24392 10934 24404
rect 14826 24392 14832 24404
rect 10928 24364 14832 24392
rect 10928 24352 10934 24364
rect 14826 24352 14832 24364
rect 14884 24352 14890 24404
rect 20438 24352 20444 24404
rect 20496 24392 20502 24404
rect 21177 24395 21235 24401
rect 21177 24392 21189 24395
rect 20496 24364 21189 24392
rect 20496 24352 20502 24364
rect 21177 24361 21189 24364
rect 21223 24361 21235 24395
rect 21177 24355 21235 24361
rect 25314 24352 25320 24404
rect 25372 24352 25378 24404
rect 13538 24284 13544 24336
rect 13596 24324 13602 24336
rect 14185 24327 14243 24333
rect 14185 24324 14197 24327
rect 13596 24296 14197 24324
rect 13596 24284 13602 24296
rect 14185 24293 14197 24296
rect 14231 24324 14243 24327
rect 14734 24324 14740 24336
rect 14231 24296 14740 24324
rect 14231 24293 14243 24296
rect 14185 24287 14243 24293
rect 14734 24284 14740 24296
rect 14792 24284 14798 24336
rect 25133 24327 25191 24333
rect 25133 24293 25145 24327
rect 25179 24324 25191 24327
rect 25590 24324 25596 24336
rect 25179 24296 25596 24324
rect 25179 24293 25191 24296
rect 25133 24287 25191 24293
rect 25590 24284 25596 24296
rect 25648 24284 25654 24336
rect 10134 24216 10140 24268
rect 10192 24256 10198 24268
rect 10192 24228 11008 24256
rect 10192 24216 10198 24228
rect 7834 24148 7840 24200
rect 7892 24188 7898 24200
rect 9125 24191 9183 24197
rect 9125 24188 9137 24191
rect 7892 24160 9137 24188
rect 7892 24148 7898 24160
rect 9125 24157 9137 24160
rect 9171 24157 9183 24191
rect 10980 24188 11008 24228
rect 11054 24216 11060 24268
rect 11112 24256 11118 24268
rect 11977 24259 12035 24265
rect 11977 24256 11989 24259
rect 11112 24228 11989 24256
rect 11112 24216 11118 24228
rect 11977 24225 11989 24228
rect 12023 24256 12035 24259
rect 12342 24256 12348 24268
rect 12023 24228 12348 24256
rect 12023 24225 12035 24228
rect 11977 24219 12035 24225
rect 12342 24216 12348 24228
rect 12400 24216 12406 24268
rect 11241 24191 11299 24197
rect 11241 24188 11253 24191
rect 10980 24160 11253 24188
rect 9125 24151 9183 24157
rect 11241 24157 11253 24160
rect 11287 24188 11299 24191
rect 11425 24191 11483 24197
rect 11425 24188 11437 24191
rect 11287 24160 11437 24188
rect 11287 24157 11299 24160
rect 11241 24151 11299 24157
rect 11425 24157 11437 24160
rect 11471 24157 11483 24191
rect 13556 24188 13584 24284
rect 18785 24259 18843 24265
rect 18785 24225 18797 24259
rect 18831 24256 18843 24259
rect 18966 24256 18972 24268
rect 18831 24228 18972 24256
rect 18831 24225 18843 24228
rect 18785 24219 18843 24225
rect 18966 24216 18972 24228
rect 19024 24216 19030 24268
rect 19426 24216 19432 24268
rect 19484 24216 19490 24268
rect 21913 24259 21971 24265
rect 21913 24225 21925 24259
rect 21959 24256 21971 24259
rect 22186 24256 22192 24268
rect 21959 24228 22192 24256
rect 21959 24225 21971 24228
rect 21913 24219 21971 24225
rect 22186 24216 22192 24228
rect 22244 24216 22250 24268
rect 24118 24216 24124 24268
rect 24176 24256 24182 24268
rect 24581 24259 24639 24265
rect 24581 24256 24593 24259
rect 24176 24228 24593 24256
rect 24176 24216 24182 24228
rect 24581 24225 24593 24228
rect 24627 24225 24639 24259
rect 24581 24219 24639 24225
rect 13386 24160 13584 24188
rect 11425 24151 11483 24157
rect 17678 24148 17684 24200
rect 17736 24148 17742 24200
rect 18506 24148 18512 24200
rect 18564 24148 18570 24200
rect 9306 24080 9312 24132
rect 9364 24120 9370 24132
rect 9401 24123 9459 24129
rect 9401 24120 9413 24123
rect 9364 24092 9413 24120
rect 9364 24080 9370 24092
rect 9401 24089 9413 24092
rect 9447 24089 9459 24123
rect 9401 24083 9459 24089
rect 9416 24052 9444 24083
rect 10134 24080 10140 24132
rect 10192 24080 10198 24132
rect 10796 24092 11928 24120
rect 10796 24052 10824 24092
rect 9416 24024 10824 24052
rect 10873 24055 10931 24061
rect 10873 24021 10885 24055
rect 10919 24052 10931 24055
rect 11054 24052 11060 24064
rect 10919 24024 11060 24052
rect 10919 24021 10931 24024
rect 10873 24015 10931 24021
rect 11054 24012 11060 24024
rect 11112 24012 11118 24064
rect 11900 24052 11928 24092
rect 11974 24080 11980 24132
rect 12032 24120 12038 24132
rect 12253 24123 12311 24129
rect 12253 24120 12265 24123
rect 12032 24092 12265 24120
rect 12032 24080 12038 24092
rect 12253 24089 12265 24092
rect 12299 24089 12311 24123
rect 12253 24083 12311 24089
rect 15933 24123 15991 24129
rect 15933 24089 15945 24123
rect 15979 24120 15991 24123
rect 18874 24120 18880 24132
rect 15979 24092 18880 24120
rect 15979 24089 15991 24092
rect 15933 24083 15991 24089
rect 18874 24080 18880 24092
rect 18932 24080 18938 24132
rect 19702 24080 19708 24132
rect 19760 24080 19766 24132
rect 21082 24120 21088 24132
rect 20930 24092 21088 24120
rect 21082 24080 21088 24092
rect 21140 24120 21146 24132
rect 22189 24123 22247 24129
rect 21140 24092 21588 24120
rect 21140 24080 21146 24092
rect 21560 24064 21588 24092
rect 22189 24089 22201 24123
rect 22235 24120 22247 24123
rect 22278 24120 22284 24132
rect 22235 24092 22284 24120
rect 22235 24089 22247 24092
rect 22189 24083 22247 24089
rect 22278 24080 22284 24092
rect 22336 24080 22342 24132
rect 23414 24092 23980 24120
rect 12618 24052 12624 24064
rect 11900 24024 12624 24052
rect 12618 24012 12624 24024
rect 12676 24052 12682 24064
rect 12894 24052 12900 24064
rect 12676 24024 12900 24052
rect 12676 24012 12682 24024
rect 12894 24012 12900 24024
rect 12952 24012 12958 24064
rect 13725 24055 13783 24061
rect 13725 24021 13737 24055
rect 13771 24052 13783 24055
rect 13906 24052 13912 24064
rect 13771 24024 13912 24052
rect 13771 24021 13783 24024
rect 13725 24015 13783 24021
rect 13906 24012 13912 24024
rect 13964 24012 13970 24064
rect 18141 24055 18199 24061
rect 18141 24021 18153 24055
rect 18187 24052 18199 24055
rect 18414 24052 18420 24064
rect 18187 24024 18420 24052
rect 18187 24021 18199 24024
rect 18141 24015 18199 24021
rect 18414 24012 18420 24024
rect 18472 24012 18478 24064
rect 18601 24055 18659 24061
rect 18601 24021 18613 24055
rect 18647 24052 18659 24055
rect 20714 24052 20720 24064
rect 18647 24024 20720 24052
rect 18647 24021 18659 24024
rect 18601 24015 18659 24021
rect 20714 24012 20720 24024
rect 20772 24012 20778 24064
rect 21542 24012 21548 24064
rect 21600 24012 21606 24064
rect 23566 24012 23572 24064
rect 23624 24052 23630 24064
rect 23952 24061 23980 24092
rect 23661 24055 23719 24061
rect 23661 24052 23673 24055
rect 23624 24024 23673 24052
rect 23624 24012 23630 24024
rect 23661 24021 23673 24024
rect 23707 24021 23719 24055
rect 23661 24015 23719 24021
rect 23937 24055 23995 24061
rect 23937 24021 23949 24055
rect 23983 24052 23995 24055
rect 25314 24052 25320 24064
rect 23983 24024 25320 24052
rect 23983 24021 23995 24024
rect 23937 24015 23995 24021
rect 25314 24012 25320 24024
rect 25372 24052 25378 24064
rect 25409 24055 25467 24061
rect 25409 24052 25421 24055
rect 25372 24024 25421 24052
rect 25372 24012 25378 24024
rect 25409 24021 25421 24024
rect 25455 24021 25467 24055
rect 25409 24015 25467 24021
rect 1104 23962 25852 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 25852 23962
rect 1104 23888 25852 23910
rect 9766 23808 9772 23860
rect 9824 23808 9830 23860
rect 10318 23808 10324 23860
rect 10376 23848 10382 23860
rect 10413 23851 10471 23857
rect 10413 23848 10425 23851
rect 10376 23820 10425 23848
rect 10376 23808 10382 23820
rect 10413 23817 10425 23820
rect 10459 23817 10471 23851
rect 10413 23811 10471 23817
rect 10781 23851 10839 23857
rect 10781 23817 10793 23851
rect 10827 23848 10839 23851
rect 13814 23848 13820 23860
rect 10827 23820 13820 23848
rect 10827 23817 10839 23820
rect 10781 23811 10839 23817
rect 13814 23808 13820 23820
rect 13872 23808 13878 23860
rect 14461 23851 14519 23857
rect 14461 23817 14473 23851
rect 14507 23817 14519 23851
rect 14461 23811 14519 23817
rect 9784 23780 9812 23808
rect 9784 23752 11008 23780
rect 7834 23672 7840 23724
rect 7892 23712 7898 23724
rect 8021 23715 8079 23721
rect 8021 23712 8033 23715
rect 7892 23684 8033 23712
rect 7892 23672 7898 23684
rect 8021 23681 8033 23684
rect 8067 23681 8079 23715
rect 9430 23684 9996 23712
rect 8021 23675 8079 23681
rect 8297 23647 8355 23653
rect 8297 23613 8309 23647
rect 8343 23644 8355 23647
rect 9674 23644 9680 23656
rect 8343 23616 9680 23644
rect 8343 23613 8355 23616
rect 8297 23607 8355 23613
rect 9674 23604 9680 23616
rect 9732 23604 9738 23656
rect 9968 23576 9996 23684
rect 10980 23656 11008 23752
rect 13630 23740 13636 23792
rect 13688 23740 13694 23792
rect 13722 23740 13728 23792
rect 13780 23740 13786 23792
rect 14476 23780 14504 23811
rect 14918 23808 14924 23860
rect 14976 23808 14982 23860
rect 16758 23808 16764 23860
rect 16816 23848 16822 23860
rect 17221 23851 17279 23857
rect 17221 23848 17233 23851
rect 16816 23820 17233 23848
rect 16816 23808 16822 23820
rect 17221 23817 17233 23820
rect 17267 23848 17279 23851
rect 18138 23848 18144 23860
rect 17267 23820 18144 23848
rect 17267 23817 17279 23820
rect 17221 23811 17279 23817
rect 18138 23808 18144 23820
rect 18196 23808 18202 23860
rect 18230 23808 18236 23860
rect 18288 23848 18294 23860
rect 18690 23848 18696 23860
rect 18288 23820 18696 23848
rect 18288 23808 18294 23820
rect 18690 23808 18696 23820
rect 18748 23808 18754 23860
rect 18874 23808 18880 23860
rect 18932 23808 18938 23860
rect 19150 23808 19156 23860
rect 19208 23848 19214 23860
rect 24949 23851 25007 23857
rect 19208 23820 22692 23848
rect 19208 23808 19214 23820
rect 14476 23752 18276 23780
rect 13998 23672 14004 23724
rect 14056 23712 14062 23724
rect 14829 23715 14887 23721
rect 14829 23712 14841 23715
rect 14056 23684 14841 23712
rect 14056 23672 14062 23684
rect 14829 23681 14841 23684
rect 14875 23681 14887 23715
rect 14829 23675 14887 23681
rect 17310 23672 17316 23724
rect 17368 23712 17374 23724
rect 18248 23721 18276 23752
rect 19702 23740 19708 23792
rect 19760 23780 19766 23792
rect 22554 23780 22560 23792
rect 19760 23752 20944 23780
rect 19760 23740 19766 23752
rect 18233 23715 18291 23721
rect 17368 23684 17540 23712
rect 17368 23672 17374 23684
rect 10042 23604 10048 23656
rect 10100 23644 10106 23656
rect 10873 23647 10931 23653
rect 10873 23644 10885 23647
rect 10100 23616 10885 23644
rect 10100 23604 10106 23616
rect 10873 23613 10885 23616
rect 10919 23613 10931 23647
rect 10873 23607 10931 23613
rect 10962 23604 10968 23656
rect 11020 23604 11026 23656
rect 13817 23647 13875 23653
rect 13817 23613 13829 23647
rect 13863 23613 13875 23647
rect 13817 23607 13875 23613
rect 9968 23548 10180 23576
rect 10152 23520 10180 23548
rect 12894 23536 12900 23588
rect 12952 23576 12958 23588
rect 13832 23576 13860 23607
rect 13906 23604 13912 23656
rect 13964 23644 13970 23656
rect 15013 23647 15071 23653
rect 15013 23644 15025 23647
rect 13964 23616 15025 23644
rect 13964 23604 13970 23616
rect 15013 23613 15025 23616
rect 15059 23613 15071 23647
rect 15013 23607 15071 23613
rect 15654 23604 15660 23656
rect 15712 23604 15718 23656
rect 16574 23604 16580 23656
rect 16632 23644 16638 23656
rect 17328 23644 17356 23672
rect 16632 23616 17356 23644
rect 17405 23647 17463 23653
rect 16632 23604 16638 23616
rect 17405 23613 17417 23647
rect 17451 23613 17463 23647
rect 17512 23644 17540 23684
rect 18233 23681 18245 23715
rect 18279 23681 18291 23715
rect 18233 23675 18291 23681
rect 19610 23672 19616 23724
rect 19668 23672 19674 23724
rect 19904 23712 20024 23716
rect 20162 23712 20168 23724
rect 19720 23688 20168 23712
rect 19720 23684 19932 23688
rect 19996 23684 20168 23688
rect 19720 23656 19748 23684
rect 20162 23672 20168 23684
rect 20220 23672 20226 23724
rect 18785 23647 18843 23653
rect 18785 23644 18797 23647
rect 17512 23616 18797 23644
rect 17405 23607 17463 23613
rect 18785 23613 18797 23616
rect 18831 23644 18843 23647
rect 19334 23644 19340 23656
rect 18831 23616 19340 23644
rect 18831 23613 18843 23616
rect 18785 23607 18843 23613
rect 12952 23548 13860 23576
rect 12952 23536 12958 23548
rect 14550 23536 14556 23588
rect 14608 23576 14614 23588
rect 17420 23576 17448 23607
rect 19334 23604 19340 23616
rect 19392 23604 19398 23656
rect 19702 23604 19708 23656
rect 19760 23604 19766 23656
rect 19889 23647 19947 23653
rect 19889 23613 19901 23647
rect 19935 23644 19947 23647
rect 20548 23644 20576 23752
rect 20806 23672 20812 23724
rect 20864 23672 20870 23724
rect 20916 23712 20944 23752
rect 22296 23752 22560 23780
rect 22296 23724 22324 23752
rect 22554 23740 22560 23752
rect 22612 23740 22618 23792
rect 22278 23712 22284 23724
rect 20916 23684 22284 23712
rect 22278 23672 22284 23684
rect 22336 23672 22342 23724
rect 22373 23715 22431 23721
rect 22373 23681 22385 23715
rect 22419 23712 22431 23715
rect 22664 23712 22692 23820
rect 24949 23817 24961 23851
rect 24995 23848 25007 23851
rect 25222 23848 25228 23860
rect 24995 23820 25228 23848
rect 24995 23817 25007 23820
rect 24949 23811 25007 23817
rect 25222 23808 25228 23820
rect 25280 23808 25286 23860
rect 25501 23851 25559 23857
rect 25501 23817 25513 23851
rect 25547 23848 25559 23851
rect 25590 23848 25596 23860
rect 25547 23820 25596 23848
rect 25547 23817 25559 23820
rect 25501 23811 25559 23817
rect 25590 23808 25596 23820
rect 25648 23808 25654 23860
rect 25222 23712 25228 23724
rect 22419 23684 22692 23712
rect 24610 23684 25228 23712
rect 22419 23681 22431 23684
rect 22373 23675 22431 23681
rect 25222 23672 25228 23684
rect 25280 23672 25286 23724
rect 19935 23616 20576 23644
rect 19935 23613 19947 23616
rect 19889 23607 19947 23613
rect 20898 23604 20904 23656
rect 20956 23604 20962 23656
rect 20990 23604 20996 23656
rect 21048 23604 21054 23656
rect 22186 23604 22192 23656
rect 22244 23644 22250 23656
rect 23201 23647 23259 23653
rect 23201 23644 23213 23647
rect 22244 23616 23213 23644
rect 22244 23604 22250 23616
rect 23201 23613 23213 23616
rect 23247 23613 23259 23647
rect 23201 23607 23259 23613
rect 23477 23647 23535 23653
rect 23477 23613 23489 23647
rect 23523 23644 23535 23647
rect 23566 23644 23572 23656
rect 23523 23616 23572 23644
rect 23523 23613 23535 23616
rect 23477 23607 23535 23613
rect 23566 23604 23572 23616
rect 23624 23604 23630 23656
rect 14608 23548 17448 23576
rect 18049 23579 18107 23585
rect 14608 23536 14614 23548
rect 18049 23545 18061 23579
rect 18095 23576 18107 23579
rect 18095 23548 23060 23576
rect 18095 23545 18107 23548
rect 18049 23539 18107 23545
rect 10134 23468 10140 23520
rect 10192 23468 10198 23520
rect 12434 23468 12440 23520
rect 12492 23508 12498 23520
rect 13265 23511 13323 23517
rect 13265 23508 13277 23511
rect 12492 23480 13277 23508
rect 12492 23468 12498 23480
rect 13265 23477 13277 23480
rect 13311 23477 13323 23511
rect 13265 23471 13323 23477
rect 16853 23511 16911 23517
rect 16853 23477 16865 23511
rect 16899 23508 16911 23511
rect 17310 23508 17316 23520
rect 16899 23480 17316 23508
rect 16899 23477 16911 23480
rect 16853 23471 16911 23477
rect 17310 23468 17316 23480
rect 17368 23468 17374 23520
rect 18138 23468 18144 23520
rect 18196 23508 18202 23520
rect 18509 23511 18567 23517
rect 18509 23508 18521 23511
rect 18196 23480 18521 23508
rect 18196 23468 18202 23480
rect 18509 23477 18521 23480
rect 18555 23508 18567 23511
rect 19150 23508 19156 23520
rect 18555 23480 19156 23508
rect 18555 23477 18567 23480
rect 18509 23471 18567 23477
rect 19150 23468 19156 23480
rect 19208 23468 19214 23520
rect 19242 23468 19248 23520
rect 19300 23468 19306 23520
rect 19334 23468 19340 23520
rect 19392 23508 19398 23520
rect 20254 23508 20260 23520
rect 19392 23480 20260 23508
rect 19392 23468 19398 23480
rect 20254 23468 20260 23480
rect 20312 23468 20318 23520
rect 20441 23511 20499 23517
rect 20441 23477 20453 23511
rect 20487 23508 20499 23511
rect 20622 23508 20628 23520
rect 20487 23480 20628 23508
rect 20487 23477 20499 23480
rect 20441 23471 20499 23477
rect 20622 23468 20628 23480
rect 20680 23468 20686 23520
rect 21542 23468 21548 23520
rect 21600 23468 21606 23520
rect 22189 23511 22247 23517
rect 22189 23477 22201 23511
rect 22235 23508 22247 23511
rect 22830 23508 22836 23520
rect 22235 23480 22836 23508
rect 22235 23477 22247 23480
rect 22189 23471 22247 23477
rect 22830 23468 22836 23480
rect 22888 23468 22894 23520
rect 23032 23508 23060 23548
rect 23934 23508 23940 23520
rect 23032 23480 23940 23508
rect 23934 23468 23940 23480
rect 23992 23468 23998 23520
rect 25222 23468 25228 23520
rect 25280 23468 25286 23520
rect 1104 23418 25852 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 25852 23418
rect 1104 23344 25852 23366
rect 9125 23307 9183 23313
rect 9125 23273 9137 23307
rect 9171 23304 9183 23307
rect 9214 23304 9220 23316
rect 9171 23276 9220 23304
rect 9171 23273 9183 23276
rect 9125 23267 9183 23273
rect 9214 23264 9220 23276
rect 9272 23264 9278 23316
rect 14369 23307 14427 23313
rect 14369 23273 14381 23307
rect 14415 23304 14427 23307
rect 14458 23304 14464 23316
rect 14415 23276 14464 23304
rect 14415 23273 14427 23276
rect 14369 23267 14427 23273
rect 14458 23264 14464 23276
rect 14516 23264 14522 23316
rect 15841 23307 15899 23313
rect 15841 23273 15853 23307
rect 15887 23304 15899 23307
rect 16758 23304 16764 23316
rect 15887 23276 16764 23304
rect 15887 23273 15899 23276
rect 15841 23267 15899 23273
rect 9398 23196 9404 23248
rect 9456 23236 9462 23248
rect 9456 23208 11928 23236
rect 9456 23196 9462 23208
rect 8662 23128 8668 23180
rect 8720 23168 8726 23180
rect 9677 23171 9735 23177
rect 9677 23168 9689 23171
rect 8720 23140 9689 23168
rect 8720 23128 8726 23140
rect 9677 23137 9689 23140
rect 9723 23137 9735 23171
rect 9677 23131 9735 23137
rect 11698 23128 11704 23180
rect 11756 23128 11762 23180
rect 11793 23171 11851 23177
rect 11793 23137 11805 23171
rect 11839 23137 11851 23171
rect 11900 23168 11928 23208
rect 12618 23196 12624 23248
rect 12676 23236 12682 23248
rect 14737 23239 14795 23245
rect 14737 23236 14749 23239
rect 12676 23208 14749 23236
rect 12676 23196 12682 23208
rect 14737 23205 14749 23208
rect 14783 23205 14795 23239
rect 14737 23199 14795 23205
rect 13541 23171 13599 23177
rect 13541 23168 13553 23171
rect 11900 23140 13553 23168
rect 11793 23131 11851 23137
rect 13541 23137 13553 23140
rect 13587 23137 13599 23171
rect 13541 23131 13599 23137
rect 9858 23060 9864 23112
rect 9916 23100 9922 23112
rect 11808 23100 11836 23131
rect 13630 23128 13636 23180
rect 13688 23168 13694 23180
rect 15289 23171 15347 23177
rect 15289 23168 15301 23171
rect 13688 23140 15301 23168
rect 13688 23128 13694 23140
rect 15289 23137 15301 23140
rect 15335 23137 15347 23171
rect 15289 23131 15347 23137
rect 9916 23072 11836 23100
rect 13357 23103 13415 23109
rect 9916 23060 9922 23072
rect 13357 23069 13369 23103
rect 13403 23100 13415 23103
rect 14458 23100 14464 23112
rect 13403 23072 14464 23100
rect 13403 23069 13415 23072
rect 13357 23063 13415 23069
rect 14458 23060 14464 23072
rect 14516 23060 14522 23112
rect 15105 23103 15163 23109
rect 15105 23069 15117 23103
rect 15151 23100 15163 23103
rect 15654 23100 15660 23112
rect 15151 23072 15660 23100
rect 15151 23069 15163 23072
rect 15105 23063 15163 23069
rect 15654 23060 15660 23072
rect 15712 23060 15718 23112
rect 9493 23035 9551 23041
rect 9493 23001 9505 23035
rect 9539 23032 9551 23035
rect 10410 23032 10416 23044
rect 9539 23004 10416 23032
rect 9539 23001 9551 23004
rect 9493 22995 9551 23001
rect 10410 22992 10416 23004
rect 10468 22992 10474 23044
rect 11609 23035 11667 23041
rect 11609 23001 11621 23035
rect 11655 23032 11667 23035
rect 11790 23032 11796 23044
rect 11655 23004 11796 23032
rect 11655 23001 11667 23004
rect 11609 22995 11667 23001
rect 11790 22992 11796 23004
rect 11848 22992 11854 23044
rect 13449 23035 13507 23041
rect 13449 23001 13461 23035
rect 13495 23032 13507 23035
rect 14185 23035 14243 23041
rect 14185 23032 14197 23035
rect 13495 23004 14197 23032
rect 13495 23001 13507 23004
rect 13449 22995 13507 23001
rect 14185 23001 14197 23004
rect 14231 23032 14243 23035
rect 15197 23035 15255 23041
rect 14231 23004 15148 23032
rect 14231 23001 14243 23004
rect 14185 22995 14243 23001
rect 9585 22967 9643 22973
rect 9585 22933 9597 22967
rect 9631 22964 9643 22967
rect 9766 22964 9772 22976
rect 9631 22936 9772 22964
rect 9631 22933 9643 22936
rect 9585 22927 9643 22933
rect 9766 22924 9772 22936
rect 9824 22924 9830 22976
rect 10502 22924 10508 22976
rect 10560 22964 10566 22976
rect 11241 22967 11299 22973
rect 11241 22964 11253 22967
rect 10560 22936 11253 22964
rect 10560 22924 10566 22936
rect 11241 22933 11253 22936
rect 11287 22933 11299 22967
rect 11241 22927 11299 22933
rect 12158 22924 12164 22976
rect 12216 22964 12222 22976
rect 12989 22967 13047 22973
rect 12989 22964 13001 22967
rect 12216 22936 13001 22964
rect 12216 22924 12222 22936
rect 12989 22933 13001 22936
rect 13035 22933 13047 22967
rect 15120 22964 15148 23004
rect 15197 23001 15209 23035
rect 15243 23032 15255 23035
rect 15856 23032 15884 23267
rect 16758 23264 16764 23276
rect 16816 23304 16822 23316
rect 26326 23304 26332 23316
rect 16816 23276 26332 23304
rect 16816 23264 16822 23276
rect 26326 23264 26332 23276
rect 26384 23264 26390 23316
rect 17865 23239 17923 23245
rect 17865 23205 17877 23239
rect 17911 23236 17923 23239
rect 18690 23236 18696 23248
rect 17911 23208 18696 23236
rect 17911 23205 17923 23208
rect 17865 23199 17923 23205
rect 18690 23196 18696 23208
rect 18748 23196 18754 23248
rect 18969 23239 19027 23245
rect 18969 23205 18981 23239
rect 19015 23236 19027 23239
rect 19702 23236 19708 23248
rect 19015 23208 19708 23236
rect 19015 23205 19027 23208
rect 18969 23199 19027 23205
rect 19702 23196 19708 23208
rect 19760 23196 19766 23248
rect 18506 23128 18512 23180
rect 18564 23128 18570 23180
rect 18598 23128 18604 23180
rect 18656 23168 18662 23180
rect 18782 23168 18788 23180
rect 18656 23140 18788 23168
rect 18656 23128 18662 23140
rect 18782 23128 18788 23140
rect 18840 23128 18846 23180
rect 19978 23128 19984 23180
rect 20036 23128 20042 23180
rect 20165 23171 20223 23177
rect 20165 23137 20177 23171
rect 20211 23168 20223 23171
rect 20438 23168 20444 23180
rect 20211 23140 20444 23168
rect 20211 23137 20223 23140
rect 20165 23131 20223 23137
rect 20438 23128 20444 23140
rect 20496 23128 20502 23180
rect 20717 23171 20775 23177
rect 20717 23137 20729 23171
rect 20763 23168 20775 23171
rect 20806 23168 20812 23180
rect 20763 23140 20812 23168
rect 20763 23137 20775 23140
rect 20717 23131 20775 23137
rect 20806 23128 20812 23140
rect 20864 23128 20870 23180
rect 24302 23128 24308 23180
rect 24360 23168 24366 23180
rect 25041 23171 25099 23177
rect 25041 23168 25053 23171
rect 24360 23140 25053 23168
rect 24360 23128 24366 23140
rect 25041 23137 25053 23140
rect 25087 23137 25099 23171
rect 25041 23131 25099 23137
rect 25225 23171 25283 23177
rect 25225 23137 25237 23171
rect 25271 23168 25283 23171
rect 25314 23168 25320 23180
rect 25271 23140 25320 23168
rect 25271 23137 25283 23140
rect 25225 23131 25283 23137
rect 25314 23128 25320 23140
rect 25372 23128 25378 23180
rect 18233 23103 18291 23109
rect 18233 23069 18245 23103
rect 18279 23100 18291 23103
rect 18322 23100 18328 23112
rect 18279 23072 18328 23100
rect 18279 23069 18291 23072
rect 18233 23063 18291 23069
rect 18322 23060 18328 23072
rect 18380 23060 18386 23112
rect 19242 23060 19248 23112
rect 19300 23100 19306 23112
rect 19889 23103 19947 23109
rect 19889 23100 19901 23103
rect 19300 23072 19901 23100
rect 19300 23060 19306 23072
rect 19889 23069 19901 23072
rect 19935 23069 19947 23103
rect 19889 23063 19947 23069
rect 21821 23103 21879 23109
rect 21821 23069 21833 23103
rect 21867 23069 21879 23103
rect 21821 23063 21879 23069
rect 22833 23103 22891 23109
rect 22833 23069 22845 23103
rect 22879 23100 22891 23103
rect 23750 23100 23756 23112
rect 22879 23072 23756 23100
rect 22879 23069 22891 23072
rect 22833 23063 22891 23069
rect 15243 23004 15884 23032
rect 15243 23001 15255 23004
rect 15197 22995 15255 23001
rect 16850 22992 16856 23044
rect 16908 23032 16914 23044
rect 21836 23032 21864 23063
rect 23750 23060 23756 23072
rect 23808 23060 23814 23112
rect 24949 23103 25007 23109
rect 24949 23069 24961 23103
rect 24995 23100 25007 23103
rect 25590 23100 25596 23112
rect 24995 23072 25596 23100
rect 24995 23069 25007 23072
rect 24949 23063 25007 23069
rect 25590 23060 25596 23072
rect 25648 23060 25654 23112
rect 16908 23004 21864 23032
rect 23845 23035 23903 23041
rect 16908 22992 16914 23004
rect 23845 23001 23857 23035
rect 23891 23032 23903 23035
rect 24854 23032 24860 23044
rect 23891 23004 24860 23032
rect 23891 23001 23903 23004
rect 23845 22995 23903 23001
rect 24854 22992 24860 23004
rect 24912 22992 24918 23044
rect 16574 22964 16580 22976
rect 15120 22936 16580 22964
rect 12989 22927 13047 22933
rect 16574 22924 16580 22936
rect 16632 22924 16638 22976
rect 18230 22924 18236 22976
rect 18288 22964 18294 22976
rect 18325 22967 18383 22973
rect 18325 22964 18337 22967
rect 18288 22936 18337 22964
rect 18288 22924 18294 22936
rect 18325 22933 18337 22936
rect 18371 22964 18383 22967
rect 18598 22964 18604 22976
rect 18371 22936 18604 22964
rect 18371 22933 18383 22936
rect 18325 22927 18383 22933
rect 18598 22924 18604 22936
rect 18656 22924 18662 22976
rect 19242 22924 19248 22976
rect 19300 22964 19306 22976
rect 19521 22967 19579 22973
rect 19521 22964 19533 22967
rect 19300 22936 19533 22964
rect 19300 22924 19306 22936
rect 19521 22933 19533 22936
rect 19567 22933 19579 22967
rect 19521 22927 19579 22933
rect 21637 22967 21695 22973
rect 21637 22933 21649 22967
rect 21683 22964 21695 22967
rect 22094 22964 22100 22976
rect 21683 22936 22100 22964
rect 21683 22933 21695 22936
rect 21637 22927 21695 22933
rect 22094 22924 22100 22936
rect 22152 22924 22158 22976
rect 22554 22924 22560 22976
rect 22612 22964 22618 22976
rect 24581 22967 24639 22973
rect 24581 22964 24593 22967
rect 22612 22936 24593 22964
rect 22612 22924 22618 22936
rect 24581 22933 24593 22936
rect 24627 22933 24639 22967
rect 24581 22927 24639 22933
rect 1104 22874 25852 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 25852 22874
rect 1104 22800 25852 22822
rect 9306 22720 9312 22772
rect 9364 22760 9370 22772
rect 10134 22760 10140 22772
rect 9364 22732 10140 22760
rect 9364 22720 9370 22732
rect 10134 22720 10140 22732
rect 10192 22720 10198 22772
rect 14461 22763 14519 22769
rect 14461 22729 14473 22763
rect 14507 22760 14519 22763
rect 14734 22760 14740 22772
rect 14507 22732 14740 22760
rect 14507 22729 14519 22732
rect 14461 22723 14519 22729
rect 8938 22652 8944 22704
rect 8996 22652 9002 22704
rect 14476 22692 14504 22723
rect 14734 22720 14740 22732
rect 14792 22720 14798 22772
rect 16850 22720 16856 22772
rect 16908 22720 16914 22772
rect 18322 22720 18328 22772
rect 18380 22760 18386 22772
rect 18693 22763 18751 22769
rect 18693 22760 18705 22763
rect 18380 22732 18705 22760
rect 18380 22720 18386 22732
rect 18693 22729 18705 22732
rect 18739 22760 18751 22763
rect 18966 22760 18972 22772
rect 18739 22732 18972 22760
rect 18739 22729 18751 22732
rect 18693 22723 18751 22729
rect 18966 22720 18972 22732
rect 19024 22720 19030 22772
rect 19610 22720 19616 22772
rect 19668 22760 19674 22772
rect 19705 22763 19763 22769
rect 19705 22760 19717 22763
rect 19668 22732 19717 22760
rect 19668 22720 19674 22732
rect 19705 22729 19717 22732
rect 19751 22729 19763 22763
rect 19705 22723 19763 22729
rect 21177 22763 21235 22769
rect 21177 22729 21189 22763
rect 21223 22760 21235 22763
rect 25130 22760 25136 22772
rect 21223 22732 25136 22760
rect 21223 22729 21235 22732
rect 21177 22723 21235 22729
rect 25130 22720 25136 22732
rect 25188 22720 25194 22772
rect 13846 22664 14504 22692
rect 18598 22652 18604 22704
rect 18656 22692 18662 22704
rect 18877 22695 18935 22701
rect 18877 22692 18889 22695
rect 18656 22664 18889 22692
rect 18656 22652 18662 22664
rect 18877 22661 18889 22664
rect 18923 22692 18935 22695
rect 20898 22692 20904 22704
rect 18923 22664 20904 22692
rect 18923 22661 18935 22664
rect 18877 22655 18935 22661
rect 20898 22652 20904 22664
rect 20956 22652 20962 22704
rect 7834 22584 7840 22636
rect 7892 22624 7898 22636
rect 8113 22627 8171 22633
rect 8113 22624 8125 22627
rect 7892 22596 8125 22624
rect 7892 22584 7898 22596
rect 8113 22593 8125 22596
rect 8159 22593 8171 22627
rect 8113 22587 8171 22593
rect 12342 22584 12348 22636
rect 12400 22584 12406 22636
rect 17037 22627 17095 22633
rect 17037 22593 17049 22627
rect 17083 22593 17095 22627
rect 17037 22587 17095 22593
rect 8389 22559 8447 22565
rect 8389 22525 8401 22559
rect 8435 22556 8447 22559
rect 10870 22556 10876 22568
rect 8435 22528 10876 22556
rect 8435 22525 8447 22528
rect 8389 22519 8447 22525
rect 10870 22516 10876 22528
rect 10928 22516 10934 22568
rect 12621 22559 12679 22565
rect 12621 22525 12633 22559
rect 12667 22556 12679 22559
rect 13354 22556 13360 22568
rect 12667 22528 13360 22556
rect 12667 22525 12679 22528
rect 12621 22519 12679 22525
rect 13354 22516 13360 22528
rect 13412 22516 13418 22568
rect 17052 22488 17080 22587
rect 20438 22584 20444 22636
rect 20496 22624 20502 22636
rect 21085 22627 21143 22633
rect 21085 22624 21097 22627
rect 20496 22596 21097 22624
rect 20496 22584 20502 22596
rect 21085 22593 21097 22596
rect 21131 22624 21143 22627
rect 21450 22624 21456 22636
rect 21131 22596 21456 22624
rect 21131 22593 21143 22596
rect 21085 22587 21143 22593
rect 21450 22584 21456 22596
rect 21508 22584 21514 22636
rect 22094 22584 22100 22636
rect 22152 22584 22158 22636
rect 22830 22584 22836 22636
rect 22888 22624 22894 22636
rect 23937 22627 23995 22633
rect 23937 22624 23949 22627
rect 22888 22596 23949 22624
rect 22888 22584 22894 22596
rect 23937 22593 23949 22596
rect 23983 22593 23995 22627
rect 23937 22587 23995 22593
rect 18598 22516 18604 22568
rect 18656 22556 18662 22568
rect 19150 22556 19156 22568
rect 18656 22528 19156 22556
rect 18656 22516 18662 22528
rect 19150 22516 19156 22528
rect 19208 22516 19214 22568
rect 19518 22516 19524 22568
rect 19576 22556 19582 22568
rect 19794 22556 19800 22568
rect 19576 22528 19800 22556
rect 19576 22516 19582 22528
rect 19794 22516 19800 22528
rect 19852 22516 19858 22568
rect 20162 22516 20168 22568
rect 20220 22556 20226 22568
rect 21269 22559 21327 22565
rect 21269 22556 21281 22559
rect 20220 22528 21281 22556
rect 20220 22516 20226 22528
rect 21269 22525 21281 22528
rect 21315 22525 21327 22559
rect 21269 22519 21327 22525
rect 23293 22559 23351 22565
rect 23293 22525 23305 22559
rect 23339 22556 23351 22559
rect 23382 22556 23388 22568
rect 23339 22528 23388 22556
rect 23339 22525 23351 22528
rect 23293 22519 23351 22525
rect 23382 22516 23388 22528
rect 23440 22516 23446 22568
rect 24762 22516 24768 22568
rect 24820 22516 24826 22568
rect 13635 22460 17080 22488
rect 6914 22380 6920 22432
rect 6972 22420 6978 22432
rect 9858 22420 9864 22432
rect 6972 22392 9864 22420
rect 6972 22380 6978 22392
rect 9858 22380 9864 22392
rect 9916 22380 9922 22432
rect 12066 22380 12072 22432
rect 12124 22420 12130 22432
rect 13635 22420 13663 22460
rect 22278 22448 22284 22500
rect 22336 22488 22342 22500
rect 22830 22488 22836 22500
rect 22336 22460 22836 22488
rect 22336 22448 22342 22460
rect 22830 22448 22836 22460
rect 22888 22448 22894 22500
rect 12124 22392 13663 22420
rect 12124 22380 12130 22392
rect 14090 22380 14096 22432
rect 14148 22380 14154 22432
rect 20438 22380 20444 22432
rect 20496 22380 20502 22432
rect 20714 22380 20720 22432
rect 20772 22380 20778 22432
rect 1104 22330 25852 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 25852 22330
rect 1104 22256 25852 22278
rect 11054 22176 11060 22228
rect 11112 22216 11118 22228
rect 21808 22219 21866 22225
rect 11112 22188 12434 22216
rect 11112 22176 11118 22188
rect 11977 22151 12035 22157
rect 11977 22117 11989 22151
rect 12023 22148 12035 22151
rect 12066 22148 12072 22160
rect 12023 22120 12072 22148
rect 12023 22117 12035 22120
rect 11977 22111 12035 22117
rect 12066 22108 12072 22120
rect 12124 22108 12130 22160
rect 12406 22148 12434 22188
rect 21808 22185 21820 22219
rect 21854 22216 21866 22219
rect 23290 22216 23296 22228
rect 21854 22188 23296 22216
rect 21854 22185 21866 22188
rect 21808 22179 21866 22185
rect 23290 22176 23296 22188
rect 23348 22176 23354 22228
rect 23750 22176 23756 22228
rect 23808 22176 23814 22228
rect 15746 22148 15752 22160
rect 12406 22120 12572 22148
rect 8938 22040 8944 22092
rect 8996 22040 9002 22092
rect 11330 22040 11336 22092
rect 11388 22040 11394 22092
rect 12434 22040 12440 22092
rect 12492 22040 12498 22092
rect 12544 22089 12572 22120
rect 15304 22120 15752 22148
rect 15304 22089 15332 22120
rect 15746 22108 15752 22120
rect 15804 22108 15810 22160
rect 25498 22148 25504 22160
rect 25240 22120 25504 22148
rect 12529 22083 12587 22089
rect 12529 22049 12541 22083
rect 12575 22049 12587 22083
rect 12529 22043 12587 22049
rect 15289 22083 15347 22089
rect 15289 22049 15301 22083
rect 15335 22080 15347 22083
rect 15473 22083 15531 22089
rect 15335 22052 15369 22080
rect 15335 22049 15347 22052
rect 15289 22043 15347 22049
rect 15473 22049 15485 22083
rect 15519 22049 15531 22083
rect 15473 22043 15531 22049
rect 9490 21972 9496 22024
rect 9548 22012 9554 22024
rect 9548 21984 11284 22012
rect 9548 21972 9554 21984
rect 11149 21947 11207 21953
rect 11149 21944 11161 21947
rect 10336 21916 11161 21944
rect 10336 21888 10364 21916
rect 11149 21913 11161 21916
rect 11195 21913 11207 21947
rect 11149 21907 11207 21913
rect 10318 21836 10324 21888
rect 10376 21836 10382 21888
rect 10686 21836 10692 21888
rect 10744 21836 10750 21888
rect 11054 21836 11060 21888
rect 11112 21836 11118 21888
rect 11256 21876 11284 21984
rect 14090 21972 14096 22024
rect 14148 22012 14154 22024
rect 15488 22012 15516 22043
rect 18782 22040 18788 22092
rect 18840 22080 18846 22092
rect 20165 22083 20223 22089
rect 20165 22080 20177 22083
rect 18840 22052 20177 22080
rect 18840 22040 18846 22052
rect 20165 22049 20177 22052
rect 20211 22049 20223 22083
rect 20165 22043 20223 22049
rect 14148 21984 15516 22012
rect 16117 22015 16175 22021
rect 14148 21972 14154 21984
rect 16117 21981 16129 22015
rect 16163 21981 16175 22015
rect 20180 22012 20208 22043
rect 20346 22040 20352 22092
rect 20404 22040 20410 22092
rect 21545 22083 21603 22089
rect 21545 22049 21557 22083
rect 21591 22080 21603 22083
rect 22186 22080 22192 22092
rect 21591 22052 22192 22080
rect 21591 22049 21603 22052
rect 21545 22043 21603 22049
rect 22186 22040 22192 22052
rect 22244 22040 22250 22092
rect 22830 22040 22836 22092
rect 22888 22080 22894 22092
rect 23293 22083 23351 22089
rect 23293 22080 23305 22083
rect 22888 22052 23305 22080
rect 22888 22040 22894 22052
rect 23293 22049 23305 22052
rect 23339 22049 23351 22083
rect 23293 22043 23351 22049
rect 25038 22040 25044 22092
rect 25096 22040 25102 22092
rect 25240 22089 25268 22120
rect 25498 22108 25504 22120
rect 25556 22108 25562 22160
rect 25225 22083 25283 22089
rect 25225 22049 25237 22083
rect 25271 22049 25283 22083
rect 25225 22043 25283 22049
rect 21358 22012 21364 22024
rect 20180 21984 21364 22012
rect 16117 21975 16175 21981
rect 12345 21879 12403 21885
rect 12345 21876 12357 21879
rect 11256 21848 12357 21876
rect 12345 21845 12357 21848
rect 12391 21845 12403 21879
rect 12345 21839 12403 21845
rect 14826 21836 14832 21888
rect 14884 21836 14890 21888
rect 15194 21836 15200 21888
rect 15252 21836 15258 21888
rect 16132 21876 16160 21975
rect 21358 21972 21364 21984
rect 21416 21972 21422 22024
rect 23934 21972 23940 22024
rect 23992 21972 23998 22024
rect 16390 21904 16396 21956
rect 16448 21944 16454 21956
rect 17770 21944 17776 21956
rect 16448 21916 16804 21944
rect 17618 21916 17776 21944
rect 16448 21904 16454 21916
rect 16574 21876 16580 21888
rect 16132 21848 16580 21876
rect 16574 21836 16580 21848
rect 16632 21836 16638 21888
rect 16776 21876 16804 21916
rect 17770 21904 17776 21916
rect 17828 21944 17834 21956
rect 18141 21947 18199 21953
rect 18141 21944 18153 21947
rect 17828 21916 18153 21944
rect 17828 21904 17834 21916
rect 18141 21913 18153 21916
rect 18187 21913 18199 21947
rect 18141 21907 18199 21913
rect 21542 21904 21548 21956
rect 21600 21944 21606 21956
rect 24949 21947 25007 21953
rect 24949 21944 24961 21947
rect 21600 21916 22310 21944
rect 23124 21916 24961 21944
rect 21600 21904 21606 21916
rect 17034 21876 17040 21888
rect 16776 21848 17040 21876
rect 17034 21836 17040 21848
rect 17092 21836 17098 21888
rect 17126 21836 17132 21888
rect 17184 21876 17190 21888
rect 17865 21879 17923 21885
rect 17865 21876 17877 21879
rect 17184 21848 17877 21876
rect 17184 21836 17190 21848
rect 17865 21845 17877 21848
rect 17911 21845 17923 21879
rect 17865 21839 17923 21845
rect 19705 21879 19763 21885
rect 19705 21845 19717 21879
rect 19751 21876 19763 21879
rect 19886 21876 19892 21888
rect 19751 21848 19892 21876
rect 19751 21845 19763 21848
rect 19705 21839 19763 21845
rect 19886 21836 19892 21848
rect 19944 21836 19950 21888
rect 20070 21836 20076 21888
rect 20128 21836 20134 21888
rect 20901 21879 20959 21885
rect 20901 21845 20913 21879
rect 20947 21876 20959 21879
rect 23124 21876 23152 21916
rect 24949 21913 24961 21916
rect 24995 21913 25007 21947
rect 24949 21907 25007 21913
rect 20947 21848 23152 21876
rect 20947 21845 20959 21848
rect 20901 21839 20959 21845
rect 24026 21836 24032 21888
rect 24084 21876 24090 21888
rect 24581 21879 24639 21885
rect 24581 21876 24593 21879
rect 24084 21848 24593 21876
rect 24084 21836 24090 21848
rect 24581 21845 24593 21848
rect 24627 21845 24639 21879
rect 24581 21839 24639 21845
rect 1104 21786 25852 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 25852 21786
rect 1104 21712 25852 21734
rect 9217 21675 9275 21681
rect 9217 21641 9229 21675
rect 9263 21641 9275 21675
rect 9217 21635 9275 21641
rect 8938 21604 8944 21616
rect 8418 21576 8944 21604
rect 8938 21564 8944 21576
rect 8996 21564 9002 21616
rect 9232 21604 9260 21635
rect 10226 21632 10232 21684
rect 10284 21672 10290 21684
rect 10413 21675 10471 21681
rect 10413 21672 10425 21675
rect 10284 21644 10425 21672
rect 10284 21632 10290 21644
rect 10413 21641 10425 21644
rect 10459 21641 10471 21675
rect 10413 21635 10471 21641
rect 11054 21632 11060 21684
rect 11112 21672 11118 21684
rect 11701 21675 11759 21681
rect 11701 21672 11713 21675
rect 11112 21644 11713 21672
rect 11112 21632 11118 21644
rect 11701 21641 11713 21644
rect 11747 21641 11759 21675
rect 14090 21672 14096 21684
rect 11701 21635 11759 21641
rect 13372 21644 14096 21672
rect 9232 21576 10640 21604
rect 9585 21539 9643 21545
rect 9585 21505 9597 21539
rect 9631 21536 9643 21539
rect 9950 21536 9956 21548
rect 9631 21508 9956 21536
rect 9631 21505 9643 21508
rect 9585 21499 9643 21505
rect 9950 21496 9956 21508
rect 10008 21496 10014 21548
rect 6917 21471 6975 21477
rect 6917 21437 6929 21471
rect 6963 21437 6975 21471
rect 6917 21431 6975 21437
rect 7193 21471 7251 21477
rect 7193 21437 7205 21471
rect 7239 21468 7251 21471
rect 8846 21468 8852 21480
rect 7239 21440 8852 21468
rect 7239 21437 7251 21440
rect 7193 21431 7251 21437
rect 6932 21332 6960 21431
rect 8846 21428 8852 21440
rect 8904 21428 8910 21480
rect 8938 21428 8944 21480
rect 8996 21468 9002 21480
rect 9677 21471 9735 21477
rect 9677 21468 9689 21471
rect 8996 21440 9689 21468
rect 8996 21428 9002 21440
rect 9677 21437 9689 21440
rect 9723 21437 9735 21471
rect 9677 21431 9735 21437
rect 9769 21471 9827 21477
rect 9769 21437 9781 21471
rect 9815 21437 9827 21471
rect 9769 21431 9827 21437
rect 7742 21332 7748 21344
rect 6932 21304 7748 21332
rect 7742 21292 7748 21304
rect 7800 21292 7806 21344
rect 8294 21292 8300 21344
rect 8352 21332 8358 21344
rect 8662 21332 8668 21344
rect 8352 21304 8668 21332
rect 8352 21292 8358 21304
rect 8662 21292 8668 21304
rect 8720 21292 8726 21344
rect 9582 21292 9588 21344
rect 9640 21332 9646 21344
rect 9784 21332 9812 21431
rect 9640 21304 9812 21332
rect 10612 21332 10640 21576
rect 10686 21564 10692 21616
rect 10744 21604 10750 21616
rect 13372 21613 13400 21644
rect 14090 21632 14096 21644
rect 14148 21632 14154 21684
rect 15102 21632 15108 21684
rect 15160 21672 15166 21684
rect 15749 21675 15807 21681
rect 15749 21672 15761 21675
rect 15160 21644 15761 21672
rect 15160 21632 15166 21644
rect 15749 21641 15761 21644
rect 15795 21641 15807 21675
rect 15749 21635 15807 21641
rect 20070 21632 20076 21684
rect 20128 21672 20134 21684
rect 21177 21675 21235 21681
rect 21177 21672 21189 21675
rect 20128 21644 21189 21672
rect 20128 21632 20134 21644
rect 21177 21641 21189 21644
rect 21223 21641 21235 21675
rect 21177 21635 21235 21641
rect 21358 21632 21364 21684
rect 21416 21632 21422 21684
rect 22462 21632 22468 21684
rect 22520 21632 22526 21684
rect 22646 21632 22652 21684
rect 22704 21672 22710 21684
rect 22830 21672 22836 21684
rect 22704 21644 22836 21672
rect 22704 21632 22710 21644
rect 22830 21632 22836 21644
rect 22888 21632 22894 21684
rect 23290 21632 23296 21684
rect 23348 21672 23354 21684
rect 25041 21675 25099 21681
rect 25041 21672 25053 21675
rect 23348 21644 25053 21672
rect 23348 21632 23354 21644
rect 25041 21641 25053 21644
rect 25087 21641 25099 21675
rect 25041 21635 25099 21641
rect 13357 21607 13415 21613
rect 10744 21576 11652 21604
rect 10744 21564 10750 21576
rect 10781 21539 10839 21545
rect 10781 21505 10793 21539
rect 10827 21536 10839 21539
rect 11514 21536 11520 21548
rect 10827 21508 11520 21536
rect 10827 21505 10839 21508
rect 10781 21499 10839 21505
rect 11514 21496 11520 21508
rect 11572 21496 11578 21548
rect 10870 21428 10876 21480
rect 10928 21428 10934 21480
rect 10962 21428 10968 21480
rect 11020 21428 11026 21480
rect 11624 21400 11652 21576
rect 13357 21573 13369 21607
rect 13403 21573 13415 21607
rect 13357 21567 13415 21573
rect 14826 21564 14832 21616
rect 14884 21604 14890 21616
rect 14884 21576 18920 21604
rect 14884 21564 14890 21576
rect 18892 21545 18920 21576
rect 22186 21564 22192 21616
rect 22244 21604 22250 21616
rect 22244 21576 23336 21604
rect 22244 21564 22250 21576
rect 15657 21539 15715 21545
rect 14490 21508 14688 21536
rect 12342 21428 12348 21480
rect 12400 21468 12406 21480
rect 12710 21468 12716 21480
rect 12400 21440 12716 21468
rect 12400 21428 12406 21440
rect 12710 21428 12716 21440
rect 12768 21468 12774 21480
rect 13081 21471 13139 21477
rect 13081 21468 13093 21471
rect 12768 21440 13093 21468
rect 12768 21428 12774 21440
rect 13081 21437 13093 21440
rect 13127 21437 13139 21471
rect 13081 21431 13139 21437
rect 14660 21412 14688 21508
rect 15657 21505 15669 21539
rect 15703 21505 15715 21539
rect 15657 21499 15715 21505
rect 18877 21539 18935 21545
rect 18877 21505 18889 21539
rect 18923 21505 18935 21539
rect 18877 21499 18935 21505
rect 19889 21539 19947 21545
rect 19889 21505 19901 21539
rect 19935 21536 19947 21539
rect 20717 21539 20775 21545
rect 20717 21536 20729 21539
rect 19935 21508 20729 21536
rect 19935 21505 19947 21508
rect 19889 21499 19947 21505
rect 20717 21505 20729 21508
rect 20763 21505 20775 21539
rect 20717 21499 20775 21505
rect 15672 21468 15700 21499
rect 22002 21496 22008 21548
rect 22060 21536 22066 21548
rect 23308 21545 23336 21576
rect 24118 21564 24124 21616
rect 24176 21564 24182 21616
rect 22373 21539 22431 21545
rect 22373 21536 22385 21539
rect 22060 21508 22385 21536
rect 22060 21496 22066 21508
rect 22373 21505 22385 21508
rect 22419 21505 22431 21539
rect 22373 21499 22431 21505
rect 23293 21539 23351 21545
rect 23293 21505 23305 21539
rect 23339 21505 23351 21539
rect 23293 21499 23351 21505
rect 19058 21468 19064 21480
rect 15672 21440 19064 21468
rect 19058 21428 19064 21440
rect 19116 21428 19122 21480
rect 19150 21428 19156 21480
rect 19208 21468 19214 21480
rect 19981 21471 20039 21477
rect 19981 21468 19993 21471
rect 19208 21440 19993 21468
rect 19208 21428 19214 21440
rect 19981 21437 19993 21440
rect 20027 21437 20039 21471
rect 19981 21431 20039 21437
rect 20162 21428 20168 21480
rect 20220 21428 20226 21480
rect 22649 21471 22707 21477
rect 22649 21437 22661 21471
rect 22695 21437 22707 21471
rect 22649 21431 22707 21437
rect 23569 21471 23627 21477
rect 23569 21437 23581 21471
rect 23615 21468 23627 21471
rect 25314 21468 25320 21480
rect 23615 21440 25320 21468
rect 23615 21437 23627 21440
rect 23569 21431 23627 21437
rect 11624 21372 13216 21400
rect 12526 21332 12532 21344
rect 10612 21304 12532 21332
rect 9640 21292 9646 21304
rect 12526 21292 12532 21304
rect 12584 21292 12590 21344
rect 13188 21332 13216 21372
rect 14642 21360 14648 21412
rect 14700 21400 14706 21412
rect 15105 21403 15163 21409
rect 15105 21400 15117 21403
rect 14700 21372 15117 21400
rect 14700 21360 14706 21372
rect 15105 21369 15117 21372
rect 15151 21369 15163 21403
rect 15105 21363 15163 21369
rect 15286 21360 15292 21412
rect 15344 21400 15350 21412
rect 18693 21403 18751 21409
rect 15344 21372 17724 21400
rect 15344 21360 15350 21372
rect 14090 21332 14096 21344
rect 13188 21304 14096 21332
rect 14090 21292 14096 21304
rect 14148 21292 14154 21344
rect 14366 21292 14372 21344
rect 14424 21332 14430 21344
rect 14829 21335 14887 21341
rect 14829 21332 14841 21335
rect 14424 21304 14841 21332
rect 14424 21292 14430 21304
rect 14829 21301 14841 21304
rect 14875 21332 14887 21335
rect 15010 21332 15016 21344
rect 14875 21304 15016 21332
rect 14875 21301 14887 21304
rect 14829 21295 14887 21301
rect 15010 21292 15016 21304
rect 15068 21292 15074 21344
rect 17696 21332 17724 21372
rect 18693 21369 18705 21403
rect 18739 21400 18751 21403
rect 21082 21400 21088 21412
rect 18739 21372 21088 21400
rect 18739 21369 18751 21372
rect 18693 21363 18751 21369
rect 21082 21360 21088 21372
rect 21140 21360 21146 21412
rect 19150 21332 19156 21344
rect 17696 21304 19156 21332
rect 19150 21292 19156 21304
rect 19208 21292 19214 21344
rect 19521 21335 19579 21341
rect 19521 21301 19533 21335
rect 19567 21332 19579 21335
rect 20438 21332 20444 21344
rect 19567 21304 20444 21332
rect 19567 21301 19579 21304
rect 19521 21295 19579 21301
rect 20438 21292 20444 21304
rect 20496 21292 20502 21344
rect 21542 21292 21548 21344
rect 21600 21292 21606 21344
rect 21726 21292 21732 21344
rect 21784 21332 21790 21344
rect 22005 21335 22063 21341
rect 22005 21332 22017 21335
rect 21784 21304 22017 21332
rect 21784 21292 21790 21304
rect 22005 21301 22017 21304
rect 22051 21301 22063 21335
rect 22664 21332 22692 21431
rect 25314 21428 25320 21440
rect 25372 21428 25378 21480
rect 23566 21332 23572 21344
rect 22664 21304 23572 21332
rect 22005 21295 22063 21301
rect 23566 21292 23572 21304
rect 23624 21292 23630 21344
rect 24118 21292 24124 21344
rect 24176 21332 24182 21344
rect 25130 21332 25136 21344
rect 24176 21304 25136 21332
rect 24176 21292 24182 21304
rect 25130 21292 25136 21304
rect 25188 21332 25194 21344
rect 25317 21335 25375 21341
rect 25317 21332 25329 21335
rect 25188 21304 25329 21332
rect 25188 21292 25194 21304
rect 25317 21301 25329 21304
rect 25363 21301 25375 21335
rect 25317 21295 25375 21301
rect 1104 21242 25852 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 25852 21242
rect 1104 21168 25852 21190
rect 3510 21088 3516 21140
rect 3568 21128 3574 21140
rect 15286 21128 15292 21140
rect 3568 21100 15292 21128
rect 3568 21088 3574 21100
rect 15286 21088 15292 21100
rect 15344 21088 15350 21140
rect 15562 21088 15568 21140
rect 15620 21128 15626 21140
rect 15620 21100 20208 21128
rect 15620 21088 15626 21100
rect 12437 21063 12495 21069
rect 12437 21029 12449 21063
rect 12483 21060 12495 21063
rect 13354 21060 13360 21072
rect 12483 21032 13360 21060
rect 12483 21029 12495 21032
rect 12437 21023 12495 21029
rect 13354 21020 13360 21032
rect 13412 21020 13418 21072
rect 16574 21020 16580 21072
rect 16632 21020 16638 21072
rect 19429 21063 19487 21069
rect 19429 21029 19441 21063
rect 19475 21060 19487 21063
rect 20070 21060 20076 21072
rect 19475 21032 20076 21060
rect 19475 21029 19487 21032
rect 19429 21023 19487 21029
rect 20070 21020 20076 21032
rect 20128 21020 20134 21072
rect 9950 20952 9956 21004
rect 10008 20952 10014 21004
rect 15197 20995 15255 21001
rect 15197 20961 15209 20995
rect 15243 20992 15255 20995
rect 16592 20992 16620 21020
rect 15243 20964 16620 20992
rect 15243 20961 15255 20964
rect 15197 20955 15255 20961
rect 19702 20952 19708 21004
rect 19760 20992 19766 21004
rect 19981 20995 20039 21001
rect 19981 20992 19993 20995
rect 19760 20964 19993 20992
rect 19760 20952 19766 20964
rect 19981 20961 19993 20964
rect 20027 20961 20039 20995
rect 20180 20992 20208 21100
rect 20898 21088 20904 21140
rect 20956 21128 20962 21140
rect 21453 21131 21511 21137
rect 21453 21128 21465 21131
rect 20956 21100 21465 21128
rect 20956 21088 20962 21100
rect 21453 21097 21465 21100
rect 21499 21097 21511 21131
rect 21453 21091 21511 21097
rect 20809 21063 20867 21069
rect 20809 21029 20821 21063
rect 20855 21060 20867 21063
rect 20855 21032 22140 21060
rect 20855 21029 20867 21032
rect 20809 21023 20867 21029
rect 20180 20964 21036 20992
rect 19981 20955 20039 20961
rect 10686 20884 10692 20936
rect 10744 20884 10750 20936
rect 18598 20884 18604 20936
rect 18656 20924 18662 20936
rect 21008 20933 21036 20964
rect 22002 20952 22008 21004
rect 22060 20952 22066 21004
rect 19797 20927 19855 20933
rect 19797 20924 19809 20927
rect 18656 20896 19809 20924
rect 18656 20884 18662 20896
rect 19797 20893 19809 20896
rect 19843 20924 19855 20927
rect 20441 20927 20499 20933
rect 20441 20924 20453 20927
rect 19843 20896 20453 20924
rect 19843 20893 19855 20896
rect 19797 20887 19855 20893
rect 20441 20893 20453 20896
rect 20487 20893 20499 20927
rect 20441 20887 20499 20893
rect 20993 20927 21051 20933
rect 20993 20893 21005 20927
rect 21039 20893 21051 20927
rect 22112 20924 22140 21032
rect 23845 20995 23903 21001
rect 23845 20961 23857 20995
rect 23891 20992 23903 20995
rect 24854 20992 24860 21004
rect 23891 20964 24860 20992
rect 23891 20961 23903 20964
rect 23845 20955 23903 20961
rect 24854 20952 24860 20964
rect 24912 20952 24918 21004
rect 24946 20952 24952 21004
rect 25004 20992 25010 21004
rect 25041 20995 25099 21001
rect 25041 20992 25053 20995
rect 25004 20964 25053 20992
rect 25004 20952 25010 20964
rect 25041 20961 25053 20964
rect 25087 20961 25099 20995
rect 25041 20955 25099 20961
rect 25133 20995 25191 21001
rect 25133 20961 25145 20995
rect 25179 20961 25191 20995
rect 25133 20955 25191 20961
rect 22649 20927 22707 20933
rect 22649 20924 22661 20927
rect 22112 20896 22661 20924
rect 20993 20887 21051 20893
rect 22649 20893 22661 20896
rect 22695 20893 22707 20927
rect 22649 20887 22707 20893
rect 23934 20884 23940 20936
rect 23992 20924 23998 20936
rect 25148 20924 25176 20955
rect 23992 20896 25176 20924
rect 23992 20884 23998 20896
rect 10870 20816 10876 20868
rect 10928 20856 10934 20868
rect 10965 20859 11023 20865
rect 10965 20856 10977 20859
rect 10928 20828 10977 20856
rect 10928 20816 10934 20828
rect 10965 20825 10977 20828
rect 11011 20825 11023 20859
rect 15473 20859 15531 20865
rect 12190 20828 12434 20856
rect 10965 20819 11023 20825
rect 8938 20748 8944 20800
rect 8996 20788 9002 20800
rect 9033 20791 9091 20797
rect 9033 20788 9045 20791
rect 8996 20760 9045 20788
rect 8996 20748 9002 20760
rect 9033 20757 9045 20760
rect 9079 20757 9091 20791
rect 12406 20788 12434 20828
rect 15473 20825 15485 20859
rect 15519 20856 15531 20859
rect 15746 20856 15752 20868
rect 15519 20828 15752 20856
rect 15519 20825 15531 20828
rect 15473 20819 15531 20825
rect 15746 20816 15752 20828
rect 15804 20816 15810 20868
rect 19889 20859 19947 20865
rect 16698 20828 17356 20856
rect 12805 20791 12863 20797
rect 12805 20788 12817 20791
rect 12406 20760 12817 20788
rect 9033 20751 9091 20757
rect 12805 20757 12817 20760
rect 12851 20788 12863 20791
rect 14642 20788 14648 20800
rect 12851 20760 14648 20788
rect 12851 20757 12863 20760
rect 12805 20751 12863 20757
rect 14642 20748 14648 20760
rect 14700 20748 14706 20800
rect 16390 20748 16396 20800
rect 16448 20788 16454 20800
rect 17328 20797 17356 20828
rect 19889 20825 19901 20859
rect 19935 20856 19947 20859
rect 20254 20856 20260 20868
rect 19935 20828 20260 20856
rect 19935 20825 19947 20828
rect 19889 20819 19947 20825
rect 20254 20816 20260 20828
rect 20312 20856 20318 20868
rect 21269 20859 21327 20865
rect 21269 20856 21281 20859
rect 20312 20828 21281 20856
rect 20312 20816 20318 20828
rect 21269 20825 21281 20828
rect 21315 20825 21327 20859
rect 21269 20819 21327 20825
rect 16945 20791 17003 20797
rect 16945 20788 16957 20791
rect 16448 20760 16957 20788
rect 16448 20748 16454 20760
rect 16945 20757 16957 20760
rect 16991 20757 17003 20791
rect 16945 20751 17003 20757
rect 17313 20791 17371 20797
rect 17313 20757 17325 20791
rect 17359 20788 17371 20791
rect 17770 20788 17776 20800
rect 17359 20760 17776 20788
rect 17359 20757 17371 20760
rect 17313 20751 17371 20757
rect 17770 20748 17776 20760
rect 17828 20788 17834 20800
rect 18693 20791 18751 20797
rect 18693 20788 18705 20791
rect 17828 20760 18705 20788
rect 17828 20748 17834 20760
rect 18693 20757 18705 20760
rect 18739 20757 18751 20791
rect 18693 20751 18751 20757
rect 18782 20748 18788 20800
rect 18840 20788 18846 20800
rect 18966 20788 18972 20800
rect 18840 20760 18972 20788
rect 18840 20748 18846 20760
rect 18966 20748 18972 20760
rect 19024 20748 19030 20800
rect 24578 20748 24584 20800
rect 24636 20748 24642 20800
rect 24854 20748 24860 20800
rect 24912 20788 24918 20800
rect 24949 20791 25007 20797
rect 24949 20788 24961 20791
rect 24912 20760 24961 20788
rect 24912 20748 24918 20760
rect 24949 20757 24961 20760
rect 24995 20757 25007 20791
rect 24949 20751 25007 20757
rect 1104 20698 25852 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 25852 20698
rect 1104 20624 25852 20646
rect 8846 20544 8852 20596
rect 8904 20584 8910 20596
rect 8904 20556 10364 20584
rect 8904 20544 8910 20556
rect 8021 20519 8079 20525
rect 8021 20485 8033 20519
rect 8067 20516 8079 20519
rect 8294 20516 8300 20528
rect 8067 20488 8300 20516
rect 8067 20485 8079 20488
rect 8021 20479 8079 20485
rect 8294 20476 8300 20488
rect 8352 20476 8358 20528
rect 9030 20476 9036 20528
rect 9088 20476 9094 20528
rect 9306 20476 9312 20528
rect 9364 20516 9370 20528
rect 9582 20516 9588 20528
rect 9364 20488 9588 20516
rect 9364 20476 9370 20488
rect 9582 20476 9588 20488
rect 9640 20516 9646 20528
rect 10045 20519 10103 20525
rect 10045 20516 10057 20519
rect 9640 20488 10057 20516
rect 9640 20476 9646 20488
rect 10045 20485 10057 20488
rect 10091 20485 10103 20519
rect 10045 20479 10103 20485
rect 10336 20448 10364 20556
rect 10410 20544 10416 20596
rect 10468 20544 10474 20596
rect 10781 20587 10839 20593
rect 10781 20553 10793 20587
rect 10827 20584 10839 20587
rect 12618 20584 12624 20596
rect 10827 20556 12624 20584
rect 10827 20553 10839 20556
rect 10781 20547 10839 20553
rect 12618 20544 12624 20556
rect 12676 20544 12682 20596
rect 13630 20544 13636 20596
rect 13688 20584 13694 20596
rect 15381 20587 15439 20593
rect 15381 20584 15393 20587
rect 13688 20556 15393 20584
rect 13688 20544 13694 20556
rect 15381 20553 15393 20556
rect 15427 20553 15439 20587
rect 15381 20547 15439 20553
rect 15470 20544 15476 20596
rect 15528 20544 15534 20596
rect 19426 20584 19432 20596
rect 16868 20556 19432 20584
rect 14642 20516 14648 20528
rect 14214 20488 14648 20516
rect 14642 20476 14648 20488
rect 14700 20476 14706 20528
rect 16868 20457 16896 20556
rect 19426 20544 19432 20556
rect 19484 20544 19490 20596
rect 20898 20544 20904 20596
rect 20956 20544 20962 20596
rect 21453 20587 21511 20593
rect 21453 20584 21465 20587
rect 21008 20556 21465 20584
rect 17126 20476 17132 20528
rect 17184 20476 17190 20528
rect 17770 20476 17776 20528
rect 17828 20476 17834 20528
rect 18782 20476 18788 20528
rect 18840 20516 18846 20528
rect 20809 20519 20867 20525
rect 20809 20516 20821 20519
rect 18840 20488 20821 20516
rect 18840 20476 18846 20488
rect 20809 20485 20821 20488
rect 20855 20516 20867 20519
rect 21008 20516 21036 20556
rect 21453 20553 21465 20556
rect 21499 20553 21511 20587
rect 21453 20547 21511 20553
rect 25314 20544 25320 20596
rect 25372 20544 25378 20596
rect 20855 20488 21036 20516
rect 20855 20485 20867 20488
rect 20809 20479 20867 20485
rect 21082 20476 21088 20528
rect 21140 20516 21146 20528
rect 21140 20488 22968 20516
rect 21140 20476 21146 20488
rect 16853 20451 16911 20457
rect 10336 20420 11008 20448
rect 7742 20340 7748 20392
rect 7800 20340 7806 20392
rect 9766 20340 9772 20392
rect 9824 20340 9830 20392
rect 10226 20340 10232 20392
rect 10284 20380 10290 20392
rect 10980 20389 11008 20420
rect 16853 20417 16865 20451
rect 16899 20417 16911 20451
rect 16853 20411 16911 20417
rect 19245 20451 19303 20457
rect 19245 20417 19257 20451
rect 19291 20448 19303 20451
rect 19518 20448 19524 20460
rect 19291 20420 19524 20448
rect 19291 20417 19303 20420
rect 19245 20411 19303 20417
rect 19518 20408 19524 20420
rect 19576 20408 19582 20460
rect 19889 20451 19947 20457
rect 19889 20417 19901 20451
rect 19935 20417 19947 20451
rect 21818 20448 21824 20460
rect 19889 20411 19947 20417
rect 21008 20420 21824 20448
rect 10873 20383 10931 20389
rect 10873 20380 10885 20383
rect 10284 20352 10885 20380
rect 10284 20340 10290 20352
rect 10873 20349 10885 20352
rect 10919 20349 10931 20383
rect 10873 20343 10931 20349
rect 10965 20383 11023 20389
rect 10965 20349 10977 20383
rect 11011 20349 11023 20383
rect 10965 20343 11023 20349
rect 12710 20340 12716 20392
rect 12768 20340 12774 20392
rect 12989 20383 13047 20389
rect 12989 20349 13001 20383
rect 13035 20380 13047 20383
rect 13446 20380 13452 20392
rect 13035 20352 13452 20380
rect 13035 20349 13047 20352
rect 12989 20343 13047 20349
rect 13446 20340 13452 20352
rect 13504 20380 13510 20392
rect 14366 20380 14372 20392
rect 13504 20352 14372 20380
rect 13504 20340 13510 20352
rect 14366 20340 14372 20352
rect 14424 20340 14430 20392
rect 15565 20383 15623 20389
rect 15565 20380 15577 20383
rect 14476 20352 15577 20380
rect 14476 20256 14504 20352
rect 15565 20349 15577 20352
rect 15611 20349 15623 20383
rect 15565 20343 15623 20349
rect 17218 20340 17224 20392
rect 17276 20380 17282 20392
rect 18506 20380 18512 20392
rect 17276 20352 18512 20380
rect 17276 20340 17282 20352
rect 18506 20340 18512 20352
rect 18564 20380 18570 20392
rect 18601 20383 18659 20389
rect 18601 20380 18613 20383
rect 18564 20352 18613 20380
rect 18564 20340 18570 20352
rect 18601 20349 18613 20352
rect 18647 20349 18659 20383
rect 19904 20380 19932 20411
rect 21008 20380 21036 20420
rect 21818 20408 21824 20420
rect 21876 20408 21882 20460
rect 22186 20408 22192 20460
rect 22244 20408 22250 20460
rect 22940 20457 22968 20488
rect 24118 20476 24124 20528
rect 24176 20516 24182 20528
rect 24176 20488 24334 20516
rect 24176 20476 24182 20488
rect 22925 20451 22983 20457
rect 22925 20417 22937 20451
rect 22971 20417 22983 20451
rect 22925 20411 22983 20417
rect 19904 20352 21036 20380
rect 21085 20383 21143 20389
rect 18601 20343 18659 20349
rect 21085 20349 21097 20383
rect 21131 20380 21143 20383
rect 23382 20380 23388 20392
rect 21131 20352 23388 20380
rect 21131 20349 21143 20352
rect 21085 20343 21143 20349
rect 23382 20340 23388 20352
rect 23440 20340 23446 20392
rect 23566 20340 23572 20392
rect 23624 20340 23630 20392
rect 23845 20383 23903 20389
rect 23845 20349 23857 20383
rect 23891 20380 23903 20383
rect 25130 20380 25136 20392
rect 23891 20352 25136 20380
rect 23891 20349 23903 20352
rect 23845 20343 23903 20349
rect 25130 20340 25136 20352
rect 25188 20340 25194 20392
rect 19150 20312 19156 20324
rect 18524 20284 19156 20312
rect 14458 20204 14464 20256
rect 14516 20204 14522 20256
rect 15013 20247 15071 20253
rect 15013 20213 15025 20247
rect 15059 20244 15071 20247
rect 18524 20244 18552 20284
rect 19150 20272 19156 20284
rect 19208 20272 19214 20324
rect 22005 20315 22063 20321
rect 22005 20281 22017 20315
rect 22051 20312 22063 20315
rect 22051 20284 23704 20312
rect 22051 20281 22063 20284
rect 22005 20275 22063 20281
rect 23676 20256 23704 20284
rect 15059 20216 18552 20244
rect 15059 20213 15071 20216
rect 15013 20207 15071 20213
rect 19058 20204 19064 20256
rect 19116 20204 19122 20256
rect 19518 20204 19524 20256
rect 19576 20244 19582 20256
rect 19705 20247 19763 20253
rect 19705 20244 19717 20247
rect 19576 20216 19717 20244
rect 19576 20204 19582 20216
rect 19705 20213 19717 20216
rect 19751 20213 19763 20247
rect 19705 20207 19763 20213
rect 20441 20247 20499 20253
rect 20441 20213 20453 20247
rect 20487 20244 20499 20247
rect 21266 20244 21272 20256
rect 20487 20216 21272 20244
rect 20487 20213 20499 20216
rect 20441 20207 20499 20213
rect 21266 20204 21272 20216
rect 21324 20204 21330 20256
rect 22738 20204 22744 20256
rect 22796 20204 22802 20256
rect 23658 20204 23664 20256
rect 23716 20204 23722 20256
rect 1104 20154 25852 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 25852 20154
rect 1104 20080 25852 20102
rect 8386 20000 8392 20052
rect 8444 20040 8450 20052
rect 8481 20043 8539 20049
rect 8481 20040 8493 20043
rect 8444 20012 8493 20040
rect 8444 20000 8450 20012
rect 8481 20009 8493 20012
rect 8527 20040 8539 20043
rect 9030 20040 9036 20052
rect 8527 20012 9036 20040
rect 8527 20009 8539 20012
rect 8481 20003 8539 20009
rect 9030 20000 9036 20012
rect 9088 20000 9094 20052
rect 11333 20043 11391 20049
rect 11333 20009 11345 20043
rect 11379 20040 11391 20043
rect 13998 20040 14004 20052
rect 11379 20012 14004 20040
rect 11379 20009 11391 20012
rect 11333 20003 11391 20009
rect 13998 20000 14004 20012
rect 14056 20000 14062 20052
rect 15746 20000 15752 20052
rect 15804 20040 15810 20052
rect 16025 20043 16083 20049
rect 16025 20040 16037 20043
rect 15804 20012 16037 20040
rect 15804 20000 15810 20012
rect 16025 20009 16037 20012
rect 16071 20009 16083 20043
rect 16025 20003 16083 20009
rect 16485 20043 16543 20049
rect 16485 20009 16497 20043
rect 16531 20040 16543 20043
rect 22186 20040 22192 20052
rect 16531 20012 22192 20040
rect 16531 20009 16543 20012
rect 16485 20003 16543 20009
rect 22186 20000 22192 20012
rect 22244 20000 22250 20052
rect 23845 20043 23903 20049
rect 23845 20009 23857 20043
rect 23891 20040 23903 20043
rect 23934 20040 23940 20052
rect 23891 20012 23940 20040
rect 23891 20009 23903 20012
rect 23845 20003 23903 20009
rect 23934 20000 23940 20012
rect 23992 20000 23998 20052
rect 17126 19932 17132 19984
rect 17184 19972 17190 19984
rect 17184 19944 18092 19972
rect 17184 19932 17190 19944
rect 10686 19904 10692 19916
rect 9140 19876 10692 19904
rect 7742 19796 7748 19848
rect 7800 19836 7806 19848
rect 9030 19836 9036 19848
rect 7800 19808 9036 19836
rect 7800 19796 7806 19808
rect 9030 19796 9036 19808
rect 9088 19836 9094 19848
rect 9140 19845 9168 19876
rect 10686 19864 10692 19876
rect 10744 19864 10750 19916
rect 11974 19864 11980 19916
rect 12032 19864 12038 19916
rect 14550 19864 14556 19916
rect 14608 19864 14614 19916
rect 14642 19864 14648 19916
rect 14700 19904 14706 19916
rect 16945 19907 17003 19913
rect 16945 19904 16957 19907
rect 14700 19876 16957 19904
rect 14700 19864 14706 19876
rect 16945 19873 16957 19876
rect 16991 19904 17003 19907
rect 17770 19904 17776 19916
rect 16991 19876 17776 19904
rect 16991 19873 17003 19876
rect 16945 19867 17003 19873
rect 17770 19864 17776 19876
rect 17828 19864 17834 19916
rect 17954 19864 17960 19916
rect 18012 19864 18018 19916
rect 18064 19913 18092 19944
rect 18049 19907 18107 19913
rect 18049 19873 18061 19907
rect 18095 19873 18107 19907
rect 18049 19867 18107 19873
rect 19889 19907 19947 19913
rect 19889 19873 19901 19907
rect 19935 19904 19947 19907
rect 20254 19904 20260 19916
rect 19935 19876 20260 19904
rect 19935 19873 19947 19876
rect 19889 19867 19947 19873
rect 20254 19864 20260 19876
rect 20312 19904 20318 19916
rect 22097 19907 22155 19913
rect 22097 19904 22109 19907
rect 20312 19876 22109 19904
rect 20312 19864 20318 19876
rect 22097 19873 22109 19876
rect 22143 19873 22155 19907
rect 22097 19867 22155 19873
rect 22830 19864 22836 19916
rect 22888 19904 22894 19916
rect 23106 19904 23112 19916
rect 22888 19876 23112 19904
rect 22888 19864 22894 19876
rect 23106 19864 23112 19876
rect 23164 19904 23170 19916
rect 24397 19907 24455 19913
rect 24397 19904 24409 19907
rect 23164 19876 24409 19904
rect 23164 19864 23170 19876
rect 24397 19873 24409 19876
rect 24443 19904 24455 19907
rect 24854 19904 24860 19916
rect 24443 19876 24860 19904
rect 24443 19873 24455 19876
rect 24397 19867 24455 19873
rect 24854 19864 24860 19876
rect 24912 19864 24918 19916
rect 9125 19839 9183 19845
rect 9125 19836 9137 19839
rect 9088 19808 9137 19836
rect 9088 19796 9094 19808
rect 9125 19805 9137 19808
rect 9171 19805 9183 19839
rect 9125 19799 9183 19805
rect 12710 19796 12716 19848
rect 12768 19836 12774 19848
rect 14277 19839 14335 19845
rect 14277 19836 14289 19839
rect 12768 19808 14289 19836
rect 12768 19796 12774 19808
rect 14277 19805 14289 19808
rect 14323 19805 14335 19839
rect 14277 19799 14335 19805
rect 15838 19796 15844 19848
rect 15896 19836 15902 19848
rect 16669 19839 16727 19845
rect 16669 19836 16681 19839
rect 15896 19808 16681 19836
rect 15896 19796 15902 19808
rect 16669 19805 16681 19808
rect 16715 19805 16727 19839
rect 17865 19839 17923 19845
rect 17865 19836 17877 19839
rect 16669 19799 16727 19805
rect 16776 19808 17877 19836
rect 8294 19728 8300 19780
rect 8352 19768 8358 19780
rect 9398 19768 9404 19780
rect 8352 19740 9404 19768
rect 8352 19728 8358 19740
rect 9398 19728 9404 19740
rect 9456 19728 9462 19780
rect 9600 19740 9890 19768
rect 9600 19712 9628 19740
rect 11238 19728 11244 19780
rect 11296 19768 11302 19780
rect 11793 19771 11851 19777
rect 11793 19768 11805 19771
rect 11296 19740 11805 19768
rect 11296 19728 11302 19740
rect 11793 19737 11805 19740
rect 11839 19737 11851 19771
rect 11793 19731 11851 19737
rect 14642 19728 14648 19780
rect 14700 19768 14706 19780
rect 14700 19740 15042 19768
rect 14700 19728 14706 19740
rect 15930 19728 15936 19780
rect 15988 19768 15994 19780
rect 16776 19768 16804 19808
rect 17865 19805 17877 19808
rect 17911 19805 17923 19839
rect 17865 19799 17923 19805
rect 18877 19839 18935 19845
rect 18877 19805 18889 19839
rect 18923 19836 18935 19839
rect 19610 19836 19616 19848
rect 18923 19808 19616 19836
rect 18923 19805 18935 19808
rect 18877 19799 18935 19805
rect 19610 19796 19616 19808
rect 19668 19796 19674 19848
rect 21542 19836 21548 19848
rect 21298 19808 21548 19836
rect 21542 19796 21548 19808
rect 21600 19836 21606 19848
rect 21818 19836 21824 19848
rect 21600 19808 21824 19836
rect 21600 19796 21606 19808
rect 21818 19796 21824 19808
rect 21876 19796 21882 19848
rect 19794 19768 19800 19780
rect 15988 19740 16804 19768
rect 18432 19740 19800 19768
rect 15988 19728 15994 19740
rect 9582 19660 9588 19712
rect 9640 19660 9646 19712
rect 10870 19660 10876 19712
rect 10928 19660 10934 19712
rect 11698 19660 11704 19712
rect 11756 19660 11762 19712
rect 14550 19660 14556 19712
rect 14608 19700 14614 19712
rect 15378 19700 15384 19712
rect 14608 19672 15384 19700
rect 14608 19660 14614 19672
rect 15378 19660 15384 19672
rect 15436 19660 15442 19712
rect 17497 19703 17555 19709
rect 17497 19669 17509 19703
rect 17543 19700 17555 19703
rect 18432 19700 18460 19740
rect 19794 19728 19800 19740
rect 19852 19728 19858 19780
rect 20162 19728 20168 19780
rect 20220 19728 20226 19780
rect 22373 19771 22431 19777
rect 22373 19768 22385 19771
rect 21652 19740 22385 19768
rect 21652 19712 21680 19740
rect 22373 19737 22385 19740
rect 22419 19737 22431 19771
rect 22373 19731 22431 19737
rect 22572 19740 22862 19768
rect 17543 19672 18460 19700
rect 17543 19669 17555 19672
rect 17497 19663 17555 19669
rect 18506 19660 18512 19712
rect 18564 19700 18570 19712
rect 18693 19703 18751 19709
rect 18693 19700 18705 19703
rect 18564 19672 18705 19700
rect 18564 19660 18570 19672
rect 18693 19669 18705 19672
rect 18739 19669 18751 19703
rect 18693 19663 18751 19669
rect 21634 19660 21640 19712
rect 21692 19660 21698 19712
rect 21818 19660 21824 19712
rect 21876 19700 21882 19712
rect 22572 19700 22600 19740
rect 21876 19672 22600 19700
rect 22756 19700 22784 19740
rect 24118 19700 24124 19712
rect 22756 19672 24124 19700
rect 21876 19660 21882 19672
rect 24118 19660 24124 19672
rect 24176 19700 24182 19712
rect 25406 19700 25412 19712
rect 24176 19672 25412 19700
rect 24176 19660 24182 19672
rect 25406 19660 25412 19672
rect 25464 19660 25470 19712
rect 1104 19610 25852 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 25852 19610
rect 1104 19536 25852 19558
rect 8754 19456 8760 19508
rect 8812 19456 8818 19508
rect 9582 19456 9588 19508
rect 9640 19496 9646 19508
rect 10965 19499 11023 19505
rect 10965 19496 10977 19499
rect 9640 19468 10977 19496
rect 9640 19456 9646 19468
rect 10965 19465 10977 19468
rect 11011 19465 11023 19499
rect 10965 19459 11023 19465
rect 8386 19428 8392 19440
rect 8050 19400 8392 19428
rect 8386 19388 8392 19400
rect 8444 19428 8450 19440
rect 8662 19428 8668 19440
rect 8444 19400 8668 19428
rect 8444 19388 8450 19400
rect 8662 19388 8668 19400
rect 8720 19388 8726 19440
rect 9125 19431 9183 19437
rect 9125 19397 9137 19431
rect 9171 19428 9183 19431
rect 9214 19428 9220 19440
rect 9171 19400 9220 19428
rect 9171 19397 9183 19400
rect 9125 19391 9183 19397
rect 9214 19388 9220 19400
rect 9272 19388 9278 19440
rect 10134 19360 10140 19372
rect 9232 19332 10140 19360
rect 6546 19252 6552 19304
rect 6604 19252 6610 19304
rect 6825 19295 6883 19301
rect 6825 19261 6837 19295
rect 6871 19292 6883 19295
rect 6914 19292 6920 19304
rect 6871 19264 6920 19292
rect 6871 19261 6883 19264
rect 6825 19255 6883 19261
rect 6914 19252 6920 19264
rect 6972 19252 6978 19304
rect 9232 19301 9260 19332
rect 10134 19320 10140 19332
rect 10192 19320 10198 19372
rect 10980 19360 11008 19459
rect 11698 19456 11704 19508
rect 11756 19456 11762 19508
rect 11790 19456 11796 19508
rect 11848 19496 11854 19508
rect 11848 19468 15240 19496
rect 11848 19456 11854 19468
rect 14642 19428 14648 19440
rect 14030 19400 14648 19428
rect 14642 19388 14648 19400
rect 14700 19388 14706 19440
rect 15212 19369 15240 19468
rect 15286 19456 15292 19508
rect 15344 19496 15350 19508
rect 15933 19499 15991 19505
rect 15933 19496 15945 19499
rect 15344 19468 15945 19496
rect 15344 19456 15350 19468
rect 15933 19465 15945 19468
rect 15979 19465 15991 19499
rect 15933 19459 15991 19465
rect 16853 19499 16911 19505
rect 16853 19465 16865 19499
rect 16899 19465 16911 19499
rect 16853 19459 16911 19465
rect 16868 19428 16896 19459
rect 17310 19456 17316 19508
rect 17368 19456 17374 19508
rect 18969 19499 19027 19505
rect 18969 19465 18981 19499
rect 19015 19465 19027 19499
rect 18969 19459 19027 19465
rect 18984 19428 19012 19459
rect 19242 19456 19248 19508
rect 19300 19496 19306 19508
rect 20073 19499 20131 19505
rect 20073 19496 20085 19499
rect 19300 19468 20085 19496
rect 19300 19456 19306 19468
rect 20073 19465 20085 19468
rect 20119 19465 20131 19499
rect 20073 19459 20131 19465
rect 20438 19456 20444 19508
rect 20496 19456 20502 19508
rect 20533 19499 20591 19505
rect 20533 19465 20545 19499
rect 20579 19496 20591 19499
rect 20714 19496 20720 19508
rect 20579 19468 20720 19496
rect 20579 19465 20591 19468
rect 20533 19459 20591 19465
rect 20714 19456 20720 19468
rect 20772 19456 20778 19508
rect 22189 19499 22247 19505
rect 22189 19465 22201 19499
rect 22235 19496 22247 19499
rect 22462 19496 22468 19508
rect 22235 19468 22468 19496
rect 22235 19465 22247 19468
rect 22189 19459 22247 19465
rect 22462 19456 22468 19468
rect 22520 19456 22526 19508
rect 22554 19456 22560 19508
rect 22612 19496 22618 19508
rect 22649 19499 22707 19505
rect 22649 19496 22661 19499
rect 22612 19468 22661 19496
rect 22612 19456 22618 19468
rect 22649 19465 22661 19468
rect 22695 19465 22707 19499
rect 22649 19459 22707 19465
rect 25130 19456 25136 19508
rect 25188 19456 25194 19508
rect 25406 19456 25412 19508
rect 25464 19456 25470 19508
rect 21542 19428 21548 19440
rect 16868 19400 18920 19428
rect 18984 19400 21548 19428
rect 15197 19363 15255 19369
rect 10980 19332 11100 19360
rect 9217 19295 9275 19301
rect 9217 19261 9229 19295
rect 9263 19261 9275 19295
rect 9217 19255 9275 19261
rect 9309 19295 9367 19301
rect 9309 19261 9321 19295
rect 9355 19261 9367 19295
rect 11072 19292 11100 19332
rect 15197 19329 15209 19363
rect 15243 19329 15255 19363
rect 15562 19360 15568 19372
rect 15197 19323 15255 19329
rect 15304 19332 15568 19360
rect 11422 19292 11428 19304
rect 11072 19264 11428 19292
rect 9309 19255 9367 19261
rect 8570 19184 8576 19236
rect 8628 19224 8634 19236
rect 9324 19224 9352 19255
rect 11422 19252 11428 19264
rect 11480 19252 11486 19304
rect 12529 19295 12587 19301
rect 12529 19261 12541 19295
rect 12575 19261 12587 19295
rect 12529 19255 12587 19261
rect 12805 19295 12863 19301
rect 12805 19261 12817 19295
rect 12851 19292 12863 19295
rect 14458 19292 14464 19304
rect 12851 19264 14464 19292
rect 12851 19261 12863 19264
rect 12805 19255 12863 19261
rect 8628 19196 9352 19224
rect 8628 19184 8634 19196
rect 8297 19159 8355 19165
rect 8297 19125 8309 19159
rect 8343 19156 8355 19159
rect 8386 19156 8392 19168
rect 8343 19128 8392 19156
rect 8343 19125 8355 19128
rect 8297 19119 8355 19125
rect 8386 19116 8392 19128
rect 8444 19116 8450 19168
rect 11238 19116 11244 19168
rect 11296 19116 11302 19168
rect 12544 19156 12572 19255
rect 14458 19252 14464 19264
rect 14516 19252 14522 19304
rect 15013 19227 15071 19233
rect 15013 19193 15025 19227
rect 15059 19224 15071 19227
rect 15304 19224 15332 19332
rect 15562 19320 15568 19332
rect 15620 19320 15626 19372
rect 16117 19363 16175 19369
rect 16117 19329 16129 19363
rect 16163 19360 16175 19363
rect 16482 19360 16488 19372
rect 16163 19332 16488 19360
rect 16163 19329 16175 19332
rect 16117 19323 16175 19329
rect 16482 19320 16488 19332
rect 16540 19320 16546 19372
rect 16666 19320 16672 19372
rect 16724 19360 16730 19372
rect 17221 19363 17279 19369
rect 17221 19360 17233 19363
rect 16724 19332 17233 19360
rect 16724 19320 16730 19332
rect 17221 19329 17233 19332
rect 17267 19329 17279 19363
rect 18892 19360 18920 19400
rect 21542 19388 21548 19400
rect 21600 19388 21606 19440
rect 23566 19428 23572 19440
rect 23400 19400 23572 19428
rect 18892 19332 19104 19360
rect 17221 19323 17279 19329
rect 15746 19252 15752 19304
rect 15804 19292 15810 19304
rect 17405 19295 17463 19301
rect 17405 19292 17417 19295
rect 15804 19264 17417 19292
rect 15804 19252 15810 19264
rect 17405 19261 17417 19264
rect 17451 19261 17463 19295
rect 19076 19292 19104 19332
rect 19150 19320 19156 19372
rect 19208 19320 19214 19372
rect 23400 19369 23428 19400
rect 23566 19388 23572 19400
rect 23624 19388 23630 19440
rect 23661 19431 23719 19437
rect 23661 19397 23673 19431
rect 23707 19428 23719 19431
rect 23934 19428 23940 19440
rect 23707 19400 23940 19428
rect 23707 19397 23719 19400
rect 23661 19391 23719 19397
rect 23934 19388 23940 19400
rect 23992 19388 23998 19440
rect 24118 19388 24124 19440
rect 24176 19388 24182 19440
rect 21269 19363 21327 19369
rect 21269 19329 21281 19363
rect 21315 19360 21327 19363
rect 22557 19363 22615 19369
rect 22557 19360 22569 19363
rect 21315 19332 22569 19360
rect 21315 19329 21327 19332
rect 21269 19323 21327 19329
rect 22557 19329 22569 19332
rect 22603 19329 22615 19363
rect 22557 19323 22615 19329
rect 23385 19363 23443 19369
rect 23385 19329 23397 19363
rect 23431 19329 23443 19363
rect 23385 19323 23443 19329
rect 19334 19292 19340 19304
rect 19076 19264 19340 19292
rect 17405 19255 17463 19261
rect 19334 19252 19340 19264
rect 19392 19252 19398 19304
rect 20717 19295 20775 19301
rect 20717 19261 20729 19295
rect 20763 19292 20775 19295
rect 21634 19292 21640 19304
rect 20763 19264 21640 19292
rect 20763 19261 20775 19264
rect 20717 19255 20775 19261
rect 21634 19252 21640 19264
rect 21692 19252 21698 19304
rect 22833 19295 22891 19301
rect 22833 19261 22845 19295
rect 22879 19292 22891 19295
rect 23290 19292 23296 19304
rect 22879 19264 23296 19292
rect 22879 19261 22891 19264
rect 22833 19255 22891 19261
rect 23290 19252 23296 19264
rect 23348 19252 23354 19304
rect 15059 19196 15332 19224
rect 15059 19193 15071 19196
rect 15013 19187 15071 19193
rect 12802 19156 12808 19168
rect 12544 19128 12808 19156
rect 12802 19116 12808 19128
rect 12860 19116 12866 19168
rect 14277 19159 14335 19165
rect 14277 19125 14289 19159
rect 14323 19156 14335 19159
rect 14366 19156 14372 19168
rect 14323 19128 14372 19156
rect 14323 19125 14335 19128
rect 14277 19119 14335 19125
rect 14366 19116 14372 19128
rect 14424 19116 14430 19168
rect 14642 19116 14648 19168
rect 14700 19116 14706 19168
rect 20990 19116 20996 19168
rect 21048 19156 21054 19168
rect 21818 19156 21824 19168
rect 21048 19128 21824 19156
rect 21048 19116 21054 19128
rect 21818 19116 21824 19128
rect 21876 19116 21882 19168
rect 1104 19066 25852 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 25852 19066
rect 1104 18992 25852 19014
rect 8662 18912 8668 18964
rect 8720 18912 8726 18964
rect 10042 18912 10048 18964
rect 10100 18912 10106 18964
rect 11517 18955 11575 18961
rect 11517 18921 11529 18955
rect 11563 18952 11575 18955
rect 15838 18952 15844 18964
rect 11563 18924 15844 18952
rect 11563 18921 11575 18924
rect 11517 18915 11575 18921
rect 15838 18912 15844 18924
rect 15896 18912 15902 18964
rect 16850 18912 16856 18964
rect 16908 18952 16914 18964
rect 25958 18952 25964 18964
rect 16908 18924 25964 18952
rect 16908 18912 16914 18924
rect 25958 18912 25964 18924
rect 26016 18912 26022 18964
rect 9950 18844 9956 18896
rect 10008 18884 10014 18896
rect 12713 18887 12771 18893
rect 12713 18884 12725 18887
rect 10008 18856 12725 18884
rect 10008 18844 10014 18856
rect 12713 18853 12725 18856
rect 12759 18853 12771 18887
rect 24486 18884 24492 18896
rect 12713 18847 12771 18853
rect 21468 18856 24492 18884
rect 6917 18819 6975 18825
rect 6917 18785 6929 18819
rect 6963 18816 6975 18819
rect 8386 18816 8392 18828
rect 6963 18788 8392 18816
rect 6963 18785 6975 18788
rect 6917 18779 6975 18785
rect 8386 18776 8392 18788
rect 8444 18776 8450 18828
rect 9674 18776 9680 18828
rect 9732 18816 9738 18828
rect 10594 18816 10600 18828
rect 9732 18788 10600 18816
rect 9732 18776 9738 18788
rect 10594 18776 10600 18788
rect 10652 18776 10658 18828
rect 10870 18776 10876 18828
rect 10928 18816 10934 18828
rect 12069 18819 12127 18825
rect 12069 18816 12081 18819
rect 10928 18788 12081 18816
rect 10928 18776 10934 18788
rect 12069 18785 12081 18788
rect 12115 18785 12127 18819
rect 13265 18819 13323 18825
rect 13265 18816 13277 18819
rect 12069 18779 12127 18785
rect 12268 18788 13277 18816
rect 6638 18708 6644 18760
rect 6696 18708 6702 18760
rect 8662 18748 8668 18760
rect 8050 18720 8668 18748
rect 8662 18708 8668 18720
rect 8720 18708 8726 18760
rect 8846 18708 8852 18760
rect 8904 18748 8910 18760
rect 9398 18748 9404 18760
rect 8904 18720 9404 18748
rect 8904 18708 8910 18720
rect 9398 18708 9404 18720
rect 9456 18748 9462 18760
rect 11977 18751 12035 18757
rect 9456 18720 11928 18748
rect 9456 18708 9462 18720
rect 9582 18680 9588 18692
rect 8220 18652 9588 18680
rect 7006 18572 7012 18624
rect 7064 18612 7070 18624
rect 8220 18612 8248 18652
rect 9582 18640 9588 18652
rect 9640 18640 9646 18692
rect 10594 18640 10600 18692
rect 10652 18680 10658 18692
rect 11698 18680 11704 18692
rect 10652 18652 11704 18680
rect 10652 18640 10658 18652
rect 11698 18640 11704 18652
rect 11756 18640 11762 18692
rect 11900 18680 11928 18720
rect 11977 18717 11989 18751
rect 12023 18748 12035 18751
rect 12158 18748 12164 18760
rect 12023 18720 12164 18748
rect 12023 18717 12035 18720
rect 11977 18711 12035 18717
rect 12158 18708 12164 18720
rect 12216 18708 12222 18760
rect 12268 18680 12296 18788
rect 13265 18785 13277 18788
rect 13311 18785 13323 18819
rect 13265 18779 13323 18785
rect 16942 18776 16948 18828
rect 17000 18816 17006 18828
rect 17497 18819 17555 18825
rect 17000 18788 17264 18816
rect 17000 18776 17006 18788
rect 12526 18708 12532 18760
rect 12584 18748 12590 18760
rect 17236 18757 17264 18788
rect 17497 18785 17509 18819
rect 17543 18816 17555 18819
rect 17770 18816 17776 18828
rect 17543 18788 17776 18816
rect 17543 18785 17555 18788
rect 17497 18779 17555 18785
rect 17770 18776 17776 18788
rect 17828 18776 17834 18828
rect 13173 18751 13231 18757
rect 13173 18748 13185 18751
rect 12584 18720 13185 18748
rect 12584 18708 12590 18720
rect 13173 18717 13185 18720
rect 13219 18717 13231 18751
rect 13173 18711 13231 18717
rect 17221 18751 17279 18757
rect 17221 18717 17233 18751
rect 17267 18748 17279 18751
rect 17310 18748 17316 18760
rect 17267 18720 17316 18748
rect 17267 18717 17279 18720
rect 17221 18711 17279 18717
rect 17310 18708 17316 18720
rect 17368 18748 17374 18760
rect 21468 18757 21496 18856
rect 24486 18844 24492 18856
rect 24544 18844 24550 18896
rect 23842 18776 23848 18828
rect 23900 18776 23906 18828
rect 17865 18751 17923 18757
rect 17865 18748 17877 18751
rect 17368 18720 17877 18748
rect 17368 18708 17374 18720
rect 17865 18717 17877 18720
rect 17911 18717 17923 18751
rect 17865 18711 17923 18717
rect 21453 18751 21511 18757
rect 21453 18717 21465 18751
rect 21499 18717 21511 18751
rect 21453 18711 21511 18717
rect 21542 18708 21548 18760
rect 21600 18748 21606 18760
rect 22189 18751 22247 18757
rect 22189 18748 22201 18751
rect 21600 18720 22201 18748
rect 21600 18708 21606 18720
rect 22189 18717 22201 18720
rect 22235 18717 22247 18751
rect 22189 18711 22247 18717
rect 22738 18708 22744 18760
rect 22796 18708 22802 18760
rect 24673 18751 24731 18757
rect 24673 18717 24685 18751
rect 24719 18748 24731 18751
rect 26602 18748 26608 18760
rect 24719 18720 26608 18748
rect 24719 18717 24731 18720
rect 24673 18711 24731 18717
rect 26602 18708 26608 18720
rect 26660 18708 26666 18760
rect 11900 18652 12296 18680
rect 12434 18640 12440 18692
rect 12492 18680 12498 18692
rect 13817 18683 13875 18689
rect 13817 18680 13829 18683
rect 12492 18652 13829 18680
rect 12492 18640 12498 18652
rect 13817 18649 13829 18652
rect 13863 18680 13875 18683
rect 16942 18680 16948 18692
rect 13863 18652 16948 18680
rect 13863 18649 13875 18652
rect 13817 18643 13875 18649
rect 16942 18640 16948 18652
rect 17000 18680 17006 18692
rect 17678 18680 17684 18692
rect 17000 18652 17684 18680
rect 17000 18640 17006 18652
rect 17678 18640 17684 18652
rect 17736 18640 17742 18692
rect 24857 18683 24915 18689
rect 24857 18649 24869 18683
rect 24903 18680 24915 18683
rect 25406 18680 25412 18692
rect 24903 18652 25412 18680
rect 24903 18649 24915 18652
rect 24857 18643 24915 18649
rect 25406 18640 25412 18652
rect 25464 18640 25470 18692
rect 7064 18584 8248 18612
rect 7064 18572 7070 18584
rect 8294 18572 8300 18624
rect 8352 18612 8358 18624
rect 8389 18615 8447 18621
rect 8389 18612 8401 18615
rect 8352 18584 8401 18612
rect 8352 18572 8358 18584
rect 8389 18581 8401 18584
rect 8435 18581 8447 18615
rect 8389 18575 8447 18581
rect 8938 18572 8944 18624
rect 8996 18612 9002 18624
rect 9677 18615 9735 18621
rect 9677 18612 9689 18615
rect 8996 18584 9689 18612
rect 8996 18572 9002 18584
rect 9677 18581 9689 18584
rect 9723 18612 9735 18615
rect 10413 18615 10471 18621
rect 10413 18612 10425 18615
rect 9723 18584 10425 18612
rect 9723 18581 9735 18584
rect 9677 18575 9735 18581
rect 10413 18581 10425 18584
rect 10459 18581 10471 18615
rect 10413 18575 10471 18581
rect 10502 18572 10508 18624
rect 10560 18572 10566 18624
rect 11330 18572 11336 18624
rect 11388 18612 11394 18624
rect 11885 18615 11943 18621
rect 11885 18612 11897 18615
rect 11388 18584 11897 18612
rect 11388 18572 11394 18584
rect 11885 18581 11897 18584
rect 11931 18581 11943 18615
rect 11885 18575 11943 18581
rect 12618 18572 12624 18624
rect 12676 18612 12682 18624
rect 13081 18615 13139 18621
rect 13081 18612 13093 18615
rect 12676 18584 13093 18612
rect 12676 18572 12682 18584
rect 13081 18581 13093 18584
rect 13127 18581 13139 18615
rect 13081 18575 13139 18581
rect 14274 18572 14280 18624
rect 14332 18572 14338 18624
rect 16758 18572 16764 18624
rect 16816 18612 16822 18624
rect 16853 18615 16911 18621
rect 16853 18612 16865 18615
rect 16816 18584 16865 18612
rect 16816 18572 16822 18584
rect 16853 18581 16865 18584
rect 16899 18581 16911 18615
rect 16853 18575 16911 18581
rect 17313 18615 17371 18621
rect 17313 18581 17325 18615
rect 17359 18612 17371 18615
rect 17586 18612 17592 18624
rect 17359 18584 17592 18612
rect 17359 18581 17371 18584
rect 17313 18575 17371 18581
rect 17586 18572 17592 18584
rect 17644 18612 17650 18624
rect 18049 18615 18107 18621
rect 18049 18612 18061 18615
rect 17644 18584 18061 18612
rect 17644 18572 17650 18584
rect 18049 18581 18061 18584
rect 18095 18581 18107 18615
rect 18049 18575 18107 18581
rect 21269 18615 21327 18621
rect 21269 18581 21281 18615
rect 21315 18612 21327 18615
rect 21358 18612 21364 18624
rect 21315 18584 21364 18612
rect 21315 18581 21327 18584
rect 21269 18575 21327 18581
rect 21358 18572 21364 18584
rect 21416 18572 21422 18624
rect 22005 18615 22063 18621
rect 22005 18581 22017 18615
rect 22051 18612 22063 18615
rect 22094 18612 22100 18624
rect 22051 18584 22100 18612
rect 22051 18581 22063 18584
rect 22005 18575 22063 18581
rect 22094 18572 22100 18584
rect 22152 18572 22158 18624
rect 1104 18522 25852 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 25852 18522
rect 1104 18448 25852 18470
rect 10042 18408 10048 18420
rect 8036 18380 10048 18408
rect 8036 18349 8064 18380
rect 10042 18368 10048 18380
rect 10100 18368 10106 18420
rect 10410 18368 10416 18420
rect 10468 18368 10474 18420
rect 10502 18368 10508 18420
rect 10560 18408 10566 18420
rect 13817 18411 13875 18417
rect 13817 18408 13829 18411
rect 10560 18380 13829 18408
rect 10560 18368 10566 18380
rect 13817 18377 13829 18380
rect 13863 18377 13875 18411
rect 13817 18371 13875 18377
rect 14185 18411 14243 18417
rect 14185 18377 14197 18411
rect 14231 18408 14243 18411
rect 14921 18411 14979 18417
rect 14921 18408 14933 18411
rect 14231 18380 14933 18408
rect 14231 18377 14243 18380
rect 14185 18371 14243 18377
rect 14921 18377 14933 18380
rect 14967 18408 14979 18411
rect 16850 18408 16856 18420
rect 14967 18380 16856 18408
rect 14967 18377 14979 18380
rect 14921 18371 14979 18377
rect 16850 18368 16856 18380
rect 16908 18368 16914 18420
rect 8021 18343 8079 18349
rect 8021 18309 8033 18343
rect 8067 18309 8079 18343
rect 8021 18303 8079 18309
rect 8662 18300 8668 18352
rect 8720 18300 8726 18352
rect 10060 18340 10088 18368
rect 11057 18343 11115 18349
rect 10060 18312 11008 18340
rect 9582 18232 9588 18284
rect 9640 18272 9646 18284
rect 10321 18275 10379 18281
rect 10321 18272 10333 18275
rect 9640 18244 10333 18272
rect 9640 18232 9646 18244
rect 10321 18241 10333 18244
rect 10367 18241 10379 18275
rect 10321 18235 10379 18241
rect 6638 18164 6644 18216
rect 6696 18204 6702 18216
rect 7745 18207 7803 18213
rect 7745 18204 7757 18207
rect 6696 18176 7757 18204
rect 6696 18164 6702 18176
rect 7745 18173 7757 18176
rect 7791 18204 7803 18207
rect 7791 18176 7880 18204
rect 7791 18173 7803 18176
rect 7745 18167 7803 18173
rect 7852 18068 7880 18176
rect 8386 18164 8392 18216
rect 8444 18204 8450 18216
rect 10505 18207 10563 18213
rect 10505 18204 10517 18207
rect 8444 18176 10517 18204
rect 8444 18164 8450 18176
rect 10505 18173 10517 18176
rect 10551 18173 10563 18207
rect 10980 18204 11008 18312
rect 11057 18309 11069 18343
rect 11103 18340 11115 18343
rect 11422 18340 11428 18352
rect 11103 18312 11428 18340
rect 11103 18309 11115 18312
rect 11057 18303 11115 18309
rect 11422 18300 11428 18312
rect 11480 18300 11486 18352
rect 11606 18300 11612 18352
rect 11664 18340 11670 18352
rect 12434 18340 12440 18352
rect 11664 18312 12440 18340
rect 11664 18300 11670 18312
rect 12434 18300 12440 18312
rect 12492 18300 12498 18352
rect 17034 18300 17040 18352
rect 17092 18340 17098 18352
rect 17129 18343 17187 18349
rect 17129 18340 17141 18343
rect 17092 18312 17141 18340
rect 17092 18300 17098 18312
rect 17129 18309 17141 18312
rect 17175 18340 17187 18343
rect 17218 18340 17224 18352
rect 17175 18312 17224 18340
rect 17175 18309 17187 18312
rect 17129 18303 17187 18309
rect 17218 18300 17224 18312
rect 17276 18300 17282 18352
rect 22186 18340 22192 18352
rect 21284 18312 22192 18340
rect 13538 18272 13544 18284
rect 12728 18244 13544 18272
rect 12728 18204 12756 18244
rect 13538 18232 13544 18244
rect 13596 18232 13602 18284
rect 16298 18232 16304 18284
rect 16356 18232 16362 18284
rect 16574 18232 16580 18284
rect 16632 18272 16638 18284
rect 21284 18281 21312 18312
rect 22186 18300 22192 18312
rect 22244 18300 22250 18352
rect 23293 18343 23351 18349
rect 23293 18309 23305 18343
rect 23339 18340 23351 18343
rect 24854 18340 24860 18352
rect 23339 18312 24860 18340
rect 23339 18309 23351 18312
rect 23293 18303 23351 18309
rect 24854 18300 24860 18312
rect 24912 18300 24918 18352
rect 16853 18275 16911 18281
rect 16853 18272 16865 18275
rect 16632 18244 16865 18272
rect 16632 18232 16638 18244
rect 16853 18241 16865 18244
rect 16899 18241 16911 18275
rect 21269 18275 21327 18281
rect 18262 18244 19012 18272
rect 16853 18235 16911 18241
rect 10980 18176 12756 18204
rect 10505 18167 10563 18173
rect 12802 18164 12808 18216
rect 12860 18204 12866 18216
rect 13173 18207 13231 18213
rect 13173 18204 13185 18207
rect 12860 18176 13185 18204
rect 12860 18164 12866 18176
rect 13173 18173 13185 18176
rect 13219 18173 13231 18207
rect 13173 18167 13231 18173
rect 14090 18164 14096 18216
rect 14148 18204 14154 18216
rect 14277 18207 14335 18213
rect 14277 18204 14289 18207
rect 14148 18176 14289 18204
rect 14148 18164 14154 18176
rect 14277 18173 14289 18176
rect 14323 18173 14335 18207
rect 14277 18167 14335 18173
rect 14458 18164 14464 18216
rect 14516 18164 14522 18216
rect 9030 18096 9036 18148
rect 9088 18136 9094 18148
rect 9582 18136 9588 18148
rect 9088 18108 9588 18136
rect 9088 18096 9094 18108
rect 9582 18096 9588 18108
rect 9640 18096 9646 18148
rect 9953 18139 10011 18145
rect 9953 18105 9965 18139
rect 9999 18136 10011 18139
rect 11790 18136 11796 18148
rect 9999 18108 11796 18136
rect 9999 18105 10011 18108
rect 9953 18099 10011 18105
rect 11790 18096 11796 18108
rect 11848 18096 11854 18148
rect 9048 18068 9076 18096
rect 7852 18040 9076 18068
rect 9398 18028 9404 18080
rect 9456 18068 9462 18080
rect 9493 18071 9551 18077
rect 9493 18068 9505 18071
rect 9456 18040 9505 18068
rect 9456 18028 9462 18040
rect 9493 18037 9505 18040
rect 9539 18037 9551 18071
rect 9493 18031 9551 18037
rect 16117 18071 16175 18077
rect 16117 18037 16129 18071
rect 16163 18068 16175 18071
rect 17586 18068 17592 18080
rect 16163 18040 17592 18068
rect 16163 18037 16175 18040
rect 16117 18031 16175 18037
rect 17586 18028 17592 18040
rect 17644 18028 17650 18080
rect 18322 18028 18328 18080
rect 18380 18068 18386 18080
rect 18984 18077 19012 18244
rect 21269 18241 21281 18275
rect 21315 18241 21327 18275
rect 21269 18235 21327 18241
rect 22094 18232 22100 18284
rect 22152 18232 22158 18284
rect 23658 18232 23664 18284
rect 23716 18272 23722 18284
rect 23937 18275 23995 18281
rect 23937 18272 23949 18275
rect 23716 18244 23949 18272
rect 23716 18232 23722 18244
rect 23937 18241 23949 18244
rect 23983 18241 23995 18275
rect 23937 18235 23995 18241
rect 24670 18164 24676 18216
rect 24728 18164 24734 18216
rect 18601 18071 18659 18077
rect 18601 18068 18613 18071
rect 18380 18040 18613 18068
rect 18380 18028 18386 18040
rect 18601 18037 18613 18040
rect 18647 18037 18659 18071
rect 18601 18031 18659 18037
rect 18969 18071 19027 18077
rect 18969 18037 18981 18071
rect 19015 18068 19027 18071
rect 19150 18068 19156 18080
rect 19015 18040 19156 18068
rect 19015 18037 19027 18040
rect 18969 18031 19027 18037
rect 19150 18028 19156 18040
rect 19208 18028 19214 18080
rect 21085 18071 21143 18077
rect 21085 18037 21097 18071
rect 21131 18068 21143 18071
rect 21542 18068 21548 18080
rect 21131 18040 21548 18068
rect 21131 18037 21143 18040
rect 21085 18031 21143 18037
rect 21542 18028 21548 18040
rect 21600 18028 21606 18080
rect 1104 17978 25852 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 25852 17978
rect 1104 17904 25852 17926
rect 7837 17867 7895 17873
rect 7837 17833 7849 17867
rect 7883 17864 7895 17867
rect 8478 17864 8484 17876
rect 7883 17836 8484 17864
rect 7883 17833 7895 17836
rect 7837 17827 7895 17833
rect 8478 17824 8484 17836
rect 8536 17824 8542 17876
rect 12253 17867 12311 17873
rect 12253 17833 12265 17867
rect 12299 17864 12311 17867
rect 15194 17864 15200 17876
rect 12299 17836 15200 17864
rect 12299 17833 12311 17836
rect 12253 17827 12311 17833
rect 15194 17824 15200 17836
rect 15252 17824 15258 17876
rect 18141 17867 18199 17873
rect 18141 17833 18153 17867
rect 18187 17864 18199 17867
rect 21818 17864 21824 17876
rect 18187 17836 21824 17864
rect 18187 17833 18199 17836
rect 18141 17827 18199 17833
rect 21818 17824 21824 17836
rect 21876 17824 21882 17876
rect 21910 17824 21916 17876
rect 21968 17864 21974 17876
rect 26050 17864 26056 17876
rect 21968 17836 26056 17864
rect 21968 17824 21974 17836
rect 26050 17824 26056 17836
rect 26108 17824 26114 17876
rect 9766 17756 9772 17808
rect 9824 17756 9830 17808
rect 19337 17799 19395 17805
rect 19337 17796 19349 17799
rect 17420 17768 19349 17796
rect 7834 17688 7840 17740
rect 7892 17728 7898 17740
rect 8389 17731 8447 17737
rect 8389 17728 8401 17731
rect 7892 17700 8401 17728
rect 7892 17688 7898 17700
rect 8389 17697 8401 17700
rect 8435 17697 8447 17731
rect 9784 17728 9812 17756
rect 17420 17740 17448 17768
rect 19337 17765 19349 17768
rect 19383 17765 19395 17799
rect 19337 17759 19395 17765
rect 20809 17799 20867 17805
rect 20809 17765 20821 17799
rect 20855 17796 20867 17799
rect 24302 17796 24308 17808
rect 20855 17768 24308 17796
rect 20855 17765 20867 17768
rect 20809 17759 20867 17765
rect 24302 17756 24308 17768
rect 24360 17756 24366 17808
rect 24578 17756 24584 17808
rect 24636 17796 24642 17808
rect 24636 17768 25084 17796
rect 24636 17756 24642 17768
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 9784 17700 10057 17728
rect 8389 17691 8447 17697
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 10045 17691 10103 17697
rect 11698 17688 11704 17740
rect 11756 17728 11762 17740
rect 11793 17731 11851 17737
rect 11793 17728 11805 17731
rect 11756 17700 11805 17728
rect 11756 17688 11762 17700
rect 11793 17697 11805 17700
rect 11839 17697 11851 17731
rect 11793 17691 11851 17697
rect 12897 17731 12955 17737
rect 12897 17697 12909 17731
rect 12943 17728 12955 17731
rect 13354 17728 13360 17740
rect 12943 17700 13360 17728
rect 12943 17697 12955 17700
rect 12897 17691 12955 17697
rect 13354 17688 13360 17700
rect 13412 17688 13418 17740
rect 13906 17688 13912 17740
rect 13964 17728 13970 17740
rect 14642 17728 14648 17740
rect 13964 17700 14648 17728
rect 13964 17688 13970 17700
rect 14642 17688 14648 17700
rect 14700 17728 14706 17740
rect 16206 17728 16212 17740
rect 14700 17700 16212 17728
rect 14700 17688 14706 17700
rect 16206 17688 16212 17700
rect 16264 17688 16270 17740
rect 17402 17688 17408 17740
rect 17460 17688 17466 17740
rect 17494 17688 17500 17740
rect 17552 17688 17558 17740
rect 18322 17688 18328 17740
rect 18380 17728 18386 17740
rect 18693 17731 18751 17737
rect 18693 17728 18705 17731
rect 18380 17700 18705 17728
rect 18380 17688 18386 17700
rect 18693 17697 18705 17700
rect 18739 17697 18751 17731
rect 18693 17691 18751 17697
rect 19794 17688 19800 17740
rect 19852 17728 19858 17740
rect 23845 17731 23903 17737
rect 19852 17700 21036 17728
rect 19852 17688 19858 17700
rect 9582 17620 9588 17672
rect 9640 17660 9646 17672
rect 9769 17663 9827 17669
rect 9769 17660 9781 17663
rect 9640 17632 9781 17660
rect 9640 17620 9646 17632
rect 9769 17629 9781 17632
rect 9815 17629 9827 17663
rect 9769 17623 9827 17629
rect 12621 17663 12679 17669
rect 12621 17629 12633 17663
rect 12667 17660 12679 17663
rect 14274 17660 14280 17672
rect 12667 17632 14280 17660
rect 12667 17629 12679 17632
rect 12621 17623 12679 17629
rect 14274 17620 14280 17632
rect 14332 17620 14338 17672
rect 17310 17620 17316 17672
rect 17368 17660 17374 17672
rect 17368 17632 18828 17660
rect 17368 17620 17374 17632
rect 8205 17595 8263 17601
rect 8205 17561 8217 17595
rect 8251 17592 8263 17595
rect 8846 17592 8852 17604
rect 8251 17564 8852 17592
rect 8251 17561 8263 17564
rect 8205 17555 8263 17561
rect 8846 17552 8852 17564
rect 8904 17552 8910 17604
rect 11422 17592 11428 17604
rect 11270 17564 11428 17592
rect 11422 17552 11428 17564
rect 11480 17552 11486 17604
rect 14090 17592 14096 17604
rect 12728 17564 14096 17592
rect 12728 17536 12756 17564
rect 14090 17552 14096 17564
rect 14148 17552 14154 17604
rect 15562 17552 15568 17604
rect 15620 17592 15626 17604
rect 18509 17595 18567 17601
rect 18509 17592 18521 17595
rect 15620 17564 18521 17592
rect 15620 17552 15626 17564
rect 18509 17561 18521 17564
rect 18555 17561 18567 17595
rect 18509 17555 18567 17561
rect 18601 17595 18659 17601
rect 18601 17561 18613 17595
rect 18647 17592 18659 17595
rect 18690 17592 18696 17604
rect 18647 17564 18696 17592
rect 18647 17561 18659 17564
rect 18601 17555 18659 17561
rect 18690 17552 18696 17564
rect 18748 17552 18754 17604
rect 18800 17592 18828 17632
rect 19334 17620 19340 17672
rect 19392 17660 19398 17672
rect 21008 17669 21036 17700
rect 23845 17697 23857 17731
rect 23891 17728 23903 17731
rect 24946 17728 24952 17740
rect 23891 17700 24952 17728
rect 23891 17697 23903 17700
rect 23845 17691 23903 17697
rect 24946 17688 24952 17700
rect 25004 17688 25010 17740
rect 25056 17737 25084 17768
rect 25041 17731 25099 17737
rect 25041 17697 25053 17731
rect 25087 17697 25099 17731
rect 25041 17691 25099 17697
rect 25130 17688 25136 17740
rect 25188 17688 25194 17740
rect 19981 17663 20039 17669
rect 19981 17660 19993 17663
rect 19392 17632 19993 17660
rect 19392 17620 19398 17632
rect 19981 17629 19993 17632
rect 20027 17629 20039 17663
rect 19981 17623 20039 17629
rect 20993 17663 21051 17669
rect 20993 17629 21005 17663
rect 21039 17629 21051 17663
rect 20993 17623 21051 17629
rect 22005 17663 22063 17669
rect 22005 17629 22017 17663
rect 22051 17660 22063 17663
rect 22833 17663 22891 17669
rect 22051 17632 22784 17660
rect 22051 17629 22063 17632
rect 22005 17623 22063 17629
rect 19429 17595 19487 17601
rect 19429 17592 19441 17595
rect 18800 17564 19441 17592
rect 19429 17561 19441 17564
rect 19475 17561 19487 17595
rect 19429 17555 19487 17561
rect 22186 17552 22192 17604
rect 22244 17552 22250 17604
rect 22756 17592 22784 17632
rect 22833 17629 22845 17663
rect 22879 17660 22891 17663
rect 24578 17660 24584 17672
rect 22879 17632 24584 17660
rect 22879 17629 22891 17632
rect 22833 17623 22891 17629
rect 24578 17620 24584 17632
rect 24636 17620 24642 17672
rect 25866 17592 25872 17604
rect 22756 17564 25872 17592
rect 25866 17552 25872 17564
rect 25924 17552 25930 17604
rect 7190 17484 7196 17536
rect 7248 17484 7254 17536
rect 7742 17484 7748 17536
rect 7800 17524 7806 17536
rect 8297 17527 8355 17533
rect 8297 17524 8309 17527
rect 7800 17496 8309 17524
rect 7800 17484 7806 17496
rect 8297 17493 8309 17496
rect 8343 17493 8355 17527
rect 8297 17487 8355 17493
rect 9125 17527 9183 17533
rect 9125 17493 9137 17527
rect 9171 17524 9183 17527
rect 9398 17524 9404 17536
rect 9171 17496 9404 17524
rect 9171 17493 9183 17496
rect 9125 17487 9183 17493
rect 9398 17484 9404 17496
rect 9456 17484 9462 17536
rect 12710 17484 12716 17536
rect 12768 17484 12774 17536
rect 13170 17484 13176 17536
rect 13228 17524 13234 17536
rect 13449 17527 13507 17533
rect 13449 17524 13461 17527
rect 13228 17496 13461 17524
rect 13228 17484 13234 17496
rect 13449 17493 13461 17496
rect 13495 17493 13507 17527
rect 13449 17487 13507 17493
rect 15746 17484 15752 17536
rect 15804 17484 15810 17536
rect 16206 17484 16212 17536
rect 16264 17524 16270 17536
rect 16393 17527 16451 17533
rect 16393 17524 16405 17527
rect 16264 17496 16405 17524
rect 16264 17484 16270 17496
rect 16393 17493 16405 17496
rect 16439 17493 16451 17527
rect 16393 17487 16451 17493
rect 16945 17527 17003 17533
rect 16945 17493 16957 17527
rect 16991 17524 17003 17527
rect 17218 17524 17224 17536
rect 16991 17496 17224 17524
rect 16991 17493 17003 17496
rect 16945 17487 17003 17493
rect 17218 17484 17224 17496
rect 17276 17484 17282 17536
rect 19797 17527 19855 17533
rect 19797 17493 19809 17527
rect 19843 17524 19855 17527
rect 20898 17524 20904 17536
rect 19843 17496 20904 17524
rect 19843 17493 19855 17496
rect 19797 17487 19855 17493
rect 20898 17484 20904 17496
rect 20956 17484 20962 17536
rect 23566 17484 23572 17536
rect 23624 17524 23630 17536
rect 24581 17527 24639 17533
rect 24581 17524 24593 17527
rect 23624 17496 24593 17524
rect 23624 17484 23630 17496
rect 24581 17493 24593 17496
rect 24627 17493 24639 17527
rect 24581 17487 24639 17493
rect 24670 17484 24676 17536
rect 24728 17524 24734 17536
rect 24949 17527 25007 17533
rect 24949 17524 24961 17527
rect 24728 17496 24961 17524
rect 24728 17484 24734 17496
rect 24949 17493 24961 17496
rect 24995 17493 25007 17527
rect 24949 17487 25007 17493
rect 1104 17434 25852 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 25852 17434
rect 1104 17360 25852 17382
rect 7190 17280 7196 17332
rect 7248 17320 7254 17332
rect 8021 17323 8079 17329
rect 8021 17320 8033 17323
rect 7248 17292 8033 17320
rect 7248 17280 7254 17292
rect 8021 17289 8033 17292
rect 8067 17289 8079 17323
rect 8021 17283 8079 17289
rect 9033 17323 9091 17329
rect 9033 17289 9045 17323
rect 9079 17289 9091 17323
rect 9033 17283 9091 17289
rect 9048 17252 9076 17283
rect 9398 17280 9404 17332
rect 9456 17280 9462 17332
rect 11606 17320 11612 17332
rect 10244 17292 11612 17320
rect 9490 17252 9496 17264
rect 9048 17224 9496 17252
rect 9490 17212 9496 17224
rect 9548 17212 9554 17264
rect 9582 17212 9588 17264
rect 9640 17212 9646 17264
rect 10244 17261 10272 17292
rect 11606 17280 11612 17292
rect 11664 17280 11670 17332
rect 13170 17280 13176 17332
rect 13228 17280 13234 17332
rect 13354 17280 13360 17332
rect 13412 17320 13418 17332
rect 14458 17320 14464 17332
rect 13412 17292 14464 17320
rect 13412 17280 13418 17292
rect 14458 17280 14464 17292
rect 14516 17280 14522 17332
rect 16390 17320 16396 17332
rect 14660 17292 16396 17320
rect 10229 17255 10287 17261
rect 10229 17221 10241 17255
rect 10275 17221 10287 17255
rect 10229 17215 10287 17221
rect 11422 17212 11428 17264
rect 11480 17252 11486 17264
rect 11882 17252 11888 17264
rect 11480 17224 11888 17252
rect 11480 17212 11486 17224
rect 11882 17212 11888 17224
rect 11940 17212 11946 17264
rect 14660 17252 14688 17292
rect 16390 17280 16396 17292
rect 16448 17320 16454 17332
rect 16574 17320 16580 17332
rect 16448 17292 16580 17320
rect 16448 17280 16454 17292
rect 16574 17280 16580 17292
rect 16632 17280 16638 17332
rect 17402 17280 17408 17332
rect 17460 17280 17466 17332
rect 18966 17320 18972 17332
rect 17972 17292 18972 17320
rect 16206 17252 16212 17264
rect 14568 17224 14688 17252
rect 16054 17224 16212 17252
rect 7650 17144 7656 17196
rect 7708 17184 7714 17196
rect 9600 17184 9628 17212
rect 10965 17187 11023 17193
rect 10965 17184 10977 17187
rect 7708 17156 8248 17184
rect 9600 17156 10977 17184
rect 7708 17144 7714 17156
rect 3326 17076 3332 17128
rect 3384 17116 3390 17128
rect 8220 17125 8248 17156
rect 10965 17153 10977 17156
rect 11011 17153 11023 17187
rect 10965 17147 11023 17153
rect 13265 17187 13323 17193
rect 13265 17153 13277 17187
rect 13311 17184 13323 17187
rect 13722 17184 13728 17196
rect 13311 17156 13728 17184
rect 13311 17153 13323 17156
rect 13265 17147 13323 17153
rect 13722 17144 13728 17156
rect 13780 17144 13786 17196
rect 14568 17193 14596 17224
rect 16206 17212 16212 17224
rect 16264 17212 16270 17264
rect 16945 17255 17003 17261
rect 16945 17221 16957 17255
rect 16991 17252 17003 17255
rect 17420 17252 17448 17280
rect 17972 17261 18000 17292
rect 18966 17280 18972 17292
rect 19024 17280 19030 17332
rect 20162 17280 20168 17332
rect 20220 17320 20226 17332
rect 20349 17323 20407 17329
rect 20349 17320 20361 17323
rect 20220 17292 20361 17320
rect 20220 17280 20226 17292
rect 20349 17289 20361 17292
rect 20395 17289 20407 17323
rect 20349 17283 20407 17289
rect 22741 17323 22799 17329
rect 22741 17289 22753 17323
rect 22787 17320 22799 17323
rect 24394 17320 24400 17332
rect 22787 17292 24400 17320
rect 22787 17289 22799 17292
rect 22741 17283 22799 17289
rect 24394 17280 24400 17292
rect 24452 17280 24458 17332
rect 16991 17224 17448 17252
rect 17957 17255 18015 17261
rect 16991 17221 17003 17224
rect 16945 17215 17003 17221
rect 17957 17221 17969 17255
rect 18003 17221 18015 17255
rect 17957 17215 18015 17221
rect 18598 17212 18604 17264
rect 18656 17252 18662 17264
rect 18877 17255 18935 17261
rect 18877 17252 18889 17255
rect 18656 17224 18889 17252
rect 18656 17212 18662 17224
rect 18877 17221 18889 17224
rect 18923 17221 18935 17255
rect 20717 17255 20775 17261
rect 20717 17252 20729 17255
rect 20102 17224 20729 17252
rect 18877 17215 18935 17221
rect 20717 17221 20729 17224
rect 20763 17252 20775 17255
rect 20990 17252 20996 17264
rect 20763 17224 20996 17252
rect 20763 17221 20775 17224
rect 20717 17215 20775 17221
rect 20990 17212 20996 17224
rect 21048 17212 21054 17264
rect 14553 17187 14611 17193
rect 14553 17153 14565 17187
rect 14599 17153 14611 17187
rect 18141 17187 18199 17193
rect 18141 17184 18153 17187
rect 14553 17147 14611 17153
rect 16040 17156 18153 17184
rect 8113 17119 8171 17125
rect 8113 17116 8125 17119
rect 3384 17088 8125 17116
rect 3384 17076 3390 17088
rect 8113 17085 8125 17088
rect 8159 17085 8171 17119
rect 8113 17079 8171 17085
rect 8205 17119 8263 17125
rect 8205 17085 8217 17119
rect 8251 17085 8263 17119
rect 8205 17079 8263 17085
rect 9490 17076 9496 17128
rect 9548 17076 9554 17128
rect 9585 17119 9643 17125
rect 9585 17085 9597 17119
rect 9631 17085 9643 17119
rect 9585 17079 9643 17085
rect 9306 17008 9312 17060
rect 9364 17048 9370 17060
rect 9600 17048 9628 17079
rect 9766 17076 9772 17128
rect 9824 17116 9830 17128
rect 13354 17116 13360 17128
rect 9824 17088 13360 17116
rect 9824 17076 9830 17088
rect 13354 17076 13360 17088
rect 13412 17076 13418 17128
rect 13446 17076 13452 17128
rect 13504 17076 13510 17128
rect 14826 17076 14832 17128
rect 14884 17076 14890 17128
rect 14918 17076 14924 17128
rect 14976 17116 14982 17128
rect 16040 17116 16068 17156
rect 18141 17153 18153 17156
rect 18187 17153 18199 17187
rect 18141 17147 18199 17153
rect 21269 17187 21327 17193
rect 21269 17153 21281 17187
rect 21315 17184 21327 17187
rect 22649 17187 22707 17193
rect 22649 17184 22661 17187
rect 21315 17156 22661 17184
rect 21315 17153 21327 17156
rect 21269 17147 21327 17153
rect 22649 17153 22661 17156
rect 22695 17153 22707 17187
rect 22649 17147 22707 17153
rect 23474 17144 23480 17196
rect 23532 17144 23538 17196
rect 24854 17144 24860 17196
rect 24912 17144 24918 17196
rect 14976 17088 16068 17116
rect 14976 17076 14982 17088
rect 17862 17076 17868 17128
rect 17920 17116 17926 17128
rect 18601 17119 18659 17125
rect 18601 17116 18613 17119
rect 17920 17088 18613 17116
rect 17920 17076 17926 17088
rect 18601 17085 18613 17088
rect 18647 17085 18659 17119
rect 18601 17079 18659 17085
rect 18966 17076 18972 17128
rect 19024 17116 19030 17128
rect 21910 17116 21916 17128
rect 19024 17088 21916 17116
rect 19024 17076 19030 17088
rect 21910 17076 21916 17088
rect 21968 17076 21974 17128
rect 22830 17076 22836 17128
rect 22888 17116 22894 17128
rect 22925 17119 22983 17125
rect 22925 17116 22937 17119
rect 22888 17088 22937 17116
rect 22888 17076 22894 17088
rect 22925 17085 22937 17088
rect 22971 17116 22983 17119
rect 23753 17119 23811 17125
rect 22971 17088 23612 17116
rect 22971 17085 22983 17088
rect 22925 17079 22983 17085
rect 9364 17020 9628 17048
rect 12805 17051 12863 17057
rect 9364 17008 9370 17020
rect 12805 17017 12817 17051
rect 12851 17048 12863 17051
rect 13630 17048 13636 17060
rect 12851 17020 13636 17048
rect 12851 17017 12863 17020
rect 12805 17011 12863 17017
rect 13630 17008 13636 17020
rect 13688 17008 13694 17060
rect 17126 17008 17132 17060
rect 17184 17008 17190 17060
rect 7653 16983 7711 16989
rect 7653 16949 7665 16983
rect 7699 16980 7711 16983
rect 11146 16980 11152 16992
rect 7699 16952 11152 16980
rect 7699 16949 7711 16952
rect 7653 16943 7711 16949
rect 11146 16940 11152 16952
rect 11204 16940 11210 16992
rect 11882 16940 11888 16992
rect 11940 16980 11946 16992
rect 13906 16980 13912 16992
rect 11940 16952 13912 16980
rect 11940 16940 11946 16952
rect 13906 16940 13912 16952
rect 13964 16940 13970 16992
rect 15378 16940 15384 16992
rect 15436 16980 15442 16992
rect 16301 16983 16359 16989
rect 16301 16980 16313 16983
rect 15436 16952 16313 16980
rect 15436 16940 15442 16952
rect 16301 16949 16313 16952
rect 16347 16949 16359 16983
rect 16301 16943 16359 16949
rect 22281 16983 22339 16989
rect 22281 16949 22293 16983
rect 22327 16980 22339 16983
rect 22554 16980 22560 16992
rect 22327 16952 22560 16980
rect 22327 16949 22339 16952
rect 22281 16943 22339 16949
rect 22554 16940 22560 16952
rect 22612 16940 22618 16992
rect 23584 16980 23612 17088
rect 23753 17085 23765 17119
rect 23799 17116 23811 17119
rect 24210 17116 24216 17128
rect 23799 17088 24216 17116
rect 23799 17085 23811 17088
rect 23753 17079 23811 17085
rect 24210 17076 24216 17088
rect 24268 17076 24274 17128
rect 25225 16983 25283 16989
rect 25225 16980 25237 16983
rect 23584 16952 25237 16980
rect 25225 16949 25237 16952
rect 25271 16949 25283 16983
rect 25225 16943 25283 16949
rect 1104 16890 25852 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 25852 16890
rect 1104 16816 25852 16838
rect 12802 16776 12808 16788
rect 11808 16748 12808 16776
rect 10042 16600 10048 16652
rect 10100 16640 10106 16652
rect 10781 16643 10839 16649
rect 10781 16640 10793 16643
rect 10100 16612 10793 16640
rect 10100 16600 10106 16612
rect 10781 16609 10793 16612
rect 10827 16640 10839 16643
rect 10962 16640 10968 16652
rect 10827 16612 10968 16640
rect 10827 16609 10839 16612
rect 10781 16603 10839 16609
rect 10962 16600 10968 16612
rect 11020 16600 11026 16652
rect 11422 16640 11428 16652
rect 11072 16612 11428 16640
rect 10410 16532 10416 16584
rect 10468 16572 10474 16584
rect 11072 16572 11100 16612
rect 11422 16600 11428 16612
rect 11480 16600 11486 16652
rect 11808 16649 11836 16748
rect 12802 16736 12808 16748
rect 12860 16736 12866 16788
rect 13906 16736 13912 16788
rect 13964 16736 13970 16788
rect 14274 16736 14280 16788
rect 14332 16776 14338 16788
rect 18966 16776 18972 16788
rect 14332 16748 18972 16776
rect 14332 16736 14338 16748
rect 18966 16736 18972 16748
rect 19024 16736 19030 16788
rect 20990 16736 20996 16788
rect 21048 16776 21054 16788
rect 22278 16776 22284 16788
rect 21048 16748 22284 16776
rect 21048 16736 21054 16748
rect 22278 16736 22284 16748
rect 22336 16736 22342 16788
rect 24578 16736 24584 16788
rect 24636 16736 24642 16788
rect 14366 16708 14372 16720
rect 13556 16680 14372 16708
rect 11793 16643 11851 16649
rect 11793 16609 11805 16643
rect 11839 16609 11851 16643
rect 11793 16603 11851 16609
rect 12069 16643 12127 16649
rect 12069 16609 12081 16643
rect 12115 16640 12127 16643
rect 13556 16640 13584 16680
rect 14366 16668 14372 16680
rect 14424 16668 14430 16720
rect 12115 16612 13584 16640
rect 12115 16609 12127 16612
rect 12069 16603 12127 16609
rect 13630 16600 13636 16652
rect 13688 16640 13694 16652
rect 15105 16643 15163 16649
rect 15105 16640 15117 16643
rect 13688 16612 15117 16640
rect 13688 16600 13694 16612
rect 15105 16609 15117 16612
rect 15151 16609 15163 16643
rect 15105 16603 15163 16609
rect 15838 16600 15844 16652
rect 15896 16640 15902 16652
rect 16209 16643 16267 16649
rect 16209 16640 16221 16643
rect 15896 16612 16221 16640
rect 15896 16600 15902 16612
rect 16209 16609 16221 16612
rect 16255 16609 16267 16643
rect 16209 16603 16267 16609
rect 16298 16600 16304 16652
rect 16356 16600 16362 16652
rect 16390 16600 16396 16652
rect 16448 16640 16454 16652
rect 17862 16640 17868 16652
rect 16448 16612 17868 16640
rect 16448 16600 16454 16612
rect 17862 16600 17868 16612
rect 17920 16640 17926 16652
rect 17957 16643 18015 16649
rect 17957 16640 17969 16643
rect 17920 16612 17969 16640
rect 17920 16600 17926 16612
rect 17957 16609 17969 16612
rect 18003 16609 18015 16643
rect 19334 16640 19340 16652
rect 17957 16603 18015 16609
rect 18064 16612 19340 16640
rect 10468 16544 11100 16572
rect 14568 16544 15700 16572
rect 10468 16532 10474 16544
rect 10318 16504 10324 16516
rect 9876 16476 10324 16504
rect 9876 16448 9904 16476
rect 10318 16464 10324 16476
rect 10376 16504 10382 16516
rect 10597 16507 10655 16513
rect 10597 16504 10609 16507
rect 10376 16476 10609 16504
rect 10376 16464 10382 16476
rect 10597 16473 10609 16476
rect 10643 16473 10655 16507
rect 13906 16504 13912 16516
rect 13294 16476 13912 16504
rect 10597 16467 10655 16473
rect 13906 16464 13912 16476
rect 13964 16464 13970 16516
rect 9858 16396 9864 16448
rect 9916 16396 9922 16448
rect 10226 16396 10232 16448
rect 10284 16396 10290 16448
rect 10689 16439 10747 16445
rect 10689 16405 10701 16439
rect 10735 16436 10747 16439
rect 12250 16436 12256 16448
rect 10735 16408 12256 16436
rect 10735 16405 10747 16408
rect 10689 16399 10747 16405
rect 12250 16396 12256 16408
rect 12308 16396 12314 16448
rect 13541 16439 13599 16445
rect 13541 16405 13553 16439
rect 13587 16436 13599 16439
rect 13630 16436 13636 16448
rect 13587 16408 13636 16436
rect 13587 16405 13599 16408
rect 13541 16399 13599 16405
rect 13630 16396 13636 16408
rect 13688 16396 13694 16448
rect 14568 16445 14596 16544
rect 14921 16507 14979 16513
rect 14921 16473 14933 16507
rect 14967 16504 14979 16507
rect 15470 16504 15476 16516
rect 14967 16476 15476 16504
rect 14967 16473 14979 16476
rect 14921 16467 14979 16473
rect 15470 16464 15476 16476
rect 15528 16464 15534 16516
rect 15672 16504 15700 16544
rect 15746 16532 15752 16584
rect 15804 16572 15810 16584
rect 16117 16575 16175 16581
rect 16117 16572 16129 16575
rect 15804 16544 16129 16572
rect 15804 16532 15810 16544
rect 16117 16541 16129 16544
rect 16163 16541 16175 16575
rect 16117 16535 16175 16541
rect 16942 16532 16948 16584
rect 17000 16572 17006 16584
rect 17221 16575 17279 16581
rect 17221 16572 17233 16575
rect 17000 16544 17233 16572
rect 17000 16532 17006 16544
rect 17221 16541 17233 16544
rect 17267 16572 17279 16575
rect 18064 16572 18092 16612
rect 19334 16600 19340 16612
rect 19392 16600 19398 16652
rect 20254 16600 20260 16652
rect 20312 16600 20318 16652
rect 18877 16575 18935 16581
rect 18877 16572 18889 16575
rect 17267 16544 18092 16572
rect 18156 16544 18889 16572
rect 17267 16541 17279 16544
rect 17221 16535 17279 16541
rect 18156 16504 18184 16544
rect 18877 16541 18889 16544
rect 18923 16541 18935 16575
rect 18877 16535 18935 16541
rect 19794 16532 19800 16584
rect 19852 16532 19858 16584
rect 22370 16532 22376 16584
rect 22428 16572 22434 16584
rect 22649 16575 22707 16581
rect 22649 16572 22661 16575
rect 22428 16544 22661 16572
rect 22428 16532 22434 16544
rect 22649 16541 22661 16544
rect 22695 16541 22707 16575
rect 22649 16535 22707 16541
rect 23842 16532 23848 16584
rect 23900 16532 23906 16584
rect 24765 16575 24823 16581
rect 24765 16541 24777 16575
rect 24811 16541 24823 16575
rect 24765 16535 24823 16541
rect 15672 16476 18184 16504
rect 18708 16476 20484 16504
rect 14553 16439 14611 16445
rect 14553 16405 14565 16439
rect 14599 16405 14611 16439
rect 14553 16399 14611 16405
rect 15010 16396 15016 16448
rect 15068 16396 15074 16448
rect 15749 16439 15807 16445
rect 15749 16405 15761 16439
rect 15795 16436 15807 16439
rect 15930 16436 15936 16448
rect 15795 16408 15936 16436
rect 15795 16405 15807 16408
rect 15749 16399 15807 16405
rect 15930 16396 15936 16408
rect 15988 16396 15994 16448
rect 18708 16445 18736 16476
rect 18693 16439 18751 16445
rect 18693 16405 18705 16439
rect 18739 16405 18751 16439
rect 18693 16399 18751 16405
rect 19610 16396 19616 16448
rect 19668 16396 19674 16448
rect 20456 16436 20484 16476
rect 20530 16464 20536 16516
rect 20588 16464 20594 16516
rect 20990 16464 20996 16516
rect 21048 16464 21054 16516
rect 24780 16504 24808 16535
rect 21823 16476 24808 16504
rect 21823 16436 21851 16476
rect 20456 16408 21851 16436
rect 21910 16396 21916 16448
rect 21968 16436 21974 16448
rect 22005 16439 22063 16445
rect 22005 16436 22017 16439
rect 21968 16408 22017 16436
rect 21968 16396 21974 16408
rect 22005 16405 22017 16408
rect 22051 16405 22063 16439
rect 22005 16399 22063 16405
rect 22278 16396 22284 16448
rect 22336 16436 22342 16448
rect 22373 16439 22431 16445
rect 22373 16436 22385 16439
rect 22336 16408 22385 16436
rect 22336 16396 22342 16408
rect 22373 16405 22385 16408
rect 22419 16436 22431 16439
rect 23658 16436 23664 16448
rect 22419 16408 23664 16436
rect 22419 16405 22431 16408
rect 22373 16399 22431 16405
rect 23658 16396 23664 16408
rect 23716 16396 23722 16448
rect 24854 16396 24860 16448
rect 24912 16436 24918 16448
rect 25130 16436 25136 16448
rect 24912 16408 25136 16436
rect 24912 16396 24918 16408
rect 25130 16396 25136 16408
rect 25188 16436 25194 16448
rect 25409 16439 25467 16445
rect 25409 16436 25421 16439
rect 25188 16408 25421 16436
rect 25188 16396 25194 16408
rect 25409 16405 25421 16408
rect 25455 16405 25467 16439
rect 25409 16399 25467 16405
rect 1104 16346 25852 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 25852 16346
rect 1104 16272 25852 16294
rect 8297 16235 8355 16241
rect 8297 16201 8309 16235
rect 8343 16232 8355 16235
rect 8570 16232 8576 16244
rect 8343 16204 8576 16232
rect 8343 16201 8355 16204
rect 8297 16195 8355 16201
rect 8570 16192 8576 16204
rect 8628 16192 8634 16244
rect 8662 16192 8668 16244
rect 8720 16192 8726 16244
rect 11054 16192 11060 16244
rect 11112 16232 11118 16244
rect 12161 16235 12219 16241
rect 12161 16232 12173 16235
rect 11112 16204 12173 16232
rect 11112 16192 11118 16204
rect 12161 16201 12173 16204
rect 12207 16201 12219 16235
rect 12161 16195 12219 16201
rect 12529 16235 12587 16241
rect 12529 16201 12541 16235
rect 12575 16232 12587 16235
rect 14182 16232 14188 16244
rect 12575 16204 14188 16232
rect 12575 16201 12587 16204
rect 12529 16195 12587 16201
rect 14182 16192 14188 16204
rect 14240 16192 14246 16244
rect 14553 16235 14611 16241
rect 14553 16201 14565 16235
rect 14599 16232 14611 16235
rect 15010 16232 15016 16244
rect 14599 16204 15016 16232
rect 14599 16201 14611 16204
rect 14553 16195 14611 16201
rect 15010 16192 15016 16204
rect 15068 16192 15074 16244
rect 15470 16192 15476 16244
rect 15528 16232 15534 16244
rect 15749 16235 15807 16241
rect 15749 16232 15761 16235
rect 15528 16204 15761 16232
rect 15528 16192 15534 16204
rect 15749 16201 15761 16204
rect 15795 16201 15807 16235
rect 15749 16195 15807 16201
rect 16850 16192 16856 16244
rect 16908 16232 16914 16244
rect 20254 16232 20260 16244
rect 16908 16204 17264 16232
rect 16908 16192 16914 16204
rect 8680 16164 8708 16192
rect 8050 16136 8708 16164
rect 13725 16167 13783 16173
rect 13725 16133 13737 16167
rect 13771 16164 13783 16167
rect 14274 16164 14280 16176
rect 13771 16136 14280 16164
rect 13771 16133 13783 16136
rect 13725 16127 13783 16133
rect 14274 16124 14280 16136
rect 14332 16124 14338 16176
rect 17236 16173 17264 16204
rect 20088 16204 20260 16232
rect 20088 16173 20116 16204
rect 20254 16192 20260 16204
rect 20312 16232 20318 16244
rect 22278 16232 22284 16244
rect 20312 16204 22284 16232
rect 20312 16192 20318 16204
rect 17221 16167 17279 16173
rect 17221 16133 17233 16167
rect 17267 16133 17279 16167
rect 20073 16167 20131 16173
rect 17221 16127 17279 16133
rect 18708 16136 20024 16164
rect 6546 16056 6552 16108
rect 6604 16056 6610 16108
rect 11698 16056 11704 16108
rect 11756 16096 11762 16108
rect 12158 16096 12164 16108
rect 11756 16068 12164 16096
rect 11756 16056 11762 16068
rect 12158 16056 12164 16068
rect 12216 16096 12222 16108
rect 12621 16099 12679 16105
rect 12216 16068 12434 16096
rect 12216 16056 12222 16068
rect 6825 16031 6883 16037
rect 6825 15997 6837 16031
rect 6871 16028 6883 16031
rect 8478 16028 8484 16040
rect 6871 16000 8484 16028
rect 6871 15997 6883 16000
rect 6825 15991 6883 15997
rect 8478 15988 8484 16000
rect 8536 16028 8542 16040
rect 9582 16028 9588 16040
rect 8536 16000 9588 16028
rect 8536 15988 8542 16000
rect 9582 15988 9588 16000
rect 9640 15988 9646 16040
rect 12406 16028 12434 16068
rect 12621 16065 12633 16099
rect 12667 16096 12679 16099
rect 12667 16068 14320 16096
rect 12667 16065 12679 16068
rect 12621 16059 12679 16065
rect 14292 16040 14320 16068
rect 14734 16056 14740 16108
rect 14792 16096 14798 16108
rect 14921 16099 14979 16105
rect 14921 16096 14933 16099
rect 14792 16068 14933 16096
rect 14792 16056 14798 16068
rect 14921 16065 14933 16068
rect 14967 16065 14979 16099
rect 14921 16059 14979 16065
rect 15013 16099 15071 16105
rect 15013 16065 15025 16099
rect 15059 16096 15071 16099
rect 18049 16099 18107 16105
rect 15059 16068 16344 16096
rect 15059 16065 15071 16068
rect 15013 16059 15071 16065
rect 12713 16031 12771 16037
rect 12713 16028 12725 16031
rect 12406 16000 12725 16028
rect 12713 15997 12725 16000
rect 12759 15997 12771 16031
rect 12713 15991 12771 15997
rect 13814 15988 13820 16040
rect 13872 15988 13878 16040
rect 13909 16031 13967 16037
rect 13909 15997 13921 16031
rect 13955 15997 13967 16031
rect 13909 15991 13967 15997
rect 11698 15920 11704 15972
rect 11756 15960 11762 15972
rect 13924 15960 13952 15991
rect 14274 15988 14280 16040
rect 14332 15988 14338 16040
rect 15105 16031 15163 16037
rect 15105 15997 15117 16031
rect 15151 15997 15163 16031
rect 15105 15991 15163 15997
rect 11756 15932 13952 15960
rect 11756 15920 11762 15932
rect 14366 15920 14372 15972
rect 14424 15960 14430 15972
rect 15120 15960 15148 15991
rect 16316 15969 16344 16068
rect 18049 16065 18061 16099
rect 18095 16096 18107 16099
rect 18414 16096 18420 16108
rect 18095 16068 18420 16096
rect 18095 16065 18107 16068
rect 18049 16059 18107 16065
rect 18414 16056 18420 16068
rect 18472 16056 18478 16108
rect 18708 16105 18736 16136
rect 18693 16099 18751 16105
rect 18693 16065 18705 16099
rect 18739 16065 18751 16099
rect 18693 16059 18751 16065
rect 19245 16099 19303 16105
rect 19245 16065 19257 16099
rect 19291 16096 19303 16099
rect 19334 16096 19340 16108
rect 19291 16068 19340 16096
rect 19291 16065 19303 16068
rect 19245 16059 19303 16065
rect 19334 16056 19340 16068
rect 19392 16056 19398 16108
rect 19996 16096 20024 16136
rect 20073 16133 20085 16167
rect 20119 16133 20131 16167
rect 20073 16127 20131 16133
rect 20346 16124 20352 16176
rect 20404 16164 20410 16176
rect 20622 16164 20628 16176
rect 20404 16136 20628 16164
rect 20404 16124 20410 16136
rect 20622 16124 20628 16136
rect 20680 16164 20686 16176
rect 21910 16164 21916 16176
rect 20680 16136 21916 16164
rect 20680 16124 20686 16136
rect 21910 16124 21916 16136
rect 21968 16124 21974 16176
rect 20438 16096 20444 16108
rect 19996 16068 20444 16096
rect 20438 16056 20444 16068
rect 20496 16056 20502 16108
rect 20806 16056 20812 16108
rect 20864 16096 20870 16108
rect 22020 16105 22048 16204
rect 22278 16192 22284 16204
rect 22336 16232 22342 16244
rect 23290 16232 23296 16244
rect 22336 16204 23296 16232
rect 22336 16192 22342 16204
rect 23290 16192 23296 16204
rect 23348 16192 23354 16244
rect 24121 16235 24179 16241
rect 24121 16232 24133 16235
rect 23768 16204 24133 16232
rect 23658 16164 23664 16176
rect 23506 16136 23664 16164
rect 23658 16124 23664 16136
rect 23716 16164 23722 16176
rect 23768 16164 23796 16204
rect 24121 16201 24133 16204
rect 24167 16232 24179 16235
rect 24854 16232 24860 16244
rect 24167 16204 24860 16232
rect 24167 16201 24179 16204
rect 24121 16195 24179 16201
rect 24854 16192 24860 16204
rect 24912 16192 24918 16244
rect 23716 16136 23796 16164
rect 23716 16124 23722 16136
rect 21085 16099 21143 16105
rect 21085 16096 21097 16099
rect 20864 16068 21097 16096
rect 20864 16056 20870 16068
rect 21085 16065 21097 16068
rect 21131 16065 21143 16099
rect 21085 16059 21143 16065
rect 22005 16099 22063 16105
rect 22005 16065 22017 16099
rect 22051 16065 22063 16099
rect 22005 16059 22063 16065
rect 23290 16056 23296 16108
rect 23348 16056 23354 16108
rect 23842 16056 23848 16108
rect 23900 16096 23906 16108
rect 24765 16099 24823 16105
rect 24765 16096 24777 16099
rect 23900 16068 24777 16096
rect 23900 16056 23906 16068
rect 24765 16065 24777 16068
rect 24811 16065 24823 16099
rect 24765 16059 24823 16065
rect 19886 15988 19892 16040
rect 19944 16028 19950 16040
rect 21177 16031 21235 16037
rect 21177 16028 21189 16031
rect 19944 16000 21189 16028
rect 19944 15988 19950 16000
rect 21177 15997 21189 16000
rect 21223 15997 21235 16031
rect 21177 15991 21235 15997
rect 21361 16031 21419 16037
rect 21361 15997 21373 16031
rect 21407 16028 21419 16031
rect 22281 16031 22339 16037
rect 21407 16000 22140 16028
rect 21407 15997 21419 16000
rect 21361 15991 21419 15997
rect 14424 15932 15148 15960
rect 16301 15963 16359 15969
rect 14424 15920 14430 15932
rect 16301 15929 16313 15963
rect 16347 15960 16359 15963
rect 17678 15960 17684 15972
rect 16347 15932 17684 15960
rect 16347 15929 16359 15932
rect 16301 15923 16359 15929
rect 17678 15920 17684 15932
rect 17736 15960 17742 15972
rect 18230 15960 18236 15972
rect 17736 15932 18236 15960
rect 17736 15920 17742 15932
rect 18230 15920 18236 15932
rect 18288 15920 18294 15972
rect 19794 15920 19800 15972
rect 19852 15960 19858 15972
rect 22002 15960 22008 15972
rect 19852 15932 22008 15960
rect 19852 15920 19858 15932
rect 22002 15920 22008 15932
rect 22060 15920 22066 15972
rect 12250 15852 12256 15904
rect 12308 15892 12314 15904
rect 13357 15895 13415 15901
rect 13357 15892 13369 15895
rect 12308 15864 13369 15892
rect 12308 15852 12314 15864
rect 13357 15861 13369 15864
rect 13403 15861 13415 15895
rect 13357 15855 13415 15861
rect 17310 15852 17316 15904
rect 17368 15852 17374 15904
rect 17770 15852 17776 15904
rect 17828 15892 17834 15904
rect 17865 15895 17923 15901
rect 17865 15892 17877 15895
rect 17828 15864 17877 15892
rect 17828 15852 17834 15864
rect 17865 15861 17877 15864
rect 17911 15861 17923 15895
rect 17865 15855 17923 15861
rect 18506 15852 18512 15904
rect 18564 15852 18570 15904
rect 20717 15895 20775 15901
rect 20717 15861 20729 15895
rect 20763 15892 20775 15895
rect 21450 15892 21456 15904
rect 20763 15864 21456 15892
rect 20763 15861 20775 15864
rect 20717 15855 20775 15861
rect 21450 15852 21456 15864
rect 21508 15852 21514 15904
rect 22112 15892 22140 16000
rect 22281 15997 22293 16031
rect 22327 16028 22339 16031
rect 22738 16028 22744 16040
rect 22327 16000 22744 16028
rect 22327 15997 22339 16000
rect 22281 15991 22339 15997
rect 22738 15988 22744 16000
rect 22796 15988 22802 16040
rect 22830 15988 22836 16040
rect 22888 16028 22894 16040
rect 23308 16028 23336 16056
rect 22888 16000 23336 16028
rect 24489 16031 24547 16037
rect 22888 15988 22894 16000
rect 24489 15997 24501 16031
rect 24535 16028 24547 16031
rect 24578 16028 24584 16040
rect 24535 16000 24584 16028
rect 24535 15997 24547 16000
rect 24489 15991 24547 15997
rect 24578 15988 24584 16000
rect 24636 15988 24642 16040
rect 23750 15892 23756 15904
rect 22112 15864 23756 15892
rect 23750 15852 23756 15864
rect 23808 15852 23814 15904
rect 1104 15802 25852 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 25852 15802
rect 1104 15728 25852 15750
rect 9125 15691 9183 15697
rect 9125 15657 9137 15691
rect 9171 15688 9183 15691
rect 9214 15688 9220 15700
rect 9171 15660 9220 15688
rect 9171 15657 9183 15660
rect 9125 15651 9183 15657
rect 9214 15648 9220 15660
rect 9272 15648 9278 15700
rect 10229 15691 10287 15697
rect 10229 15657 10241 15691
rect 10275 15688 10287 15691
rect 10410 15688 10416 15700
rect 10275 15660 10416 15688
rect 10275 15657 10287 15660
rect 10229 15651 10287 15657
rect 10410 15648 10416 15660
rect 10468 15648 10474 15700
rect 11514 15648 11520 15700
rect 11572 15688 11578 15700
rect 11609 15691 11667 15697
rect 11609 15688 11621 15691
rect 11572 15660 11621 15688
rect 11572 15648 11578 15660
rect 11609 15657 11621 15660
rect 11655 15657 11667 15691
rect 11609 15651 11667 15657
rect 17678 15648 17684 15700
rect 17736 15688 17742 15700
rect 17862 15688 17868 15700
rect 17736 15660 17868 15688
rect 17736 15648 17742 15660
rect 17862 15648 17868 15660
rect 17920 15688 17926 15700
rect 18141 15691 18199 15697
rect 18141 15688 18153 15691
rect 17920 15660 18153 15688
rect 17920 15648 17926 15660
rect 18141 15657 18153 15660
rect 18187 15657 18199 15691
rect 18141 15651 18199 15657
rect 18509 15691 18567 15697
rect 18509 15657 18521 15691
rect 18555 15688 18567 15691
rect 19150 15688 19156 15700
rect 18555 15660 19156 15688
rect 18555 15657 18567 15660
rect 18509 15651 18567 15657
rect 9582 15512 9588 15564
rect 9640 15552 9646 15564
rect 9677 15555 9735 15561
rect 9677 15552 9689 15555
rect 9640 15524 9689 15552
rect 9640 15512 9646 15524
rect 9677 15521 9689 15524
rect 9723 15521 9735 15555
rect 9677 15515 9735 15521
rect 12158 15512 12164 15564
rect 12216 15512 12222 15564
rect 16390 15512 16396 15564
rect 16448 15512 16454 15564
rect 16669 15555 16727 15561
rect 16669 15521 16681 15555
rect 16715 15552 16727 15555
rect 18322 15552 18328 15564
rect 16715 15524 18328 15552
rect 16715 15521 16727 15524
rect 16669 15515 16727 15521
rect 18322 15512 18328 15524
rect 18380 15512 18386 15564
rect 18524 15484 18552 15651
rect 19150 15648 19156 15660
rect 19208 15688 19214 15700
rect 19208 15660 20760 15688
rect 19208 15648 19214 15660
rect 20732 15620 20760 15660
rect 21450 15648 21456 15700
rect 21508 15688 21514 15700
rect 22738 15688 22744 15700
rect 21508 15660 22744 15688
rect 21508 15648 21514 15660
rect 22738 15648 22744 15660
rect 22796 15648 22802 15700
rect 22922 15648 22928 15700
rect 22980 15688 22986 15700
rect 24029 15691 24087 15697
rect 24029 15688 24041 15691
rect 22980 15660 24041 15688
rect 22980 15648 22986 15660
rect 24029 15657 24041 15660
rect 24075 15657 24087 15691
rect 24029 15651 24087 15657
rect 25130 15648 25136 15700
rect 25188 15648 25194 15700
rect 20732 15592 20944 15620
rect 19429 15555 19487 15561
rect 19429 15521 19441 15555
rect 19475 15552 19487 15555
rect 20254 15552 20260 15564
rect 19475 15524 20260 15552
rect 19475 15521 19487 15524
rect 19429 15515 19487 15521
rect 20254 15512 20260 15524
rect 20312 15512 20318 15564
rect 17802 15470 18552 15484
rect 17788 15456 18552 15470
rect 9214 15376 9220 15428
rect 9272 15416 9278 15428
rect 9585 15419 9643 15425
rect 9585 15416 9597 15419
rect 9272 15388 9597 15416
rect 9272 15376 9278 15388
rect 9585 15385 9597 15388
rect 9631 15385 9643 15419
rect 9585 15379 9643 15385
rect 11977 15419 12035 15425
rect 11977 15385 11989 15419
rect 12023 15416 12035 15419
rect 12526 15416 12532 15428
rect 12023 15388 12532 15416
rect 12023 15385 12035 15388
rect 11977 15379 12035 15385
rect 12526 15376 12532 15388
rect 12584 15376 12590 15428
rect 9493 15351 9551 15357
rect 9493 15317 9505 15351
rect 9539 15348 9551 15351
rect 10042 15348 10048 15360
rect 9539 15320 10048 15348
rect 9539 15317 9551 15320
rect 9493 15311 9551 15317
rect 10042 15308 10048 15320
rect 10100 15308 10106 15360
rect 12066 15308 12072 15360
rect 12124 15308 12130 15360
rect 14274 15308 14280 15360
rect 14332 15308 14338 15360
rect 15746 15308 15752 15360
rect 15804 15308 15810 15360
rect 16390 15308 16396 15360
rect 16448 15348 16454 15360
rect 17788 15348 17816 15456
rect 19702 15376 19708 15428
rect 19760 15376 19766 15428
rect 20916 15416 20944 15592
rect 22278 15512 22284 15564
rect 22336 15512 22342 15564
rect 22557 15555 22615 15561
rect 22557 15521 22569 15555
rect 22603 15552 22615 15555
rect 23750 15552 23756 15564
rect 22603 15524 23756 15552
rect 22603 15521 22615 15524
rect 22557 15515 22615 15521
rect 23750 15512 23756 15524
rect 23808 15512 23814 15564
rect 24581 15555 24639 15561
rect 24581 15521 24593 15555
rect 24627 15552 24639 15555
rect 24670 15552 24676 15564
rect 24627 15524 24676 15552
rect 24627 15521 24639 15524
rect 24581 15515 24639 15521
rect 24670 15512 24676 15524
rect 24728 15512 24734 15564
rect 21818 15444 21824 15496
rect 21876 15444 21882 15496
rect 23658 15444 23664 15496
rect 23716 15444 23722 15496
rect 21082 15416 21088 15428
rect 20916 15402 21088 15416
rect 20930 15388 21088 15402
rect 21082 15376 21088 15388
rect 21140 15376 21146 15428
rect 25222 15416 25228 15428
rect 23952 15388 25228 15416
rect 16448 15320 17816 15348
rect 16448 15308 16454 15320
rect 20530 15308 20536 15360
rect 20588 15348 20594 15360
rect 21177 15351 21235 15357
rect 21177 15348 21189 15351
rect 20588 15320 21189 15348
rect 20588 15308 20594 15320
rect 21177 15317 21189 15320
rect 21223 15317 21235 15351
rect 21177 15311 21235 15317
rect 21637 15351 21695 15357
rect 21637 15317 21649 15351
rect 21683 15348 21695 15351
rect 23952 15348 23980 15388
rect 25222 15376 25228 15388
rect 25280 15376 25286 15428
rect 21683 15320 23980 15348
rect 21683 15317 21695 15320
rect 21637 15311 21695 15317
rect 1104 15258 25852 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 25852 15258
rect 1104 15184 25852 15206
rect 10134 15104 10140 15156
rect 10192 15104 10198 15156
rect 10410 15104 10416 15156
rect 10468 15144 10474 15156
rect 10870 15144 10876 15156
rect 10468 15116 10876 15144
rect 10468 15104 10474 15116
rect 10870 15104 10876 15116
rect 10928 15144 10934 15156
rect 12069 15147 12127 15153
rect 12069 15144 12081 15147
rect 10928 15116 12081 15144
rect 10928 15104 10934 15116
rect 12069 15113 12081 15116
rect 12115 15113 12127 15147
rect 12069 15107 12127 15113
rect 14093 15147 14151 15153
rect 14093 15113 14105 15147
rect 14139 15144 14151 15147
rect 14274 15144 14280 15156
rect 14139 15116 14280 15144
rect 14139 15113 14151 15116
rect 14093 15107 14151 15113
rect 14274 15104 14280 15116
rect 14332 15104 14338 15156
rect 15562 15104 15568 15156
rect 15620 15104 15626 15156
rect 15746 15104 15752 15156
rect 15804 15144 15810 15156
rect 15933 15147 15991 15153
rect 15933 15144 15945 15147
rect 15804 15116 15945 15144
rect 15804 15104 15810 15116
rect 15933 15113 15945 15116
rect 15979 15113 15991 15147
rect 15933 15107 15991 15113
rect 20070 15104 20076 15156
rect 20128 15104 20134 15156
rect 20162 15104 20168 15156
rect 20220 15144 20226 15156
rect 25682 15144 25688 15156
rect 20220 15116 25688 15144
rect 20220 15104 20226 15116
rect 25682 15104 25688 15116
rect 25740 15104 25746 15156
rect 8662 15036 8668 15088
rect 8720 15036 8726 15088
rect 10597 15079 10655 15085
rect 10597 15045 10609 15079
rect 10643 15076 10655 15079
rect 11514 15076 11520 15088
rect 10643 15048 11520 15076
rect 10643 15045 10655 15048
rect 10597 15039 10655 15045
rect 11514 15036 11520 15048
rect 11572 15036 11578 15088
rect 18693 15079 18751 15085
rect 18693 15045 18705 15079
rect 18739 15076 18751 15079
rect 19242 15076 19248 15088
rect 18739 15048 19248 15076
rect 18739 15045 18751 15048
rect 18693 15039 18751 15045
rect 19242 15036 19248 15048
rect 19300 15036 19306 15088
rect 21082 15036 21088 15088
rect 21140 15076 21146 15088
rect 21269 15079 21327 15085
rect 21269 15076 21281 15079
rect 21140 15048 21281 15076
rect 21140 15036 21146 15048
rect 21269 15045 21281 15048
rect 21315 15045 21327 15079
rect 21269 15039 21327 15045
rect 23290 15036 23296 15088
rect 23348 15036 23354 15088
rect 9582 14968 9588 15020
rect 9640 15008 9646 15020
rect 10505 15011 10563 15017
rect 9640 14980 9812 15008
rect 9640 14968 9646 14980
rect 7653 14943 7711 14949
rect 7653 14909 7665 14943
rect 7699 14940 7711 14943
rect 7929 14943 7987 14949
rect 7699 14912 7788 14940
rect 7699 14909 7711 14912
rect 7653 14903 7711 14909
rect 7760 14804 7788 14912
rect 7929 14909 7941 14943
rect 7975 14940 7987 14943
rect 8570 14940 8576 14952
rect 7975 14912 8576 14940
rect 7975 14909 7987 14912
rect 7929 14903 7987 14909
rect 8570 14900 8576 14912
rect 8628 14900 8634 14952
rect 9306 14900 9312 14952
rect 9364 14940 9370 14952
rect 9677 14943 9735 14949
rect 9677 14940 9689 14943
rect 9364 14912 9689 14940
rect 9364 14900 9370 14912
rect 9677 14909 9689 14912
rect 9723 14909 9735 14943
rect 9784 14940 9812 14980
rect 10505 14977 10517 15011
rect 10551 15008 10563 15011
rect 11422 15008 11428 15020
rect 10551 14980 11428 15008
rect 10551 14977 10563 14980
rect 10505 14971 10563 14977
rect 11422 14968 11428 14980
rect 11480 14968 11486 15020
rect 19426 14968 19432 15020
rect 19484 15008 19490 15020
rect 19981 15011 20039 15017
rect 19981 15008 19993 15011
rect 19484 14980 19993 15008
rect 19484 14968 19490 14980
rect 19981 14977 19993 14980
rect 20027 14977 20039 15011
rect 19981 14971 20039 14977
rect 20993 15011 21051 15017
rect 20993 14977 21005 15011
rect 21039 14977 21051 15011
rect 20993 14971 21051 14977
rect 10689 14943 10747 14949
rect 10689 14940 10701 14943
rect 9784 14912 10701 14940
rect 9677 14903 9735 14909
rect 10689 14909 10701 14912
rect 10735 14909 10747 14943
rect 10689 14903 10747 14909
rect 11882 14900 11888 14952
rect 11940 14940 11946 14952
rect 14185 14943 14243 14949
rect 14185 14940 14197 14943
rect 11940 14912 14197 14940
rect 11940 14900 11946 14912
rect 14185 14909 14197 14912
rect 14231 14909 14243 14943
rect 14185 14903 14243 14909
rect 14369 14943 14427 14949
rect 14369 14909 14381 14943
rect 14415 14940 14427 14943
rect 15378 14940 15384 14952
rect 14415 14912 15384 14940
rect 14415 14909 14427 14912
rect 14369 14903 14427 14909
rect 15378 14900 15384 14912
rect 15436 14900 15442 14952
rect 15470 14900 15476 14952
rect 15528 14940 15534 14952
rect 16025 14943 16083 14949
rect 16025 14940 16037 14943
rect 15528 14912 16037 14940
rect 15528 14900 15534 14912
rect 16025 14909 16037 14912
rect 16071 14909 16083 14943
rect 16025 14903 16083 14909
rect 16209 14943 16267 14949
rect 16209 14909 16221 14943
rect 16255 14940 16267 14943
rect 17034 14940 17040 14952
rect 16255 14912 17040 14940
rect 16255 14909 16267 14912
rect 16209 14903 16267 14909
rect 17034 14900 17040 14912
rect 17092 14900 17098 14952
rect 20257 14943 20315 14949
rect 20257 14909 20269 14943
rect 20303 14940 20315 14943
rect 20530 14940 20536 14952
rect 20303 14912 20536 14940
rect 20303 14909 20315 14912
rect 20257 14903 20315 14909
rect 20530 14900 20536 14912
rect 20588 14900 20594 14952
rect 21008 14940 21036 14971
rect 22094 14968 22100 15020
rect 22152 14968 22158 15020
rect 24118 14968 24124 15020
rect 24176 14968 24182 15020
rect 24026 14940 24032 14952
rect 21008 14912 24032 14940
rect 24026 14900 24032 14912
rect 24084 14900 24090 14952
rect 24762 14900 24768 14952
rect 24820 14900 24826 14952
rect 13725 14875 13783 14881
rect 13725 14841 13737 14875
rect 13771 14872 13783 14875
rect 16666 14872 16672 14884
rect 13771 14844 16672 14872
rect 13771 14841 13783 14844
rect 13725 14835 13783 14841
rect 16666 14832 16672 14844
rect 16724 14832 16730 14884
rect 18874 14832 18880 14884
rect 18932 14832 18938 14884
rect 19613 14875 19671 14881
rect 19613 14841 19625 14875
rect 19659 14872 19671 14875
rect 19659 14844 24072 14872
rect 19659 14841 19671 14844
rect 19613 14835 19671 14841
rect 24044 14816 24072 14844
rect 8294 14804 8300 14816
rect 7760 14776 8300 14804
rect 8294 14764 8300 14776
rect 8352 14764 8358 14816
rect 20714 14764 20720 14816
rect 20772 14804 20778 14816
rect 20809 14807 20867 14813
rect 20809 14804 20821 14807
rect 20772 14776 20821 14804
rect 20772 14764 20778 14776
rect 20809 14773 20821 14776
rect 20855 14773 20867 14807
rect 20809 14767 20867 14773
rect 24026 14764 24032 14816
rect 24084 14764 24090 14816
rect 1104 14714 25852 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 25852 14714
rect 1104 14640 25852 14662
rect 7834 14560 7840 14612
rect 7892 14600 7898 14612
rect 8205 14603 8263 14609
rect 8205 14600 8217 14603
rect 7892 14572 8217 14600
rect 7892 14560 7898 14572
rect 8205 14569 8217 14572
rect 8251 14569 8263 14603
rect 8205 14563 8263 14569
rect 8573 14603 8631 14609
rect 8573 14569 8585 14603
rect 8619 14600 8631 14603
rect 8662 14600 8668 14612
rect 8619 14572 8668 14600
rect 8619 14569 8631 14572
rect 8573 14563 8631 14569
rect 8588 14532 8616 14563
rect 8662 14560 8668 14572
rect 8720 14560 8726 14612
rect 9306 14560 9312 14612
rect 9364 14600 9370 14612
rect 12437 14603 12495 14609
rect 9364 14572 11284 14600
rect 9364 14560 9370 14572
rect 9585 14535 9643 14541
rect 9585 14532 9597 14535
rect 8588 14504 9597 14532
rect 6454 14424 6460 14476
rect 6512 14464 6518 14476
rect 8294 14464 8300 14476
rect 6512 14436 8300 14464
rect 6512 14424 6518 14436
rect 8294 14424 8300 14436
rect 8352 14424 8358 14476
rect 8588 14396 8616 14504
rect 9585 14501 9597 14504
rect 9631 14501 9643 14535
rect 11256 14532 11284 14572
rect 12437 14569 12449 14603
rect 12483 14600 12495 14603
rect 12618 14600 12624 14612
rect 12483 14572 12624 14600
rect 12483 14569 12495 14572
rect 12437 14563 12495 14569
rect 12618 14560 12624 14572
rect 12676 14560 12682 14612
rect 21453 14603 21511 14609
rect 21453 14569 21465 14603
rect 21499 14600 21511 14603
rect 25038 14600 25044 14612
rect 21499 14572 25044 14600
rect 21499 14569 21511 14572
rect 21453 14563 21511 14569
rect 25038 14560 25044 14572
rect 25096 14560 25102 14612
rect 15746 14532 15752 14544
rect 11256 14504 15752 14532
rect 9585 14495 9643 14501
rect 9766 14424 9772 14476
rect 9824 14464 9830 14476
rect 10229 14467 10287 14473
rect 10229 14464 10241 14467
rect 9824 14436 10241 14464
rect 9824 14424 9830 14436
rect 10229 14433 10241 14436
rect 10275 14464 10287 14467
rect 11698 14464 11704 14476
rect 10275 14436 11704 14464
rect 10275 14433 10287 14436
rect 10229 14427 10287 14433
rect 11698 14424 11704 14436
rect 11756 14424 11762 14476
rect 13081 14467 13139 14473
rect 13081 14464 13093 14467
rect 12406 14436 13093 14464
rect 7866 14368 8616 14396
rect 9582 14356 9588 14408
rect 9640 14396 9646 14408
rect 9953 14399 10011 14405
rect 9953 14396 9965 14399
rect 9640 14368 9965 14396
rect 9640 14356 9646 14368
rect 9953 14365 9965 14368
rect 9999 14365 10011 14399
rect 9953 14359 10011 14365
rect 6733 14331 6791 14337
rect 6733 14297 6745 14331
rect 6779 14297 6791 14331
rect 9398 14328 9404 14340
rect 6733 14291 6791 14297
rect 8404 14300 9404 14328
rect 6748 14260 6776 14291
rect 8404 14260 8432 14300
rect 9398 14288 9404 14300
rect 9456 14288 9462 14340
rect 10870 14288 10876 14340
rect 10928 14288 10934 14340
rect 11977 14331 12035 14337
rect 11977 14297 11989 14331
rect 12023 14328 12035 14331
rect 12406 14328 12434 14436
rect 13081 14433 13093 14436
rect 13127 14464 13139 14467
rect 13446 14464 13452 14476
rect 13127 14436 13452 14464
rect 13127 14433 13139 14436
rect 13081 14427 13139 14433
rect 13446 14424 13452 14436
rect 13504 14424 13510 14476
rect 14844 14473 14872 14504
rect 15746 14492 15752 14504
rect 15804 14492 15810 14544
rect 16485 14535 16543 14541
rect 16485 14501 16497 14535
rect 16531 14532 16543 14535
rect 20346 14532 20352 14544
rect 16531 14504 20352 14532
rect 16531 14501 16543 14504
rect 16485 14495 16543 14501
rect 20346 14492 20352 14504
rect 20404 14492 20410 14544
rect 24302 14492 24308 14544
rect 24360 14532 24366 14544
rect 24360 14504 25084 14532
rect 24360 14492 24366 14504
rect 14829 14467 14887 14473
rect 14829 14433 14841 14467
rect 14875 14433 14887 14467
rect 14829 14427 14887 14433
rect 14918 14424 14924 14476
rect 14976 14464 14982 14476
rect 17037 14467 17095 14473
rect 17037 14464 17049 14467
rect 14976 14436 17049 14464
rect 14976 14424 14982 14436
rect 17037 14433 17049 14436
rect 17083 14433 17095 14467
rect 17037 14427 17095 14433
rect 21266 14424 21272 14476
rect 21324 14464 21330 14476
rect 21913 14467 21971 14473
rect 21913 14464 21925 14467
rect 21324 14436 21925 14464
rect 21324 14424 21330 14436
rect 21913 14433 21925 14436
rect 21959 14433 21971 14467
rect 21913 14427 21971 14433
rect 22097 14467 22155 14473
rect 22097 14433 22109 14467
rect 22143 14464 22155 14467
rect 23198 14464 23204 14476
rect 22143 14436 23204 14464
rect 22143 14433 22155 14436
rect 22097 14427 22155 14433
rect 23198 14424 23204 14436
rect 23256 14464 23262 14476
rect 23382 14464 23388 14476
rect 23256 14436 23388 14464
rect 23256 14424 23262 14436
rect 23382 14424 23388 14436
rect 23440 14424 23446 14476
rect 23845 14467 23903 14473
rect 23845 14433 23857 14467
rect 23891 14464 23903 14467
rect 24854 14464 24860 14476
rect 23891 14436 24860 14464
rect 23891 14433 23903 14436
rect 23845 14427 23903 14433
rect 24854 14424 24860 14436
rect 24912 14424 24918 14476
rect 14645 14399 14703 14405
rect 14645 14365 14657 14399
rect 14691 14396 14703 14399
rect 15381 14399 15439 14405
rect 15381 14396 15393 14399
rect 14691 14368 15393 14396
rect 14691 14365 14703 14368
rect 14645 14359 14703 14365
rect 15381 14365 15393 14368
rect 15427 14396 15439 14399
rect 20162 14396 20168 14408
rect 15427 14368 20168 14396
rect 15427 14365 15439 14368
rect 15381 14359 15439 14365
rect 20162 14356 20168 14368
rect 20220 14356 20226 14408
rect 20441 14399 20499 14405
rect 20441 14365 20453 14399
rect 20487 14396 20499 14399
rect 21726 14396 21732 14408
rect 20487 14368 21732 14396
rect 20487 14365 20499 14368
rect 20441 14359 20499 14365
rect 21726 14356 21732 14368
rect 21784 14356 21790 14408
rect 22833 14399 22891 14405
rect 22833 14365 22845 14399
rect 22879 14396 22891 14399
rect 24486 14396 24492 14408
rect 22879 14368 24492 14396
rect 22879 14365 22891 14368
rect 22833 14359 22891 14365
rect 24486 14356 24492 14368
rect 24544 14356 24550 14408
rect 25056 14405 25084 14504
rect 25041 14399 25099 14405
rect 25041 14365 25053 14399
rect 25087 14365 25099 14399
rect 25041 14359 25099 14365
rect 12023 14300 12434 14328
rect 16853 14331 16911 14337
rect 12023 14297 12035 14300
rect 11977 14291 12035 14297
rect 16853 14297 16865 14331
rect 16899 14328 16911 14331
rect 17681 14331 17739 14337
rect 17681 14328 17693 14331
rect 16899 14300 17693 14328
rect 16899 14297 16911 14300
rect 16853 14291 16911 14297
rect 17681 14297 17693 14300
rect 17727 14297 17739 14331
rect 17681 14291 17739 14297
rect 6748 14232 8432 14260
rect 10962 14220 10968 14272
rect 11020 14260 11026 14272
rect 11992 14260 12020 14291
rect 20898 14288 20904 14340
rect 20956 14328 20962 14340
rect 24394 14328 24400 14340
rect 20956 14300 24400 14328
rect 20956 14288 20962 14300
rect 24394 14288 24400 14300
rect 24452 14288 24458 14340
rect 11020 14232 12020 14260
rect 11020 14220 11026 14232
rect 12802 14220 12808 14272
rect 12860 14220 12866 14272
rect 12897 14263 12955 14269
rect 12897 14229 12909 14263
rect 12943 14260 12955 14263
rect 13354 14260 13360 14272
rect 12943 14232 13360 14260
rect 12943 14229 12955 14232
rect 12897 14223 12955 14229
rect 13354 14220 13360 14232
rect 13412 14220 13418 14272
rect 13538 14220 13544 14272
rect 13596 14220 13602 14272
rect 14277 14263 14335 14269
rect 14277 14229 14289 14263
rect 14323 14260 14335 14263
rect 14458 14260 14464 14272
rect 14323 14232 14464 14260
rect 14323 14229 14335 14232
rect 14277 14223 14335 14229
rect 14458 14220 14464 14232
rect 14516 14220 14522 14272
rect 14734 14220 14740 14272
rect 14792 14220 14798 14272
rect 16574 14220 16580 14272
rect 16632 14260 16638 14272
rect 16945 14263 17003 14269
rect 16945 14260 16957 14263
rect 16632 14232 16957 14260
rect 16632 14220 16638 14232
rect 16945 14229 16957 14232
rect 16991 14229 17003 14263
rect 16945 14223 17003 14229
rect 20254 14220 20260 14272
rect 20312 14220 20318 14272
rect 21818 14220 21824 14272
rect 21876 14220 21882 14272
rect 22002 14220 22008 14272
rect 22060 14260 22066 14272
rect 22462 14260 22468 14272
rect 22060 14232 22468 14260
rect 22060 14220 22066 14232
rect 22462 14220 22468 14232
rect 22520 14220 22526 14272
rect 24854 14220 24860 14272
rect 24912 14220 24918 14272
rect 1104 14170 25852 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 25852 14170
rect 1104 14096 25852 14118
rect 8294 14056 8300 14068
rect 7852 14028 8300 14056
rect 7852 13988 7880 14028
rect 8294 14016 8300 14028
rect 8352 14056 8358 14068
rect 9582 14056 9588 14068
rect 8352 14028 9588 14056
rect 8352 14016 8358 14028
rect 9582 14016 9588 14028
rect 9640 14016 9646 14068
rect 11606 14056 11612 14068
rect 10244 14028 11612 14056
rect 7760 13960 7880 13988
rect 7760 13929 7788 13960
rect 7926 13948 7932 14000
rect 7984 13988 7990 14000
rect 8021 13991 8079 13997
rect 8021 13988 8033 13991
rect 7984 13960 8033 13988
rect 7984 13948 7990 13960
rect 8021 13957 8033 13960
rect 8067 13957 8079 13991
rect 8021 13951 8079 13957
rect 8662 13948 8668 14000
rect 8720 13948 8726 14000
rect 9766 13948 9772 14000
rect 9824 13948 9830 14000
rect 10244 13997 10272 14028
rect 11606 14016 11612 14028
rect 11664 14056 11670 14068
rect 12161 14059 12219 14065
rect 12161 14056 12173 14059
rect 11664 14028 12173 14056
rect 11664 14016 11670 14028
rect 12161 14025 12173 14028
rect 12207 14056 12219 14059
rect 12342 14056 12348 14068
rect 12207 14028 12348 14056
rect 12207 14025 12219 14028
rect 12161 14019 12219 14025
rect 12342 14016 12348 14028
rect 12400 14016 12406 14068
rect 12989 14059 13047 14065
rect 12989 14025 13001 14059
rect 13035 14056 13047 14059
rect 13538 14056 13544 14068
rect 13035 14028 13544 14056
rect 13035 14025 13047 14028
rect 12989 14019 13047 14025
rect 13538 14016 13544 14028
rect 13596 14016 13602 14068
rect 14826 14016 14832 14068
rect 14884 14056 14890 14068
rect 15565 14059 15623 14065
rect 15565 14056 15577 14059
rect 14884 14028 15577 14056
rect 14884 14016 14890 14028
rect 15565 14025 15577 14028
rect 15611 14025 15623 14059
rect 15565 14019 15623 14025
rect 15933 14059 15991 14065
rect 15933 14025 15945 14059
rect 15979 14056 15991 14059
rect 16390 14056 16396 14068
rect 15979 14028 16396 14056
rect 15979 14025 15991 14028
rect 15933 14019 15991 14025
rect 10229 13991 10287 13997
rect 10229 13957 10241 13991
rect 10275 13957 10287 13991
rect 10229 13951 10287 13957
rect 13262 13948 13268 14000
rect 13320 13988 13326 14000
rect 15948 13988 15976 14019
rect 16390 14016 16396 14028
rect 16448 14016 16454 14068
rect 18598 14016 18604 14068
rect 18656 14056 18662 14068
rect 18782 14056 18788 14068
rect 18656 14028 18788 14056
rect 18656 14016 18662 14028
rect 18782 14016 18788 14028
rect 18840 14016 18846 14068
rect 18966 14016 18972 14068
rect 19024 14056 19030 14068
rect 19061 14059 19119 14065
rect 19061 14056 19073 14059
rect 19024 14028 19073 14056
rect 19024 14016 19030 14028
rect 19061 14025 19073 14028
rect 19107 14056 19119 14059
rect 19150 14056 19156 14068
rect 19107 14028 19156 14056
rect 19107 14025 19119 14028
rect 19061 14019 19119 14025
rect 19150 14016 19156 14028
rect 19208 14016 19214 14068
rect 20165 14059 20223 14065
rect 20165 14025 20177 14059
rect 20211 14056 20223 14059
rect 21082 14056 21088 14068
rect 20211 14028 21088 14056
rect 20211 14025 20223 14028
rect 20165 14019 20223 14025
rect 21082 14016 21088 14028
rect 21140 14016 21146 14068
rect 23474 14016 23480 14068
rect 23532 14056 23538 14068
rect 25041 14059 25099 14065
rect 25041 14056 25053 14059
rect 23532 14028 25053 14056
rect 23532 14016 23538 14028
rect 25041 14025 25053 14028
rect 25087 14025 25099 14059
rect 25041 14019 25099 14025
rect 18877 13991 18935 13997
rect 18877 13988 18889 13991
rect 13320 13960 13584 13988
rect 15318 13960 15976 13988
rect 18354 13960 18889 13988
rect 13320 13948 13326 13960
rect 13556 13932 13584 13960
rect 18877 13957 18889 13960
rect 18923 13988 18935 13991
rect 19242 13988 19248 14000
rect 18923 13960 19248 13988
rect 18923 13957 18935 13960
rect 18877 13951 18935 13957
rect 19242 13948 19248 13960
rect 19300 13948 19306 14000
rect 19521 13991 19579 13997
rect 19521 13957 19533 13991
rect 19567 13988 19579 13991
rect 22646 13988 22652 14000
rect 19567 13960 22048 13988
rect 19567 13957 19579 13960
rect 19521 13951 19579 13957
rect 7745 13923 7803 13929
rect 7745 13889 7757 13923
rect 7791 13889 7803 13923
rect 7745 13883 7803 13889
rect 9582 13880 9588 13932
rect 9640 13920 9646 13932
rect 10965 13923 11023 13929
rect 10965 13920 10977 13923
rect 9640 13892 10977 13920
rect 9640 13880 9646 13892
rect 10965 13889 10977 13892
rect 11011 13889 11023 13923
rect 10965 13883 11023 13889
rect 13538 13880 13544 13932
rect 13596 13880 13602 13932
rect 20346 13880 20352 13932
rect 20404 13880 20410 13932
rect 21085 13923 21143 13929
rect 21085 13889 21097 13923
rect 21131 13920 21143 13923
rect 21910 13920 21916 13932
rect 21131 13892 21916 13920
rect 21131 13889 21143 13892
rect 21085 13883 21143 13889
rect 21910 13880 21916 13892
rect 21968 13880 21974 13932
rect 22020 13920 22048 13960
rect 22112 13960 22652 13988
rect 22112 13920 22140 13960
rect 22646 13948 22652 13960
rect 22704 13948 22710 14000
rect 23658 13948 23664 14000
rect 23716 13948 23722 14000
rect 22020 13892 22140 13920
rect 22189 13923 22247 13929
rect 22189 13889 22201 13923
rect 22235 13920 22247 13923
rect 22278 13920 22284 13932
rect 22235 13892 22284 13920
rect 22235 13889 22247 13892
rect 22189 13883 22247 13889
rect 22278 13880 22284 13892
rect 22336 13880 22342 13932
rect 24394 13880 24400 13932
rect 24452 13920 24458 13932
rect 25225 13923 25283 13929
rect 25225 13920 25237 13923
rect 24452 13892 25237 13920
rect 24452 13880 24458 13892
rect 25225 13889 25237 13892
rect 25271 13889 25283 13923
rect 25225 13883 25283 13889
rect 11054 13812 11060 13864
rect 11112 13852 11118 13864
rect 11701 13855 11759 13861
rect 11701 13852 11713 13855
rect 11112 13824 11713 13852
rect 11112 13812 11118 13824
rect 11701 13821 11713 13824
rect 11747 13821 11759 13855
rect 11701 13815 11759 13821
rect 12710 13812 12716 13864
rect 12768 13852 12774 13864
rect 13081 13855 13139 13861
rect 13081 13852 13093 13855
rect 12768 13824 13093 13852
rect 12768 13812 12774 13824
rect 13081 13821 13093 13824
rect 13127 13821 13139 13855
rect 13081 13815 13139 13821
rect 13265 13855 13323 13861
rect 13265 13821 13277 13855
rect 13311 13821 13323 13855
rect 13265 13815 13323 13821
rect 11146 13676 11152 13728
rect 11204 13716 11210 13728
rect 12250 13716 12256 13728
rect 11204 13688 12256 13716
rect 11204 13676 11210 13688
rect 12250 13676 12256 13688
rect 12308 13676 12314 13728
rect 12618 13676 12624 13728
rect 12676 13676 12682 13728
rect 13280 13716 13308 13815
rect 13814 13812 13820 13864
rect 13872 13812 13878 13864
rect 16850 13812 16856 13864
rect 16908 13812 16914 13864
rect 19705 13855 19763 13861
rect 19705 13821 19717 13855
rect 19751 13852 19763 13855
rect 19886 13852 19892 13864
rect 19751 13824 19892 13852
rect 19751 13821 19763 13824
rect 19705 13815 19763 13821
rect 19886 13812 19892 13824
rect 19944 13812 19950 13864
rect 22370 13852 22376 13864
rect 20916 13824 21956 13852
rect 15102 13744 15108 13796
rect 15160 13784 15166 13796
rect 15654 13784 15660 13796
rect 15160 13756 15660 13784
rect 15160 13744 15166 13756
rect 15654 13744 15660 13756
rect 15712 13744 15718 13796
rect 20916 13793 20944 13824
rect 21928 13796 21956 13824
rect 22020 13824 22376 13852
rect 20901 13787 20959 13793
rect 20901 13753 20913 13787
rect 20947 13753 20959 13787
rect 20901 13747 20959 13753
rect 21910 13744 21916 13796
rect 21968 13744 21974 13796
rect 22020 13793 22048 13824
rect 22370 13812 22376 13824
rect 22428 13812 22434 13864
rect 22646 13812 22652 13864
rect 22704 13852 22710 13864
rect 22833 13855 22891 13861
rect 22833 13852 22845 13855
rect 22704 13824 22845 13852
rect 22704 13812 22710 13824
rect 22833 13821 22845 13824
rect 22879 13821 22891 13855
rect 22833 13815 22891 13821
rect 23198 13812 23204 13864
rect 23256 13852 23262 13864
rect 24581 13855 24639 13861
rect 24581 13852 24593 13855
rect 23256 13824 24593 13852
rect 23256 13812 23262 13824
rect 24581 13821 24593 13824
rect 24627 13821 24639 13855
rect 24581 13815 24639 13821
rect 22005 13787 22063 13793
rect 22005 13753 22017 13787
rect 22051 13753 22063 13787
rect 22005 13747 22063 13753
rect 13906 13716 13912 13728
rect 13280 13688 13912 13716
rect 13906 13676 13912 13688
rect 13964 13676 13970 13728
rect 14090 13725 14096 13728
rect 14080 13719 14096 13725
rect 14080 13685 14092 13719
rect 14080 13679 14096 13685
rect 14090 13676 14096 13679
rect 14148 13676 14154 13728
rect 17126 13725 17132 13728
rect 17116 13719 17132 13725
rect 17116 13685 17128 13719
rect 17184 13716 17190 13728
rect 17494 13716 17500 13728
rect 17184 13688 17500 13716
rect 17116 13679 17132 13685
rect 17126 13676 17132 13679
rect 17184 13676 17190 13688
rect 17494 13676 17500 13688
rect 17552 13676 17558 13728
rect 22462 13676 22468 13728
rect 22520 13716 22526 13728
rect 22830 13716 22836 13728
rect 22520 13688 22836 13716
rect 22520 13676 22526 13688
rect 22830 13676 22836 13688
rect 22888 13716 22894 13728
rect 23090 13719 23148 13725
rect 23090 13716 23102 13719
rect 22888 13688 23102 13716
rect 22888 13676 22894 13688
rect 23090 13685 23102 13688
rect 23136 13685 23148 13719
rect 23090 13679 23148 13685
rect 1104 13626 25852 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 25852 13626
rect 1104 13552 25852 13574
rect 8297 13515 8355 13521
rect 8297 13481 8309 13515
rect 8343 13512 8355 13515
rect 8478 13512 8484 13524
rect 8343 13484 8484 13512
rect 8343 13481 8355 13484
rect 8297 13475 8355 13481
rect 8478 13472 8484 13484
rect 8536 13472 8542 13524
rect 8662 13472 8668 13524
rect 8720 13472 8726 13524
rect 8846 13472 8852 13524
rect 8904 13512 8910 13524
rect 9217 13515 9275 13521
rect 9217 13512 9229 13515
rect 8904 13484 9229 13512
rect 8904 13472 8910 13484
rect 9217 13481 9229 13484
rect 9263 13481 9275 13515
rect 9217 13475 9275 13481
rect 10676 13515 10734 13521
rect 10676 13481 10688 13515
rect 10722 13512 10734 13515
rect 13630 13512 13636 13524
rect 10722 13484 13636 13512
rect 10722 13481 10734 13484
rect 10676 13475 10734 13481
rect 13630 13472 13636 13484
rect 13688 13472 13694 13524
rect 14274 13472 14280 13524
rect 14332 13512 14338 13524
rect 14737 13515 14795 13521
rect 14737 13512 14749 13515
rect 14332 13484 14749 13512
rect 14332 13472 14338 13484
rect 14737 13481 14749 13484
rect 14783 13512 14795 13515
rect 17310 13512 17316 13524
rect 14783 13484 17316 13512
rect 14783 13481 14795 13484
rect 14737 13475 14795 13481
rect 17310 13472 17316 13484
rect 17368 13472 17374 13524
rect 17402 13472 17408 13524
rect 17460 13472 17466 13524
rect 18322 13472 18328 13524
rect 18380 13512 18386 13524
rect 21174 13512 21180 13524
rect 18380 13484 21180 13512
rect 18380 13472 18386 13484
rect 21174 13472 21180 13484
rect 21232 13472 21238 13524
rect 24486 13472 24492 13524
rect 24544 13512 24550 13524
rect 24581 13515 24639 13521
rect 24581 13512 24593 13515
rect 24544 13484 24593 13512
rect 24544 13472 24550 13484
rect 24581 13481 24593 13484
rect 24627 13481 24639 13515
rect 24581 13475 24639 13481
rect 9398 13404 9404 13456
rect 9456 13444 9462 13456
rect 9582 13444 9588 13456
rect 9456 13416 9588 13444
rect 9456 13404 9462 13416
rect 9582 13404 9588 13416
rect 9640 13444 9646 13456
rect 9640 13416 9812 13444
rect 9640 13404 9646 13416
rect 6454 13336 6460 13388
rect 6512 13376 6518 13388
rect 6549 13379 6607 13385
rect 6549 13376 6561 13379
rect 6512 13348 6561 13376
rect 6512 13336 6518 13348
rect 6549 13345 6561 13348
rect 6595 13345 6607 13379
rect 6549 13339 6607 13345
rect 6825 13379 6883 13385
rect 6825 13345 6837 13379
rect 6871 13376 6883 13379
rect 9674 13376 9680 13388
rect 6871 13348 9680 13376
rect 6871 13345 6883 13348
rect 6825 13339 6883 13345
rect 9674 13336 9680 13348
rect 9732 13336 9738 13388
rect 9784 13385 9812 13416
rect 13170 13404 13176 13456
rect 13228 13444 13234 13456
rect 15102 13444 15108 13456
rect 13228 13416 15108 13444
rect 13228 13404 13234 13416
rect 15102 13404 15108 13416
rect 15160 13404 15166 13456
rect 16482 13404 16488 13456
rect 16540 13444 16546 13456
rect 19794 13444 19800 13456
rect 16540 13416 19800 13444
rect 16540 13404 16546 13416
rect 19794 13404 19800 13416
rect 19852 13404 19858 13456
rect 20898 13404 20904 13456
rect 20956 13444 20962 13456
rect 21591 13447 21649 13453
rect 21591 13444 21603 13447
rect 20956 13416 21603 13444
rect 20956 13404 20962 13416
rect 21591 13413 21603 13416
rect 21637 13413 21649 13447
rect 21591 13407 21649 13413
rect 22094 13404 22100 13456
rect 22152 13444 22158 13456
rect 22830 13444 22836 13456
rect 22152 13416 22836 13444
rect 22152 13404 22158 13416
rect 22830 13404 22836 13416
rect 22888 13404 22894 13456
rect 23658 13404 23664 13456
rect 23716 13444 23722 13456
rect 25041 13447 25099 13453
rect 25041 13444 25053 13447
rect 23716 13416 25053 13444
rect 23716 13404 23722 13416
rect 25041 13413 25053 13416
rect 25087 13413 25099 13447
rect 25041 13407 25099 13413
rect 9769 13379 9827 13385
rect 9769 13345 9781 13379
rect 9815 13345 9827 13379
rect 9769 13339 9827 13345
rect 10413 13379 10471 13385
rect 10413 13345 10425 13379
rect 10459 13376 10471 13379
rect 11698 13376 11704 13388
rect 10459 13348 11704 13376
rect 10459 13345 10471 13348
rect 10413 13339 10471 13345
rect 11698 13336 11704 13348
rect 11756 13376 11762 13388
rect 13449 13379 13507 13385
rect 13449 13376 13461 13379
rect 11756 13348 13461 13376
rect 11756 13336 11762 13348
rect 13449 13345 13461 13348
rect 13495 13376 13507 13379
rect 13814 13376 13820 13388
rect 13495 13348 13820 13376
rect 13495 13345 13507 13348
rect 13449 13339 13507 13345
rect 13814 13336 13820 13348
rect 13872 13336 13878 13388
rect 15746 13336 15752 13388
rect 15804 13376 15810 13388
rect 16206 13376 16212 13388
rect 15804 13348 16212 13376
rect 15804 13336 15810 13348
rect 16206 13336 16212 13348
rect 16264 13336 16270 13388
rect 17310 13336 17316 13388
rect 17368 13376 17374 13388
rect 17862 13376 17868 13388
rect 17368 13348 17868 13376
rect 17368 13336 17374 13348
rect 17862 13336 17868 13348
rect 17920 13336 17926 13388
rect 18049 13379 18107 13385
rect 18049 13345 18061 13379
rect 18095 13376 18107 13379
rect 18598 13376 18604 13388
rect 18095 13348 18604 13376
rect 18095 13345 18107 13348
rect 18049 13339 18107 13345
rect 18598 13336 18604 13348
rect 18656 13336 18662 13388
rect 20990 13376 20996 13388
rect 18708 13348 20996 13376
rect 13906 13268 13912 13320
rect 13964 13308 13970 13320
rect 15102 13308 15108 13320
rect 13964 13280 15108 13308
rect 13964 13268 13970 13280
rect 15102 13268 15108 13280
rect 15160 13268 15166 13320
rect 15657 13311 15715 13317
rect 15657 13308 15669 13311
rect 15212 13280 15669 13308
rect 8662 13240 8668 13252
rect 8050 13212 8668 13240
rect 8662 13200 8668 13212
rect 8720 13200 8726 13252
rect 9585 13243 9643 13249
rect 9585 13209 9597 13243
rect 9631 13240 9643 13243
rect 9631 13212 11100 13240
rect 9631 13209 9643 13212
rect 9585 13203 9643 13209
rect 9674 13132 9680 13184
rect 9732 13132 9738 13184
rect 11072 13172 11100 13212
rect 11146 13200 11152 13252
rect 11204 13200 11210 13252
rect 12342 13200 12348 13252
rect 12400 13240 12406 13252
rect 12621 13243 12679 13249
rect 12621 13240 12633 13243
rect 12400 13212 12633 13240
rect 12400 13200 12406 13212
rect 12621 13209 12633 13212
rect 12667 13209 12679 13243
rect 12621 13203 12679 13209
rect 11974 13172 11980 13184
rect 11072 13144 11980 13172
rect 11974 13132 11980 13144
rect 12032 13132 12038 13184
rect 12158 13132 12164 13184
rect 12216 13132 12222 13184
rect 12636 13172 12664 13203
rect 12894 13200 12900 13252
rect 12952 13240 12958 13252
rect 15212 13240 15240 13280
rect 15657 13277 15669 13280
rect 15703 13308 15715 13311
rect 15838 13308 15844 13320
rect 15703 13280 15844 13308
rect 15703 13277 15715 13280
rect 15657 13271 15715 13277
rect 15838 13268 15844 13280
rect 15896 13268 15902 13320
rect 16114 13268 16120 13320
rect 16172 13308 16178 13320
rect 18708 13308 18736 13348
rect 20990 13336 20996 13348
rect 21048 13336 21054 13388
rect 21082 13336 21088 13388
rect 21140 13376 21146 13388
rect 21140 13348 23612 13376
rect 21140 13336 21146 13348
rect 16172 13280 18736 13308
rect 16172 13268 16178 13280
rect 19334 13268 19340 13320
rect 19392 13308 19398 13320
rect 19429 13311 19487 13317
rect 19429 13308 19441 13311
rect 19392 13280 19441 13308
rect 19392 13268 19398 13280
rect 19429 13277 19441 13280
rect 19475 13308 19487 13311
rect 20625 13311 20683 13317
rect 20625 13308 20637 13311
rect 19475 13280 20637 13308
rect 19475 13277 19487 13280
rect 19429 13271 19487 13277
rect 20625 13277 20637 13280
rect 20671 13277 20683 13311
rect 20625 13271 20683 13277
rect 21361 13311 21419 13317
rect 21361 13277 21373 13311
rect 21407 13277 21419 13311
rect 21361 13271 21419 13277
rect 22833 13311 22891 13317
rect 22833 13277 22845 13311
rect 22879 13308 22891 13311
rect 23474 13308 23480 13320
rect 22879 13280 23480 13308
rect 22879 13277 22891 13280
rect 22833 13271 22891 13277
rect 12952 13212 15240 13240
rect 15565 13243 15623 13249
rect 12952 13200 12958 13212
rect 15565 13209 15577 13243
rect 15611 13240 15623 13243
rect 15611 13212 16344 13240
rect 15611 13209 15623 13212
rect 15565 13203 15623 13209
rect 16316 13184 16344 13212
rect 17402 13200 17408 13252
rect 17460 13240 17466 13252
rect 17865 13243 17923 13249
rect 17865 13240 17877 13243
rect 17460 13212 17877 13240
rect 17460 13200 17466 13212
rect 17865 13209 17877 13212
rect 17911 13209 17923 13243
rect 17865 13203 17923 13209
rect 18601 13243 18659 13249
rect 18601 13209 18613 13243
rect 18647 13209 18659 13243
rect 18601 13203 18659 13209
rect 18785 13243 18843 13249
rect 18785 13209 18797 13243
rect 18831 13240 18843 13243
rect 18966 13240 18972 13252
rect 18831 13212 18972 13240
rect 18831 13209 18843 13212
rect 18785 13203 18843 13209
rect 13906 13172 13912 13184
rect 12636 13144 13912 13172
rect 13906 13132 13912 13144
rect 13964 13132 13970 13184
rect 15194 13132 15200 13184
rect 15252 13132 15258 13184
rect 16298 13132 16304 13184
rect 16356 13132 16362 13184
rect 18616 13172 18644 13203
rect 18966 13200 18972 13212
rect 19024 13200 19030 13252
rect 20257 13243 20315 13249
rect 20257 13209 20269 13243
rect 20303 13240 20315 13243
rect 20438 13240 20444 13252
rect 20303 13212 20444 13240
rect 20303 13209 20315 13212
rect 20257 13203 20315 13209
rect 20438 13200 20444 13212
rect 20496 13200 20502 13252
rect 21376 13240 21404 13271
rect 23474 13268 23480 13280
rect 23532 13268 23538 13320
rect 23584 13308 23612 13348
rect 23842 13336 23848 13388
rect 23900 13336 23906 13388
rect 24765 13311 24823 13317
rect 24765 13308 24777 13311
rect 23584 13280 24777 13308
rect 24765 13277 24777 13280
rect 24811 13277 24823 13311
rect 24765 13271 24823 13277
rect 25130 13240 25136 13252
rect 21376 13212 25136 13240
rect 25130 13200 25136 13212
rect 25188 13200 25194 13252
rect 19150 13172 19156 13184
rect 18616 13144 19156 13172
rect 19150 13132 19156 13144
rect 19208 13132 19214 13184
rect 20162 13132 20168 13184
rect 20220 13172 20226 13184
rect 22554 13172 22560 13184
rect 20220 13144 22560 13172
rect 20220 13132 20226 13144
rect 22554 13132 22560 13144
rect 22612 13132 22618 13184
rect 1104 13082 25852 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 25852 13082
rect 1104 13008 25852 13030
rect 6641 12971 6699 12977
rect 6641 12937 6653 12971
rect 6687 12968 6699 12971
rect 7006 12968 7012 12980
rect 6687 12940 7012 12968
rect 6687 12937 6699 12940
rect 6641 12931 6699 12937
rect 7006 12928 7012 12940
rect 7064 12928 7070 12980
rect 9033 12971 9091 12977
rect 9033 12937 9045 12971
rect 9079 12968 9091 12971
rect 9214 12968 9220 12980
rect 9079 12940 9220 12968
rect 9079 12937 9091 12940
rect 9033 12931 9091 12937
rect 9214 12928 9220 12940
rect 9272 12928 9278 12980
rect 9398 12928 9404 12980
rect 9456 12928 9462 12980
rect 10042 12928 10048 12980
rect 10100 12968 10106 12980
rect 10413 12971 10471 12977
rect 10413 12968 10425 12971
rect 10100 12940 10425 12968
rect 10100 12928 10106 12940
rect 10413 12937 10425 12940
rect 10459 12937 10471 12971
rect 10413 12931 10471 12937
rect 10781 12971 10839 12977
rect 10781 12937 10793 12971
rect 10827 12968 10839 12971
rect 11054 12968 11060 12980
rect 10827 12940 11060 12968
rect 10827 12937 10839 12940
rect 10781 12931 10839 12937
rect 11054 12928 11060 12940
rect 11112 12928 11118 12980
rect 12250 12928 12256 12980
rect 12308 12928 12314 12980
rect 13078 12928 13084 12980
rect 13136 12968 13142 12980
rect 15013 12971 15071 12977
rect 15013 12968 15025 12971
rect 13136 12940 15025 12968
rect 13136 12928 13142 12940
rect 15013 12937 15025 12940
rect 15059 12937 15071 12971
rect 15013 12931 15071 12937
rect 15470 12928 15476 12980
rect 15528 12928 15534 12980
rect 16114 12968 16120 12980
rect 15856 12940 16120 12968
rect 6914 12860 6920 12912
rect 6972 12900 6978 12912
rect 12618 12900 12624 12912
rect 6972 12872 7236 12900
rect 6972 12860 6978 12872
rect 7006 12792 7012 12844
rect 7064 12792 7070 12844
rect 6914 12724 6920 12776
rect 6972 12764 6978 12776
rect 7208 12773 7236 12872
rect 9508 12872 12624 12900
rect 8202 12792 8208 12844
rect 8260 12792 8266 12844
rect 9508 12841 9536 12872
rect 12618 12860 12624 12872
rect 12676 12860 12682 12912
rect 12989 12903 13047 12909
rect 12989 12869 13001 12903
rect 13035 12900 13047 12903
rect 13998 12900 14004 12912
rect 13035 12872 14004 12900
rect 13035 12869 13047 12872
rect 12989 12863 13047 12869
rect 13998 12860 14004 12872
rect 14056 12860 14062 12912
rect 14274 12860 14280 12912
rect 14332 12860 14338 12912
rect 15381 12903 15439 12909
rect 15381 12869 15393 12903
rect 15427 12900 15439 12903
rect 15856 12900 15884 12940
rect 16114 12928 16120 12940
rect 16172 12928 16178 12980
rect 17218 12928 17224 12980
rect 17276 12968 17282 12980
rect 17313 12971 17371 12977
rect 17313 12968 17325 12971
rect 17276 12940 17325 12968
rect 17276 12928 17282 12940
rect 17313 12937 17325 12940
rect 17359 12937 17371 12971
rect 19245 12971 19303 12977
rect 19245 12968 19257 12971
rect 17313 12931 17371 12937
rect 17420 12940 19257 12968
rect 15427 12872 15884 12900
rect 15427 12869 15439 12872
rect 15381 12863 15439 12869
rect 15930 12860 15936 12912
rect 15988 12900 15994 12912
rect 17420 12900 17448 12940
rect 19245 12937 19257 12940
rect 19291 12937 19303 12971
rect 19245 12931 19303 12937
rect 19794 12928 19800 12980
rect 19852 12968 19858 12980
rect 21085 12971 21143 12977
rect 21085 12968 21097 12971
rect 19852 12940 21097 12968
rect 19852 12928 19858 12940
rect 21085 12937 21097 12940
rect 21131 12937 21143 12971
rect 21085 12931 21143 12937
rect 21174 12928 21180 12980
rect 21232 12968 21238 12980
rect 22465 12971 22523 12977
rect 22465 12968 22477 12971
rect 21232 12940 22477 12968
rect 21232 12928 21238 12940
rect 22465 12937 22477 12940
rect 22511 12937 22523 12971
rect 22465 12931 22523 12937
rect 22741 12971 22799 12977
rect 22741 12937 22753 12971
rect 22787 12968 22799 12971
rect 23658 12968 23664 12980
rect 22787 12940 23664 12968
rect 22787 12937 22799 12940
rect 22741 12931 22799 12937
rect 15988 12872 17448 12900
rect 15988 12860 15994 12872
rect 18046 12860 18052 12912
rect 18104 12900 18110 12912
rect 22278 12900 22284 12912
rect 18104 12872 22284 12900
rect 18104 12860 18110 12872
rect 22278 12860 22284 12872
rect 22336 12860 22342 12912
rect 22370 12860 22376 12912
rect 22428 12900 22434 12912
rect 22756 12900 22784 12931
rect 23658 12928 23664 12940
rect 23716 12968 23722 12980
rect 25133 12971 25191 12977
rect 25133 12968 25145 12971
rect 23716 12940 25145 12968
rect 23716 12928 23722 12940
rect 22428 12872 22784 12900
rect 22428 12860 22434 12872
rect 23382 12860 23388 12912
rect 23440 12860 23446 12912
rect 23768 12900 23796 12940
rect 25133 12937 25145 12940
rect 25179 12937 25191 12971
rect 25133 12931 25191 12937
rect 23768 12872 23874 12900
rect 9493 12835 9551 12841
rect 9493 12801 9505 12835
rect 9539 12801 9551 12835
rect 9493 12795 9551 12801
rect 10873 12835 10931 12841
rect 10873 12801 10885 12835
rect 10919 12832 10931 12835
rect 10919 12804 11652 12832
rect 10919 12801 10931 12804
rect 10873 12795 10931 12801
rect 7101 12767 7159 12773
rect 7101 12764 7113 12767
rect 6972 12736 7113 12764
rect 6972 12724 6978 12736
rect 7101 12733 7113 12736
rect 7147 12733 7159 12767
rect 7101 12727 7159 12733
rect 7193 12767 7251 12773
rect 7193 12733 7205 12767
rect 7239 12733 7251 12767
rect 7193 12727 7251 12733
rect 7650 12724 7656 12776
rect 7708 12764 7714 12776
rect 8297 12767 8355 12773
rect 8297 12764 8309 12767
rect 7708 12736 8309 12764
rect 7708 12724 7714 12736
rect 8297 12733 8309 12736
rect 8343 12733 8355 12767
rect 8297 12727 8355 12733
rect 8386 12724 8392 12776
rect 8444 12724 8450 12776
rect 9677 12767 9735 12773
rect 9677 12733 9689 12767
rect 9723 12764 9735 12767
rect 9766 12764 9772 12776
rect 9723 12736 9772 12764
rect 9723 12733 9735 12736
rect 9677 12727 9735 12733
rect 9766 12724 9772 12736
rect 9824 12764 9830 12776
rect 9950 12764 9956 12776
rect 9824 12736 9956 12764
rect 9824 12724 9830 12736
rect 9950 12724 9956 12736
rect 10008 12764 10014 12776
rect 10962 12764 10968 12776
rect 10008 12736 10968 12764
rect 10008 12724 10014 12736
rect 10962 12724 10968 12736
rect 11020 12724 11026 12776
rect 11624 12764 11652 12804
rect 11790 12792 11796 12844
rect 11848 12832 11854 12844
rect 12894 12832 12900 12844
rect 11848 12804 12900 12832
rect 11848 12792 11854 12804
rect 12894 12792 12900 12804
rect 12952 12792 12958 12844
rect 13081 12835 13139 12841
rect 13081 12801 13093 12835
rect 13127 12832 13139 12835
rect 13538 12832 13544 12844
rect 13127 12804 13544 12832
rect 13127 12801 13139 12804
rect 13081 12795 13139 12801
rect 13538 12792 13544 12804
rect 13596 12792 13602 12844
rect 13722 12792 13728 12844
rect 13780 12832 13786 12844
rect 14185 12835 14243 12841
rect 14185 12832 14197 12835
rect 13780 12804 14197 12832
rect 13780 12792 13786 12804
rect 14185 12801 14197 12804
rect 14231 12801 14243 12835
rect 14185 12795 14243 12801
rect 14918 12792 14924 12844
rect 14976 12832 14982 12844
rect 16482 12832 16488 12844
rect 14976 12804 16488 12832
rect 14976 12792 14982 12804
rect 16482 12792 16488 12804
rect 16540 12792 16546 12844
rect 17218 12792 17224 12844
rect 17276 12792 17282 12844
rect 18233 12835 18291 12841
rect 18233 12832 18245 12835
rect 17328 12804 18245 12832
rect 13170 12764 13176 12776
rect 11624 12736 13176 12764
rect 13170 12724 13176 12736
rect 13228 12724 13234 12776
rect 13265 12767 13323 12773
rect 13265 12733 13277 12767
rect 13311 12764 13323 12767
rect 13446 12764 13452 12776
rect 13311 12736 13452 12764
rect 13311 12733 13323 12736
rect 13265 12727 13323 12733
rect 13446 12724 13452 12736
rect 13504 12724 13510 12776
rect 14274 12724 14280 12776
rect 14332 12764 14338 12776
rect 14369 12767 14427 12773
rect 14369 12764 14381 12767
rect 14332 12736 14381 12764
rect 14332 12724 14338 12736
rect 14369 12733 14381 12736
rect 14415 12733 14427 12767
rect 14369 12727 14427 12733
rect 14826 12724 14832 12776
rect 14884 12764 14890 12776
rect 15102 12764 15108 12776
rect 14884 12736 15108 12764
rect 14884 12724 14890 12736
rect 15102 12724 15108 12736
rect 15160 12764 15166 12776
rect 15565 12767 15623 12773
rect 15565 12764 15577 12767
rect 15160 12736 15577 12764
rect 15160 12724 15166 12736
rect 15565 12733 15577 12736
rect 15611 12733 15623 12767
rect 15565 12727 15623 12733
rect 15654 12724 15660 12776
rect 15712 12764 15718 12776
rect 17328 12764 17356 12804
rect 18233 12801 18245 12804
rect 18279 12801 18291 12835
rect 18233 12795 18291 12801
rect 19150 12792 19156 12844
rect 19208 12792 19214 12844
rect 20162 12792 20168 12844
rect 20220 12792 20226 12844
rect 20346 12792 20352 12844
rect 20404 12832 20410 12844
rect 22189 12835 22247 12841
rect 22189 12832 22201 12835
rect 20404 12804 22201 12832
rect 20404 12792 20410 12804
rect 22189 12801 22201 12804
rect 22235 12801 22247 12835
rect 22189 12795 22247 12801
rect 15712 12736 17356 12764
rect 17497 12767 17555 12773
rect 15712 12724 15718 12736
rect 17497 12733 17509 12767
rect 17543 12764 17555 12767
rect 18782 12764 18788 12776
rect 17543 12736 18788 12764
rect 17543 12733 17555 12736
rect 17497 12727 17555 12733
rect 18782 12724 18788 12736
rect 18840 12724 18846 12776
rect 19429 12767 19487 12773
rect 19429 12733 19441 12767
rect 19475 12764 19487 12767
rect 20622 12764 20628 12776
rect 19475 12736 20628 12764
rect 19475 12733 19487 12736
rect 19429 12727 19487 12733
rect 20622 12724 20628 12736
rect 20680 12724 20686 12776
rect 21361 12767 21419 12773
rect 21361 12733 21373 12767
rect 21407 12733 21419 12767
rect 21361 12727 21419 12733
rect 7837 12699 7895 12705
rect 7837 12665 7849 12699
rect 7883 12696 7895 12699
rect 11330 12696 11336 12708
rect 7883 12668 11336 12696
rect 7883 12665 7895 12668
rect 7837 12659 7895 12665
rect 11330 12656 11336 12668
rect 11388 12656 11394 12708
rect 12342 12656 12348 12708
rect 12400 12696 12406 12708
rect 19981 12699 20039 12705
rect 19981 12696 19993 12699
rect 12400 12668 19993 12696
rect 12400 12656 12406 12668
rect 19981 12665 19993 12668
rect 20027 12665 20039 12699
rect 20806 12696 20812 12708
rect 19981 12659 20039 12665
rect 20088 12668 20812 12696
rect 11238 12588 11244 12640
rect 11296 12628 11302 12640
rect 11790 12628 11796 12640
rect 11296 12600 11796 12628
rect 11296 12588 11302 12600
rect 11790 12588 11796 12600
rect 11848 12588 11854 12640
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 12621 12631 12679 12637
rect 12621 12628 12633 12631
rect 12492 12600 12633 12628
rect 12492 12588 12498 12600
rect 12621 12597 12633 12600
rect 12667 12597 12679 12631
rect 12621 12591 12679 12597
rect 13817 12631 13875 12637
rect 13817 12597 13829 12631
rect 13863 12628 13875 12631
rect 16574 12628 16580 12640
rect 13863 12600 16580 12628
rect 13863 12597 13875 12600
rect 13817 12591 13875 12597
rect 16574 12588 16580 12600
rect 16632 12588 16638 12640
rect 16853 12631 16911 12637
rect 16853 12597 16865 12631
rect 16899 12628 16911 12631
rect 17402 12628 17408 12640
rect 16899 12600 17408 12628
rect 16899 12597 16911 12600
rect 16853 12591 16911 12597
rect 17402 12588 17408 12600
rect 17460 12588 17466 12640
rect 18046 12588 18052 12640
rect 18104 12588 18110 12640
rect 18785 12631 18843 12637
rect 18785 12597 18797 12631
rect 18831 12628 18843 12631
rect 20088 12628 20116 12668
rect 20806 12656 20812 12668
rect 20864 12656 20870 12708
rect 21376 12696 21404 12727
rect 22646 12724 22652 12776
rect 22704 12764 22710 12776
rect 23109 12767 23167 12773
rect 23109 12764 23121 12767
rect 22704 12736 23121 12764
rect 22704 12724 22710 12736
rect 23109 12733 23121 12736
rect 23155 12733 23167 12767
rect 23109 12727 23167 12733
rect 21376 12668 23244 12696
rect 18831 12600 20116 12628
rect 20717 12631 20775 12637
rect 18831 12597 18843 12600
rect 18785 12591 18843 12597
rect 20717 12597 20729 12631
rect 20763 12628 20775 12631
rect 21910 12628 21916 12640
rect 20763 12600 21916 12628
rect 20763 12597 20775 12600
rect 20717 12591 20775 12597
rect 21910 12588 21916 12600
rect 21968 12588 21974 12640
rect 22005 12631 22063 12637
rect 22005 12597 22017 12631
rect 22051 12628 22063 12631
rect 22830 12628 22836 12640
rect 22051 12600 22836 12628
rect 22051 12597 22063 12600
rect 22005 12591 22063 12597
rect 22830 12588 22836 12600
rect 22888 12588 22894 12640
rect 23216 12628 23244 12668
rect 23382 12628 23388 12640
rect 23216 12600 23388 12628
rect 23382 12588 23388 12600
rect 23440 12628 23446 12640
rect 24857 12631 24915 12637
rect 24857 12628 24869 12631
rect 23440 12600 24869 12628
rect 23440 12588 23446 12600
rect 24857 12597 24869 12600
rect 24903 12597 24915 12631
rect 24857 12591 24915 12597
rect 1104 12538 25852 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 25852 12538
rect 1104 12464 25852 12486
rect 7742 12384 7748 12436
rect 7800 12424 7806 12436
rect 10229 12427 10287 12433
rect 10229 12424 10241 12427
rect 7800 12396 10241 12424
rect 7800 12384 7806 12396
rect 10229 12393 10241 12396
rect 10275 12393 10287 12427
rect 10229 12387 10287 12393
rect 11422 12384 11428 12436
rect 11480 12384 11486 12436
rect 12526 12384 12532 12436
rect 12584 12424 12590 12436
rect 12621 12427 12679 12433
rect 12621 12424 12633 12427
rect 12584 12396 12633 12424
rect 12584 12384 12590 12396
rect 12621 12393 12633 12396
rect 12667 12393 12679 12427
rect 12621 12387 12679 12393
rect 13906 12384 13912 12436
rect 13964 12424 13970 12436
rect 16301 12427 16359 12433
rect 16301 12424 16313 12427
rect 13964 12396 16313 12424
rect 13964 12384 13970 12396
rect 16301 12393 16313 12396
rect 16347 12424 16359 12427
rect 17310 12424 17316 12436
rect 16347 12396 17316 12424
rect 16347 12393 16359 12396
rect 16301 12387 16359 12393
rect 17310 12384 17316 12396
rect 17368 12384 17374 12436
rect 18874 12424 18880 12436
rect 17512 12396 18880 12424
rect 12066 12316 12072 12368
rect 12124 12356 12130 12368
rect 13078 12356 13084 12368
rect 12124 12328 13084 12356
rect 12124 12316 12130 12328
rect 13078 12316 13084 12328
rect 13136 12316 13142 12368
rect 14182 12316 14188 12368
rect 14240 12356 14246 12368
rect 14277 12359 14335 12365
rect 14277 12356 14289 12359
rect 14240 12328 14289 12356
rect 14240 12316 14246 12328
rect 14277 12325 14289 12328
rect 14323 12325 14335 12359
rect 14277 12319 14335 12325
rect 14642 12316 14648 12368
rect 14700 12356 14706 12368
rect 17512 12356 17540 12396
rect 18874 12384 18880 12396
rect 18932 12424 18938 12436
rect 19242 12424 19248 12436
rect 18932 12396 19248 12424
rect 18932 12384 18938 12396
rect 19242 12384 19248 12396
rect 19300 12384 19306 12436
rect 20070 12384 20076 12436
rect 20128 12384 20134 12436
rect 22189 12427 22247 12433
rect 22189 12424 22201 12427
rect 20548 12396 22201 12424
rect 14700 12328 17540 12356
rect 14700 12316 14706 12328
rect 17586 12316 17592 12368
rect 17644 12356 17650 12368
rect 19518 12356 19524 12368
rect 17644 12328 19524 12356
rect 17644 12316 17650 12328
rect 19518 12316 19524 12328
rect 19576 12316 19582 12368
rect 19702 12316 19708 12368
rect 19760 12356 19766 12368
rect 20548 12356 20576 12396
rect 22189 12393 22201 12396
rect 22235 12393 22247 12427
rect 22189 12387 22247 12393
rect 24118 12384 24124 12436
rect 24176 12424 24182 12436
rect 24581 12427 24639 12433
rect 24581 12424 24593 12427
rect 24176 12396 24593 12424
rect 24176 12384 24182 12396
rect 24581 12393 24593 12396
rect 24627 12393 24639 12427
rect 24581 12387 24639 12393
rect 19760 12328 20576 12356
rect 19760 12316 19766 12328
rect 7006 12248 7012 12300
rect 7064 12288 7070 12300
rect 7377 12291 7435 12297
rect 7377 12288 7389 12291
rect 7064 12260 7389 12288
rect 7064 12248 7070 12260
rect 7377 12257 7389 12260
rect 7423 12257 7435 12291
rect 7377 12251 7435 12257
rect 8202 12248 8208 12300
rect 8260 12248 8266 12300
rect 9582 12248 9588 12300
rect 9640 12288 9646 12300
rect 10781 12291 10839 12297
rect 10781 12288 10793 12291
rect 9640 12260 10793 12288
rect 9640 12248 9646 12260
rect 10781 12257 10793 12260
rect 10827 12257 10839 12291
rect 10781 12251 10839 12257
rect 10962 12248 10968 12300
rect 11020 12288 11026 12300
rect 11977 12291 12035 12297
rect 11977 12288 11989 12291
rect 11020 12260 11989 12288
rect 11020 12248 11026 12260
rect 11977 12257 11989 12260
rect 12023 12288 12035 12291
rect 12158 12288 12164 12300
rect 12023 12260 12164 12288
rect 12023 12257 12035 12260
rect 11977 12251 12035 12257
rect 12158 12248 12164 12260
rect 12216 12248 12222 12300
rect 13265 12291 13323 12297
rect 13265 12257 13277 12291
rect 13311 12288 13323 12291
rect 13630 12288 13636 12300
rect 13311 12260 13636 12288
rect 13311 12257 13323 12260
rect 13265 12251 13323 12257
rect 13630 12248 13636 12260
rect 13688 12248 13694 12300
rect 13906 12248 13912 12300
rect 13964 12288 13970 12300
rect 14550 12288 14556 12300
rect 13964 12260 14556 12288
rect 13964 12248 13970 12260
rect 14550 12248 14556 12260
rect 14608 12288 14614 12300
rect 14737 12291 14795 12297
rect 14737 12288 14749 12291
rect 14608 12260 14749 12288
rect 14608 12248 14614 12260
rect 14737 12257 14749 12260
rect 14783 12257 14795 12291
rect 14737 12251 14795 12257
rect 14921 12291 14979 12297
rect 14921 12257 14933 12291
rect 14967 12288 14979 12291
rect 15102 12288 15108 12300
rect 14967 12260 15108 12288
rect 14967 12257 14979 12260
rect 14921 12251 14979 12257
rect 15102 12248 15108 12260
rect 15160 12248 15166 12300
rect 16390 12248 16396 12300
rect 16448 12288 16454 12300
rect 18414 12288 18420 12300
rect 16448 12260 18420 12288
rect 16448 12248 16454 12260
rect 18414 12248 18420 12260
rect 18472 12248 18478 12300
rect 18693 12291 18751 12297
rect 18693 12257 18705 12291
rect 18739 12288 18751 12291
rect 19150 12288 19156 12300
rect 18739 12260 19156 12288
rect 18739 12257 18751 12260
rect 18693 12251 18751 12257
rect 19150 12248 19156 12260
rect 19208 12248 19214 12300
rect 20438 12248 20444 12300
rect 20496 12248 20502 12300
rect 20717 12291 20775 12297
rect 20717 12257 20729 12291
rect 20763 12288 20775 12291
rect 21266 12288 21272 12300
rect 20763 12260 21272 12288
rect 20763 12257 20775 12260
rect 20717 12251 20775 12257
rect 21266 12248 21272 12260
rect 21324 12248 21330 12300
rect 11793 12223 11851 12229
rect 11793 12189 11805 12223
rect 11839 12220 11851 12223
rect 12434 12220 12440 12232
rect 11839 12192 12440 12220
rect 11839 12189 11851 12192
rect 11793 12183 11851 12189
rect 12434 12180 12440 12192
rect 12492 12180 12498 12232
rect 12526 12180 12532 12232
rect 12584 12220 12590 12232
rect 13081 12223 13139 12229
rect 13081 12220 13093 12223
rect 12584 12192 13093 12220
rect 12584 12180 12590 12192
rect 13081 12189 13093 12192
rect 13127 12220 13139 12223
rect 13722 12220 13728 12232
rect 13127 12192 13728 12220
rect 13127 12189 13139 12192
rect 13081 12183 13139 12189
rect 13722 12180 13728 12192
rect 13780 12180 13786 12232
rect 17310 12180 17316 12232
rect 17368 12180 17374 12232
rect 19521 12223 19579 12229
rect 19521 12189 19533 12223
rect 19567 12220 19579 12223
rect 20070 12220 20076 12232
rect 19567 12192 20076 12220
rect 19567 12189 19579 12192
rect 19521 12183 19579 12189
rect 20070 12180 20076 12192
rect 20128 12180 20134 12232
rect 21818 12180 21824 12232
rect 21876 12220 21882 12232
rect 22370 12220 22376 12232
rect 21876 12192 22376 12220
rect 21876 12180 21882 12192
rect 22370 12180 22376 12192
rect 22428 12180 22434 12232
rect 22830 12180 22836 12232
rect 22888 12180 22894 12232
rect 24765 12223 24823 12229
rect 24765 12220 24777 12223
rect 22940 12192 24777 12220
rect 10689 12155 10747 12161
rect 10689 12121 10701 12155
rect 10735 12152 10747 12155
rect 12618 12152 12624 12164
rect 10735 12124 12624 12152
rect 10735 12121 10747 12124
rect 10689 12115 10747 12121
rect 12618 12112 12624 12124
rect 12676 12112 12682 12164
rect 13446 12152 13452 12164
rect 12912 12124 13452 12152
rect 10594 12044 10600 12096
rect 10652 12044 10658 12096
rect 11885 12087 11943 12093
rect 11885 12053 11897 12087
rect 11931 12084 11943 12087
rect 12912 12084 12940 12124
rect 13446 12112 13452 12124
rect 13504 12112 13510 12164
rect 16390 12152 16396 12164
rect 14568 12124 16396 12152
rect 11931 12056 12940 12084
rect 12989 12087 13047 12093
rect 11931 12053 11943 12056
rect 11885 12047 11943 12053
rect 12989 12053 13001 12087
rect 13035 12084 13047 12087
rect 14568 12084 14596 12124
rect 16390 12112 16396 12124
rect 16448 12112 16454 12164
rect 16942 12112 16948 12164
rect 17000 12152 17006 12164
rect 18049 12155 18107 12161
rect 18049 12152 18061 12155
rect 17000 12124 18061 12152
rect 17000 12112 17006 12124
rect 18049 12121 18061 12124
rect 18095 12121 18107 12155
rect 18049 12115 18107 12121
rect 13035 12056 14596 12084
rect 14645 12087 14703 12093
rect 13035 12053 13047 12056
rect 12989 12047 13047 12053
rect 14645 12053 14657 12087
rect 14691 12084 14703 12087
rect 15010 12084 15016 12096
rect 14691 12056 15016 12084
rect 14691 12053 14703 12056
rect 14645 12047 14703 12053
rect 15010 12044 15016 12056
rect 15068 12044 15074 12096
rect 15286 12044 15292 12096
rect 15344 12084 15350 12096
rect 15838 12084 15844 12096
rect 15344 12056 15844 12084
rect 15344 12044 15350 12056
rect 15838 12044 15844 12056
rect 15896 12044 15902 12096
rect 16669 12087 16727 12093
rect 16669 12053 16681 12087
rect 16715 12084 16727 12087
rect 18414 12084 18420 12096
rect 16715 12056 18420 12084
rect 16715 12053 16727 12056
rect 16669 12047 16727 12053
rect 18414 12044 18420 12056
rect 18472 12044 18478 12096
rect 18966 12044 18972 12096
rect 19024 12084 19030 12096
rect 19613 12087 19671 12093
rect 19613 12084 19625 12087
rect 19024 12056 19625 12084
rect 19024 12044 19030 12056
rect 19613 12053 19625 12056
rect 19659 12053 19671 12087
rect 19613 12047 19671 12053
rect 20990 12044 20996 12096
rect 21048 12084 21054 12096
rect 22940 12084 22968 12192
rect 24765 12189 24777 12192
rect 24811 12189 24823 12223
rect 24765 12183 24823 12189
rect 23845 12155 23903 12161
rect 23845 12121 23857 12155
rect 23891 12152 23903 12155
rect 24946 12152 24952 12164
rect 23891 12124 24952 12152
rect 23891 12121 23903 12124
rect 23845 12115 23903 12121
rect 24946 12112 24952 12124
rect 25004 12112 25010 12164
rect 21048 12056 22968 12084
rect 21048 12044 21054 12056
rect 1104 11994 25852 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 25852 11994
rect 1104 11920 25852 11942
rect 5258 11840 5264 11892
rect 5316 11880 5322 11892
rect 9033 11883 9091 11889
rect 5316 11852 8892 11880
rect 5316 11840 5322 11852
rect 8864 11812 8892 11852
rect 9033 11849 9045 11883
rect 9079 11880 9091 11883
rect 9582 11880 9588 11892
rect 9079 11852 9588 11880
rect 9079 11849 9091 11852
rect 9033 11843 9091 11849
rect 9582 11840 9588 11852
rect 9640 11840 9646 11892
rect 9674 11840 9680 11892
rect 9732 11880 9738 11892
rect 9861 11883 9919 11889
rect 9861 11880 9873 11883
rect 9732 11852 9873 11880
rect 9732 11840 9738 11852
rect 9861 11849 9873 11852
rect 9907 11849 9919 11883
rect 11146 11880 11152 11892
rect 9861 11843 9919 11849
rect 10244 11852 11152 11880
rect 10244 11821 10272 11852
rect 11146 11840 11152 11852
rect 11204 11840 11210 11892
rect 11885 11883 11943 11889
rect 11885 11849 11897 11883
rect 11931 11880 11943 11883
rect 12802 11880 12808 11892
rect 11931 11852 12808 11880
rect 11931 11849 11943 11852
rect 11885 11843 11943 11849
rect 12802 11840 12808 11852
rect 12860 11840 12866 11892
rect 13078 11840 13084 11892
rect 13136 11840 13142 11892
rect 13446 11840 13452 11892
rect 13504 11880 13510 11892
rect 14182 11880 14188 11892
rect 13504 11852 14188 11880
rect 13504 11840 13510 11852
rect 14182 11840 14188 11852
rect 14240 11840 14246 11892
rect 14277 11883 14335 11889
rect 14277 11849 14289 11883
rect 14323 11880 14335 11883
rect 14366 11880 14372 11892
rect 14323 11852 14372 11880
rect 14323 11849 14335 11852
rect 14277 11843 14335 11849
rect 14366 11840 14372 11852
rect 14424 11840 14430 11892
rect 16758 11840 16764 11892
rect 16816 11880 16822 11892
rect 17313 11883 17371 11889
rect 17313 11880 17325 11883
rect 16816 11852 17325 11880
rect 16816 11840 16822 11852
rect 17313 11849 17325 11852
rect 17359 11849 17371 11883
rect 17313 11843 17371 11849
rect 18049 11883 18107 11889
rect 18049 11849 18061 11883
rect 18095 11849 18107 11883
rect 18049 11843 18107 11849
rect 9493 11815 9551 11821
rect 9493 11812 9505 11815
rect 8864 11784 9505 11812
rect 9493 11781 9505 11784
rect 9539 11812 9551 11815
rect 10229 11815 10287 11821
rect 10229 11812 10241 11815
rect 9539 11784 10241 11812
rect 9539 11781 9551 11784
rect 9493 11775 9551 11781
rect 10229 11781 10241 11784
rect 10275 11781 10287 11815
rect 10229 11775 10287 11781
rect 10321 11815 10379 11821
rect 10321 11781 10333 11815
rect 10367 11781 10379 11815
rect 10321 11775 10379 11781
rect 8662 11704 8668 11756
rect 8720 11744 8726 11756
rect 9309 11747 9367 11753
rect 9309 11744 9321 11747
rect 8720 11716 9321 11744
rect 8720 11704 8726 11716
rect 9309 11713 9321 11716
rect 9355 11713 9367 11747
rect 10336 11744 10364 11775
rect 11790 11772 11796 11824
rect 11848 11812 11854 11824
rect 12253 11815 12311 11821
rect 12253 11812 12265 11815
rect 11848 11784 12265 11812
rect 11848 11772 11854 11784
rect 12253 11781 12265 11784
rect 12299 11781 12311 11815
rect 12253 11775 12311 11781
rect 12342 11772 12348 11824
rect 12400 11812 12406 11824
rect 14458 11812 14464 11824
rect 12400 11784 14464 11812
rect 12400 11772 12406 11784
rect 14458 11772 14464 11784
rect 14516 11772 14522 11824
rect 17494 11812 17500 11824
rect 14568 11784 17500 11812
rect 12066 11744 12072 11756
rect 10336 11716 12072 11744
rect 9309 11707 9367 11713
rect 12066 11704 12072 11716
rect 12124 11704 12130 11756
rect 13449 11747 13507 11753
rect 13449 11713 13461 11747
rect 13495 11744 13507 11747
rect 14568 11744 14596 11784
rect 17494 11772 17500 11784
rect 17552 11772 17558 11824
rect 18064 11812 18092 11843
rect 18414 11840 18420 11892
rect 18472 11840 18478 11892
rect 25774 11880 25780 11892
rect 21376 11852 25780 11880
rect 19426 11812 19432 11824
rect 18064 11784 19432 11812
rect 19426 11772 19432 11784
rect 19484 11772 19490 11824
rect 19978 11772 19984 11824
rect 20036 11812 20042 11824
rect 21376 11821 21404 11852
rect 25774 11840 25780 11852
rect 25832 11840 25838 11892
rect 20073 11815 20131 11821
rect 20073 11812 20085 11815
rect 20036 11784 20085 11812
rect 20036 11772 20042 11784
rect 20073 11781 20085 11784
rect 20119 11812 20131 11815
rect 21361 11815 21419 11821
rect 21361 11812 21373 11815
rect 20119 11784 21373 11812
rect 20119 11781 20131 11784
rect 20073 11775 20131 11781
rect 21361 11781 21373 11784
rect 21407 11781 21419 11815
rect 21361 11775 21419 11781
rect 23293 11815 23351 11821
rect 23293 11781 23305 11815
rect 23339 11812 23351 11815
rect 24854 11812 24860 11824
rect 23339 11784 24860 11812
rect 23339 11781 23351 11784
rect 23293 11775 23351 11781
rect 24854 11772 24860 11784
rect 24912 11772 24918 11824
rect 13495 11716 14596 11744
rect 13495 11713 13507 11716
rect 13449 11707 13507 11713
rect 14642 11704 14648 11756
rect 14700 11704 14706 11756
rect 16114 11704 16120 11756
rect 16172 11744 16178 11756
rect 17221 11747 17279 11753
rect 17221 11744 17233 11747
rect 16172 11716 17233 11744
rect 16172 11704 16178 11716
rect 17221 11713 17233 11716
rect 17267 11713 17279 11747
rect 17221 11707 17279 11713
rect 19334 11704 19340 11756
rect 19392 11744 19398 11756
rect 21177 11747 21235 11753
rect 21177 11744 21189 11747
rect 19392 11716 21189 11744
rect 19392 11704 19398 11716
rect 21177 11713 21189 11716
rect 21223 11744 21235 11747
rect 22281 11747 22339 11753
rect 21223 11716 22094 11744
rect 21223 11713 21235 11716
rect 21177 11707 21235 11713
rect 7285 11679 7343 11685
rect 7285 11645 7297 11679
rect 7331 11645 7343 11679
rect 7285 11639 7343 11645
rect 7561 11679 7619 11685
rect 7561 11645 7573 11679
rect 7607 11676 7619 11679
rect 10413 11679 10471 11685
rect 10413 11676 10425 11679
rect 7607 11648 10425 11676
rect 7607 11645 7619 11648
rect 7561 11639 7619 11645
rect 10413 11645 10425 11648
rect 10459 11676 10471 11679
rect 11054 11676 11060 11688
rect 10459 11648 11060 11676
rect 10459 11645 10471 11648
rect 10413 11639 10471 11645
rect 7300 11540 7328 11639
rect 11054 11636 11060 11648
rect 11112 11636 11118 11688
rect 12345 11679 12403 11685
rect 12345 11645 12357 11679
rect 12391 11645 12403 11679
rect 12345 11639 12403 11645
rect 12437 11679 12495 11685
rect 12437 11645 12449 11679
rect 12483 11645 12495 11679
rect 12437 11639 12495 11645
rect 13541 11679 13599 11685
rect 13541 11645 13553 11679
rect 13587 11645 13599 11679
rect 13541 11639 13599 11645
rect 10502 11568 10508 11620
rect 10560 11608 10566 11620
rect 11882 11608 11888 11620
rect 10560 11580 11888 11608
rect 10560 11568 10566 11580
rect 11882 11568 11888 11580
rect 11940 11608 11946 11620
rect 12360 11608 12388 11639
rect 11940 11580 12388 11608
rect 11940 11568 11946 11580
rect 8294 11540 8300 11552
rect 7300 11512 8300 11540
rect 8294 11500 8300 11512
rect 8352 11500 8358 11552
rect 11606 11500 11612 11552
rect 11664 11540 11670 11552
rect 12342 11540 12348 11552
rect 11664 11512 12348 11540
rect 11664 11500 11670 11512
rect 12342 11500 12348 11512
rect 12400 11540 12406 11552
rect 12452 11540 12480 11639
rect 13446 11568 13452 11620
rect 13504 11608 13510 11620
rect 13556 11608 13584 11639
rect 13630 11636 13636 11688
rect 13688 11676 13694 11688
rect 13725 11679 13783 11685
rect 13725 11676 13737 11679
rect 13688 11648 13737 11676
rect 13688 11636 13694 11648
rect 13725 11645 13737 11648
rect 13771 11645 13783 11679
rect 13725 11639 13783 11645
rect 13504 11580 13584 11608
rect 13740 11608 13768 11639
rect 14366 11636 14372 11688
rect 14424 11676 14430 11688
rect 14737 11679 14795 11685
rect 14737 11676 14749 11679
rect 14424 11648 14749 11676
rect 14424 11636 14430 11648
rect 14737 11645 14749 11648
rect 14783 11645 14795 11679
rect 14737 11639 14795 11645
rect 14921 11679 14979 11685
rect 14921 11645 14933 11679
rect 14967 11676 14979 11679
rect 15102 11676 15108 11688
rect 14967 11648 15108 11676
rect 14967 11645 14979 11648
rect 14921 11639 14979 11645
rect 14936 11608 14964 11639
rect 15102 11636 15108 11648
rect 15160 11636 15166 11688
rect 16666 11636 16672 11688
rect 16724 11676 16730 11688
rect 17405 11679 17463 11685
rect 17405 11676 17417 11679
rect 16724 11648 17417 11676
rect 16724 11636 16730 11648
rect 17405 11645 17417 11648
rect 17451 11645 17463 11679
rect 17405 11639 17463 11645
rect 18230 11636 18236 11688
rect 18288 11676 18294 11688
rect 18509 11679 18567 11685
rect 18509 11676 18521 11679
rect 18288 11648 18521 11676
rect 18288 11636 18294 11648
rect 18509 11645 18521 11648
rect 18555 11645 18567 11679
rect 18509 11639 18567 11645
rect 18693 11679 18751 11685
rect 18693 11645 18705 11679
rect 18739 11676 18751 11679
rect 19702 11676 19708 11688
rect 18739 11648 19708 11676
rect 18739 11645 18751 11648
rect 18693 11639 18751 11645
rect 19702 11636 19708 11648
rect 19760 11636 19766 11688
rect 19978 11636 19984 11688
rect 20036 11676 20042 11688
rect 20717 11679 20775 11685
rect 20717 11676 20729 11679
rect 20036 11648 20729 11676
rect 20036 11636 20042 11648
rect 20717 11645 20729 11648
rect 20763 11645 20775 11679
rect 20717 11639 20775 11645
rect 13740 11580 14964 11608
rect 13504 11568 13510 11580
rect 15470 11568 15476 11620
rect 15528 11608 15534 11620
rect 16482 11608 16488 11620
rect 15528 11580 16488 11608
rect 15528 11568 15534 11580
rect 16482 11568 16488 11580
rect 16540 11608 16546 11620
rect 16758 11608 16764 11620
rect 16540 11580 16764 11608
rect 16540 11568 16546 11580
rect 16758 11568 16764 11580
rect 16816 11568 16822 11620
rect 16853 11611 16911 11617
rect 16853 11577 16865 11611
rect 16899 11608 16911 11611
rect 21726 11608 21732 11620
rect 16899 11580 21732 11608
rect 16899 11577 16911 11580
rect 16853 11571 16911 11577
rect 21726 11568 21732 11580
rect 21784 11568 21790 11620
rect 22066 11608 22094 11716
rect 22281 11713 22293 11747
rect 22327 11744 22339 11747
rect 23934 11744 23940 11756
rect 22327 11716 23940 11744
rect 22327 11713 22339 11716
rect 22281 11707 22339 11713
rect 23934 11704 23940 11716
rect 23992 11704 23998 11756
rect 24121 11747 24179 11753
rect 24121 11713 24133 11747
rect 24167 11744 24179 11747
rect 24946 11744 24952 11756
rect 24167 11716 24952 11744
rect 24167 11713 24179 11716
rect 24121 11707 24179 11713
rect 24946 11704 24952 11716
rect 25004 11704 25010 11756
rect 24762 11636 24768 11688
rect 24820 11636 24826 11688
rect 26142 11608 26148 11620
rect 22066 11580 26148 11608
rect 26142 11568 26148 11580
rect 26200 11568 26206 11620
rect 12400 11512 12480 11540
rect 12400 11500 12406 11512
rect 14826 11500 14832 11552
rect 14884 11540 14890 11552
rect 15010 11540 15016 11552
rect 14884 11512 15016 11540
rect 14884 11500 14890 11512
rect 15010 11500 15016 11512
rect 15068 11500 15074 11552
rect 15378 11500 15384 11552
rect 15436 11540 15442 11552
rect 17678 11540 17684 11552
rect 15436 11512 17684 11540
rect 15436 11500 15442 11512
rect 17678 11500 17684 11512
rect 17736 11500 17742 11552
rect 19429 11543 19487 11549
rect 19429 11509 19441 11543
rect 19475 11540 19487 11543
rect 19702 11540 19708 11552
rect 19475 11512 19708 11540
rect 19475 11509 19487 11512
rect 19429 11503 19487 11509
rect 19702 11500 19708 11512
rect 19760 11500 19766 11552
rect 20165 11543 20223 11549
rect 20165 11509 20177 11543
rect 20211 11540 20223 11543
rect 20714 11540 20720 11552
rect 20211 11512 20720 11540
rect 20211 11509 20223 11512
rect 20165 11503 20223 11509
rect 20714 11500 20720 11512
rect 20772 11500 20778 11552
rect 23750 11500 23756 11552
rect 23808 11540 23814 11552
rect 24118 11540 24124 11552
rect 23808 11512 24124 11540
rect 23808 11500 23814 11512
rect 24118 11500 24124 11512
rect 24176 11500 24182 11552
rect 1104 11450 25852 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 25852 11450
rect 1104 11376 25852 11398
rect 7190 11296 7196 11348
rect 7248 11336 7254 11348
rect 10502 11336 10508 11348
rect 7248 11308 10508 11336
rect 7248 11296 7254 11308
rect 10502 11296 10508 11308
rect 10560 11296 10566 11348
rect 10594 11296 10600 11348
rect 10652 11336 10658 11348
rect 12621 11339 12679 11345
rect 12621 11336 12633 11339
rect 10652 11308 12633 11336
rect 10652 11296 10658 11308
rect 12621 11305 12633 11308
rect 12667 11305 12679 11339
rect 12621 11299 12679 11305
rect 13262 11296 13268 11348
rect 13320 11336 13326 11348
rect 13446 11336 13452 11348
rect 13320 11308 13452 11336
rect 13320 11296 13326 11308
rect 13446 11296 13452 11308
rect 13504 11296 13510 11348
rect 15194 11336 15200 11348
rect 14108 11308 15200 11336
rect 11425 11271 11483 11277
rect 11425 11237 11437 11271
rect 11471 11268 11483 11271
rect 12802 11268 12808 11280
rect 11471 11240 12808 11268
rect 11471 11237 11483 11240
rect 11425 11231 11483 11237
rect 12802 11228 12808 11240
rect 12860 11228 12866 11280
rect 13170 11228 13176 11280
rect 13228 11268 13234 11280
rect 13633 11271 13691 11277
rect 13633 11268 13645 11271
rect 13228 11240 13645 11268
rect 13228 11228 13234 11240
rect 13633 11237 13645 11240
rect 13679 11268 13691 11271
rect 13814 11268 13820 11280
rect 13679 11240 13820 11268
rect 13679 11237 13691 11240
rect 13633 11231 13691 11237
rect 13814 11228 13820 11240
rect 13872 11228 13878 11280
rect 9401 11203 9459 11209
rect 9401 11169 9413 11203
rect 9447 11200 9459 11203
rect 9447 11172 11836 11200
rect 9447 11169 9459 11172
rect 9401 11163 9459 11169
rect 9122 11092 9128 11144
rect 9180 11092 9186 11144
rect 11808 11132 11836 11172
rect 11882 11160 11888 11212
rect 11940 11160 11946 11212
rect 11977 11203 12035 11209
rect 11977 11169 11989 11203
rect 12023 11200 12035 11203
rect 12250 11200 12256 11212
rect 12023 11172 12256 11200
rect 12023 11169 12035 11172
rect 11977 11163 12035 11169
rect 11992 11132 12020 11163
rect 12250 11160 12256 11172
rect 12308 11160 12314 11212
rect 13265 11203 13323 11209
rect 13265 11200 13277 11203
rect 12820 11172 13277 11200
rect 11808 11104 12020 11132
rect 12066 11092 12072 11144
rect 12124 11132 12130 11144
rect 12710 11132 12716 11144
rect 12124 11104 12716 11132
rect 12124 11092 12130 11104
rect 12710 11092 12716 11104
rect 12768 11092 12774 11144
rect 8662 11024 8668 11076
rect 8720 11064 8726 11076
rect 9858 11064 9864 11076
rect 8720 11036 9864 11064
rect 8720 11024 8726 11036
rect 9858 11024 9864 11036
rect 9916 11024 9922 11076
rect 11054 11024 11060 11076
rect 11112 11064 11118 11076
rect 12820 11064 12848 11172
rect 13265 11169 13277 11172
rect 13311 11200 13323 11203
rect 13538 11200 13544 11212
rect 13311 11172 13544 11200
rect 13311 11169 13323 11172
rect 13265 11163 13323 11169
rect 13538 11160 13544 11172
rect 13596 11160 13602 11212
rect 12989 11135 13047 11141
rect 12989 11101 13001 11135
rect 13035 11132 13047 11135
rect 14108 11132 14136 11308
rect 15194 11296 15200 11308
rect 15252 11296 15258 11348
rect 16298 11296 16304 11348
rect 16356 11336 16362 11348
rect 19426 11336 19432 11348
rect 16356 11308 19432 11336
rect 16356 11296 16362 11308
rect 19426 11296 19432 11308
rect 19484 11296 19490 11348
rect 19613 11339 19671 11345
rect 19613 11305 19625 11339
rect 19659 11336 19671 11339
rect 21634 11336 21640 11348
rect 19659 11308 21640 11336
rect 19659 11305 19671 11308
rect 19613 11299 19671 11305
rect 21634 11296 21640 11308
rect 21692 11296 21698 11348
rect 22830 11296 22836 11348
rect 22888 11336 22894 11348
rect 25041 11339 25099 11345
rect 25041 11336 25053 11339
rect 22888 11308 25053 11336
rect 22888 11296 22894 11308
rect 25041 11305 25053 11308
rect 25087 11305 25099 11339
rect 25041 11299 25099 11305
rect 14458 11228 14464 11280
rect 14516 11268 14522 11280
rect 14826 11268 14832 11280
rect 14516 11240 14832 11268
rect 14516 11228 14522 11240
rect 14826 11228 14832 11240
rect 14884 11228 14890 11280
rect 16666 11228 16672 11280
rect 16724 11228 16730 11280
rect 16758 11228 16764 11280
rect 16816 11268 16822 11280
rect 17037 11271 17095 11277
rect 17037 11268 17049 11271
rect 16816 11240 17049 11268
rect 16816 11228 16822 11240
rect 17037 11237 17049 11240
rect 17083 11237 17095 11271
rect 17037 11231 17095 11237
rect 18141 11271 18199 11277
rect 18141 11237 18153 11271
rect 18187 11268 18199 11271
rect 21358 11268 21364 11280
rect 18187 11240 21364 11268
rect 18187 11237 18199 11240
rect 18141 11231 18199 11237
rect 21358 11228 21364 11240
rect 21416 11228 21422 11280
rect 21545 11271 21603 11277
rect 21545 11237 21557 11271
rect 21591 11268 21603 11271
rect 23750 11268 23756 11280
rect 21591 11240 23756 11268
rect 21591 11237 21603 11240
rect 21545 11231 21603 11237
rect 23750 11228 23756 11240
rect 23808 11228 23814 11280
rect 14366 11160 14372 11212
rect 14424 11200 14430 11212
rect 14734 11200 14740 11212
rect 14424 11172 14740 11200
rect 14424 11160 14430 11172
rect 14734 11160 14740 11172
rect 14792 11160 14798 11212
rect 14921 11203 14979 11209
rect 14921 11169 14933 11203
rect 14967 11200 14979 11203
rect 16942 11200 16948 11212
rect 14967 11172 16948 11200
rect 14967 11169 14979 11172
rect 14921 11163 14979 11169
rect 16942 11160 16948 11172
rect 17000 11160 17006 11212
rect 17310 11160 17316 11212
rect 17368 11200 17374 11212
rect 17494 11200 17500 11212
rect 17368 11172 17500 11200
rect 17368 11160 17374 11172
rect 17494 11160 17500 11172
rect 17552 11160 17558 11212
rect 17954 11160 17960 11212
rect 18012 11200 18018 11212
rect 18601 11203 18659 11209
rect 18601 11200 18613 11203
rect 18012 11172 18613 11200
rect 18012 11160 18018 11172
rect 18601 11169 18613 11172
rect 18647 11169 18659 11203
rect 18601 11163 18659 11169
rect 18785 11203 18843 11209
rect 18785 11169 18797 11203
rect 18831 11200 18843 11203
rect 20257 11203 20315 11209
rect 18831 11172 20208 11200
rect 18831 11169 18843 11172
rect 18785 11163 18843 11169
rect 13035 11104 14136 11132
rect 13035 11101 13047 11104
rect 12989 11095 13047 11101
rect 14182 11092 14188 11144
rect 14240 11132 14246 11144
rect 14550 11132 14556 11144
rect 14240 11104 14556 11132
rect 14240 11092 14246 11104
rect 14550 11092 14556 11104
rect 14608 11092 14614 11144
rect 18616 11132 18644 11163
rect 19245 11135 19303 11141
rect 19245 11132 19257 11135
rect 18616 11104 19257 11132
rect 19245 11101 19257 11104
rect 19291 11101 19303 11135
rect 19245 11095 19303 11101
rect 19978 11092 19984 11144
rect 20036 11092 20042 11144
rect 20180 11132 20208 11172
rect 20257 11169 20269 11203
rect 20303 11200 20315 11203
rect 22462 11200 22468 11212
rect 20303 11172 22468 11200
rect 20303 11169 20315 11172
rect 20257 11163 20315 11169
rect 22462 11160 22468 11172
rect 22520 11160 22526 11212
rect 26694 11200 26700 11212
rect 23584 11172 26700 11200
rect 20806 11132 20812 11144
rect 20180 11104 20812 11132
rect 20806 11092 20812 11104
rect 20864 11092 20870 11144
rect 20901 11135 20959 11141
rect 20901 11101 20913 11135
rect 20947 11132 20959 11135
rect 21082 11132 21088 11144
rect 20947 11104 21088 11132
rect 20947 11101 20959 11104
rect 20901 11095 20959 11101
rect 21082 11092 21088 11104
rect 21140 11092 21146 11144
rect 21726 11092 21732 11144
rect 21784 11092 21790 11144
rect 22833 11135 22891 11141
rect 22833 11101 22845 11135
rect 22879 11132 22891 11135
rect 23474 11132 23480 11144
rect 22879 11104 23480 11132
rect 22879 11101 22891 11104
rect 22833 11095 22891 11101
rect 23474 11092 23480 11104
rect 23532 11092 23538 11144
rect 11112 11036 12848 11064
rect 13081 11067 13139 11073
rect 11112 11024 11118 11036
rect 13081 11033 13093 11067
rect 13127 11064 13139 11067
rect 15102 11064 15108 11076
rect 13127 11036 15108 11064
rect 13127 11033 13139 11036
rect 13081 11027 13139 11033
rect 15102 11024 15108 11036
rect 15160 11024 15166 11076
rect 15194 11024 15200 11076
rect 15252 11024 15258 11076
rect 15470 11064 15476 11076
rect 15304 11036 15476 11064
rect 9674 10956 9680 11008
rect 9732 10996 9738 11008
rect 10870 10996 10876 11008
rect 9732 10968 10876 10996
rect 9732 10956 9738 10968
rect 10870 10956 10876 10968
rect 10928 10956 10934 11008
rect 11793 10999 11851 11005
rect 11793 10965 11805 10999
rect 11839 10996 11851 10999
rect 11882 10996 11888 11008
rect 11839 10968 11888 10996
rect 11839 10965 11851 10968
rect 11793 10959 11851 10965
rect 11882 10956 11888 10968
rect 11940 10996 11946 11008
rect 12066 10996 12072 11008
rect 11940 10968 12072 10996
rect 11940 10956 11946 10968
rect 12066 10956 12072 10968
rect 12124 10956 12130 11008
rect 12434 10956 12440 11008
rect 12492 10996 12498 11008
rect 13446 10996 13452 11008
rect 12492 10968 13452 10996
rect 12492 10956 12498 10968
rect 13446 10956 13452 10968
rect 13504 10956 13510 11008
rect 14274 10956 14280 11008
rect 14332 10956 14338 11008
rect 14826 10956 14832 11008
rect 14884 10996 14890 11008
rect 15304 10996 15332 11036
rect 15470 11024 15476 11036
rect 15528 11064 15534 11076
rect 15528 11036 15686 11064
rect 16868 11036 17080 11064
rect 15528 11024 15534 11036
rect 14884 10968 15332 10996
rect 14884 10956 14890 10968
rect 15378 10956 15384 11008
rect 15436 10996 15442 11008
rect 16868 10996 16896 11036
rect 15436 10968 16896 10996
rect 17052 10996 17080 11036
rect 17678 11024 17684 11076
rect 17736 11064 17742 11076
rect 17736 11036 18460 11064
rect 17736 11024 17742 11036
rect 18230 10996 18236 11008
rect 17052 10968 18236 10996
rect 15436 10956 15442 10968
rect 18230 10956 18236 10968
rect 18288 10956 18294 11008
rect 18432 10996 18460 11036
rect 18506 11024 18512 11076
rect 18564 11024 18570 11076
rect 18616 11036 19564 11064
rect 18616 10996 18644 11036
rect 18432 10968 18644 10996
rect 19536 10996 19564 11036
rect 19610 11024 19616 11076
rect 19668 11064 19674 11076
rect 21100 11064 21128 11092
rect 23584 11064 23612 11172
rect 26694 11160 26700 11172
rect 26752 11160 26758 11212
rect 25222 11092 25228 11144
rect 25280 11092 25286 11144
rect 19668 11036 21036 11064
rect 21100 11036 23612 11064
rect 19668 11024 19674 11036
rect 21008 11005 21036 11036
rect 22112 11005 22140 11036
rect 23842 11024 23848 11076
rect 23900 11024 23906 11076
rect 20073 10999 20131 11005
rect 20073 10996 20085 10999
rect 19536 10968 20085 10996
rect 20073 10965 20085 10968
rect 20119 10965 20131 10999
rect 20073 10959 20131 10965
rect 20993 10999 21051 11005
rect 20993 10965 21005 10999
rect 21039 10965 21051 10999
rect 20993 10959 21051 10965
rect 22097 10999 22155 11005
rect 22097 10965 22109 10999
rect 22143 10996 22155 10999
rect 22143 10968 22177 10996
rect 22143 10965 22155 10968
rect 22097 10959 22155 10965
rect 1104 10906 25852 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 25852 10906
rect 1104 10832 25852 10854
rect 8662 10752 8668 10804
rect 8720 10752 8726 10804
rect 9950 10752 9956 10804
rect 10008 10752 10014 10804
rect 12713 10795 12771 10801
rect 12713 10761 12725 10795
rect 12759 10792 12771 10795
rect 14274 10792 14280 10804
rect 12759 10764 14280 10792
rect 12759 10761 12771 10764
rect 12713 10755 12771 10761
rect 14274 10752 14280 10764
rect 14332 10752 14338 10804
rect 14366 10752 14372 10804
rect 14424 10792 14430 10804
rect 20622 10792 20628 10804
rect 14424 10764 17080 10792
rect 14424 10752 14430 10764
rect 7098 10684 7104 10736
rect 7156 10724 7162 10736
rect 8481 10727 8539 10733
rect 8481 10724 8493 10727
rect 7156 10696 8493 10724
rect 7156 10684 7162 10696
rect 8481 10693 8493 10696
rect 8527 10693 8539 10727
rect 8680 10724 8708 10752
rect 8680 10696 8970 10724
rect 8481 10687 8539 10693
rect 9858 10684 9864 10736
rect 9916 10724 9922 10736
rect 10321 10727 10379 10733
rect 10321 10724 10333 10727
rect 9916 10696 10333 10724
rect 9916 10684 9922 10696
rect 10321 10693 10333 10696
rect 10367 10724 10379 10727
rect 10965 10727 11023 10733
rect 10965 10724 10977 10727
rect 10367 10696 10977 10724
rect 10367 10693 10379 10696
rect 10321 10687 10379 10693
rect 10965 10693 10977 10696
rect 11011 10693 11023 10727
rect 10965 10687 11023 10693
rect 12342 10684 12348 10736
rect 12400 10724 12406 10736
rect 12400 10696 12756 10724
rect 12400 10684 12406 10696
rect 10870 10616 10876 10668
rect 10928 10656 10934 10668
rect 12728 10656 12756 10696
rect 12802 10684 12808 10736
rect 12860 10684 12866 10736
rect 15286 10724 15292 10736
rect 12912 10696 15292 10724
rect 12912 10656 12940 10696
rect 15286 10684 15292 10696
rect 15344 10724 15350 10736
rect 15344 10696 16252 10724
rect 15344 10684 15350 10696
rect 10928 10628 12664 10656
rect 12728 10628 12940 10656
rect 10928 10616 10934 10628
rect 8205 10591 8263 10597
rect 8205 10557 8217 10591
rect 8251 10557 8263 10591
rect 8205 10551 8263 10557
rect 11701 10591 11759 10597
rect 11701 10557 11713 10591
rect 11747 10588 11759 10591
rect 12066 10588 12072 10600
rect 11747 10560 12072 10588
rect 11747 10557 11759 10560
rect 11701 10551 11759 10557
rect 8220 10452 8248 10551
rect 12066 10548 12072 10560
rect 12124 10548 12130 10600
rect 12636 10520 12664 10628
rect 13354 10616 13360 10668
rect 13412 10616 13418 10668
rect 14182 10616 14188 10668
rect 14240 10616 14246 10668
rect 14274 10616 14280 10668
rect 14332 10616 14338 10668
rect 15933 10659 15991 10665
rect 15933 10625 15945 10659
rect 15979 10625 15991 10659
rect 15933 10619 15991 10625
rect 12897 10591 12955 10597
rect 12897 10557 12909 10591
rect 12943 10557 12955 10591
rect 12897 10551 12955 10557
rect 12912 10520 12940 10551
rect 12636 10492 12940 10520
rect 13372 10520 13400 10616
rect 14461 10591 14519 10597
rect 14461 10557 14473 10591
rect 14507 10588 14519 10591
rect 15286 10588 15292 10600
rect 14507 10560 15292 10588
rect 14507 10557 14519 10560
rect 14461 10551 14519 10557
rect 15286 10548 15292 10560
rect 15344 10548 15350 10600
rect 13817 10523 13875 10529
rect 13817 10520 13829 10523
rect 13372 10492 13829 10520
rect 13817 10489 13829 10492
rect 13863 10489 13875 10523
rect 13817 10483 13875 10489
rect 13998 10480 14004 10532
rect 14056 10520 14062 10532
rect 15565 10523 15623 10529
rect 15565 10520 15577 10523
rect 14056 10492 15577 10520
rect 14056 10480 14062 10492
rect 15565 10489 15577 10492
rect 15611 10489 15623 10523
rect 15948 10520 15976 10619
rect 16022 10548 16028 10600
rect 16080 10548 16086 10600
rect 16224 10597 16252 10696
rect 17052 10665 17080 10764
rect 18156 10764 20628 10792
rect 17586 10684 17592 10736
rect 17644 10684 17650 10736
rect 17037 10659 17095 10665
rect 17037 10625 17049 10659
rect 17083 10625 17095 10659
rect 17037 10619 17095 10625
rect 16209 10591 16267 10597
rect 16209 10557 16221 10591
rect 16255 10588 16267 10591
rect 16482 10588 16488 10600
rect 16255 10560 16488 10588
rect 16255 10557 16267 10560
rect 16209 10551 16267 10557
rect 16482 10548 16488 10560
rect 16540 10548 16546 10600
rect 18156 10520 18184 10764
rect 20622 10752 20628 10764
rect 20680 10752 20686 10804
rect 20717 10795 20775 10801
rect 20717 10761 20729 10795
rect 20763 10761 20775 10795
rect 23566 10792 23572 10804
rect 20717 10755 20775 10761
rect 22204 10764 23572 10792
rect 20732 10724 20760 10755
rect 19076 10696 20760 10724
rect 21177 10727 21235 10733
rect 18414 10616 18420 10668
rect 18472 10616 18478 10668
rect 19076 10665 19104 10696
rect 21177 10693 21189 10727
rect 21223 10724 21235 10727
rect 21358 10724 21364 10736
rect 21223 10696 21364 10724
rect 21223 10693 21235 10696
rect 21177 10687 21235 10693
rect 21358 10684 21364 10696
rect 21416 10684 21422 10736
rect 19061 10659 19119 10665
rect 19061 10625 19073 10659
rect 19107 10625 19119 10659
rect 19061 10619 19119 10625
rect 19242 10616 19248 10668
rect 19300 10656 19306 10668
rect 19889 10659 19947 10665
rect 19889 10656 19901 10659
rect 19300 10628 19901 10656
rect 19300 10616 19306 10628
rect 19889 10625 19901 10628
rect 19935 10625 19947 10659
rect 19889 10619 19947 10625
rect 21082 10616 21088 10668
rect 21140 10616 21146 10668
rect 22204 10665 22232 10764
rect 23566 10752 23572 10764
rect 23624 10752 23630 10804
rect 23382 10684 23388 10736
rect 23440 10684 23446 10736
rect 22189 10659 22247 10665
rect 22189 10625 22201 10659
rect 22235 10625 22247 10659
rect 22189 10619 22247 10625
rect 22646 10616 22652 10668
rect 22704 10656 22710 10668
rect 23109 10659 23167 10665
rect 23109 10656 23121 10659
rect 22704 10628 23121 10656
rect 22704 10616 22710 10628
rect 23109 10625 23121 10628
rect 23155 10625 23167 10659
rect 23109 10619 23167 10625
rect 19426 10548 19432 10600
rect 19484 10588 19490 10600
rect 19978 10588 19984 10600
rect 19484 10560 19984 10588
rect 19484 10548 19490 10560
rect 19978 10548 19984 10560
rect 20036 10548 20042 10600
rect 20162 10548 20168 10600
rect 20220 10548 20226 10600
rect 21266 10548 21272 10600
rect 21324 10548 21330 10600
rect 21910 10548 21916 10600
rect 21968 10588 21974 10600
rect 22557 10591 22615 10597
rect 22557 10588 22569 10591
rect 21968 10560 22569 10588
rect 21968 10548 21974 10560
rect 22557 10557 22569 10560
rect 22603 10588 22615 10591
rect 24394 10588 24400 10600
rect 22603 10560 24400 10588
rect 22603 10557 22615 10560
rect 22557 10551 22615 10557
rect 24394 10548 24400 10560
rect 24452 10588 24458 10600
rect 24504 10588 24532 10642
rect 25133 10591 25191 10597
rect 25133 10588 25145 10591
rect 24452 10560 25145 10588
rect 24452 10548 24458 10560
rect 25133 10557 25145 10560
rect 25179 10557 25191 10591
rect 25133 10551 25191 10557
rect 15948 10492 18184 10520
rect 18233 10523 18291 10529
rect 15565 10483 15623 10489
rect 18233 10489 18245 10523
rect 18279 10520 18291 10523
rect 20346 10520 20352 10532
rect 18279 10492 20352 10520
rect 18279 10489 18291 10492
rect 18233 10483 18291 10489
rect 20346 10480 20352 10492
rect 20404 10480 20410 10532
rect 8294 10452 8300 10464
rect 8220 10424 8300 10452
rect 8294 10412 8300 10424
rect 8352 10452 8358 10464
rect 9122 10452 9128 10464
rect 8352 10424 9128 10452
rect 8352 10412 8358 10424
rect 9122 10412 9128 10424
rect 9180 10452 9186 10464
rect 9582 10452 9588 10464
rect 9180 10424 9588 10452
rect 9180 10412 9186 10424
rect 9582 10412 9588 10424
rect 9640 10412 9646 10464
rect 12345 10455 12403 10461
rect 12345 10421 12357 10455
rect 12391 10452 12403 10455
rect 15654 10452 15660 10464
rect 12391 10424 15660 10452
rect 12391 10421 12403 10424
rect 12345 10415 12403 10421
rect 15654 10412 15660 10424
rect 15712 10412 15718 10464
rect 16850 10412 16856 10464
rect 16908 10412 16914 10464
rect 17034 10412 17040 10464
rect 17092 10452 17098 10464
rect 17681 10455 17739 10461
rect 17681 10452 17693 10455
rect 17092 10424 17693 10452
rect 17092 10412 17098 10424
rect 17681 10421 17693 10424
rect 17727 10421 17739 10455
rect 17681 10415 17739 10421
rect 18874 10412 18880 10464
rect 18932 10412 18938 10464
rect 19521 10455 19579 10461
rect 19521 10421 19533 10455
rect 19567 10452 19579 10455
rect 21358 10452 21364 10464
rect 19567 10424 21364 10452
rect 19567 10421 19579 10424
rect 19521 10415 19579 10421
rect 21358 10412 21364 10424
rect 21416 10412 21422 10464
rect 21818 10412 21824 10464
rect 21876 10452 21882 10464
rect 22005 10455 22063 10461
rect 22005 10452 22017 10455
rect 21876 10424 22017 10452
rect 21876 10412 21882 10424
rect 22005 10421 22017 10424
rect 22051 10421 22063 10455
rect 22005 10415 22063 10421
rect 23382 10412 23388 10464
rect 23440 10452 23446 10464
rect 24857 10455 24915 10461
rect 24857 10452 24869 10455
rect 23440 10424 24869 10452
rect 23440 10412 23446 10424
rect 24857 10421 24869 10424
rect 24903 10421 24915 10455
rect 24857 10415 24915 10421
rect 1104 10362 25852 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 25852 10362
rect 1104 10288 25852 10310
rect 11054 10208 11060 10260
rect 11112 10208 11118 10260
rect 11514 10208 11520 10260
rect 11572 10248 11578 10260
rect 11609 10251 11667 10257
rect 11609 10248 11621 10251
rect 11572 10220 11621 10248
rect 11572 10208 11578 10220
rect 11609 10217 11621 10220
rect 11655 10217 11667 10251
rect 11609 10211 11667 10217
rect 11974 10208 11980 10260
rect 12032 10248 12038 10260
rect 12805 10251 12863 10257
rect 12805 10248 12817 10251
rect 12032 10220 12817 10248
rect 12032 10208 12038 10220
rect 12805 10217 12817 10220
rect 12851 10217 12863 10251
rect 12805 10211 12863 10217
rect 14550 10208 14556 10260
rect 14608 10208 14614 10260
rect 14734 10208 14740 10260
rect 14792 10248 14798 10260
rect 14792 10220 16804 10248
rect 14792 10208 14798 10220
rect 12710 10140 12716 10192
rect 12768 10180 12774 10192
rect 13722 10180 13728 10192
rect 12768 10152 13728 10180
rect 12768 10140 12774 10152
rect 13722 10140 13728 10152
rect 13780 10140 13786 10192
rect 16022 10140 16028 10192
rect 16080 10180 16086 10192
rect 16298 10180 16304 10192
rect 16080 10152 16304 10180
rect 16080 10140 16086 10152
rect 16298 10140 16304 10152
rect 16356 10140 16362 10192
rect 9309 10115 9367 10121
rect 9309 10081 9321 10115
rect 9355 10112 9367 10115
rect 9582 10112 9588 10124
rect 9355 10084 9588 10112
rect 9355 10081 9367 10084
rect 9309 10075 9367 10081
rect 9582 10072 9588 10084
rect 9640 10072 9646 10124
rect 12158 10072 12164 10124
rect 12216 10072 12222 10124
rect 13449 10115 13507 10121
rect 13449 10081 13461 10115
rect 13495 10112 13507 10115
rect 13538 10112 13544 10124
rect 13495 10084 13544 10112
rect 13495 10081 13507 10084
rect 13449 10075 13507 10081
rect 13538 10072 13544 10084
rect 13596 10072 13602 10124
rect 14918 10072 14924 10124
rect 14976 10112 14982 10124
rect 15105 10115 15163 10121
rect 15105 10112 15117 10115
rect 14976 10084 15117 10112
rect 14976 10072 14982 10084
rect 15105 10081 15117 10084
rect 15151 10081 15163 10115
rect 16776 10112 16804 10220
rect 16850 10208 16856 10260
rect 16908 10248 16914 10260
rect 20990 10248 20996 10260
rect 16908 10220 20996 10248
rect 16908 10208 16914 10220
rect 20990 10208 20996 10220
rect 21048 10208 21054 10260
rect 24578 10208 24584 10260
rect 24636 10208 24642 10260
rect 17957 10183 18015 10189
rect 17957 10149 17969 10183
rect 18003 10180 18015 10183
rect 18322 10180 18328 10192
rect 18003 10152 18328 10180
rect 18003 10149 18015 10152
rect 17957 10143 18015 10149
rect 18322 10140 18328 10152
rect 18380 10140 18386 10192
rect 19794 10180 19800 10192
rect 18432 10152 19800 10180
rect 17678 10112 17684 10124
rect 16776 10084 17684 10112
rect 15105 10075 15163 10081
rect 17678 10072 17684 10084
rect 17736 10072 17742 10124
rect 17770 10072 17776 10124
rect 17828 10112 17834 10124
rect 18432 10112 18460 10152
rect 19794 10140 19800 10152
rect 19852 10140 19858 10192
rect 19978 10140 19984 10192
rect 20036 10180 20042 10192
rect 20165 10183 20223 10189
rect 20165 10180 20177 10183
rect 20036 10152 20177 10180
rect 20036 10140 20042 10152
rect 20165 10149 20177 10152
rect 20211 10149 20223 10183
rect 20165 10143 20223 10149
rect 22278 10140 22284 10192
rect 22336 10140 22342 10192
rect 17828 10084 18460 10112
rect 18601 10115 18659 10121
rect 17828 10072 17834 10084
rect 18601 10081 18613 10115
rect 18647 10112 18659 10115
rect 18874 10112 18880 10124
rect 18647 10084 18880 10112
rect 18647 10081 18659 10084
rect 18601 10075 18659 10081
rect 18874 10072 18880 10084
rect 18932 10072 18938 10124
rect 19518 10072 19524 10124
rect 19576 10112 19582 10124
rect 19705 10115 19763 10121
rect 19705 10112 19717 10115
rect 19576 10084 19717 10112
rect 19576 10072 19582 10084
rect 19705 10081 19717 10084
rect 19751 10081 19763 10115
rect 19705 10075 19763 10081
rect 20806 10072 20812 10124
rect 20864 10072 20870 10124
rect 22002 10072 22008 10124
rect 22060 10112 22066 10124
rect 23293 10115 23351 10121
rect 23293 10112 23305 10115
rect 22060 10084 23305 10112
rect 22060 10072 22066 10084
rect 23293 10081 23305 10084
rect 23339 10081 23351 10115
rect 23293 10075 23351 10081
rect 23382 10072 23388 10124
rect 23440 10072 23446 10124
rect 12066 10004 12072 10056
rect 12124 10044 12130 10056
rect 13173 10047 13231 10053
rect 13173 10044 13185 10047
rect 12124 10016 13185 10044
rect 12124 10004 12130 10016
rect 13173 10013 13185 10016
rect 13219 10013 13231 10047
rect 15010 10044 15016 10056
rect 13173 10007 13231 10013
rect 14936 10016 15016 10044
rect 9306 9936 9312 9988
rect 9364 9976 9370 9988
rect 9585 9979 9643 9985
rect 9585 9976 9597 9979
rect 9364 9948 9597 9976
rect 9364 9936 9370 9948
rect 9585 9945 9597 9948
rect 9631 9945 9643 9979
rect 9585 9939 9643 9945
rect 9858 9936 9864 9988
rect 9916 9976 9922 9988
rect 11977 9979 12035 9985
rect 9916 9948 10074 9976
rect 9916 9936 9922 9948
rect 11977 9945 11989 9979
rect 12023 9976 12035 9979
rect 13722 9976 13728 9988
rect 12023 9948 13728 9976
rect 12023 9945 12035 9948
rect 11977 9939 12035 9945
rect 13722 9936 13728 9948
rect 13780 9936 13786 9988
rect 14936 9985 14964 10016
rect 15010 10004 15016 10016
rect 15068 10004 15074 10056
rect 16942 10004 16948 10056
rect 17000 10044 17006 10056
rect 20533 10047 20591 10053
rect 20533 10044 20545 10047
rect 17000 10016 20545 10044
rect 17000 10004 17006 10016
rect 20533 10013 20545 10016
rect 20579 10013 20591 10047
rect 20533 10007 20591 10013
rect 21910 10004 21916 10056
rect 21968 10004 21974 10056
rect 24026 10004 24032 10056
rect 24084 10044 24090 10056
rect 24765 10047 24823 10053
rect 24765 10044 24777 10047
rect 24084 10016 24777 10044
rect 24084 10004 24090 10016
rect 24765 10013 24777 10016
rect 24811 10013 24823 10047
rect 24765 10007 24823 10013
rect 14921 9979 14979 9985
rect 14921 9945 14933 9979
rect 14967 9945 14979 9979
rect 14921 9939 14979 9945
rect 16853 9979 16911 9985
rect 16853 9945 16865 9979
rect 16899 9976 16911 9979
rect 19058 9976 19064 9988
rect 16899 9948 19064 9976
rect 16899 9945 16911 9948
rect 16853 9939 16911 9945
rect 19058 9936 19064 9948
rect 19116 9936 19122 9988
rect 19521 9979 19579 9985
rect 19521 9945 19533 9979
rect 19567 9976 19579 9979
rect 23290 9976 23296 9988
rect 19567 9948 21220 9976
rect 19567 9945 19579 9948
rect 19521 9939 19579 9945
rect 21192 9920 21220 9948
rect 22848 9948 23296 9976
rect 12069 9911 12127 9917
rect 12069 9877 12081 9911
rect 12115 9908 12127 9911
rect 12802 9908 12808 9920
rect 12115 9880 12808 9908
rect 12115 9877 12127 9880
rect 12069 9871 12127 9877
rect 12802 9868 12808 9880
rect 12860 9868 12866 9920
rect 13265 9911 13323 9917
rect 13265 9877 13277 9911
rect 13311 9908 13323 9911
rect 13446 9908 13452 9920
rect 13311 9880 13452 9908
rect 13311 9877 13323 9880
rect 13265 9871 13323 9877
rect 13446 9868 13452 9880
rect 13504 9868 13510 9920
rect 13906 9868 13912 9920
rect 13964 9908 13970 9920
rect 14826 9908 14832 9920
rect 13964 9880 14832 9908
rect 13964 9868 13970 9880
rect 14826 9868 14832 9880
rect 14884 9868 14890 9920
rect 15013 9911 15071 9917
rect 15013 9877 15025 9911
rect 15059 9908 15071 9911
rect 15378 9908 15384 9920
rect 15059 9880 15384 9908
rect 15059 9877 15071 9880
rect 15013 9871 15071 9877
rect 15378 9868 15384 9880
rect 15436 9868 15442 9920
rect 16114 9868 16120 9920
rect 16172 9868 16178 9920
rect 16758 9868 16764 9920
rect 16816 9908 16822 9920
rect 16945 9911 17003 9917
rect 16945 9908 16957 9911
rect 16816 9880 16957 9908
rect 16816 9868 16822 9880
rect 16945 9877 16957 9880
rect 16991 9877 17003 9911
rect 16945 9871 17003 9877
rect 17678 9868 17684 9920
rect 17736 9908 17742 9920
rect 18325 9911 18383 9917
rect 18325 9908 18337 9911
rect 17736 9880 18337 9908
rect 17736 9868 17742 9880
rect 18325 9877 18337 9880
rect 18371 9877 18383 9911
rect 18325 9871 18383 9877
rect 18417 9911 18475 9917
rect 18417 9877 18429 9911
rect 18463 9908 18475 9911
rect 18690 9908 18696 9920
rect 18463 9880 18696 9908
rect 18463 9877 18475 9880
rect 18417 9871 18475 9877
rect 18690 9868 18696 9880
rect 18748 9908 18754 9920
rect 18969 9911 19027 9917
rect 18969 9908 18981 9911
rect 18748 9880 18981 9908
rect 18748 9868 18754 9880
rect 18969 9877 18981 9880
rect 19015 9877 19027 9911
rect 18969 9871 19027 9877
rect 21174 9868 21180 9920
rect 21232 9868 21238 9920
rect 22848 9917 22876 9948
rect 23290 9936 23296 9948
rect 23348 9936 23354 9988
rect 22833 9911 22891 9917
rect 22833 9877 22845 9911
rect 22879 9877 22891 9911
rect 22833 9871 22891 9877
rect 23201 9911 23259 9917
rect 23201 9877 23213 9911
rect 23247 9908 23259 9911
rect 24210 9908 24216 9920
rect 23247 9880 24216 9908
rect 23247 9877 23259 9880
rect 23201 9871 23259 9877
rect 24210 9868 24216 9880
rect 24268 9868 24274 9920
rect 1104 9818 25852 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 25852 9818
rect 1104 9744 25852 9766
rect 7098 9664 7104 9716
rect 7156 9704 7162 9716
rect 7156 9676 14596 9704
rect 7156 9664 7162 9676
rect 9858 9596 9864 9648
rect 9916 9636 9922 9648
rect 11146 9636 11152 9648
rect 9916 9608 11152 9636
rect 9916 9596 9922 9608
rect 11146 9596 11152 9608
rect 11204 9636 11210 9648
rect 11241 9639 11299 9645
rect 11241 9636 11253 9639
rect 11204 9608 11253 9636
rect 11204 9596 11210 9608
rect 11241 9605 11253 9608
rect 11287 9605 11299 9639
rect 13906 9636 13912 9648
rect 13202 9622 13912 9636
rect 11241 9599 11299 9605
rect 13188 9608 13912 9622
rect 11698 9528 11704 9580
rect 11756 9528 11762 9580
rect 11977 9503 12035 9509
rect 11977 9469 11989 9503
rect 12023 9500 12035 9503
rect 12526 9500 12532 9512
rect 12023 9472 12532 9500
rect 12023 9469 12035 9472
rect 11977 9463 12035 9469
rect 12526 9460 12532 9472
rect 12584 9460 12590 9512
rect 11146 9324 11152 9376
rect 11204 9364 11210 9376
rect 13188 9364 13216 9608
rect 13906 9596 13912 9608
rect 13964 9596 13970 9648
rect 13998 9596 14004 9648
rect 14056 9636 14062 9648
rect 14369 9639 14427 9645
rect 14369 9636 14381 9639
rect 14056 9608 14381 9636
rect 14056 9596 14062 9608
rect 14369 9605 14381 9608
rect 14415 9605 14427 9639
rect 14369 9599 14427 9605
rect 14277 9571 14335 9577
rect 14277 9537 14289 9571
rect 14323 9568 14335 9571
rect 14458 9568 14464 9580
rect 14323 9540 14464 9568
rect 14323 9537 14335 9540
rect 14277 9531 14335 9537
rect 14458 9528 14464 9540
rect 14516 9528 14522 9580
rect 13449 9503 13507 9509
rect 13449 9469 13461 9503
rect 13495 9500 13507 9503
rect 14090 9500 14096 9512
rect 13495 9472 14096 9500
rect 13495 9469 13507 9472
rect 13449 9463 13507 9469
rect 14090 9460 14096 9472
rect 14148 9460 14154 9512
rect 14568 9509 14596 9676
rect 16114 9664 16120 9716
rect 16172 9704 16178 9716
rect 20990 9704 20996 9716
rect 16172 9676 20996 9704
rect 16172 9664 16178 9676
rect 20990 9664 20996 9676
rect 21048 9664 21054 9716
rect 21082 9664 21088 9716
rect 21140 9704 21146 9716
rect 22005 9707 22063 9713
rect 22005 9704 22017 9707
rect 21140 9676 22017 9704
rect 21140 9664 21146 9676
rect 22005 9673 22017 9676
rect 22051 9673 22063 9707
rect 22005 9667 22063 9673
rect 22370 9664 22376 9716
rect 22428 9704 22434 9716
rect 24397 9707 24455 9713
rect 24397 9704 24409 9707
rect 22428 9676 24409 9704
rect 22428 9664 22434 9676
rect 24397 9673 24409 9676
rect 24443 9673 24455 9707
rect 24397 9667 24455 9673
rect 15473 9639 15531 9645
rect 15473 9605 15485 9639
rect 15519 9636 15531 9639
rect 17862 9636 17868 9648
rect 15519 9608 17868 9636
rect 15519 9605 15531 9608
rect 15473 9599 15531 9605
rect 17862 9596 17868 9608
rect 17920 9596 17926 9648
rect 19426 9636 19432 9648
rect 18814 9608 19432 9636
rect 19426 9596 19432 9608
rect 19484 9596 19490 9648
rect 19334 9528 19340 9580
rect 19392 9568 19398 9580
rect 20073 9571 20131 9577
rect 20073 9568 20085 9571
rect 19392 9540 20085 9568
rect 19392 9528 19398 9540
rect 20073 9537 20085 9540
rect 20119 9537 20131 9571
rect 20073 9531 20131 9537
rect 21269 9571 21327 9577
rect 21269 9537 21281 9571
rect 21315 9568 21327 9571
rect 22462 9568 22468 9580
rect 21315 9540 22468 9568
rect 21315 9537 21327 9540
rect 21269 9531 21327 9537
rect 22462 9528 22468 9540
rect 22520 9528 22526 9580
rect 24026 9528 24032 9580
rect 24084 9528 24090 9580
rect 25041 9571 25099 9577
rect 25041 9537 25053 9571
rect 25087 9537 25099 9571
rect 25041 9531 25099 9537
rect 14553 9503 14611 9509
rect 14553 9469 14565 9503
rect 14599 9500 14611 9503
rect 14918 9500 14924 9512
rect 14599 9472 14924 9500
rect 14599 9469 14611 9472
rect 14553 9463 14611 9469
rect 14918 9460 14924 9472
rect 14976 9460 14982 9512
rect 15565 9503 15623 9509
rect 15565 9469 15577 9503
rect 15611 9500 15623 9503
rect 15654 9500 15660 9512
rect 15611 9472 15660 9500
rect 15611 9469 15623 9472
rect 15565 9463 15623 9469
rect 15654 9460 15660 9472
rect 15712 9460 15718 9512
rect 15749 9503 15807 9509
rect 15749 9469 15761 9503
rect 15795 9500 15807 9503
rect 16206 9500 16212 9512
rect 15795 9472 16212 9500
rect 15795 9469 15807 9472
rect 15749 9463 15807 9469
rect 16206 9460 16212 9472
rect 16264 9460 16270 9512
rect 16942 9460 16948 9512
rect 17000 9500 17006 9512
rect 17313 9503 17371 9509
rect 17313 9500 17325 9503
rect 17000 9472 17325 9500
rect 17000 9460 17006 9472
rect 17313 9469 17325 9472
rect 17359 9469 17371 9503
rect 17313 9463 17371 9469
rect 17586 9460 17592 9512
rect 17644 9460 17650 9512
rect 17954 9460 17960 9512
rect 18012 9500 18018 9512
rect 19058 9500 19064 9512
rect 18012 9472 19064 9500
rect 18012 9460 18018 9472
rect 19058 9460 19064 9472
rect 19116 9460 19122 9512
rect 22002 9500 22008 9512
rect 19168 9472 22008 9500
rect 13722 9392 13728 9444
rect 13780 9432 13786 9444
rect 13909 9435 13967 9441
rect 13909 9432 13921 9435
rect 13780 9404 13921 9432
rect 13780 9392 13786 9404
rect 13909 9401 13921 9404
rect 13955 9401 13967 9435
rect 13909 9395 13967 9401
rect 15102 9392 15108 9444
rect 15160 9392 15166 9444
rect 19168 9432 19196 9472
rect 22002 9460 22008 9472
rect 22060 9460 22066 9512
rect 22646 9460 22652 9512
rect 22704 9460 22710 9512
rect 22925 9503 22983 9509
rect 22925 9469 22937 9503
rect 22971 9500 22983 9503
rect 23382 9500 23388 9512
rect 22971 9472 23388 9500
rect 22971 9469 22983 9472
rect 22925 9463 22983 9469
rect 23382 9460 23388 9472
rect 23440 9460 23446 9512
rect 25056 9500 25084 9531
rect 23952 9472 25084 9500
rect 18616 9404 19196 9432
rect 11204 9336 13216 9364
rect 11204 9324 11210 9336
rect 17402 9324 17408 9376
rect 17460 9364 17466 9376
rect 18616 9364 18644 9404
rect 20438 9392 20444 9444
rect 20496 9432 20502 9444
rect 21726 9432 21732 9444
rect 20496 9404 21732 9432
rect 20496 9392 20502 9404
rect 21726 9392 21732 9404
rect 21784 9432 21790 9444
rect 22664 9432 22692 9460
rect 21784 9404 22692 9432
rect 21784 9392 21790 9404
rect 17460 9336 18644 9364
rect 19061 9367 19119 9373
rect 17460 9324 17466 9336
rect 19061 9333 19073 9367
rect 19107 9364 19119 9367
rect 19150 9364 19156 9376
rect 19107 9336 19156 9364
rect 19107 9333 19119 9336
rect 19061 9327 19119 9333
rect 19150 9324 19156 9336
rect 19208 9324 19214 9376
rect 19426 9324 19432 9376
rect 19484 9364 19490 9376
rect 20346 9364 20352 9376
rect 19484 9336 20352 9364
rect 19484 9324 19490 9336
rect 20346 9324 20352 9336
rect 20404 9364 20410 9376
rect 21634 9364 21640 9376
rect 20404 9336 21640 9364
rect 20404 9324 20410 9336
rect 21634 9324 21640 9336
rect 21692 9324 21698 9376
rect 22738 9324 22744 9376
rect 22796 9364 22802 9376
rect 23952 9364 23980 9472
rect 24026 9392 24032 9444
rect 24084 9432 24090 9444
rect 24394 9432 24400 9444
rect 24084 9404 24400 9432
rect 24084 9392 24090 9404
rect 24394 9392 24400 9404
rect 24452 9432 24458 9444
rect 25317 9435 25375 9441
rect 25317 9432 25329 9435
rect 24452 9404 25329 9432
rect 24452 9392 24458 9404
rect 25317 9401 25329 9404
rect 25363 9401 25375 9435
rect 25317 9395 25375 9401
rect 22796 9336 23980 9364
rect 22796 9324 22802 9336
rect 24854 9324 24860 9376
rect 24912 9324 24918 9376
rect 1104 9274 25852 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 25852 9274
rect 1104 9200 25852 9222
rect 11146 9120 11152 9172
rect 11204 9120 11210 9172
rect 12802 9120 12808 9172
rect 12860 9160 12866 9172
rect 14277 9163 14335 9169
rect 14277 9160 14289 9163
rect 12860 9132 14289 9160
rect 12860 9120 12866 9132
rect 14277 9129 14289 9132
rect 14323 9129 14335 9163
rect 14277 9123 14335 9129
rect 15654 9120 15660 9172
rect 15712 9160 15718 9172
rect 18506 9160 18512 9172
rect 15712 9132 18512 9160
rect 15712 9120 15718 9132
rect 18506 9120 18512 9132
rect 18564 9120 18570 9172
rect 18690 9120 18696 9172
rect 18748 9160 18754 9172
rect 21542 9160 21548 9172
rect 18748 9132 21548 9160
rect 18748 9120 18754 9132
rect 21542 9120 21548 9132
rect 21600 9120 21606 9172
rect 21634 9120 21640 9172
rect 21692 9160 21698 9172
rect 22738 9160 22744 9172
rect 21692 9132 22744 9160
rect 21692 9120 21698 9132
rect 22738 9120 22744 9132
rect 22796 9120 22802 9172
rect 23934 9120 23940 9172
rect 23992 9160 23998 9172
rect 24581 9163 24639 9169
rect 24581 9160 24593 9163
rect 23992 9132 24593 9160
rect 23992 9120 23998 9132
rect 24581 9129 24593 9132
rect 24627 9129 24639 9163
rect 24581 9123 24639 9129
rect 12618 9052 12624 9104
rect 12676 9092 12682 9104
rect 12989 9095 13047 9101
rect 12989 9092 13001 9095
rect 12676 9064 13001 9092
rect 12676 9052 12682 9064
rect 12989 9061 13001 9064
rect 13035 9061 13047 9095
rect 12989 9055 13047 9061
rect 13630 9052 13636 9104
rect 13688 9092 13694 9104
rect 15933 9095 15991 9101
rect 15933 9092 15945 9095
rect 13688 9064 15945 9092
rect 13688 9052 13694 9064
rect 15933 9061 15945 9064
rect 15979 9061 15991 9095
rect 15933 9055 15991 9061
rect 17862 9052 17868 9104
rect 17920 9092 17926 9104
rect 19150 9092 19156 9104
rect 17920 9064 19156 9092
rect 17920 9052 17926 9064
rect 19150 9052 19156 9064
rect 19208 9052 19214 9104
rect 9125 9027 9183 9033
rect 9125 8993 9137 9027
rect 9171 9024 9183 9027
rect 11054 9024 11060 9036
rect 9171 8996 11060 9024
rect 9171 8993 9183 8996
rect 9125 8987 9183 8993
rect 11054 8984 11060 8996
rect 11112 9024 11118 9036
rect 11698 9024 11704 9036
rect 11112 8996 11704 9024
rect 11112 8984 11118 8996
rect 11698 8984 11704 8996
rect 11756 8984 11762 9036
rect 13538 8984 13544 9036
rect 13596 8984 13602 9036
rect 14918 8984 14924 9036
rect 14976 8984 14982 9036
rect 16482 8984 16488 9036
rect 16540 8984 16546 9036
rect 17052 8996 17264 9024
rect 14642 8916 14648 8968
rect 14700 8916 14706 8968
rect 16301 8959 16359 8965
rect 16301 8925 16313 8959
rect 16347 8956 16359 8959
rect 17052 8956 17080 8996
rect 16347 8928 17080 8956
rect 17236 8956 17264 8996
rect 17402 8984 17408 9036
rect 17460 9024 17466 9036
rect 17681 9027 17739 9033
rect 17681 9024 17693 9027
rect 17460 8996 17693 9024
rect 17460 8984 17466 8996
rect 17681 8993 17693 8996
rect 17727 8993 17739 9027
rect 17681 8987 17739 8993
rect 18506 8984 18512 9036
rect 18564 9024 18570 9036
rect 19613 9027 19671 9033
rect 19613 9024 19625 9027
rect 18564 8996 19625 9024
rect 18564 8984 18570 8996
rect 19613 8993 19625 8996
rect 19659 9024 19671 9027
rect 20438 9024 20444 9036
rect 19659 8996 20444 9024
rect 19659 8993 19671 8996
rect 19613 8987 19671 8993
rect 20438 8984 20444 8996
rect 20496 8984 20502 9036
rect 21634 8956 21640 8968
rect 17236 8928 19656 8956
rect 21022 8928 21640 8956
rect 16347 8925 16359 8928
rect 16301 8919 16359 8925
rect 9401 8891 9459 8897
rect 9401 8857 9413 8891
rect 9447 8888 9459 8891
rect 9674 8888 9680 8900
rect 9447 8860 9680 8888
rect 9447 8857 9459 8860
rect 9401 8851 9459 8857
rect 9674 8848 9680 8860
rect 9732 8848 9738 8900
rect 9858 8848 9864 8900
rect 9916 8848 9922 8900
rect 13357 8891 13415 8897
rect 13357 8857 13369 8891
rect 13403 8888 13415 8891
rect 13403 8860 17172 8888
rect 13403 8857 13415 8860
rect 13357 8851 13415 8857
rect 10873 8823 10931 8829
rect 10873 8789 10885 8823
rect 10919 8820 10931 8823
rect 10962 8820 10968 8832
rect 10919 8792 10968 8820
rect 10919 8789 10931 8792
rect 10873 8783 10931 8789
rect 10962 8780 10968 8792
rect 11020 8780 11026 8832
rect 13449 8823 13507 8829
rect 13449 8789 13461 8823
rect 13495 8820 13507 8823
rect 14182 8820 14188 8832
rect 13495 8792 14188 8820
rect 13495 8789 13507 8792
rect 13449 8783 13507 8789
rect 14182 8780 14188 8792
rect 14240 8780 14246 8832
rect 14642 8780 14648 8832
rect 14700 8820 14706 8832
rect 14737 8823 14795 8829
rect 14737 8820 14749 8823
rect 14700 8792 14749 8820
rect 14700 8780 14706 8792
rect 14737 8789 14749 8792
rect 14783 8789 14795 8823
rect 14737 8783 14795 8789
rect 15930 8780 15936 8832
rect 15988 8820 15994 8832
rect 16393 8823 16451 8829
rect 16393 8820 16405 8823
rect 15988 8792 16405 8820
rect 15988 8780 15994 8792
rect 16393 8789 16405 8792
rect 16439 8820 16451 8823
rect 16850 8820 16856 8832
rect 16439 8792 16856 8820
rect 16439 8789 16451 8792
rect 16393 8783 16451 8789
rect 16850 8780 16856 8792
rect 16908 8780 16914 8832
rect 17144 8829 17172 8860
rect 18690 8848 18696 8900
rect 18748 8848 18754 8900
rect 18877 8891 18935 8897
rect 18877 8857 18889 8891
rect 18923 8888 18935 8891
rect 19426 8888 19432 8900
rect 18923 8860 19432 8888
rect 18923 8857 18935 8860
rect 18877 8851 18935 8857
rect 19426 8848 19432 8860
rect 19484 8848 19490 8900
rect 17129 8823 17187 8829
rect 17129 8789 17141 8823
rect 17175 8789 17187 8823
rect 17129 8783 17187 8789
rect 17494 8780 17500 8832
rect 17552 8780 17558 8832
rect 17589 8823 17647 8829
rect 17589 8789 17601 8823
rect 17635 8820 17647 8823
rect 17678 8820 17684 8832
rect 17635 8792 17684 8820
rect 17635 8789 17647 8792
rect 17589 8783 17647 8789
rect 17678 8780 17684 8792
rect 17736 8780 17742 8832
rect 19628 8820 19656 8928
rect 21634 8916 21640 8928
rect 21692 8916 21698 8968
rect 22002 8916 22008 8968
rect 22060 8916 22066 8968
rect 22646 8916 22652 8968
rect 22704 8916 22710 8968
rect 23750 8916 23756 8968
rect 23808 8956 23814 8968
rect 24765 8959 24823 8965
rect 24765 8956 24777 8959
rect 23808 8928 24777 8956
rect 23808 8916 23814 8928
rect 24765 8925 24777 8928
rect 24811 8925 24823 8959
rect 24765 8919 24823 8925
rect 19889 8891 19947 8897
rect 19889 8857 19901 8891
rect 19935 8888 19947 8891
rect 19978 8888 19984 8900
rect 19935 8860 19984 8888
rect 19935 8857 19947 8860
rect 19889 8851 19947 8857
rect 19978 8848 19984 8860
rect 20036 8848 20042 8900
rect 23566 8888 23572 8900
rect 22066 8860 23572 8888
rect 20622 8820 20628 8832
rect 19628 8792 20628 8820
rect 20622 8780 20628 8792
rect 20680 8780 20686 8832
rect 20806 8780 20812 8832
rect 20864 8820 20870 8832
rect 21361 8823 21419 8829
rect 21361 8820 21373 8823
rect 20864 8792 21373 8820
rect 20864 8780 20870 8792
rect 21361 8789 21373 8792
rect 21407 8789 21419 8823
rect 21361 8783 21419 8789
rect 21821 8823 21879 8829
rect 21821 8789 21833 8823
rect 21867 8820 21879 8823
rect 22066 8820 22094 8860
rect 23566 8848 23572 8860
rect 23624 8848 23630 8900
rect 23845 8891 23903 8897
rect 23845 8857 23857 8891
rect 23891 8888 23903 8891
rect 24946 8888 24952 8900
rect 23891 8860 24952 8888
rect 23891 8857 23903 8860
rect 23845 8851 23903 8857
rect 24946 8848 24952 8860
rect 25004 8848 25010 8900
rect 21867 8792 22094 8820
rect 22373 8823 22431 8829
rect 21867 8789 21879 8792
rect 21821 8783 21879 8789
rect 22373 8789 22385 8823
rect 22419 8820 22431 8823
rect 22738 8820 22744 8832
rect 22419 8792 22744 8820
rect 22419 8789 22431 8792
rect 22373 8783 22431 8789
rect 22738 8780 22744 8792
rect 22796 8820 22802 8832
rect 23934 8820 23940 8832
rect 22796 8792 23940 8820
rect 22796 8780 22802 8792
rect 23934 8780 23940 8792
rect 23992 8780 23998 8832
rect 1104 8730 25852 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 25852 8730
rect 1104 8656 25852 8678
rect 15746 8616 15752 8628
rect 13924 8588 15752 8616
rect 13924 8557 13952 8588
rect 15746 8576 15752 8588
rect 15804 8576 15810 8628
rect 16850 8576 16856 8628
rect 16908 8616 16914 8628
rect 17313 8619 17371 8625
rect 17313 8616 17325 8619
rect 16908 8588 17325 8616
rect 16908 8576 16914 8588
rect 17313 8585 17325 8588
rect 17359 8585 17371 8619
rect 17313 8579 17371 8585
rect 17494 8576 17500 8628
rect 17552 8616 17558 8628
rect 20254 8616 20260 8628
rect 17552 8588 20260 8616
rect 17552 8576 17558 8588
rect 20254 8576 20260 8588
rect 20312 8616 20318 8628
rect 21266 8616 21272 8628
rect 20312 8588 21272 8616
rect 20312 8576 20318 8588
rect 21266 8576 21272 8588
rect 21324 8576 21330 8628
rect 22462 8576 22468 8628
rect 22520 8616 22526 8628
rect 24394 8616 24400 8628
rect 22520 8588 24400 8616
rect 22520 8576 22526 8588
rect 24394 8576 24400 8588
rect 24452 8576 24458 8628
rect 13909 8551 13967 8557
rect 13909 8517 13921 8551
rect 13955 8517 13967 8551
rect 13909 8511 13967 8517
rect 15120 8520 21772 8548
rect 14274 8440 14280 8492
rect 14332 8480 14338 8492
rect 15120 8489 15148 8520
rect 15105 8483 15163 8489
rect 14332 8452 15056 8480
rect 14332 8440 14338 8452
rect 11698 8372 11704 8424
rect 11756 8372 11762 8424
rect 13173 8415 13231 8421
rect 13173 8381 13185 8415
rect 13219 8412 13231 8415
rect 13354 8412 13360 8424
rect 13219 8384 13360 8412
rect 13219 8381 13231 8384
rect 13173 8375 13231 8381
rect 13354 8372 13360 8384
rect 13412 8372 13418 8424
rect 14016 8384 14780 8412
rect 10502 8304 10508 8356
rect 10560 8344 10566 8356
rect 14016 8344 14044 8384
rect 10560 8316 14044 8344
rect 10560 8304 10566 8316
rect 14090 8304 14096 8356
rect 14148 8304 14154 8356
rect 14752 8344 14780 8384
rect 14826 8372 14832 8424
rect 14884 8372 14890 8424
rect 15028 8412 15056 8452
rect 15105 8449 15117 8483
rect 15151 8449 15163 8483
rect 17221 8483 17279 8489
rect 17221 8480 17233 8483
rect 15105 8443 15163 8449
rect 15212 8452 17233 8480
rect 15212 8412 15240 8452
rect 17221 8449 17233 8452
rect 17267 8449 17279 8483
rect 17221 8443 17279 8449
rect 17328 8452 17540 8480
rect 15028 8384 15240 8412
rect 16114 8372 16120 8424
rect 16172 8372 16178 8424
rect 17328 8412 17356 8452
rect 16776 8384 17356 8412
rect 16776 8344 16804 8384
rect 17402 8372 17408 8424
rect 17460 8372 17466 8424
rect 17512 8412 17540 8452
rect 17770 8440 17776 8492
rect 17828 8480 17834 8492
rect 17865 8483 17923 8489
rect 17865 8480 17877 8483
rect 17828 8452 17877 8480
rect 17828 8440 17834 8452
rect 17865 8449 17877 8452
rect 17911 8449 17923 8483
rect 17865 8443 17923 8449
rect 18230 8440 18236 8492
rect 18288 8440 18294 8492
rect 20070 8440 20076 8492
rect 20128 8440 20134 8492
rect 17678 8412 17684 8424
rect 17512 8384 17684 8412
rect 17678 8372 17684 8384
rect 17736 8372 17742 8424
rect 19429 8415 19487 8421
rect 19429 8381 19441 8415
rect 19475 8412 19487 8415
rect 20530 8412 20536 8424
rect 19475 8384 20536 8412
rect 19475 8381 19487 8384
rect 19429 8375 19487 8381
rect 20530 8372 20536 8384
rect 20588 8372 20594 8424
rect 21269 8415 21327 8421
rect 21269 8381 21281 8415
rect 21315 8412 21327 8415
rect 21634 8412 21640 8424
rect 21315 8384 21640 8412
rect 21315 8381 21327 8384
rect 21269 8375 21327 8381
rect 21634 8372 21640 8384
rect 21692 8372 21698 8424
rect 21744 8412 21772 8520
rect 22278 8440 22284 8492
rect 22336 8440 22342 8492
rect 23937 8483 23995 8489
rect 23937 8480 23949 8483
rect 22388 8452 23949 8480
rect 22388 8412 22416 8452
rect 23937 8449 23949 8452
rect 23983 8449 23995 8483
rect 23937 8443 23995 8449
rect 21744 8384 22416 8412
rect 22462 8372 22468 8424
rect 22520 8412 22526 8424
rect 22557 8415 22615 8421
rect 22557 8412 22569 8415
rect 22520 8384 22569 8412
rect 22520 8372 22526 8384
rect 22557 8381 22569 8384
rect 22603 8381 22615 8415
rect 22557 8375 22615 8381
rect 24762 8372 24768 8424
rect 24820 8372 24826 8424
rect 14752 8316 16804 8344
rect 16853 8347 16911 8353
rect 16853 8313 16865 8347
rect 16899 8344 16911 8347
rect 19242 8344 19248 8356
rect 16899 8316 19248 8344
rect 16899 8313 16911 8316
rect 16853 8307 16911 8313
rect 19242 8304 19248 8316
rect 19300 8304 19306 8356
rect 11146 8236 11152 8288
rect 11204 8276 11210 8288
rect 17218 8276 17224 8288
rect 11204 8248 17224 8276
rect 11204 8236 11210 8248
rect 17218 8236 17224 8248
rect 17276 8236 17282 8288
rect 17954 8236 17960 8288
rect 18012 8276 18018 8288
rect 22830 8276 22836 8288
rect 18012 8248 22836 8276
rect 18012 8236 18018 8248
rect 22830 8236 22836 8248
rect 22888 8236 22894 8288
rect 1104 8186 25852 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 25852 8186
rect 1104 8112 25852 8134
rect 11057 8075 11115 8081
rect 11057 8041 11069 8075
rect 11103 8072 11115 8075
rect 11146 8072 11152 8084
rect 11103 8044 11152 8072
rect 11103 8041 11115 8044
rect 11057 8035 11115 8041
rect 11146 8032 11152 8044
rect 11204 8032 11210 8084
rect 12989 8075 13047 8081
rect 12989 8041 13001 8075
rect 13035 8072 13047 8075
rect 13538 8072 13544 8084
rect 13035 8044 13544 8072
rect 13035 8041 13047 8044
rect 12989 8035 13047 8041
rect 13538 8032 13544 8044
rect 13596 8032 13602 8084
rect 14182 8032 14188 8084
rect 14240 8072 14246 8084
rect 15841 8075 15899 8081
rect 15841 8072 15853 8075
rect 14240 8044 15853 8072
rect 14240 8032 14246 8044
rect 15841 8041 15853 8044
rect 15887 8041 15899 8075
rect 15841 8035 15899 8041
rect 16482 8032 16488 8084
rect 16540 8072 16546 8084
rect 21818 8072 21824 8084
rect 16540 8044 21824 8072
rect 16540 8032 16546 8044
rect 21818 8032 21824 8044
rect 21876 8032 21882 8084
rect 22066 8044 23428 8072
rect 12526 7964 12532 8016
rect 12584 8004 12590 8016
rect 12584 7976 14688 8004
rect 12584 7964 12590 7976
rect 11606 7896 11612 7948
rect 11664 7896 11670 7948
rect 13633 7939 13691 7945
rect 13633 7905 13645 7939
rect 13679 7936 13691 7939
rect 14550 7936 14556 7948
rect 13679 7908 14556 7936
rect 13679 7905 13691 7908
rect 13633 7899 13691 7905
rect 14550 7896 14556 7908
rect 14608 7896 14614 7948
rect 14660 7936 14688 7976
rect 15010 7964 15016 8016
rect 15068 8004 15074 8016
rect 18414 8004 18420 8016
rect 15068 7976 18420 8004
rect 15068 7964 15074 7976
rect 18414 7964 18420 7976
rect 18472 7964 18478 8016
rect 19981 8007 20039 8013
rect 19981 7973 19993 8007
rect 20027 8004 20039 8007
rect 20346 8004 20352 8016
rect 20027 7976 20352 8004
rect 20027 7973 20039 7976
rect 19981 7967 20039 7973
rect 20346 7964 20352 7976
rect 20404 7964 20410 8016
rect 22066 8004 22094 8044
rect 20456 7976 22094 8004
rect 23400 8004 23428 8044
rect 23474 8032 23480 8084
rect 23532 8072 23538 8084
rect 24765 8075 24823 8081
rect 24765 8072 24777 8075
rect 23532 8044 24777 8072
rect 23532 8032 23538 8044
rect 24765 8041 24777 8044
rect 24811 8041 24823 8075
rect 24765 8035 24823 8041
rect 24026 8004 24032 8016
rect 23400 7976 24032 8004
rect 14829 7939 14887 7945
rect 14829 7936 14841 7939
rect 14660 7908 14841 7936
rect 14829 7905 14841 7908
rect 14875 7905 14887 7939
rect 14829 7899 14887 7905
rect 16206 7896 16212 7948
rect 16264 7936 16270 7948
rect 16485 7939 16543 7945
rect 16485 7936 16497 7939
rect 16264 7908 16497 7936
rect 16264 7896 16270 7908
rect 16485 7905 16497 7908
rect 16531 7936 16543 7939
rect 17494 7936 17500 7948
rect 16531 7908 17500 7936
rect 16531 7905 16543 7908
rect 16485 7899 16543 7905
rect 17494 7896 17500 7908
rect 17552 7896 17558 7948
rect 18693 7939 18751 7945
rect 18693 7905 18705 7939
rect 18739 7936 18751 7939
rect 20254 7936 20260 7948
rect 18739 7908 20260 7936
rect 18739 7905 18751 7908
rect 18693 7899 18751 7905
rect 20254 7896 20260 7908
rect 20312 7896 20318 7948
rect 11425 7871 11483 7877
rect 11425 7837 11437 7871
rect 11471 7868 11483 7871
rect 11698 7868 11704 7880
rect 11471 7840 11704 7868
rect 11471 7837 11483 7840
rect 11425 7831 11483 7837
rect 11698 7828 11704 7840
rect 11756 7828 11762 7880
rect 13354 7828 13360 7880
rect 13412 7828 13418 7880
rect 14645 7871 14703 7877
rect 14645 7837 14657 7871
rect 14691 7868 14703 7871
rect 16114 7868 16120 7880
rect 14691 7840 16120 7868
rect 14691 7837 14703 7840
rect 14645 7831 14703 7837
rect 16114 7828 16120 7840
rect 16172 7828 16178 7880
rect 16301 7871 16359 7877
rect 16301 7868 16313 7871
rect 16211 7840 16313 7868
rect 11517 7803 11575 7809
rect 11517 7800 11529 7803
rect 2746 7772 11529 7800
rect 2222 7692 2228 7744
rect 2280 7732 2286 7744
rect 2746 7732 2774 7772
rect 11517 7769 11529 7772
rect 11563 7769 11575 7803
rect 13449 7803 13507 7809
rect 13449 7800 13461 7803
rect 11517 7763 11575 7769
rect 11624 7772 13461 7800
rect 2280 7704 2774 7732
rect 2280 7692 2286 7704
rect 11146 7692 11152 7744
rect 11204 7732 11210 7744
rect 11624 7732 11652 7772
rect 13449 7769 13461 7772
rect 13495 7769 13507 7803
rect 14737 7803 14795 7809
rect 14737 7800 14749 7803
rect 13449 7763 13507 7769
rect 13556 7772 14749 7800
rect 11204 7704 11652 7732
rect 12345 7735 12403 7741
rect 11204 7692 11210 7704
rect 12345 7701 12357 7735
rect 12391 7732 12403 7735
rect 12618 7732 12624 7744
rect 12391 7704 12624 7732
rect 12391 7701 12403 7704
rect 12345 7695 12403 7701
rect 12618 7692 12624 7704
rect 12676 7692 12682 7744
rect 13354 7692 13360 7744
rect 13412 7732 13418 7744
rect 13556 7732 13584 7772
rect 14737 7769 14749 7772
rect 14783 7769 14795 7803
rect 14737 7763 14795 7769
rect 15746 7760 15752 7812
rect 15804 7800 15810 7812
rect 16211 7800 16239 7840
rect 16301 7837 16313 7840
rect 16347 7837 16359 7871
rect 16301 7831 16359 7837
rect 17681 7871 17739 7877
rect 17681 7837 17693 7871
rect 17727 7868 17739 7871
rect 17954 7868 17960 7880
rect 17727 7840 17960 7868
rect 17727 7837 17739 7840
rect 17681 7831 17739 7837
rect 17954 7828 17960 7840
rect 18012 7828 18018 7880
rect 19613 7871 19671 7877
rect 19613 7837 19625 7871
rect 19659 7868 19671 7871
rect 19794 7868 19800 7880
rect 19659 7840 19800 7868
rect 19659 7837 19671 7840
rect 19613 7831 19671 7837
rect 19794 7828 19800 7840
rect 19852 7828 19858 7880
rect 19886 7828 19892 7880
rect 19944 7868 19950 7880
rect 20162 7868 20168 7880
rect 19944 7840 20168 7868
rect 19944 7828 19950 7840
rect 20162 7828 20168 7840
rect 20220 7828 20226 7880
rect 20456 7877 20484 7976
rect 24026 7964 24032 7976
rect 24084 7964 24090 8016
rect 22370 7896 22376 7948
rect 22428 7896 22434 7948
rect 20441 7871 20499 7877
rect 20441 7837 20453 7871
rect 20487 7837 20499 7871
rect 20441 7831 20499 7837
rect 21726 7828 21732 7880
rect 21784 7868 21790 7880
rect 22097 7871 22155 7877
rect 22097 7868 22109 7871
rect 21784 7840 22109 7868
rect 21784 7828 21790 7840
rect 22097 7837 22109 7840
rect 22143 7837 22155 7871
rect 23934 7868 23940 7880
rect 23506 7840 23940 7868
rect 22097 7831 22155 7837
rect 23934 7828 23940 7840
rect 23992 7828 23998 7880
rect 15804 7772 16239 7800
rect 15804 7760 15810 7772
rect 17770 7760 17776 7812
rect 17828 7800 17834 7812
rect 18322 7800 18328 7812
rect 17828 7772 18328 7800
rect 17828 7760 17834 7772
rect 18322 7760 18328 7772
rect 18380 7760 18386 7812
rect 21082 7800 21088 7812
rect 19444 7772 21088 7800
rect 13412 7704 13584 7732
rect 14277 7735 14335 7741
rect 13412 7692 13418 7704
rect 14277 7701 14289 7735
rect 14323 7732 14335 7735
rect 15010 7732 15016 7744
rect 14323 7704 15016 7732
rect 14323 7701 14335 7704
rect 14277 7695 14335 7701
rect 15010 7692 15016 7704
rect 15068 7692 15074 7744
rect 16209 7735 16267 7741
rect 16209 7701 16221 7735
rect 16255 7732 16267 7735
rect 16482 7732 16488 7744
rect 16255 7704 16488 7732
rect 16255 7701 16267 7704
rect 16209 7695 16267 7701
rect 16482 7692 16488 7704
rect 16540 7692 16546 7744
rect 16850 7692 16856 7744
rect 16908 7732 16914 7744
rect 17126 7732 17132 7744
rect 16908 7704 17132 7732
rect 16908 7692 16914 7704
rect 17126 7692 17132 7704
rect 17184 7732 17190 7744
rect 17862 7732 17868 7744
rect 17184 7704 17868 7732
rect 17184 7692 17190 7704
rect 17862 7692 17868 7704
rect 17920 7692 17926 7744
rect 19444 7741 19472 7772
rect 21082 7760 21088 7772
rect 21140 7760 21146 7812
rect 21450 7760 21456 7812
rect 21508 7760 21514 7812
rect 24673 7803 24731 7809
rect 24673 7800 24685 7803
rect 23676 7772 24685 7800
rect 19429 7735 19487 7741
rect 19429 7701 19441 7735
rect 19475 7701 19487 7735
rect 19429 7695 19487 7701
rect 20806 7692 20812 7744
rect 20864 7732 20870 7744
rect 23676 7732 23704 7772
rect 24673 7769 24685 7772
rect 24719 7769 24731 7803
rect 24673 7763 24731 7769
rect 20864 7704 23704 7732
rect 20864 7692 20870 7704
rect 23842 7692 23848 7744
rect 23900 7692 23906 7744
rect 23934 7692 23940 7744
rect 23992 7732 23998 7744
rect 24213 7735 24271 7741
rect 24213 7732 24225 7735
rect 23992 7704 24225 7732
rect 23992 7692 23998 7704
rect 24213 7701 24225 7704
rect 24259 7732 24271 7735
rect 24762 7732 24768 7744
rect 24259 7704 24768 7732
rect 24259 7701 24271 7704
rect 24213 7695 24271 7701
rect 24762 7692 24768 7704
rect 24820 7692 24826 7744
rect 1104 7642 25852 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 25852 7642
rect 1104 7568 25852 7590
rect 12253 7531 12311 7537
rect 12253 7497 12265 7531
rect 12299 7528 12311 7531
rect 12299 7500 12434 7528
rect 12299 7497 12311 7500
rect 12253 7491 12311 7497
rect 9582 7460 9588 7472
rect 9048 7432 9588 7460
rect 9048 7401 9076 7432
rect 9582 7420 9588 7432
rect 9640 7420 9646 7472
rect 11514 7460 11520 7472
rect 10534 7432 11520 7460
rect 11514 7420 11520 7432
rect 11572 7420 11578 7472
rect 12406 7460 12434 7500
rect 12618 7488 12624 7540
rect 12676 7488 12682 7540
rect 13630 7488 13636 7540
rect 13688 7528 13694 7540
rect 15473 7531 15531 7537
rect 15473 7528 15485 7531
rect 13688 7500 15485 7528
rect 13688 7488 13694 7500
rect 15473 7497 15485 7500
rect 15519 7497 15531 7531
rect 15473 7491 15531 7497
rect 17770 7488 17776 7540
rect 17828 7488 17834 7540
rect 19150 7488 19156 7540
rect 19208 7528 19214 7540
rect 19208 7500 20116 7528
rect 19208 7488 19214 7500
rect 14274 7460 14280 7472
rect 12406 7432 14280 7460
rect 14274 7420 14280 7432
rect 14332 7420 14338 7472
rect 15010 7420 15016 7472
rect 15068 7420 15074 7472
rect 16301 7463 16359 7469
rect 16301 7429 16313 7463
rect 16347 7460 16359 7463
rect 18782 7460 18788 7472
rect 16347 7432 18788 7460
rect 16347 7429 16359 7432
rect 16301 7423 16359 7429
rect 18782 7420 18788 7432
rect 18840 7420 18846 7472
rect 20088 7460 20116 7500
rect 20254 7488 20260 7540
rect 20312 7528 20318 7540
rect 25314 7528 25320 7540
rect 20312 7500 25320 7528
rect 20312 7488 20318 7500
rect 25314 7488 25320 7500
rect 25372 7488 25378 7540
rect 20346 7460 20352 7472
rect 20010 7432 20352 7460
rect 20346 7420 20352 7432
rect 20404 7420 20410 7472
rect 20990 7420 20996 7472
rect 21048 7460 21054 7472
rect 21085 7463 21143 7469
rect 21085 7460 21097 7463
rect 21048 7432 21097 7460
rect 21048 7420 21054 7432
rect 21085 7429 21097 7432
rect 21131 7429 21143 7463
rect 21085 7423 21143 7429
rect 21174 7420 21180 7472
rect 21232 7460 21238 7472
rect 21232 7432 23980 7460
rect 21232 7420 21238 7432
rect 9033 7395 9091 7401
rect 9033 7361 9045 7395
rect 9079 7361 9091 7395
rect 9033 7355 9091 7361
rect 16117 7395 16175 7401
rect 16117 7361 16129 7395
rect 16163 7392 16175 7395
rect 16390 7392 16396 7404
rect 16163 7364 16396 7392
rect 16163 7361 16175 7364
rect 16117 7355 16175 7361
rect 16390 7352 16396 7364
rect 16448 7352 16454 7404
rect 17678 7352 17684 7404
rect 17736 7352 17742 7404
rect 18506 7352 18512 7404
rect 18564 7352 18570 7404
rect 23952 7401 23980 7432
rect 25130 7420 25136 7472
rect 25188 7420 25194 7472
rect 22281 7395 22339 7401
rect 22281 7361 22293 7395
rect 22327 7392 22339 7395
rect 23937 7395 23995 7401
rect 22327 7364 22968 7392
rect 22327 7361 22339 7364
rect 22281 7355 22339 7361
rect 9309 7327 9367 7333
rect 9309 7293 9321 7327
rect 9355 7324 9367 7327
rect 10962 7324 10968 7336
rect 9355 7296 10968 7324
rect 9355 7293 9367 7296
rect 9309 7287 9367 7293
rect 10962 7284 10968 7296
rect 11020 7284 11026 7336
rect 11422 7284 11428 7336
rect 11480 7324 11486 7336
rect 12713 7327 12771 7333
rect 12713 7324 12725 7327
rect 11480 7296 12725 7324
rect 11480 7284 11486 7296
rect 12713 7293 12725 7296
rect 12759 7293 12771 7327
rect 12713 7287 12771 7293
rect 12805 7327 12863 7333
rect 12805 7293 12817 7327
rect 12851 7293 12863 7327
rect 12805 7287 12863 7293
rect 13725 7327 13783 7333
rect 13725 7293 13737 7327
rect 13771 7293 13783 7327
rect 13725 7287 13783 7293
rect 14001 7327 14059 7333
rect 14001 7293 14013 7327
rect 14047 7324 14059 7327
rect 16666 7324 16672 7336
rect 14047 7296 16672 7324
rect 14047 7293 14059 7296
rect 14001 7287 14059 7293
rect 12820 7256 12848 7287
rect 10796 7228 12848 7256
rect 10796 7200 10824 7228
rect 10778 7148 10784 7200
rect 10836 7148 10842 7200
rect 11149 7191 11207 7197
rect 11149 7157 11161 7191
rect 11195 7188 11207 7191
rect 11514 7188 11520 7200
rect 11195 7160 11520 7188
rect 11195 7157 11207 7160
rect 11149 7151 11207 7157
rect 11514 7148 11520 7160
rect 11572 7148 11578 7200
rect 13740 7188 13768 7287
rect 16666 7284 16672 7296
rect 16724 7284 16730 7336
rect 17586 7284 17592 7336
rect 17644 7324 17650 7336
rect 17865 7327 17923 7333
rect 17865 7324 17877 7327
rect 17644 7296 17877 7324
rect 17644 7284 17650 7296
rect 17865 7293 17877 7296
rect 17911 7293 17923 7327
rect 17865 7287 17923 7293
rect 18785 7327 18843 7333
rect 18785 7293 18797 7327
rect 18831 7324 18843 7327
rect 18874 7324 18880 7336
rect 18831 7296 18880 7324
rect 18831 7293 18843 7296
rect 18785 7287 18843 7293
rect 18874 7284 18880 7296
rect 18932 7284 18938 7336
rect 19242 7284 19248 7336
rect 19300 7324 19306 7336
rect 21177 7327 21235 7333
rect 21177 7324 21189 7327
rect 19300 7296 21189 7324
rect 19300 7284 19306 7296
rect 21177 7293 21189 7296
rect 21223 7293 21235 7327
rect 21177 7287 21235 7293
rect 21269 7327 21327 7333
rect 21269 7293 21281 7327
rect 21315 7293 21327 7327
rect 21269 7287 21327 7293
rect 18322 7256 18328 7268
rect 16684 7228 18328 7256
rect 15102 7188 15108 7200
rect 13740 7160 15108 7188
rect 15102 7148 15108 7160
rect 15160 7148 15166 7200
rect 15470 7148 15476 7200
rect 15528 7188 15534 7200
rect 16684 7197 16712 7228
rect 18322 7216 18328 7228
rect 18380 7216 18386 7268
rect 19886 7216 19892 7268
rect 19944 7256 19950 7268
rect 21284 7256 21312 7287
rect 19944 7228 21312 7256
rect 22940 7256 22968 7364
rect 23937 7361 23949 7395
rect 23983 7361 23995 7395
rect 23937 7355 23995 7361
rect 23293 7327 23351 7333
rect 23293 7293 23305 7327
rect 23339 7324 23351 7327
rect 24854 7324 24860 7336
rect 23339 7296 24860 7324
rect 23339 7293 23351 7296
rect 23293 7287 23351 7293
rect 24854 7284 24860 7296
rect 24912 7284 24918 7336
rect 24118 7256 24124 7268
rect 22940 7228 24124 7256
rect 19944 7216 19950 7228
rect 24118 7216 24124 7228
rect 24176 7216 24182 7268
rect 16669 7191 16727 7197
rect 16669 7188 16681 7191
rect 15528 7160 16681 7188
rect 15528 7148 15534 7160
rect 16669 7157 16681 7160
rect 16715 7157 16727 7191
rect 16669 7151 16727 7157
rect 17037 7191 17095 7197
rect 17037 7157 17049 7191
rect 17083 7188 17095 7191
rect 17218 7188 17224 7200
rect 17083 7160 17224 7188
rect 17083 7157 17095 7160
rect 17037 7151 17095 7157
rect 17218 7148 17224 7160
rect 17276 7148 17282 7200
rect 17313 7191 17371 7197
rect 17313 7157 17325 7191
rect 17359 7188 17371 7191
rect 17770 7188 17776 7200
rect 17359 7160 17776 7188
rect 17359 7157 17371 7160
rect 17313 7151 17371 7157
rect 17770 7148 17776 7160
rect 17828 7148 17834 7200
rect 19242 7148 19248 7200
rect 19300 7188 19306 7200
rect 20257 7191 20315 7197
rect 20257 7188 20269 7191
rect 19300 7160 20269 7188
rect 19300 7148 19306 7160
rect 20257 7157 20269 7160
rect 20303 7157 20315 7191
rect 20257 7151 20315 7157
rect 20717 7191 20775 7197
rect 20717 7157 20729 7191
rect 20763 7188 20775 7191
rect 22554 7188 22560 7200
rect 20763 7160 22560 7188
rect 20763 7157 20775 7160
rect 20717 7151 20775 7157
rect 22554 7148 22560 7160
rect 22612 7148 22618 7200
rect 1104 7098 25852 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 25852 7098
rect 1104 7024 25852 7046
rect 11606 6944 11612 6996
rect 11664 6984 11670 6996
rect 16850 6984 16856 6996
rect 11664 6956 16856 6984
rect 11664 6944 11670 6956
rect 16850 6944 16856 6956
rect 16908 6944 16914 6996
rect 17126 6944 17132 6996
rect 17184 6984 17190 6996
rect 17184 6956 18460 6984
rect 17184 6944 17190 6956
rect 15013 6919 15071 6925
rect 15013 6885 15025 6919
rect 15059 6916 15071 6919
rect 18432 6916 18460 6956
rect 19242 6944 19248 6996
rect 19300 6984 19306 6996
rect 23934 6984 23940 6996
rect 19300 6956 23940 6984
rect 19300 6944 19306 6956
rect 23934 6944 23940 6956
rect 23992 6944 23998 6996
rect 21174 6916 21180 6928
rect 15059 6888 15148 6916
rect 18432 6888 21180 6916
rect 15059 6885 15071 6888
rect 15013 6879 15071 6885
rect 10781 6851 10839 6857
rect 10781 6817 10793 6851
rect 10827 6848 10839 6851
rect 11054 6848 11060 6860
rect 10827 6820 11060 6848
rect 10827 6817 10839 6820
rect 10781 6811 10839 6817
rect 11054 6808 11060 6820
rect 11112 6808 11118 6860
rect 11514 6808 11520 6860
rect 11572 6848 11578 6860
rect 11572 6820 12434 6848
rect 11572 6808 11578 6820
rect 12406 6780 12434 6820
rect 12526 6808 12532 6860
rect 12584 6808 12590 6860
rect 12897 6851 12955 6857
rect 12897 6817 12909 6851
rect 12943 6848 12955 6851
rect 12943 6820 15056 6848
rect 12943 6817 12955 6820
rect 12897 6811 12955 6817
rect 12912 6780 12940 6811
rect 15028 6792 15056 6820
rect 12406 6752 12940 6780
rect 13722 6740 13728 6792
rect 13780 6740 13786 6792
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6780 14611 6783
rect 14734 6780 14740 6792
rect 14599 6752 14740 6780
rect 14599 6749 14611 6752
rect 14553 6743 14611 6749
rect 14734 6740 14740 6752
rect 14792 6740 14798 6792
rect 15010 6740 15016 6792
rect 15068 6740 15074 6792
rect 15120 6780 15148 6888
rect 21174 6876 21180 6888
rect 21232 6876 21238 6928
rect 23842 6876 23848 6928
rect 23900 6916 23906 6928
rect 23900 6888 25176 6916
rect 23900 6876 23906 6888
rect 15378 6808 15384 6860
rect 15436 6848 15442 6860
rect 15565 6851 15623 6857
rect 15565 6848 15577 6851
rect 15436 6820 15577 6848
rect 15436 6808 15442 6820
rect 15565 6817 15577 6820
rect 15611 6817 15623 6851
rect 15565 6811 15623 6817
rect 15746 6808 15752 6860
rect 15804 6848 15810 6860
rect 18877 6851 18935 6857
rect 15804 6820 18644 6848
rect 15804 6808 15810 6820
rect 16390 6780 16396 6792
rect 15120 6752 16396 6780
rect 16390 6740 16396 6752
rect 16448 6740 16454 6792
rect 16942 6740 16948 6792
rect 17000 6780 17006 6792
rect 17129 6783 17187 6789
rect 17129 6780 17141 6783
rect 17000 6752 17141 6780
rect 17000 6740 17006 6752
rect 17129 6749 17141 6752
rect 17175 6749 17187 6783
rect 18616 6780 18644 6820
rect 18877 6817 18889 6851
rect 18923 6848 18935 6851
rect 19886 6848 19892 6860
rect 18923 6820 19892 6848
rect 18923 6817 18935 6820
rect 18877 6811 18935 6817
rect 19886 6808 19892 6820
rect 19944 6808 19950 6860
rect 19978 6808 19984 6860
rect 20036 6848 20042 6860
rect 20073 6851 20131 6857
rect 20073 6848 20085 6851
rect 20036 6820 20085 6848
rect 20036 6808 20042 6820
rect 20073 6817 20085 6820
rect 20119 6848 20131 6851
rect 23750 6848 23756 6860
rect 20119 6820 23756 6848
rect 20119 6817 20131 6820
rect 20073 6811 20131 6817
rect 23750 6808 23756 6820
rect 23808 6808 23814 6860
rect 25148 6857 25176 6888
rect 25133 6851 25191 6857
rect 25133 6817 25145 6851
rect 25179 6817 25191 6851
rect 25133 6811 25191 6817
rect 19797 6783 19855 6789
rect 19797 6780 19809 6783
rect 18616 6752 19809 6780
rect 17129 6743 17187 6749
rect 19797 6749 19809 6752
rect 19843 6749 19855 6783
rect 19797 6743 19855 6749
rect 20346 6740 20352 6792
rect 20404 6780 20410 6792
rect 20441 6783 20499 6789
rect 20441 6780 20453 6783
rect 20404 6752 20453 6780
rect 20404 6740 20410 6752
rect 20441 6749 20453 6752
rect 20487 6749 20499 6783
rect 20441 6743 20499 6749
rect 20898 6740 20904 6792
rect 20956 6740 20962 6792
rect 22646 6740 22652 6792
rect 22704 6740 22710 6792
rect 23845 6783 23903 6789
rect 23845 6749 23857 6783
rect 23891 6780 23903 6783
rect 24946 6780 24952 6792
rect 23891 6752 24952 6780
rect 23891 6749 23903 6752
rect 23845 6743 23903 6749
rect 24946 6740 24952 6752
rect 25004 6740 25010 6792
rect 11057 6715 11115 6721
rect 11057 6681 11069 6715
rect 11103 6712 11115 6715
rect 11330 6712 11336 6724
rect 11103 6684 11336 6712
rect 11103 6681 11115 6684
rect 11057 6675 11115 6681
rect 11330 6672 11336 6684
rect 11388 6672 11394 6724
rect 11514 6672 11520 6724
rect 11572 6672 11578 6724
rect 12802 6672 12808 6724
rect 12860 6712 12866 6724
rect 15381 6715 15439 6721
rect 15381 6712 15393 6715
rect 12860 6684 15393 6712
rect 12860 6672 12866 6684
rect 15381 6681 15393 6684
rect 15427 6681 15439 6715
rect 15381 6675 15439 6681
rect 15470 6672 15476 6724
rect 15528 6672 15534 6724
rect 15838 6672 15844 6724
rect 15896 6712 15902 6724
rect 16485 6715 16543 6721
rect 16485 6712 16497 6715
rect 15896 6684 16497 6712
rect 15896 6672 15902 6684
rect 16485 6681 16497 6684
rect 16531 6681 16543 6715
rect 16485 6675 16543 6681
rect 16574 6672 16580 6724
rect 16632 6712 16638 6724
rect 16669 6715 16727 6721
rect 16669 6712 16681 6715
rect 16632 6684 16681 6712
rect 16632 6672 16638 6684
rect 16669 6681 16681 6684
rect 16715 6681 16727 6715
rect 16669 6675 16727 6681
rect 17402 6672 17408 6724
rect 17460 6672 17466 6724
rect 19150 6712 19156 6724
rect 18630 6684 19156 6712
rect 13538 6604 13544 6656
rect 13596 6604 13602 6656
rect 14366 6604 14372 6656
rect 14424 6604 14430 6656
rect 15010 6604 15016 6656
rect 15068 6644 15074 6656
rect 16117 6647 16175 6653
rect 16117 6644 16129 6647
rect 15068 6616 16129 6644
rect 15068 6604 15074 6616
rect 16117 6613 16129 6616
rect 16163 6644 16175 6647
rect 17218 6644 17224 6656
rect 16163 6616 17224 6644
rect 16163 6613 16175 6616
rect 16117 6607 16175 6613
rect 17218 6604 17224 6616
rect 17276 6644 17282 6656
rect 18708 6644 18736 6684
rect 19150 6672 19156 6684
rect 19208 6672 19214 6724
rect 20990 6712 20996 6724
rect 19812 6684 20996 6712
rect 17276 6616 18736 6644
rect 19429 6647 19487 6653
rect 17276 6604 17282 6616
rect 19429 6613 19441 6647
rect 19475 6644 19487 6647
rect 19812 6644 19840 6684
rect 20990 6672 20996 6684
rect 21048 6672 21054 6724
rect 22005 6715 22063 6721
rect 22005 6681 22017 6715
rect 22051 6712 22063 6715
rect 22830 6712 22836 6724
rect 22051 6684 22836 6712
rect 22051 6681 22063 6684
rect 22005 6675 22063 6681
rect 22830 6672 22836 6684
rect 22888 6672 22894 6724
rect 25041 6715 25099 6721
rect 25041 6712 25053 6715
rect 23676 6684 25053 6712
rect 19475 6616 19840 6644
rect 19475 6613 19487 6616
rect 19429 6607 19487 6613
rect 19886 6604 19892 6656
rect 19944 6644 19950 6656
rect 21174 6644 21180 6656
rect 19944 6616 21180 6644
rect 19944 6604 19950 6616
rect 21174 6604 21180 6616
rect 21232 6604 21238 6656
rect 21358 6604 21364 6656
rect 21416 6644 21422 6656
rect 23676 6644 23704 6684
rect 25041 6681 25053 6684
rect 25087 6681 25099 6715
rect 25041 6675 25099 6681
rect 21416 6616 23704 6644
rect 21416 6604 21422 6616
rect 24578 6604 24584 6656
rect 24636 6604 24642 6656
rect 24670 6604 24676 6656
rect 24728 6644 24734 6656
rect 24949 6647 25007 6653
rect 24949 6644 24961 6647
rect 24728 6616 24961 6644
rect 24728 6604 24734 6616
rect 24949 6613 24961 6616
rect 24995 6613 25007 6647
rect 24949 6607 25007 6613
rect 1104 6554 25852 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 25852 6554
rect 1104 6480 25852 6502
rect 10413 6443 10471 6449
rect 10413 6409 10425 6443
rect 10459 6440 10471 6443
rect 11422 6440 11428 6452
rect 10459 6412 11428 6440
rect 10459 6409 10471 6412
rect 10413 6403 10471 6409
rect 11422 6400 11428 6412
rect 11480 6400 11486 6452
rect 11701 6443 11759 6449
rect 11701 6409 11713 6443
rect 11747 6440 11759 6443
rect 13354 6440 13360 6452
rect 11747 6412 13360 6440
rect 11747 6409 11759 6412
rect 11701 6403 11759 6409
rect 13354 6400 13360 6412
rect 13412 6400 13418 6452
rect 13814 6400 13820 6452
rect 13872 6400 13878 6452
rect 14366 6400 14372 6452
rect 14424 6440 14430 6452
rect 20806 6440 20812 6452
rect 14424 6412 20812 6440
rect 14424 6400 14430 6412
rect 20806 6400 20812 6412
rect 20864 6400 20870 6452
rect 21836 6412 22048 6440
rect 12713 6375 12771 6381
rect 12713 6372 12725 6375
rect 12268 6344 12725 6372
rect 6362 6264 6368 6316
rect 6420 6304 6426 6316
rect 10781 6307 10839 6313
rect 10781 6304 10793 6307
rect 6420 6276 10793 6304
rect 6420 6264 6426 6276
rect 10781 6273 10793 6276
rect 10827 6273 10839 6307
rect 10781 6267 10839 6273
rect 12066 6264 12072 6316
rect 12124 6264 12130 6316
rect 12161 6307 12219 6313
rect 12161 6273 12173 6307
rect 12207 6304 12219 6307
rect 12268 6304 12296 6344
rect 12713 6341 12725 6344
rect 12759 6372 12771 6375
rect 13262 6372 13268 6384
rect 12759 6344 13268 6372
rect 12759 6341 12771 6344
rect 12713 6335 12771 6341
rect 13262 6332 13268 6344
rect 13320 6332 13326 6384
rect 13538 6332 13544 6384
rect 13596 6372 13602 6384
rect 13596 6344 18276 6372
rect 13596 6332 13602 6344
rect 13725 6307 13783 6313
rect 13725 6304 13737 6307
rect 12207 6276 12296 6304
rect 12636 6276 13737 6304
rect 12207 6273 12219 6276
rect 12161 6267 12219 6273
rect 10870 6196 10876 6248
rect 10928 6196 10934 6248
rect 10962 6196 10968 6248
rect 11020 6196 11026 6248
rect 12342 6196 12348 6248
rect 12400 6196 12406 6248
rect 8294 6060 8300 6112
rect 8352 6100 8358 6112
rect 12636 6100 12664 6276
rect 13725 6273 13737 6276
rect 13771 6273 13783 6307
rect 13725 6267 13783 6273
rect 13814 6264 13820 6316
rect 13872 6304 13878 6316
rect 14369 6307 14427 6313
rect 14369 6304 14381 6307
rect 13872 6276 14381 6304
rect 13872 6264 13878 6276
rect 14369 6273 14381 6276
rect 14415 6273 14427 6307
rect 14369 6267 14427 6273
rect 15105 6307 15163 6313
rect 15105 6273 15117 6307
rect 15151 6304 15163 6307
rect 15151 6276 16620 6304
rect 15151 6273 15163 6276
rect 15105 6267 15163 6273
rect 12894 6196 12900 6248
rect 12952 6196 12958 6248
rect 13909 6239 13967 6245
rect 13909 6205 13921 6239
rect 13955 6205 13967 6239
rect 13909 6199 13967 6205
rect 13630 6128 13636 6180
rect 13688 6168 13694 6180
rect 13924 6168 13952 6199
rect 16114 6196 16120 6248
rect 16172 6196 16178 6248
rect 13688 6140 13952 6168
rect 16592 6168 16620 6276
rect 17310 6264 17316 6316
rect 17368 6304 17374 6316
rect 18248 6313 18276 6344
rect 19242 6332 19248 6384
rect 19300 6372 19306 6384
rect 21836 6372 21864 6412
rect 19300 6344 21864 6372
rect 22020 6372 22048 6412
rect 22186 6400 22192 6452
rect 22244 6440 22250 6452
rect 22370 6440 22376 6452
rect 22244 6412 22376 6440
rect 22244 6400 22250 6412
rect 22370 6400 22376 6412
rect 22428 6400 22434 6452
rect 24578 6440 24584 6452
rect 22480 6412 24584 6440
rect 22480 6372 22508 6412
rect 24578 6400 24584 6412
rect 24636 6400 24642 6452
rect 24857 6443 24915 6449
rect 24857 6409 24869 6443
rect 24903 6440 24915 6443
rect 25222 6440 25228 6452
rect 24903 6412 25228 6440
rect 24903 6409 24915 6412
rect 24857 6403 24915 6409
rect 25222 6400 25228 6412
rect 25280 6400 25286 6452
rect 22020 6344 22508 6372
rect 23506 6344 23980 6372
rect 19300 6332 19306 6344
rect 17589 6307 17647 6313
rect 17589 6304 17601 6307
rect 17368 6276 17601 6304
rect 17368 6264 17374 6276
rect 17589 6273 17601 6276
rect 17635 6273 17647 6307
rect 17589 6267 17647 6273
rect 18233 6307 18291 6313
rect 18233 6273 18245 6307
rect 18279 6273 18291 6307
rect 18233 6267 18291 6273
rect 18322 6264 18328 6316
rect 18380 6304 18386 6316
rect 19886 6304 19892 6316
rect 18380 6276 19892 6304
rect 18380 6264 18386 6276
rect 19886 6264 19892 6276
rect 19944 6264 19950 6316
rect 20254 6264 20260 6316
rect 20312 6264 20318 6316
rect 21818 6264 21824 6316
rect 21876 6304 21882 6316
rect 22005 6308 22063 6313
rect 21928 6307 22063 6308
rect 21928 6304 22017 6307
rect 21876 6280 22017 6304
rect 21876 6276 21956 6280
rect 21876 6264 21882 6276
rect 22005 6273 22017 6280
rect 22051 6273 22063 6307
rect 23842 6304 23848 6316
rect 22005 6267 22063 6273
rect 23676 6276 23848 6304
rect 16850 6196 16856 6248
rect 16908 6196 16914 6248
rect 19429 6239 19487 6245
rect 19429 6205 19441 6239
rect 19475 6236 19487 6239
rect 21269 6239 21327 6245
rect 19475 6208 21220 6236
rect 19475 6205 19487 6208
rect 19429 6199 19487 6205
rect 20622 6168 20628 6180
rect 16592 6140 20628 6168
rect 13688 6128 13694 6140
rect 20622 6128 20628 6140
rect 20680 6128 20686 6180
rect 21192 6168 21220 6208
rect 21269 6205 21281 6239
rect 21315 6236 21327 6239
rect 21726 6236 21732 6248
rect 21315 6208 21732 6236
rect 21315 6205 21327 6208
rect 21269 6199 21327 6205
rect 21726 6196 21732 6208
rect 21784 6196 21790 6248
rect 22281 6239 22339 6245
rect 22281 6205 22293 6239
rect 22327 6236 22339 6239
rect 23676 6236 23704 6276
rect 23842 6264 23848 6276
rect 23900 6264 23906 6316
rect 23952 6304 23980 6344
rect 24210 6332 24216 6384
rect 24268 6332 24274 6384
rect 24762 6304 24768 6316
rect 23952 6276 24768 6304
rect 24762 6264 24768 6276
rect 24820 6264 24826 6316
rect 25038 6264 25044 6316
rect 25096 6264 25102 6316
rect 22327 6208 23704 6236
rect 22327 6205 22339 6208
rect 22281 6199 22339 6205
rect 23750 6196 23756 6248
rect 23808 6196 23814 6248
rect 22002 6168 22008 6180
rect 21192 6140 22008 6168
rect 22002 6128 22008 6140
rect 22060 6128 22066 6180
rect 8352 6072 12664 6100
rect 8352 6060 8358 6072
rect 13354 6060 13360 6112
rect 13412 6060 13418 6112
rect 16390 6060 16396 6112
rect 16448 6100 16454 6112
rect 17586 6100 17592 6112
rect 16448 6072 17592 6100
rect 16448 6060 16454 6072
rect 17586 6060 17592 6072
rect 17644 6060 17650 6112
rect 17681 6103 17739 6109
rect 17681 6069 17693 6103
rect 17727 6100 17739 6103
rect 22094 6100 22100 6112
rect 17727 6072 22100 6100
rect 17727 6069 17739 6072
rect 17681 6063 17739 6069
rect 22094 6060 22100 6072
rect 22152 6060 22158 6112
rect 24762 6060 24768 6112
rect 24820 6100 24826 6112
rect 25317 6103 25375 6109
rect 25317 6100 25329 6103
rect 24820 6072 25329 6100
rect 24820 6060 24826 6072
rect 25317 6069 25329 6072
rect 25363 6069 25375 6103
rect 25317 6063 25375 6069
rect 1104 6010 25852 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 25852 6010
rect 1104 5936 25852 5958
rect 11330 5856 11336 5908
rect 11388 5896 11394 5908
rect 11793 5899 11851 5905
rect 11793 5896 11805 5899
rect 11388 5868 11805 5896
rect 11388 5856 11394 5868
rect 11793 5865 11805 5868
rect 11839 5896 11851 5899
rect 12342 5896 12348 5908
rect 11839 5868 12348 5896
rect 11839 5865 11851 5868
rect 11793 5859 11851 5865
rect 12342 5856 12348 5868
rect 12400 5856 12406 5908
rect 14734 5856 14740 5908
rect 14792 5856 14798 5908
rect 16196 5899 16254 5905
rect 16196 5865 16208 5899
rect 16242 5896 16254 5899
rect 16242 5868 17264 5896
rect 16242 5865 16254 5868
rect 16196 5859 16254 5865
rect 14918 5788 14924 5840
rect 14976 5828 14982 5840
rect 14976 5800 15332 5828
rect 14976 5788 14982 5800
rect 10321 5763 10379 5769
rect 10321 5729 10333 5763
rect 10367 5760 10379 5763
rect 10778 5760 10784 5772
rect 10367 5732 10784 5760
rect 10367 5729 10379 5732
rect 10321 5723 10379 5729
rect 10778 5720 10784 5732
rect 10836 5720 10842 5772
rect 13354 5720 13360 5772
rect 13412 5760 13418 5772
rect 15304 5769 15332 5800
rect 17236 5772 17264 5868
rect 17402 5856 17408 5908
rect 17460 5896 17466 5908
rect 17681 5899 17739 5905
rect 17681 5896 17693 5899
rect 17460 5868 17693 5896
rect 17460 5856 17466 5868
rect 17681 5865 17693 5868
rect 17727 5865 17739 5899
rect 17681 5859 17739 5865
rect 20254 5856 20260 5908
rect 20312 5896 20318 5908
rect 23845 5899 23903 5905
rect 23845 5896 23857 5899
rect 20312 5868 23857 5896
rect 20312 5856 20318 5868
rect 23845 5865 23857 5868
rect 23891 5865 23903 5899
rect 23845 5859 23903 5865
rect 18141 5831 18199 5837
rect 18141 5797 18153 5831
rect 18187 5828 18199 5831
rect 18187 5800 20576 5828
rect 18187 5797 18199 5800
rect 18141 5791 18199 5797
rect 15197 5763 15255 5769
rect 15197 5760 15209 5763
rect 13412 5732 15209 5760
rect 13412 5720 13418 5732
rect 15197 5729 15209 5732
rect 15243 5729 15255 5763
rect 15197 5723 15255 5729
rect 15289 5763 15347 5769
rect 15289 5729 15301 5763
rect 15335 5729 15347 5763
rect 16942 5760 16948 5772
rect 15289 5723 15347 5729
rect 15948 5732 16948 5760
rect 9582 5652 9588 5704
rect 9640 5692 9646 5704
rect 10045 5695 10103 5701
rect 10045 5692 10057 5695
rect 9640 5664 10057 5692
rect 9640 5652 9646 5664
rect 10045 5661 10057 5664
rect 10091 5661 10103 5695
rect 10045 5655 10103 5661
rect 11422 5652 11428 5704
rect 11480 5692 11486 5704
rect 12069 5695 12127 5701
rect 12069 5692 12081 5695
rect 11480 5664 12081 5692
rect 11480 5652 11486 5664
rect 12069 5661 12081 5664
rect 12115 5661 12127 5695
rect 12069 5655 12127 5661
rect 13446 5652 13452 5704
rect 13504 5692 13510 5704
rect 13725 5695 13783 5701
rect 13725 5692 13737 5695
rect 13504 5664 13737 5692
rect 13504 5652 13510 5664
rect 13725 5661 13737 5664
rect 13771 5661 13783 5695
rect 13725 5655 13783 5661
rect 14461 5695 14519 5701
rect 14461 5661 14473 5695
rect 14507 5692 14519 5695
rect 15010 5692 15016 5704
rect 14507 5664 15016 5692
rect 14507 5661 14519 5664
rect 14461 5655 14519 5661
rect 15010 5652 15016 5664
rect 15068 5652 15074 5704
rect 15102 5652 15108 5704
rect 15160 5692 15166 5704
rect 15948 5701 15976 5732
rect 16942 5720 16948 5732
rect 17000 5720 17006 5772
rect 17218 5720 17224 5772
rect 17276 5760 17282 5772
rect 18693 5763 18751 5769
rect 18693 5760 18705 5763
rect 17276 5732 18705 5760
rect 17276 5720 17282 5732
rect 18693 5729 18705 5732
rect 18739 5729 18751 5763
rect 18693 5723 18751 5729
rect 19334 5720 19340 5772
rect 19392 5760 19398 5772
rect 19889 5763 19947 5769
rect 19889 5760 19901 5763
rect 19392 5732 19901 5760
rect 19392 5720 19398 5732
rect 19889 5729 19901 5732
rect 19935 5729 19947 5763
rect 19889 5723 19947 5729
rect 15933 5695 15991 5701
rect 15933 5692 15945 5695
rect 15160 5664 15945 5692
rect 15160 5652 15166 5664
rect 15933 5661 15945 5664
rect 15979 5661 15991 5695
rect 15933 5655 15991 5661
rect 17310 5652 17316 5704
rect 17368 5652 17374 5704
rect 17586 5652 17592 5704
rect 17644 5692 17650 5704
rect 18601 5695 18659 5701
rect 18601 5692 18613 5695
rect 17644 5664 18613 5692
rect 17644 5652 17650 5664
rect 18601 5661 18613 5664
rect 18647 5661 18659 5695
rect 18601 5655 18659 5661
rect 19610 5652 19616 5704
rect 19668 5652 19674 5704
rect 11698 5584 11704 5636
rect 11756 5624 11762 5636
rect 15746 5624 15752 5636
rect 11756 5596 15752 5624
rect 11756 5584 11762 5596
rect 15746 5584 15752 5596
rect 15804 5584 15810 5636
rect 20548 5624 20576 5800
rect 20622 5788 20628 5840
rect 20680 5828 20686 5840
rect 24857 5831 24915 5837
rect 24857 5828 24869 5831
rect 20680 5800 24869 5828
rect 20680 5788 20686 5800
rect 24857 5797 24869 5800
rect 24903 5797 24915 5831
rect 24857 5791 24915 5797
rect 20714 5720 20720 5772
rect 20772 5760 20778 5772
rect 21729 5763 21787 5769
rect 21729 5760 21741 5763
rect 20772 5732 21741 5760
rect 20772 5720 20778 5732
rect 21729 5729 21741 5732
rect 21775 5729 21787 5763
rect 21729 5723 21787 5729
rect 23566 5720 23572 5772
rect 23624 5760 23630 5772
rect 23624 5732 24716 5760
rect 23624 5720 23630 5732
rect 21082 5652 21088 5704
rect 21140 5692 21146 5704
rect 21269 5695 21327 5701
rect 21269 5692 21281 5695
rect 21140 5664 21281 5692
rect 21140 5652 21146 5664
rect 21269 5661 21281 5664
rect 21315 5661 21327 5695
rect 21269 5655 21327 5661
rect 22738 5652 22744 5704
rect 22796 5692 22802 5704
rect 23201 5695 23259 5701
rect 23201 5692 23213 5695
rect 22796 5664 23213 5692
rect 22796 5652 22802 5664
rect 23201 5661 23213 5664
rect 23247 5661 23259 5695
rect 23201 5655 23259 5661
rect 23658 5652 23664 5704
rect 23716 5692 23722 5704
rect 24688 5701 24716 5732
rect 24029 5695 24087 5701
rect 24029 5692 24041 5695
rect 23716 5664 24041 5692
rect 23716 5652 23722 5664
rect 24029 5661 24041 5664
rect 24075 5661 24087 5695
rect 24029 5655 24087 5661
rect 24673 5695 24731 5701
rect 24673 5661 24685 5695
rect 24719 5661 24731 5695
rect 24673 5655 24731 5661
rect 23385 5627 23443 5633
rect 20548 5596 22094 5624
rect 13538 5516 13544 5568
rect 13596 5516 13602 5568
rect 15105 5559 15163 5565
rect 15105 5525 15117 5559
rect 15151 5556 15163 5559
rect 16850 5556 16856 5568
rect 15151 5528 16856 5556
rect 15151 5525 15163 5528
rect 15105 5519 15163 5525
rect 16850 5516 16856 5528
rect 16908 5516 16914 5568
rect 18322 5516 18328 5568
rect 18380 5556 18386 5568
rect 18509 5559 18567 5565
rect 18509 5556 18521 5559
rect 18380 5528 18521 5556
rect 18380 5516 18386 5528
rect 18509 5525 18521 5528
rect 18555 5525 18567 5559
rect 22066 5556 22094 5596
rect 23385 5593 23397 5627
rect 23431 5624 23443 5627
rect 23750 5624 23756 5636
rect 23431 5596 23756 5624
rect 23431 5593 23443 5596
rect 23385 5587 23443 5593
rect 23750 5584 23756 5596
rect 23808 5584 23814 5636
rect 25130 5556 25136 5568
rect 22066 5528 25136 5556
rect 18509 5519 18567 5525
rect 25130 5516 25136 5528
rect 25188 5516 25194 5568
rect 1104 5466 25852 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 25852 5466
rect 1104 5392 25852 5414
rect 7834 5312 7840 5364
rect 7892 5352 7898 5364
rect 11238 5352 11244 5364
rect 7892 5324 11244 5352
rect 7892 5312 7898 5324
rect 11238 5312 11244 5324
rect 11296 5312 11302 5364
rect 13630 5312 13636 5364
rect 13688 5312 13694 5364
rect 18874 5312 18880 5364
rect 18932 5352 18938 5364
rect 20533 5355 20591 5361
rect 20533 5352 20545 5355
rect 18932 5324 20545 5352
rect 18932 5312 18938 5324
rect 20533 5321 20545 5324
rect 20579 5321 20591 5355
rect 20533 5315 20591 5321
rect 21174 5312 21180 5364
rect 21232 5352 21238 5364
rect 21545 5355 21603 5361
rect 21545 5352 21557 5355
rect 21232 5324 21557 5352
rect 21232 5312 21238 5324
rect 21545 5321 21557 5324
rect 21591 5321 21603 5355
rect 21545 5315 21603 5321
rect 13449 5287 13507 5293
rect 13449 5253 13461 5287
rect 13495 5284 13507 5287
rect 13648 5284 13676 5312
rect 15010 5284 15016 5296
rect 13495 5256 13676 5284
rect 14674 5256 15016 5284
rect 13495 5253 13507 5256
rect 13449 5247 13507 5253
rect 15010 5244 15016 5256
rect 15068 5284 15074 5296
rect 15470 5284 15476 5296
rect 15068 5256 15476 5284
rect 15068 5244 15074 5256
rect 15470 5244 15476 5256
rect 15528 5244 15534 5296
rect 19150 5284 19156 5296
rect 15764 5256 19156 5284
rect 15764 5225 15792 5256
rect 19150 5244 19156 5256
rect 19208 5244 19214 5296
rect 20346 5284 20352 5296
rect 20286 5256 20352 5284
rect 20346 5244 20352 5256
rect 20404 5244 20410 5296
rect 20438 5244 20444 5296
rect 20496 5284 20502 5296
rect 22925 5287 22983 5293
rect 22925 5284 22937 5287
rect 20496 5256 22937 5284
rect 20496 5244 20502 5256
rect 22925 5253 22937 5256
rect 22971 5253 22983 5287
rect 22925 5247 22983 5253
rect 15749 5219 15807 5225
rect 15749 5185 15761 5219
rect 15795 5185 15807 5219
rect 15749 5179 15807 5185
rect 17129 5219 17187 5225
rect 17129 5185 17141 5219
rect 17175 5216 17187 5219
rect 17175 5188 18460 5216
rect 17175 5185 17187 5188
rect 17129 5179 17187 5185
rect 11054 5108 11060 5160
rect 11112 5148 11118 5160
rect 13173 5151 13231 5157
rect 13173 5148 13185 5151
rect 11112 5120 13185 5148
rect 11112 5108 11118 5120
rect 13173 5117 13185 5120
rect 13219 5117 13231 5151
rect 13173 5111 13231 5117
rect 15473 5151 15531 5157
rect 15473 5117 15485 5151
rect 15519 5117 15531 5151
rect 15473 5111 15531 5117
rect 13188 5012 13216 5111
rect 15488 5080 15516 5111
rect 18138 5108 18144 5160
rect 18196 5108 18202 5160
rect 17954 5080 17960 5092
rect 15488 5052 17960 5080
rect 17954 5040 17960 5052
rect 18012 5040 18018 5092
rect 13906 5012 13912 5024
rect 13188 4984 13912 5012
rect 13906 4972 13912 4984
rect 13964 4972 13970 5024
rect 14182 4972 14188 5024
rect 14240 5012 14246 5024
rect 14918 5012 14924 5024
rect 14240 4984 14924 5012
rect 14240 4972 14246 4984
rect 14918 4972 14924 4984
rect 14976 4972 14982 5024
rect 18432 5012 18460 5188
rect 18506 5176 18512 5228
rect 18564 5216 18570 5228
rect 18785 5219 18843 5225
rect 18785 5216 18797 5219
rect 18564 5188 18797 5216
rect 18564 5176 18570 5188
rect 18785 5185 18797 5188
rect 18831 5185 18843 5219
rect 18785 5179 18843 5185
rect 21082 5176 21088 5228
rect 21140 5176 21146 5228
rect 22094 5176 22100 5228
rect 22152 5176 22158 5228
rect 23750 5176 23756 5228
rect 23808 5216 23814 5228
rect 23845 5219 23903 5225
rect 23845 5216 23857 5219
rect 23808 5188 23857 5216
rect 23808 5176 23814 5188
rect 23845 5185 23857 5188
rect 23891 5185 23903 5219
rect 23845 5179 23903 5185
rect 19061 5151 19119 5157
rect 19061 5117 19073 5151
rect 19107 5148 19119 5151
rect 21174 5148 21180 5160
rect 19107 5120 21180 5148
rect 19107 5117 19119 5120
rect 19061 5111 19119 5117
rect 21174 5108 21180 5120
rect 21232 5108 21238 5160
rect 21358 5108 21364 5160
rect 21416 5148 21422 5160
rect 24305 5151 24363 5157
rect 21416 5120 22876 5148
rect 21416 5108 21422 5120
rect 21269 5083 21327 5089
rect 21269 5049 21281 5083
rect 21315 5080 21327 5083
rect 22848 5080 22876 5120
rect 24305 5117 24317 5151
rect 24351 5117 24363 5151
rect 24305 5111 24363 5117
rect 24320 5080 24348 5111
rect 21315 5052 22094 5080
rect 22848 5052 24348 5080
rect 21315 5049 21327 5052
rect 21269 5043 21327 5049
rect 20438 5012 20444 5024
rect 18432 4984 20444 5012
rect 20438 4972 20444 4984
rect 20496 4972 20502 5024
rect 22066 5012 22094 5052
rect 23842 5012 23848 5024
rect 22066 4984 23848 5012
rect 23842 4972 23848 4984
rect 23900 4972 23906 5024
rect 1104 4922 25852 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 25852 4922
rect 1104 4848 25852 4870
rect 16853 4811 16911 4817
rect 12452 4780 16804 4808
rect 12250 4700 12256 4752
rect 12308 4700 12314 4752
rect 5077 4675 5135 4681
rect 5077 4641 5089 4675
rect 5123 4672 5135 4675
rect 9582 4672 9588 4684
rect 5123 4644 9588 4672
rect 5123 4641 5135 4644
rect 5077 4635 5135 4641
rect 9582 4632 9588 4644
rect 9640 4632 9646 4684
rect 7377 4607 7435 4613
rect 7377 4604 7389 4607
rect 6486 4576 7389 4604
rect 7377 4573 7389 4576
rect 7423 4604 7435 4607
rect 11422 4604 11428 4616
rect 7423 4576 11428 4604
rect 7423 4573 7435 4576
rect 7377 4567 7435 4573
rect 11422 4564 11428 4576
rect 11480 4564 11486 4616
rect 12452 4613 12480 4780
rect 12618 4700 12624 4752
rect 12676 4740 12682 4752
rect 14461 4743 14519 4749
rect 14461 4740 14473 4743
rect 12676 4712 14473 4740
rect 12676 4700 12682 4712
rect 14461 4709 14473 4712
rect 14507 4709 14519 4743
rect 16776 4740 16804 4780
rect 16853 4777 16865 4811
rect 16899 4808 16911 4811
rect 17218 4808 17224 4820
rect 16899 4780 17224 4808
rect 16899 4777 16911 4780
rect 16853 4771 16911 4777
rect 17218 4768 17224 4780
rect 17276 4768 17282 4820
rect 19058 4768 19064 4820
rect 19116 4808 19122 4820
rect 21082 4808 21088 4820
rect 19116 4780 21088 4808
rect 19116 4768 19122 4780
rect 21082 4768 21088 4780
rect 21140 4768 21146 4820
rect 21174 4768 21180 4820
rect 21232 4808 21238 4820
rect 21269 4811 21327 4817
rect 21269 4808 21281 4811
rect 21232 4780 21281 4808
rect 21232 4768 21238 4780
rect 21269 4777 21281 4780
rect 21315 4777 21327 4811
rect 21269 4771 21327 4777
rect 24026 4768 24032 4820
rect 24084 4808 24090 4820
rect 24765 4811 24823 4817
rect 24765 4808 24777 4811
rect 24084 4780 24777 4808
rect 24084 4768 24090 4780
rect 24765 4777 24777 4780
rect 24811 4777 24823 4811
rect 24765 4771 24823 4777
rect 17310 4740 17316 4752
rect 14461 4703 14519 4709
rect 14660 4712 15240 4740
rect 16776 4712 17316 4740
rect 13173 4675 13231 4681
rect 13173 4641 13185 4675
rect 13219 4672 13231 4675
rect 13814 4672 13820 4684
rect 13219 4644 13820 4672
rect 13219 4641 13231 4644
rect 13173 4635 13231 4641
rect 13814 4632 13820 4644
rect 13872 4632 13878 4684
rect 14660 4613 14688 4712
rect 15102 4632 15108 4684
rect 15160 4632 15166 4684
rect 15212 4672 15240 4712
rect 17310 4700 17316 4712
rect 17368 4700 17374 4752
rect 17402 4672 17408 4684
rect 15212 4644 17408 4672
rect 17402 4632 17408 4644
rect 17460 4632 17466 4684
rect 17494 4632 17500 4684
rect 17552 4672 17558 4684
rect 17865 4675 17923 4681
rect 17865 4672 17877 4675
rect 17552 4644 17877 4672
rect 17552 4632 17558 4644
rect 17865 4641 17877 4644
rect 17911 4641 17923 4675
rect 17865 4635 17923 4641
rect 18506 4632 18512 4684
rect 18564 4672 18570 4684
rect 19521 4675 19579 4681
rect 19521 4672 19533 4675
rect 18564 4644 19533 4672
rect 18564 4632 18570 4644
rect 19521 4641 19533 4644
rect 19567 4641 19579 4675
rect 19521 4635 19579 4641
rect 19794 4632 19800 4684
rect 19852 4632 19858 4684
rect 19886 4632 19892 4684
rect 19944 4672 19950 4684
rect 22189 4675 22247 4681
rect 22189 4672 22201 4675
rect 19944 4644 22201 4672
rect 19944 4632 19950 4644
rect 22189 4641 22201 4644
rect 22235 4641 22247 4675
rect 22189 4635 22247 4641
rect 22370 4632 22376 4684
rect 22428 4632 22434 4684
rect 12437 4607 12495 4613
rect 12437 4573 12449 4607
rect 12483 4573 12495 4607
rect 12437 4567 12495 4573
rect 12897 4607 12955 4613
rect 12897 4573 12909 4607
rect 12943 4573 12955 4607
rect 12897 4567 12955 4573
rect 14645 4607 14703 4613
rect 14645 4573 14657 4607
rect 14691 4573 14703 4607
rect 14645 4567 14703 4573
rect 17589 4607 17647 4613
rect 17589 4573 17601 4607
rect 17635 4573 17647 4607
rect 17589 4567 17647 4573
rect 21913 4607 21971 4613
rect 21913 4573 21925 4607
rect 21959 4604 21971 4607
rect 22388 4604 22416 4632
rect 21959 4576 22416 4604
rect 23661 4607 23719 4613
rect 21959 4573 21971 4576
rect 21913 4567 21971 4573
rect 23661 4573 23673 4607
rect 23707 4604 23719 4607
rect 24302 4604 24308 4616
rect 23707 4576 24308 4604
rect 23707 4573 23719 4576
rect 23661 4567 23719 4573
rect 5350 4496 5356 4548
rect 5408 4496 5414 4548
rect 7098 4496 7104 4548
rect 7156 4496 7162 4548
rect 12912 4536 12940 4567
rect 15102 4536 15108 4548
rect 12912 4508 15108 4536
rect 15102 4496 15108 4508
rect 15160 4496 15166 4548
rect 15378 4496 15384 4548
rect 15436 4496 15442 4548
rect 15470 4496 15476 4548
rect 15528 4536 15534 4548
rect 15838 4536 15844 4548
rect 15528 4508 15844 4536
rect 15528 4496 15534 4508
rect 15838 4496 15844 4508
rect 15896 4496 15902 4548
rect 17604 4536 17632 4567
rect 24302 4564 24308 4576
rect 24360 4564 24366 4616
rect 24486 4564 24492 4616
rect 24544 4604 24550 4616
rect 24673 4607 24731 4613
rect 24673 4604 24685 4607
rect 24544 4576 24685 4604
rect 24544 4564 24550 4576
rect 24673 4573 24685 4576
rect 24719 4573 24731 4607
rect 24673 4567 24731 4573
rect 19518 4536 19524 4548
rect 17604 4508 19524 4536
rect 19518 4496 19524 4508
rect 19576 4496 19582 4548
rect 20346 4496 20352 4548
rect 20404 4496 20410 4548
rect 1486 4428 1492 4480
rect 1544 4428 1550 4480
rect 11146 4428 11152 4480
rect 11204 4468 11210 4480
rect 11241 4471 11299 4477
rect 11241 4468 11253 4471
rect 11204 4440 11253 4468
rect 11204 4428 11210 4440
rect 11241 4437 11253 4440
rect 11287 4437 11299 4471
rect 11241 4431 11299 4437
rect 14185 4471 14243 4477
rect 14185 4437 14197 4471
rect 14231 4468 14243 4471
rect 14918 4468 14924 4480
rect 14231 4440 14924 4468
rect 14231 4437 14243 4440
rect 14185 4431 14243 4437
rect 14918 4428 14924 4440
rect 14976 4468 14982 4480
rect 15488 4468 15516 4496
rect 14976 4440 15516 4468
rect 14976 4428 14982 4440
rect 18138 4428 18144 4480
rect 18196 4468 18202 4480
rect 22278 4468 22284 4480
rect 18196 4440 22284 4468
rect 18196 4428 18202 4440
rect 22278 4428 22284 4440
rect 22336 4428 22342 4480
rect 23750 4428 23756 4480
rect 23808 4428 23814 4480
rect 24213 4471 24271 4477
rect 24213 4437 24225 4471
rect 24259 4468 24271 4471
rect 24762 4468 24768 4480
rect 24259 4440 24768 4468
rect 24259 4437 24271 4440
rect 24213 4431 24271 4437
rect 24762 4428 24768 4440
rect 24820 4428 24826 4480
rect 1104 4378 25852 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 25852 4378
rect 1104 4304 25852 4326
rect 11149 4267 11207 4273
rect 11149 4233 11161 4267
rect 11195 4264 11207 4267
rect 16117 4267 16175 4273
rect 11195 4236 15516 4264
rect 11195 4233 11207 4236
rect 11149 4227 11207 4233
rect 14182 4156 14188 4208
rect 14240 4156 14246 4208
rect 14918 4156 14924 4208
rect 14976 4156 14982 4208
rect 15488 4196 15516 4236
rect 16117 4233 16129 4267
rect 16163 4264 16175 4267
rect 18322 4264 18328 4276
rect 16163 4236 18328 4264
rect 16163 4233 16175 4236
rect 16117 4227 16175 4233
rect 18322 4224 18328 4236
rect 18380 4224 18386 4276
rect 20346 4224 20352 4276
rect 20404 4264 20410 4276
rect 21545 4267 21603 4273
rect 21545 4264 21557 4267
rect 20404 4236 21557 4264
rect 20404 4224 20410 4236
rect 21545 4233 21557 4236
rect 21591 4264 21603 4267
rect 21818 4264 21824 4276
rect 21591 4236 21824 4264
rect 21591 4233 21603 4236
rect 21545 4227 21603 4233
rect 21818 4224 21824 4236
rect 21876 4224 21882 4276
rect 21928 4236 22968 4264
rect 17126 4196 17132 4208
rect 15488 4168 17132 4196
rect 17126 4156 17132 4168
rect 17184 4156 17190 4208
rect 17402 4156 17408 4208
rect 17460 4196 17466 4208
rect 19610 4196 19616 4208
rect 17460 4168 19616 4196
rect 17460 4156 17466 4168
rect 19610 4156 19616 4168
rect 19668 4156 19674 4208
rect 21928 4196 21956 4236
rect 22940 4205 22968 4236
rect 22925 4199 22983 4205
rect 19720 4168 21956 4196
rect 22020 4168 22508 4196
rect 1486 4088 1492 4140
rect 1544 4128 1550 4140
rect 1765 4131 1823 4137
rect 1765 4128 1777 4131
rect 1544 4100 1777 4128
rect 1544 4088 1550 4100
rect 1765 4097 1777 4100
rect 1811 4097 1823 4131
rect 1765 4091 1823 4097
rect 1854 4088 1860 4140
rect 1912 4128 1918 4140
rect 2409 4131 2467 4137
rect 2409 4128 2421 4131
rect 1912 4100 2421 4128
rect 1912 4088 1918 4100
rect 2409 4097 2421 4100
rect 2455 4128 2467 4131
rect 2685 4131 2743 4137
rect 2685 4128 2697 4131
rect 2455 4100 2697 4128
rect 2455 4097 2467 4100
rect 2409 4091 2467 4097
rect 2685 4097 2697 4100
rect 2731 4097 2743 4131
rect 2685 4091 2743 4097
rect 4062 4088 4068 4140
rect 4120 4128 4126 4140
rect 4341 4131 4399 4137
rect 4341 4128 4353 4131
rect 4120 4100 4353 4128
rect 4120 4088 4126 4100
rect 4341 4097 4353 4100
rect 4387 4128 4399 4131
rect 4617 4131 4675 4137
rect 4617 4128 4629 4131
rect 4387 4100 4629 4128
rect 4387 4097 4399 4100
rect 4341 4091 4399 4097
rect 4617 4097 4629 4100
rect 4663 4097 4675 4131
rect 4617 4091 4675 4097
rect 9214 4088 9220 4140
rect 9272 4128 9278 4140
rect 9493 4131 9551 4137
rect 9493 4128 9505 4131
rect 9272 4100 9505 4128
rect 9272 4088 9278 4100
rect 9493 4097 9505 4100
rect 9539 4128 9551 4131
rect 9769 4131 9827 4137
rect 9769 4128 9781 4131
rect 9539 4100 9781 4128
rect 9539 4097 9551 4100
rect 9493 4091 9551 4097
rect 9769 4097 9781 4100
rect 9815 4097 9827 4131
rect 9769 4091 9827 4097
rect 10873 4131 10931 4137
rect 10873 4097 10885 4131
rect 10919 4128 10931 4131
rect 10962 4128 10968 4140
rect 10919 4100 10968 4128
rect 10919 4097 10931 4100
rect 10873 4091 10931 4097
rect 10962 4088 10968 4100
rect 11020 4088 11026 4140
rect 12250 4088 12256 4140
rect 12308 4088 12314 4140
rect 13906 4088 13912 4140
rect 13964 4088 13970 4140
rect 17037 4131 17095 4137
rect 17037 4097 17049 4131
rect 17083 4128 17095 4131
rect 18690 4128 18696 4140
rect 17083 4100 18696 4128
rect 17083 4097 17095 4100
rect 17037 4091 17095 4097
rect 18690 4088 18696 4100
rect 18748 4088 18754 4140
rect 18782 4088 18788 4140
rect 18840 4088 18846 4140
rect 19518 4088 19524 4140
rect 19576 4128 19582 4140
rect 19720 4128 19748 4168
rect 19576 4100 19748 4128
rect 19576 4088 19582 4100
rect 20898 4088 20904 4140
rect 20956 4088 20962 4140
rect 20990 4088 20996 4140
rect 21048 4088 21054 4140
rect 21542 4128 21548 4140
rect 21100 4100 21548 4128
rect 5350 4060 5356 4072
rect 1596 4032 5356 4060
rect 1596 4001 1624 4032
rect 5350 4020 5356 4032
rect 5408 4020 5414 4072
rect 12802 4060 12808 4072
rect 9324 4032 12808 4060
rect 1581 3995 1639 4001
rect 1581 3961 1593 3995
rect 1627 3961 1639 3995
rect 1581 3955 1639 3961
rect 2222 3952 2228 4004
rect 2280 3952 2286 4004
rect 4157 3995 4215 4001
rect 4157 3961 4169 3995
rect 4203 3992 4215 3995
rect 6914 3992 6920 4004
rect 4203 3964 6920 3992
rect 4203 3961 4215 3964
rect 4157 3955 4215 3961
rect 6914 3952 6920 3964
rect 6972 3952 6978 4004
rect 9324 4001 9352 4032
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 13265 4063 13323 4069
rect 13265 4029 13277 4063
rect 13311 4060 13323 4063
rect 16022 4060 16028 4072
rect 13311 4032 16028 4060
rect 13311 4029 13323 4032
rect 13265 4023 13323 4029
rect 16022 4020 16028 4032
rect 16080 4020 16086 4072
rect 16206 4020 16212 4072
rect 16264 4060 16270 4072
rect 17313 4063 17371 4069
rect 17313 4060 17325 4063
rect 16264 4032 17325 4060
rect 16264 4020 16270 4032
rect 17313 4029 17325 4032
rect 17359 4029 17371 4063
rect 17313 4023 17371 4029
rect 18322 4020 18328 4072
rect 18380 4060 18386 4072
rect 19153 4063 19211 4069
rect 19153 4060 19165 4063
rect 18380 4032 19165 4060
rect 18380 4020 18386 4032
rect 19153 4029 19165 4032
rect 19199 4029 19211 4063
rect 19153 4023 19211 4029
rect 20530 4020 20536 4072
rect 20588 4060 20594 4072
rect 21100 4060 21128 4100
rect 21542 4088 21548 4100
rect 21600 4088 21606 4140
rect 22020 4137 22048 4168
rect 22005 4131 22063 4137
rect 22005 4097 22017 4131
rect 22051 4097 22063 4131
rect 22005 4091 22063 4097
rect 22094 4088 22100 4140
rect 22152 4128 22158 4140
rect 22370 4128 22376 4140
rect 22152 4100 22376 4128
rect 22152 4088 22158 4100
rect 22370 4088 22376 4100
rect 22428 4088 22434 4140
rect 22480 4128 22508 4168
rect 22925 4165 22937 4199
rect 22971 4165 22983 4199
rect 22925 4159 22983 4165
rect 22480 4100 23060 4128
rect 20588 4032 21128 4060
rect 20588 4020 20594 4032
rect 21174 4020 21180 4072
rect 21232 4020 21238 4072
rect 23032 4060 23060 4100
rect 23842 4088 23848 4140
rect 23900 4088 23906 4140
rect 25406 4128 25412 4140
rect 23952 4100 25412 4128
rect 23952 4060 23980 4100
rect 25406 4088 25412 4100
rect 25464 4088 25470 4140
rect 23032 4032 23980 4060
rect 24305 4063 24363 4069
rect 24305 4029 24317 4063
rect 24351 4029 24363 4063
rect 24305 4023 24363 4029
rect 9309 3995 9367 4001
rect 9309 3961 9321 3995
rect 9355 3961 9367 3995
rect 9309 3955 9367 3961
rect 9398 3952 9404 4004
rect 9456 3992 9462 4004
rect 12434 3992 12440 4004
rect 9456 3964 12440 3992
rect 9456 3952 9462 3964
rect 12434 3952 12440 3964
rect 12492 3952 12498 4004
rect 15470 3952 15476 4004
rect 15528 3992 15534 4004
rect 15657 3995 15715 4001
rect 15657 3992 15669 3995
rect 15528 3964 15669 3992
rect 15528 3952 15534 3964
rect 15657 3961 15669 3964
rect 15703 3961 15715 3995
rect 15657 3955 15715 3961
rect 20990 3952 20996 4004
rect 21048 3992 21054 4004
rect 21048 3964 22508 3992
rect 21048 3952 21054 3964
rect 2866 3884 2872 3936
rect 2924 3884 2930 3936
rect 10594 3884 10600 3936
rect 10652 3884 10658 3936
rect 11606 3884 11612 3936
rect 11664 3884 11670 3936
rect 11793 3927 11851 3933
rect 11793 3893 11805 3927
rect 11839 3924 11851 3927
rect 12526 3924 12532 3936
rect 11839 3896 12532 3924
rect 11839 3893 11851 3896
rect 11793 3887 11851 3893
rect 12526 3884 12532 3896
rect 12584 3884 12590 3936
rect 13354 3884 13360 3936
rect 13412 3924 13418 3936
rect 20162 3924 20168 3936
rect 13412 3896 20168 3924
rect 13412 3884 13418 3896
rect 20162 3884 20168 3896
rect 20220 3884 20226 3936
rect 20530 3884 20536 3936
rect 20588 3884 20594 3936
rect 21542 3884 21548 3936
rect 21600 3924 21606 3936
rect 22370 3924 22376 3936
rect 21600 3896 22376 3924
rect 21600 3884 21606 3896
rect 22370 3884 22376 3896
rect 22428 3884 22434 3936
rect 22480 3924 22508 3964
rect 24320 3924 24348 4023
rect 22480 3896 24348 3924
rect 1104 3834 25852 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 25852 3834
rect 1104 3760 25852 3782
rect 2869 3723 2927 3729
rect 2869 3689 2881 3723
rect 2915 3720 2927 3723
rect 3326 3720 3332 3732
rect 2915 3692 3332 3720
rect 2915 3689 2927 3692
rect 2869 3683 2927 3689
rect 3326 3680 3332 3692
rect 3384 3680 3390 3732
rect 4249 3723 4307 3729
rect 4249 3689 4261 3723
rect 4295 3720 4307 3723
rect 7650 3720 7656 3732
rect 4295 3692 7656 3720
rect 4295 3689 4307 3692
rect 4249 3683 4307 3689
rect 7650 3680 7656 3692
rect 7708 3680 7714 3732
rect 8389 3723 8447 3729
rect 8389 3689 8401 3723
rect 8435 3720 8447 3723
rect 10870 3720 10876 3732
rect 8435 3692 10876 3720
rect 8435 3689 8447 3692
rect 8389 3683 8447 3689
rect 10870 3680 10876 3692
rect 10928 3680 10934 3732
rect 10962 3680 10968 3732
rect 11020 3720 11026 3732
rect 15930 3720 15936 3732
rect 11020 3692 15936 3720
rect 11020 3680 11026 3692
rect 15930 3680 15936 3692
rect 15988 3680 15994 3732
rect 17954 3680 17960 3732
rect 18012 3680 18018 3732
rect 18785 3723 18843 3729
rect 18785 3689 18797 3723
rect 18831 3720 18843 3723
rect 22094 3720 22100 3732
rect 18831 3692 22100 3720
rect 18831 3689 18843 3692
rect 18785 3683 18843 3689
rect 22094 3680 22100 3692
rect 22152 3680 22158 3732
rect 22738 3680 22744 3732
rect 22796 3720 22802 3732
rect 23109 3723 23167 3729
rect 23109 3720 23121 3723
rect 22796 3692 23121 3720
rect 22796 3680 22802 3692
rect 23109 3689 23121 3692
rect 23155 3689 23167 3723
rect 23109 3683 23167 3689
rect 6362 3612 6368 3664
rect 6420 3612 6426 3664
rect 7101 3655 7159 3661
rect 7101 3621 7113 3655
rect 7147 3652 7159 3655
rect 9398 3652 9404 3664
rect 7147 3624 9404 3652
rect 7147 3621 7159 3624
rect 7101 3615 7159 3621
rect 9398 3612 9404 3624
rect 9456 3612 9462 3664
rect 12710 3652 12716 3664
rect 9508 3624 12716 3652
rect 1581 3587 1639 3593
rect 1581 3553 1593 3587
rect 1627 3584 1639 3587
rect 2866 3584 2872 3596
rect 1627 3556 2872 3584
rect 1627 3553 1639 3556
rect 1581 3547 1639 3553
rect 2866 3544 2872 3556
rect 2924 3584 2930 3596
rect 3694 3584 3700 3596
rect 2924 3556 3700 3584
rect 2924 3544 2930 3556
rect 3694 3544 3700 3556
rect 3752 3544 3758 3596
rect 5166 3544 5172 3596
rect 5224 3544 5230 3596
rect 5442 3544 5448 3596
rect 5500 3584 5506 3596
rect 9508 3584 9536 3624
rect 12710 3612 12716 3624
rect 12768 3612 12774 3664
rect 16022 3612 16028 3664
rect 16080 3652 16086 3664
rect 23474 3652 23480 3664
rect 16080 3624 23480 3652
rect 16080 3612 16086 3624
rect 23474 3612 23480 3624
rect 23532 3612 23538 3664
rect 24946 3612 24952 3664
rect 25004 3612 25010 3664
rect 5500 3556 9536 3584
rect 11057 3587 11115 3593
rect 5500 3544 5506 3556
rect 11057 3553 11069 3587
rect 11103 3584 11115 3587
rect 12526 3584 12532 3596
rect 11103 3556 12532 3584
rect 11103 3553 11115 3556
rect 11057 3547 11115 3553
rect 12526 3544 12532 3556
rect 12584 3544 12590 3596
rect 12802 3544 12808 3596
rect 12860 3544 12866 3596
rect 13998 3544 14004 3596
rect 14056 3584 14062 3596
rect 14737 3587 14795 3593
rect 14737 3584 14749 3587
rect 14056 3556 14749 3584
rect 14056 3544 14062 3556
rect 14737 3553 14749 3556
rect 14783 3553 14795 3587
rect 14737 3547 14795 3553
rect 15470 3544 15476 3596
rect 15528 3584 15534 3596
rect 16577 3587 16635 3593
rect 16577 3584 16589 3587
rect 15528 3556 16589 3584
rect 15528 3544 15534 3556
rect 16577 3553 16589 3556
rect 16623 3553 16635 3587
rect 16577 3547 16635 3553
rect 17678 3544 17684 3596
rect 17736 3584 17742 3596
rect 19889 3587 19947 3593
rect 19889 3584 19901 3587
rect 17736 3556 19901 3584
rect 17736 3544 17742 3556
rect 19889 3553 19901 3556
rect 19935 3553 19947 3587
rect 19889 3547 19947 3553
rect 21729 3587 21787 3593
rect 21729 3553 21741 3587
rect 21775 3553 21787 3587
rect 21729 3547 21787 3553
rect 23845 3587 23903 3593
rect 23845 3553 23857 3587
rect 23891 3584 23903 3587
rect 23934 3584 23940 3596
rect 23891 3556 23940 3584
rect 23891 3553 23903 3556
rect 23845 3547 23903 3553
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3485 1915 3519
rect 1857 3479 1915 3485
rect 1872 3448 1900 3479
rect 2222 3476 2228 3528
rect 2280 3516 2286 3528
rect 3053 3519 3111 3525
rect 3053 3516 3065 3519
rect 2280 3488 3065 3516
rect 2280 3476 2286 3488
rect 3053 3485 3065 3488
rect 3099 3516 3111 3519
rect 3513 3519 3571 3525
rect 3513 3516 3525 3519
rect 3099 3488 3525 3516
rect 3099 3485 3111 3488
rect 3053 3479 3111 3485
rect 3513 3485 3525 3488
rect 3559 3485 3571 3519
rect 3513 3479 3571 3485
rect 4430 3476 4436 3528
rect 4488 3476 4494 3528
rect 4890 3476 4896 3528
rect 4948 3476 4954 3528
rect 6089 3519 6147 3525
rect 6089 3485 6101 3519
rect 6135 3516 6147 3519
rect 6270 3516 6276 3528
rect 6135 3488 6276 3516
rect 6135 3485 6147 3488
rect 6089 3479 6147 3485
rect 6270 3476 6276 3488
rect 6328 3516 6334 3528
rect 6549 3519 6607 3525
rect 6549 3516 6561 3519
rect 6328 3488 6561 3516
rect 6328 3476 6334 3488
rect 6549 3485 6561 3488
rect 6595 3485 6607 3519
rect 6549 3479 6607 3485
rect 7006 3476 7012 3528
rect 7064 3516 7070 3528
rect 7285 3519 7343 3525
rect 7285 3516 7297 3519
rect 7064 3488 7297 3516
rect 7064 3476 7070 3488
rect 7285 3485 7297 3488
rect 7331 3516 7343 3519
rect 7745 3519 7803 3525
rect 7745 3516 7757 3519
rect 7331 3488 7757 3516
rect 7331 3485 7343 3488
rect 7285 3479 7343 3485
rect 7745 3485 7757 3488
rect 7791 3485 7803 3519
rect 7745 3479 7803 3485
rect 8478 3476 8484 3528
rect 8536 3516 8542 3528
rect 8573 3519 8631 3525
rect 8573 3516 8585 3519
rect 8536 3488 8585 3516
rect 8536 3476 8542 3488
rect 8573 3485 8585 3488
rect 8619 3516 8631 3519
rect 8941 3519 8999 3525
rect 8941 3516 8953 3519
rect 8619 3488 8953 3516
rect 8619 3485 8631 3488
rect 8573 3479 8631 3485
rect 8941 3485 8953 3488
rect 8987 3485 8999 3519
rect 8941 3479 8999 3485
rect 9401 3519 9459 3525
rect 9401 3485 9413 3519
rect 9447 3516 9459 3519
rect 9582 3516 9588 3528
rect 9447 3488 9588 3516
rect 9447 3485 9459 3488
rect 9401 3479 9459 3485
rect 9582 3476 9588 3488
rect 9640 3516 9646 3528
rect 9861 3519 9919 3525
rect 9861 3516 9873 3519
rect 9640 3488 9873 3516
rect 9640 3476 9646 3488
rect 9861 3485 9873 3488
rect 9907 3485 9919 3519
rect 9861 3479 9919 3485
rect 10594 3476 10600 3528
rect 10652 3476 10658 3528
rect 11333 3519 11391 3525
rect 11333 3485 11345 3519
rect 11379 3485 11391 3519
rect 11333 3479 11391 3485
rect 12437 3519 12495 3525
rect 12437 3485 12449 3519
rect 12483 3516 12495 3519
rect 13354 3516 13360 3528
rect 12483 3488 13360 3516
rect 12483 3485 12495 3488
rect 12437 3479 12495 3485
rect 9306 3448 9312 3460
rect 1872 3420 9312 3448
rect 9306 3408 9312 3420
rect 9364 3408 9370 3460
rect 11348 3448 11376 3479
rect 13354 3476 13360 3488
rect 13412 3476 13418 3528
rect 14458 3476 14464 3528
rect 14516 3476 14522 3528
rect 16301 3519 16359 3525
rect 16301 3485 16313 3519
rect 16347 3516 16359 3519
rect 17034 3516 17040 3528
rect 16347 3488 17040 3516
rect 16347 3485 16359 3488
rect 16301 3479 16359 3485
rect 17034 3476 17040 3488
rect 17092 3476 17098 3528
rect 18141 3519 18199 3525
rect 18141 3485 18153 3519
rect 18187 3516 18199 3519
rect 19242 3516 19248 3528
rect 18187 3488 19248 3516
rect 18187 3485 18199 3488
rect 18141 3479 18199 3485
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 19426 3476 19432 3528
rect 19484 3476 19490 3528
rect 20806 3476 20812 3528
rect 20864 3516 20870 3528
rect 21269 3519 21327 3525
rect 21269 3516 21281 3519
rect 20864 3488 21281 3516
rect 20864 3476 20870 3488
rect 21269 3485 21281 3488
rect 21315 3485 21327 3519
rect 21269 3479 21327 3485
rect 9692 3420 11100 3448
rect 11348 3420 14504 3448
rect 3418 3340 3424 3392
rect 3476 3340 3482 3392
rect 7374 3340 7380 3392
rect 7432 3380 7438 3392
rect 9692 3389 9720 3420
rect 7561 3383 7619 3389
rect 7561 3380 7573 3383
rect 7432 3352 7573 3380
rect 7432 3340 7438 3352
rect 7561 3349 7573 3352
rect 7607 3349 7619 3383
rect 7561 3343 7619 3349
rect 9677 3383 9735 3389
rect 9677 3349 9689 3383
rect 9723 3349 9735 3383
rect 9677 3343 9735 3349
rect 10410 3340 10416 3392
rect 10468 3340 10474 3392
rect 11072 3380 11100 3420
rect 14274 3380 14280 3392
rect 11072 3352 14280 3380
rect 14274 3340 14280 3352
rect 14332 3340 14338 3392
rect 14476 3380 14504 3420
rect 14550 3408 14556 3460
rect 14608 3448 14614 3460
rect 18693 3451 18751 3457
rect 18693 3448 18705 3451
rect 14608 3420 18705 3448
rect 14608 3408 14614 3420
rect 18693 3417 18705 3420
rect 18739 3417 18751 3451
rect 18693 3411 18751 3417
rect 18874 3408 18880 3460
rect 18932 3448 18938 3460
rect 21744 3448 21772 3547
rect 23934 3544 23940 3556
rect 23992 3544 23998 3596
rect 22554 3476 22560 3528
rect 22612 3516 22618 3528
rect 23293 3519 23351 3525
rect 23293 3516 23305 3519
rect 22612 3488 23305 3516
rect 22612 3476 22618 3488
rect 23293 3485 23305 3488
rect 23339 3485 23351 3519
rect 23293 3479 23351 3485
rect 25130 3476 25136 3528
rect 25188 3476 25194 3528
rect 18932 3420 21772 3448
rect 18932 3408 18938 3420
rect 21818 3408 21824 3460
rect 21876 3448 21882 3460
rect 24762 3448 24768 3460
rect 21876 3420 24768 3448
rect 21876 3408 21882 3420
rect 24762 3408 24768 3420
rect 24820 3408 24826 3460
rect 14642 3380 14648 3392
rect 14476 3352 14648 3380
rect 14642 3340 14648 3352
rect 14700 3340 14706 3392
rect 20806 3340 20812 3392
rect 20864 3380 20870 3392
rect 21266 3380 21272 3392
rect 20864 3352 21272 3380
rect 20864 3340 20870 3352
rect 21266 3340 21272 3352
rect 21324 3340 21330 3392
rect 21450 3340 21456 3392
rect 21508 3380 21514 3392
rect 22830 3380 22836 3392
rect 21508 3352 22836 3380
rect 21508 3340 21514 3352
rect 22830 3340 22836 3352
rect 22888 3340 22894 3392
rect 1104 3290 25852 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 25852 3290
rect 1104 3216 25852 3238
rect 4430 3136 4436 3188
rect 4488 3176 4494 3188
rect 4525 3179 4583 3185
rect 4525 3176 4537 3179
rect 4488 3148 4537 3176
rect 4488 3136 4494 3148
rect 4525 3145 4537 3148
rect 4571 3145 4583 3179
rect 4525 3139 4583 3145
rect 4801 3179 4859 3185
rect 4801 3145 4813 3179
rect 4847 3176 4859 3179
rect 4890 3176 4896 3188
rect 4847 3148 4896 3176
rect 4847 3145 4859 3148
rect 4801 3139 4859 3145
rect 4890 3136 4896 3148
rect 4948 3136 4954 3188
rect 6549 3179 6607 3185
rect 6549 3145 6561 3179
rect 6595 3176 6607 3179
rect 6595 3148 10640 3176
rect 6595 3145 6607 3148
rect 6549 3139 6607 3145
rect 7834 3068 7840 3120
rect 7892 3068 7898 3120
rect 9401 3111 9459 3117
rect 9401 3077 9413 3111
rect 9447 3108 9459 3111
rect 10612 3108 10640 3148
rect 10962 3136 10968 3188
rect 11020 3136 11026 3188
rect 12066 3176 12072 3188
rect 11072 3148 12072 3176
rect 11072 3108 11100 3148
rect 12066 3136 12072 3148
rect 12124 3136 12130 3188
rect 20438 3136 20444 3188
rect 20496 3176 20502 3188
rect 20625 3179 20683 3185
rect 20625 3176 20637 3179
rect 20496 3148 20637 3176
rect 20496 3136 20502 3148
rect 20625 3145 20637 3148
rect 20671 3145 20683 3179
rect 20625 3139 20683 3145
rect 20898 3136 20904 3188
rect 20956 3176 20962 3188
rect 21269 3179 21327 3185
rect 21269 3176 21281 3179
rect 20956 3148 21281 3176
rect 20956 3136 20962 3148
rect 21269 3145 21281 3148
rect 21315 3145 21327 3179
rect 21269 3139 21327 3145
rect 22741 3179 22799 3185
rect 22741 3145 22753 3179
rect 22787 3176 22799 3179
rect 24670 3176 24676 3188
rect 22787 3148 24676 3176
rect 22787 3145 22799 3148
rect 22741 3139 22799 3145
rect 24670 3136 24676 3148
rect 24728 3136 24734 3188
rect 24762 3136 24768 3188
rect 24820 3176 24826 3188
rect 24857 3179 24915 3185
rect 24857 3176 24869 3179
rect 24820 3148 24869 3176
rect 24820 3136 24826 3148
rect 24857 3145 24869 3148
rect 24903 3145 24915 3179
rect 24857 3139 24915 3145
rect 11790 3108 11796 3120
rect 9447 3080 10548 3108
rect 10612 3080 11100 3108
rect 11164 3080 11796 3108
rect 9447 3077 9459 3080
rect 9401 3071 9459 3077
rect 2133 3043 2191 3049
rect 2133 3009 2145 3043
rect 2179 3040 2191 3043
rect 2590 3040 2596 3052
rect 2179 3012 2596 3040
rect 2179 3009 2191 3012
rect 2133 3003 2191 3009
rect 2590 3000 2596 3012
rect 2648 3000 2654 3052
rect 3418 3000 3424 3052
rect 3476 3000 3482 3052
rect 3697 3043 3755 3049
rect 3697 3009 3709 3043
rect 3743 3040 3755 3043
rect 5258 3040 5264 3052
rect 3743 3012 5264 3040
rect 3743 3009 3755 3012
rect 3697 3003 3755 3009
rect 5258 3000 5264 3012
rect 5316 3000 5322 3052
rect 5442 3000 5448 3052
rect 5500 3000 5506 3052
rect 6638 3000 6644 3052
rect 6696 3040 6702 3052
rect 6733 3043 6791 3049
rect 6733 3040 6745 3043
rect 6696 3012 6745 3040
rect 6696 3000 6702 3012
rect 6733 3009 6745 3012
rect 6779 3009 6791 3043
rect 6733 3003 6791 3009
rect 7374 3000 7380 3052
rect 7432 3000 7438 3052
rect 7852 3040 7880 3068
rect 8113 3043 8171 3049
rect 8113 3040 8125 3043
rect 7852 3012 8125 3040
rect 8113 3009 8125 3012
rect 8159 3009 8171 3043
rect 8113 3003 8171 3009
rect 9217 3043 9275 3049
rect 9217 3009 9229 3043
rect 9263 3040 9275 3043
rect 9861 3043 9919 3049
rect 9861 3040 9873 3043
rect 9263 3012 9873 3040
rect 9263 3009 9275 3012
rect 9217 3003 9275 3009
rect 9861 3009 9873 3012
rect 9907 3040 9919 3043
rect 10318 3040 10324 3052
rect 9907 3012 10324 3040
rect 9907 3009 9919 3012
rect 9861 3003 9919 3009
rect 10318 3000 10324 3012
rect 10376 3000 10382 3052
rect 10520 3049 10548 3080
rect 11164 3052 11192 3080
rect 11790 3068 11796 3080
rect 11848 3068 11854 3120
rect 13906 3108 13912 3120
rect 12406 3080 13912 3108
rect 10505 3043 10563 3049
rect 10505 3009 10517 3043
rect 10551 3040 10563 3043
rect 11054 3040 11060 3052
rect 10551 3012 11060 3040
rect 10551 3009 10563 3012
rect 10505 3003 10563 3009
rect 11054 3000 11060 3012
rect 11112 3000 11118 3052
rect 11146 3000 11152 3052
rect 11204 3000 11210 3052
rect 11606 3000 11612 3052
rect 11664 3040 11670 3052
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 11664 3012 11713 3040
rect 11664 3000 11670 3012
rect 11701 3009 11713 3012
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 11977 3043 12035 3049
rect 11977 3009 11989 3043
rect 12023 3040 12035 3043
rect 12406 3040 12434 3080
rect 13906 3068 13912 3080
rect 13964 3068 13970 3120
rect 16574 3068 16580 3120
rect 16632 3108 16638 3120
rect 22097 3111 22155 3117
rect 16632 3080 19196 3108
rect 16632 3068 16638 3080
rect 12023 3012 12434 3040
rect 12023 3009 12035 3012
rect 11977 3003 12035 3009
rect 13170 3000 13176 3052
rect 13228 3000 13234 3052
rect 14090 3000 14096 3052
rect 14148 3040 14154 3052
rect 14829 3043 14887 3049
rect 14829 3040 14841 3043
rect 14148 3012 14841 3040
rect 14148 3000 14154 3012
rect 14829 3009 14841 3012
rect 14875 3009 14887 3043
rect 14829 3003 14887 3009
rect 15010 3000 15016 3052
rect 15068 3040 15074 3052
rect 15378 3040 15384 3052
rect 15068 3012 15384 3040
rect 15068 3000 15074 3012
rect 15378 3000 15384 3012
rect 15436 3000 15442 3052
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3040 17095 3043
rect 18598 3040 18604 3052
rect 17083 3012 18604 3040
rect 17083 3009 17095 3012
rect 17037 3003 17095 3009
rect 18598 3000 18604 3012
rect 18656 3000 18662 3052
rect 18877 3043 18935 3049
rect 18877 3009 18889 3043
rect 18923 3040 18935 3043
rect 18966 3040 18972 3052
rect 18923 3012 18972 3040
rect 18923 3009 18935 3012
rect 18877 3003 18935 3009
rect 18966 3000 18972 3012
rect 19024 3000 19030 3052
rect 2409 2975 2467 2981
rect 2409 2941 2421 2975
rect 2455 2941 2467 2975
rect 2409 2935 2467 2941
rect 2424 2904 2452 2935
rect 5166 2932 5172 2984
rect 5224 2932 5230 2984
rect 7742 2932 7748 2984
rect 7800 2972 7806 2984
rect 7837 2975 7895 2981
rect 7837 2972 7849 2975
rect 7800 2944 7849 2972
rect 7800 2932 7806 2944
rect 7837 2941 7849 2944
rect 7883 2941 7895 2975
rect 7837 2935 7895 2941
rect 10410 2932 10416 2984
rect 10468 2972 10474 2984
rect 10468 2944 12434 2972
rect 10468 2932 10474 2944
rect 8938 2904 8944 2916
rect 2424 2876 8944 2904
rect 8938 2864 8944 2876
rect 8996 2864 9002 2916
rect 9677 2907 9735 2913
rect 9677 2873 9689 2907
rect 9723 2904 9735 2907
rect 12406 2904 12434 2944
rect 13630 2932 13636 2984
rect 13688 2932 13694 2984
rect 14734 2932 14740 2984
rect 14792 2972 14798 2984
rect 15289 2975 15347 2981
rect 15289 2972 15301 2975
rect 14792 2944 15301 2972
rect 14792 2932 14798 2944
rect 15289 2941 15301 2944
rect 15335 2941 15347 2975
rect 15289 2935 15347 2941
rect 15838 2932 15844 2984
rect 15896 2972 15902 2984
rect 19168 2981 19196 3080
rect 22097 3077 22109 3111
rect 22143 3108 22155 3111
rect 22186 3108 22192 3120
rect 22143 3080 22192 3108
rect 22143 3077 22155 3080
rect 22097 3071 22155 3077
rect 22186 3068 22192 3080
rect 22244 3068 22250 3120
rect 20806 3000 20812 3052
rect 20864 3000 20870 3052
rect 23566 3000 23572 3052
rect 23624 3000 23630 3052
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 15896 2944 17325 2972
rect 15896 2932 15902 2944
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 19153 2975 19211 2981
rect 19153 2941 19165 2975
rect 19199 2941 19211 2975
rect 19153 2935 19211 2941
rect 20070 2932 20076 2984
rect 20128 2972 20134 2984
rect 22281 2975 22339 2981
rect 22281 2972 22293 2975
rect 20128 2944 22293 2972
rect 20128 2932 20134 2944
rect 22281 2941 22293 2944
rect 22327 2941 22339 2975
rect 22281 2935 22339 2941
rect 16298 2904 16304 2916
rect 9723 2876 11100 2904
rect 12406 2876 16304 2904
rect 9723 2873 9735 2876
rect 9677 2867 9735 2873
rect 7190 2796 7196 2848
rect 7248 2796 7254 2848
rect 9030 2796 9036 2848
rect 9088 2796 9094 2848
rect 10321 2839 10379 2845
rect 10321 2805 10333 2839
rect 10367 2836 10379 2839
rect 10502 2836 10508 2848
rect 10367 2808 10508 2836
rect 10367 2805 10379 2808
rect 10321 2799 10379 2805
rect 10502 2796 10508 2808
rect 10560 2796 10566 2848
rect 11072 2836 11100 2876
rect 16298 2864 16304 2876
rect 16356 2864 16362 2916
rect 16942 2864 16948 2916
rect 17000 2904 17006 2916
rect 20346 2904 20352 2916
rect 17000 2876 20352 2904
rect 17000 2864 17006 2876
rect 20346 2864 20352 2876
rect 20404 2864 20410 2916
rect 22094 2904 22100 2916
rect 22066 2864 22100 2904
rect 22152 2864 22158 2916
rect 15010 2836 15016 2848
rect 11072 2808 15016 2836
rect 15010 2796 15016 2808
rect 15068 2796 15074 2848
rect 15102 2796 15108 2848
rect 15160 2836 15166 2848
rect 17310 2836 17316 2848
rect 15160 2808 17316 2836
rect 15160 2796 15166 2808
rect 17310 2796 17316 2808
rect 17368 2796 17374 2848
rect 18414 2796 18420 2848
rect 18472 2836 18478 2848
rect 22066 2836 22094 2864
rect 18472 2808 22094 2836
rect 18472 2796 18478 2808
rect 1104 2746 25852 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 25852 2746
rect 1104 2672 25852 2694
rect 4525 2635 4583 2641
rect 4525 2601 4537 2635
rect 4571 2632 4583 2635
rect 11882 2632 11888 2644
rect 4571 2604 11888 2632
rect 4571 2601 4583 2604
rect 4525 2595 4583 2601
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 15194 2592 15200 2644
rect 15252 2632 15258 2644
rect 18693 2635 18751 2641
rect 18693 2632 18705 2635
rect 15252 2604 18705 2632
rect 15252 2592 15258 2604
rect 18693 2601 18705 2604
rect 18739 2601 18751 2635
rect 18693 2595 18751 2601
rect 19610 2592 19616 2644
rect 19668 2632 19674 2644
rect 21269 2635 21327 2641
rect 21269 2632 21281 2635
rect 19668 2604 21281 2632
rect 19668 2592 19674 2604
rect 21269 2601 21281 2604
rect 21315 2601 21327 2635
rect 21269 2595 21327 2601
rect 23566 2592 23572 2644
rect 23624 2632 23630 2644
rect 24302 2632 24308 2644
rect 23624 2604 24308 2632
rect 23624 2592 23630 2604
rect 24302 2592 24308 2604
rect 24360 2632 24366 2644
rect 25409 2635 25467 2641
rect 25409 2632 25421 2635
rect 24360 2604 25421 2632
rect 24360 2592 24366 2604
rect 25409 2601 25421 2604
rect 25455 2601 25467 2635
rect 25409 2595 25467 2601
rect 9674 2564 9680 2576
rect 2884 2536 9680 2564
rect 2884 2505 2912 2536
rect 9674 2524 9680 2536
rect 9732 2524 9738 2576
rect 12618 2564 12624 2576
rect 9876 2536 12624 2564
rect 2869 2499 2927 2505
rect 2869 2465 2881 2499
rect 2915 2465 2927 2499
rect 2869 2459 2927 2465
rect 5442 2456 5448 2508
rect 5500 2456 5506 2508
rect 8294 2496 8300 2508
rect 7208 2468 8300 2496
rect 2593 2431 2651 2437
rect 2593 2397 2605 2431
rect 2639 2428 2651 2431
rect 2958 2428 2964 2440
rect 2639 2400 2964 2428
rect 2639 2397 2651 2400
rect 2593 2391 2651 2397
rect 2958 2388 2964 2400
rect 3016 2428 3022 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3016 2400 3985 2428
rect 3016 2388 3022 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4709 2431 4767 2437
rect 4709 2397 4721 2431
rect 4755 2397 4767 2431
rect 4709 2391 4767 2397
rect 5169 2431 5227 2437
rect 5169 2397 5181 2431
rect 5215 2428 5227 2431
rect 5534 2428 5540 2440
rect 5215 2400 5540 2428
rect 5215 2397 5227 2400
rect 5169 2391 5227 2397
rect 4249 2363 4307 2369
rect 4249 2329 4261 2363
rect 4295 2360 4307 2363
rect 4724 2360 4752 2391
rect 5534 2388 5540 2400
rect 5592 2428 5598 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 5592 2400 6561 2428
rect 5592 2388 5598 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 5902 2360 5908 2372
rect 4295 2332 5908 2360
rect 4295 2329 4307 2332
rect 4249 2323 4307 2329
rect 5902 2320 5908 2332
rect 5960 2320 5966 2372
rect 2590 2252 2596 2304
rect 2648 2292 2654 2304
rect 3789 2295 3847 2301
rect 3789 2292 3801 2295
rect 2648 2264 3801 2292
rect 2648 2252 2654 2264
rect 3789 2261 3801 2264
rect 3835 2261 3847 2295
rect 3789 2255 3847 2261
rect 5166 2252 5172 2304
rect 5224 2292 5230 2304
rect 6365 2295 6423 2301
rect 6365 2292 6377 2295
rect 5224 2264 6377 2292
rect 5224 2252 5230 2264
rect 6365 2261 6377 2264
rect 6411 2261 6423 2295
rect 6365 2255 6423 2261
rect 6638 2252 6644 2304
rect 6696 2292 6702 2304
rect 6733 2295 6791 2301
rect 6733 2292 6745 2295
rect 6696 2264 6745 2292
rect 6696 2252 6702 2264
rect 6733 2261 6745 2264
rect 6779 2261 6791 2295
rect 6733 2255 6791 2261
rect 7101 2295 7159 2301
rect 7101 2261 7113 2295
rect 7147 2292 7159 2295
rect 7208 2292 7236 2468
rect 8294 2456 8300 2468
rect 8352 2456 8358 2508
rect 7285 2431 7343 2437
rect 7285 2397 7297 2431
rect 7331 2397 7343 2431
rect 7285 2391 7343 2397
rect 7300 2360 7328 2391
rect 7834 2388 7840 2440
rect 7892 2428 7898 2440
rect 8021 2431 8079 2437
rect 8021 2428 8033 2431
rect 7892 2400 8033 2428
rect 7892 2388 7898 2400
rect 8021 2397 8033 2400
rect 8067 2428 8079 2431
rect 8573 2431 8631 2437
rect 8573 2428 8585 2431
rect 8067 2400 8585 2428
rect 8067 2397 8079 2400
rect 8021 2391 8079 2397
rect 8573 2397 8585 2400
rect 8619 2397 8631 2431
rect 8573 2391 8631 2397
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 9876 2437 9904 2536
rect 12618 2524 12624 2536
rect 12676 2524 12682 2576
rect 13538 2524 13544 2576
rect 13596 2564 13602 2576
rect 13596 2536 15056 2564
rect 13596 2524 13602 2536
rect 12158 2496 12164 2508
rect 11900 2468 12164 2496
rect 11900 2437 11928 2468
rect 12158 2456 12164 2468
rect 12216 2496 12222 2508
rect 14093 2499 14151 2505
rect 14093 2496 14105 2499
rect 12216 2468 14105 2496
rect 12216 2456 12222 2468
rect 14093 2465 14105 2468
rect 14139 2465 14151 2499
rect 14093 2459 14151 2465
rect 14366 2456 14372 2508
rect 14424 2496 14430 2508
rect 14921 2499 14979 2505
rect 14921 2496 14933 2499
rect 14424 2468 14933 2496
rect 14424 2456 14430 2468
rect 14921 2465 14933 2468
rect 14967 2465 14979 2499
rect 14921 2459 14979 2465
rect 9309 2431 9367 2437
rect 9309 2428 9321 2431
rect 9088 2400 9321 2428
rect 9088 2388 9094 2400
rect 9309 2397 9321 2400
rect 9355 2397 9367 2431
rect 9309 2391 9367 2397
rect 9861 2431 9919 2437
rect 9861 2397 9873 2431
rect 9907 2397 9919 2431
rect 9861 2391 9919 2397
rect 11885 2431 11943 2437
rect 11885 2397 11897 2431
rect 11931 2397 11943 2431
rect 11885 2391 11943 2397
rect 12529 2431 12587 2437
rect 12529 2397 12541 2431
rect 12575 2428 12587 2431
rect 14645 2431 14703 2437
rect 12575 2400 14412 2428
rect 12575 2397 12587 2400
rect 12529 2391 12587 2397
rect 7929 2363 7987 2369
rect 7929 2360 7941 2363
rect 7300 2332 7941 2360
rect 7929 2329 7941 2332
rect 7975 2360 7987 2363
rect 8846 2360 8852 2372
rect 7975 2332 8852 2360
rect 7975 2329 7987 2332
rect 7929 2323 7987 2329
rect 8846 2320 8852 2332
rect 8904 2320 8910 2372
rect 9324 2360 9352 2391
rect 9950 2360 9956 2372
rect 9324 2332 9956 2360
rect 9950 2320 9956 2332
rect 10008 2320 10014 2372
rect 10962 2320 10968 2372
rect 11020 2320 11026 2372
rect 11624 2332 12388 2360
rect 7147 2264 7236 2292
rect 7147 2261 7159 2264
rect 7101 2255 7159 2261
rect 7742 2252 7748 2304
rect 7800 2252 7806 2304
rect 8386 2252 8392 2304
rect 8444 2252 8450 2304
rect 9125 2295 9183 2301
rect 9125 2261 9137 2295
rect 9171 2292 9183 2295
rect 11624 2292 11652 2332
rect 9171 2264 11652 2292
rect 9171 2261 9183 2264
rect 9125 2255 9183 2261
rect 11698 2252 11704 2304
rect 11756 2252 11762 2304
rect 12360 2292 12388 2332
rect 13262 2320 13268 2372
rect 13320 2320 13326 2372
rect 14384 2360 14412 2400
rect 14645 2397 14657 2431
rect 14691 2428 14703 2431
rect 15028 2428 15056 2536
rect 16114 2524 16120 2576
rect 16172 2564 16178 2576
rect 22278 2564 22284 2576
rect 16172 2536 22284 2564
rect 16172 2524 16178 2536
rect 22278 2524 22284 2536
rect 22336 2524 22342 2576
rect 22646 2524 22652 2576
rect 22704 2564 22710 2576
rect 24581 2567 24639 2573
rect 24581 2564 24593 2567
rect 22704 2536 24593 2564
rect 22704 2524 22710 2536
rect 24581 2533 24593 2536
rect 24627 2533 24639 2567
rect 24581 2527 24639 2533
rect 17310 2456 17316 2508
rect 17368 2456 17374 2508
rect 20530 2496 20536 2508
rect 18892 2468 20536 2496
rect 14691 2400 15056 2428
rect 14691 2397 14703 2400
rect 14645 2391 14703 2397
rect 16022 2388 16028 2440
rect 16080 2428 16086 2440
rect 16117 2431 16175 2437
rect 16117 2428 16129 2431
rect 16080 2400 16129 2428
rect 16080 2388 16086 2400
rect 16117 2397 16129 2400
rect 16163 2397 16175 2431
rect 16117 2391 16175 2397
rect 16758 2388 16764 2440
rect 16816 2428 16822 2440
rect 18892 2437 18920 2468
rect 20530 2456 20536 2468
rect 20588 2456 20594 2508
rect 20640 2468 22048 2496
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16816 2400 16865 2428
rect 16816 2388 16822 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 18877 2431 18935 2437
rect 18877 2397 18889 2431
rect 18923 2397 18935 2431
rect 18877 2391 18935 2397
rect 19613 2431 19671 2437
rect 19613 2397 19625 2431
rect 19659 2428 19671 2431
rect 19702 2428 19708 2440
rect 19659 2400 19708 2428
rect 19659 2397 19671 2400
rect 19613 2391 19671 2397
rect 19702 2388 19708 2400
rect 19760 2388 19766 2440
rect 20346 2388 20352 2440
rect 20404 2388 20410 2440
rect 16298 2360 16304 2372
rect 14384 2332 16304 2360
rect 16298 2320 16304 2332
rect 16356 2320 16362 2372
rect 16666 2320 16672 2372
rect 16724 2360 16730 2372
rect 20640 2360 20668 2468
rect 22020 2437 22048 2468
rect 22186 2456 22192 2508
rect 22244 2496 22250 2508
rect 22465 2499 22523 2505
rect 22465 2496 22477 2499
rect 22244 2468 22477 2496
rect 22244 2456 22250 2468
rect 22465 2465 22477 2468
rect 22511 2465 22523 2499
rect 22465 2459 22523 2465
rect 21453 2431 21511 2437
rect 21453 2397 21465 2431
rect 21499 2397 21511 2431
rect 21453 2391 21511 2397
rect 22005 2431 22063 2437
rect 22005 2397 22017 2431
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 16724 2332 20668 2360
rect 16724 2320 16730 2332
rect 15654 2292 15660 2304
rect 12360 2264 15660 2292
rect 15654 2252 15660 2264
rect 15712 2252 15718 2304
rect 17770 2252 17776 2304
rect 17828 2292 17834 2304
rect 21468 2292 21496 2391
rect 23382 2388 23388 2440
rect 23440 2428 23446 2440
rect 24029 2431 24087 2437
rect 24029 2428 24041 2431
rect 23440 2400 24041 2428
rect 23440 2388 23446 2400
rect 24029 2397 24041 2400
rect 24075 2397 24087 2431
rect 24029 2391 24087 2397
rect 24765 2431 24823 2437
rect 24765 2397 24777 2431
rect 24811 2428 24823 2431
rect 24946 2428 24952 2440
rect 24811 2400 24952 2428
rect 24811 2397 24823 2400
rect 24765 2391 24823 2397
rect 24946 2388 24952 2400
rect 25004 2388 25010 2440
rect 17828 2264 21496 2292
rect 17828 2252 17834 2264
rect 23842 2252 23848 2304
rect 23900 2252 23906 2304
rect 1104 2202 25852 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 25852 2202
rect 1104 2128 25852 2150
rect 13722 1980 13728 2032
rect 13780 2020 13786 2032
rect 23842 2020 23848 2032
rect 13780 1992 23848 2020
rect 13780 1980 13786 1992
rect 23842 1980 23848 1992
rect 23900 1980 23906 2032
rect 8386 1912 8392 1964
rect 8444 1952 8450 1964
rect 15562 1952 15568 1964
rect 8444 1924 15568 1952
rect 8444 1912 8450 1924
rect 15562 1912 15568 1924
rect 15620 1912 15626 1964
rect 10962 1776 10968 1828
rect 11020 1816 11026 1828
rect 22094 1816 22100 1828
rect 11020 1788 22100 1816
rect 11020 1776 11026 1788
rect 22094 1776 22100 1788
rect 22152 1776 22158 1828
rect 21634 1232 21640 1284
rect 21692 1272 21698 1284
rect 23198 1272 23204 1284
rect 21692 1244 23204 1272
rect 21692 1232 21698 1244
rect 23198 1232 23204 1244
rect 23256 1232 23262 1284
<< via1 >>
rect 7950 54374 8002 54426
rect 8014 54374 8066 54426
rect 8078 54374 8130 54426
rect 8142 54374 8194 54426
rect 8206 54374 8258 54426
rect 17950 54374 18002 54426
rect 18014 54374 18066 54426
rect 18078 54374 18130 54426
rect 18142 54374 18194 54426
rect 18206 54374 18258 54426
rect 13820 54315 13872 54324
rect 13820 54281 13829 54315
rect 13829 54281 13863 54315
rect 13863 54281 13872 54315
rect 13820 54272 13872 54281
rect 18972 54315 19024 54324
rect 18972 54281 18981 54315
rect 18981 54281 19015 54315
rect 19015 54281 19024 54315
rect 18972 54272 19024 54281
rect 4068 54136 4120 54188
rect 4804 54179 4856 54188
rect 4804 54145 4813 54179
rect 4813 54145 4847 54179
rect 4847 54145 4856 54179
rect 4804 54136 4856 54145
rect 7380 54179 7432 54188
rect 7380 54145 7389 54179
rect 7389 54145 7423 54179
rect 7423 54145 7432 54179
rect 7380 54136 7432 54145
rect 9588 54179 9640 54188
rect 9588 54145 9597 54179
rect 9597 54145 9631 54179
rect 9631 54145 9640 54179
rect 9588 54136 9640 54145
rect 11704 54136 11756 54188
rect 2412 54068 2464 54120
rect 5172 54111 5224 54120
rect 5172 54077 5181 54111
rect 5181 54077 5215 54111
rect 5215 54077 5224 54111
rect 5172 54068 5224 54077
rect 7840 54111 7892 54120
rect 7840 54077 7849 54111
rect 7849 54077 7883 54111
rect 7883 54077 7892 54111
rect 7840 54068 7892 54077
rect 9312 54068 9364 54120
rect 12348 54068 12400 54120
rect 14832 54136 14884 54188
rect 16580 54136 16632 54188
rect 17592 54136 17644 54188
rect 8300 54000 8352 54052
rect 16672 54068 16724 54120
rect 20720 54179 20772 54188
rect 20720 54145 20729 54179
rect 20729 54145 20763 54179
rect 20763 54145 20772 54179
rect 20720 54136 20772 54145
rect 21732 54136 21784 54188
rect 23112 54136 23164 54188
rect 24492 54136 24544 54188
rect 13912 54000 13964 54052
rect 16120 54000 16172 54052
rect 25044 54000 25096 54052
rect 12716 53932 12768 53984
rect 15660 53932 15712 53984
rect 22192 53975 22244 53984
rect 22192 53941 22201 53975
rect 22201 53941 22235 53975
rect 22235 53941 22244 53975
rect 22192 53932 22244 53941
rect 22652 53932 22704 53984
rect 24676 53932 24728 53984
rect 25136 53932 25188 53984
rect 2950 53830 3002 53882
rect 3014 53830 3066 53882
rect 3078 53830 3130 53882
rect 3142 53830 3194 53882
rect 3206 53830 3258 53882
rect 12950 53830 13002 53882
rect 13014 53830 13066 53882
rect 13078 53830 13130 53882
rect 13142 53830 13194 53882
rect 13206 53830 13258 53882
rect 22950 53830 23002 53882
rect 23014 53830 23066 53882
rect 23078 53830 23130 53882
rect 23142 53830 23194 53882
rect 23206 53830 23258 53882
rect 10692 53660 10744 53712
rect 1032 53592 1084 53644
rect 3792 53592 3844 53644
rect 6552 53592 6604 53644
rect 4160 53567 4212 53576
rect 4160 53533 4169 53567
rect 4169 53533 4203 53567
rect 4203 53533 4212 53567
rect 4160 53524 4212 53533
rect 7840 53524 7892 53576
rect 10692 53524 10744 53576
rect 23388 53524 23440 53576
rect 24584 53728 24636 53780
rect 24768 53771 24820 53780
rect 24768 53737 24777 53771
rect 24777 53737 24811 53771
rect 24811 53737 24820 53771
rect 24768 53728 24820 53737
rect 25044 53567 25096 53576
rect 25044 53533 25053 53567
rect 25053 53533 25087 53567
rect 25087 53533 25096 53567
rect 25044 53524 25096 53533
rect 5540 53456 5592 53508
rect 22836 53388 22888 53440
rect 23940 53431 23992 53440
rect 23940 53397 23949 53431
rect 23949 53397 23983 53431
rect 23983 53397 23992 53431
rect 23940 53388 23992 53397
rect 26516 53388 26568 53440
rect 7950 53286 8002 53338
rect 8014 53286 8066 53338
rect 8078 53286 8130 53338
rect 8142 53286 8194 53338
rect 8206 53286 8258 53338
rect 17950 53286 18002 53338
rect 18014 53286 18066 53338
rect 18078 53286 18130 53338
rect 18142 53286 18194 53338
rect 18206 53286 18258 53338
rect 4068 53184 4120 53236
rect 23388 53227 23440 53236
rect 23388 53193 23397 53227
rect 23397 53193 23431 53227
rect 23431 53193 23440 53227
rect 23388 53184 23440 53193
rect 7748 53048 7800 53100
rect 24768 53048 24820 53100
rect 25044 53091 25096 53100
rect 25044 53057 25053 53091
rect 25053 53057 25087 53091
rect 25087 53057 25096 53091
rect 25044 53048 25096 53057
rect 15568 52912 15620 52964
rect 24492 52887 24544 52896
rect 24492 52853 24501 52887
rect 24501 52853 24535 52887
rect 24535 52853 24544 52887
rect 24492 52844 24544 52853
rect 2950 52742 3002 52794
rect 3014 52742 3066 52794
rect 3078 52742 3130 52794
rect 3142 52742 3194 52794
rect 3206 52742 3258 52794
rect 12950 52742 13002 52794
rect 13014 52742 13066 52794
rect 13078 52742 13130 52794
rect 13142 52742 13194 52794
rect 13206 52742 13258 52794
rect 22950 52742 23002 52794
rect 23014 52742 23066 52794
rect 23078 52742 23130 52794
rect 23142 52742 23194 52794
rect 23206 52742 23258 52794
rect 4160 52640 4212 52692
rect 16396 52640 16448 52692
rect 24492 52640 24544 52692
rect 9404 52436 9456 52488
rect 26792 52436 26844 52488
rect 24952 52411 25004 52420
rect 24952 52377 24961 52411
rect 24961 52377 24995 52411
rect 24995 52377 25004 52411
rect 24952 52368 25004 52377
rect 7950 52198 8002 52250
rect 8014 52198 8066 52250
rect 8078 52198 8130 52250
rect 8142 52198 8194 52250
rect 8206 52198 8258 52250
rect 17950 52198 18002 52250
rect 18014 52198 18066 52250
rect 18078 52198 18130 52250
rect 18142 52198 18194 52250
rect 18206 52198 18258 52250
rect 25872 51960 25924 52012
rect 24860 51756 24912 51808
rect 2950 51654 3002 51706
rect 3014 51654 3066 51706
rect 3078 51654 3130 51706
rect 3142 51654 3194 51706
rect 3206 51654 3258 51706
rect 12950 51654 13002 51706
rect 13014 51654 13066 51706
rect 13078 51654 13130 51706
rect 13142 51654 13194 51706
rect 13206 51654 13258 51706
rect 22950 51654 23002 51706
rect 23014 51654 23066 51706
rect 23078 51654 23130 51706
rect 23142 51654 23194 51706
rect 23206 51654 23258 51706
rect 7380 51552 7432 51604
rect 7840 51484 7892 51536
rect 4804 51348 4856 51400
rect 8484 51391 8536 51400
rect 8484 51357 8493 51391
rect 8493 51357 8527 51391
rect 8527 51357 8536 51391
rect 8484 51348 8536 51357
rect 10508 51348 10560 51400
rect 10784 51280 10836 51332
rect 24952 51323 25004 51332
rect 24952 51289 24961 51323
rect 24961 51289 24995 51323
rect 24995 51289 25004 51323
rect 24952 51280 25004 51289
rect 26884 51280 26936 51332
rect 7950 51110 8002 51162
rect 8014 51110 8066 51162
rect 8078 51110 8130 51162
rect 8142 51110 8194 51162
rect 8206 51110 8258 51162
rect 17950 51110 18002 51162
rect 18014 51110 18066 51162
rect 18078 51110 18130 51162
rect 18142 51110 18194 51162
rect 18206 51110 18258 51162
rect 24952 50915 25004 50924
rect 24952 50881 24961 50915
rect 24961 50881 24995 50915
rect 24995 50881 25004 50915
rect 24952 50872 25004 50881
rect 25044 50711 25096 50720
rect 25044 50677 25053 50711
rect 25053 50677 25087 50711
rect 25087 50677 25096 50711
rect 25044 50668 25096 50677
rect 2950 50566 3002 50618
rect 3014 50566 3066 50618
rect 3078 50566 3130 50618
rect 3142 50566 3194 50618
rect 3206 50566 3258 50618
rect 12950 50566 13002 50618
rect 13014 50566 13066 50618
rect 13078 50566 13130 50618
rect 13142 50566 13194 50618
rect 13206 50566 13258 50618
rect 22950 50566 23002 50618
rect 23014 50566 23066 50618
rect 23078 50566 23130 50618
rect 23142 50566 23194 50618
rect 23206 50566 23258 50618
rect 5540 50464 5592 50516
rect 8392 50464 8444 50516
rect 9588 50507 9640 50516
rect 9588 50473 9597 50507
rect 9597 50473 9631 50507
rect 9631 50473 9640 50507
rect 9588 50464 9640 50473
rect 16028 50464 16080 50516
rect 25044 50464 25096 50516
rect 7748 50396 7800 50448
rect 8300 50260 8352 50312
rect 9588 50260 9640 50312
rect 25504 50167 25556 50176
rect 25504 50133 25513 50167
rect 25513 50133 25547 50167
rect 25547 50133 25556 50167
rect 25504 50124 25556 50133
rect 7950 50022 8002 50074
rect 8014 50022 8066 50074
rect 8078 50022 8130 50074
rect 8142 50022 8194 50074
rect 8206 50022 8258 50074
rect 17950 50022 18002 50074
rect 18014 50022 18066 50074
rect 18078 50022 18130 50074
rect 18142 50022 18194 50074
rect 18206 50022 18258 50074
rect 25504 49784 25556 49836
rect 23664 49716 23716 49768
rect 2950 49478 3002 49530
rect 3014 49478 3066 49530
rect 3078 49478 3130 49530
rect 3142 49478 3194 49530
rect 3206 49478 3258 49530
rect 12950 49478 13002 49530
rect 13014 49478 13066 49530
rect 13078 49478 13130 49530
rect 13142 49478 13194 49530
rect 13206 49478 13258 49530
rect 22950 49478 23002 49530
rect 23014 49478 23066 49530
rect 23078 49478 23130 49530
rect 23142 49478 23194 49530
rect 23206 49478 23258 49530
rect 10692 49351 10744 49360
rect 10692 49317 10701 49351
rect 10701 49317 10735 49351
rect 10735 49317 10744 49351
rect 10692 49308 10744 49317
rect 11704 49351 11756 49360
rect 11704 49317 11713 49351
rect 11713 49317 11747 49351
rect 11747 49317 11756 49351
rect 11704 49308 11756 49317
rect 10232 49104 10284 49156
rect 10876 49104 10928 49156
rect 25136 49147 25188 49156
rect 25136 49113 25145 49147
rect 25145 49113 25179 49147
rect 25179 49113 25188 49147
rect 25136 49104 25188 49113
rect 25228 49079 25280 49088
rect 25228 49045 25237 49079
rect 25237 49045 25271 49079
rect 25271 49045 25280 49079
rect 25228 49036 25280 49045
rect 7950 48934 8002 48986
rect 8014 48934 8066 48986
rect 8078 48934 8130 48986
rect 8142 48934 8194 48986
rect 8206 48934 8258 48986
rect 17950 48934 18002 48986
rect 18014 48934 18066 48986
rect 18078 48934 18130 48986
rect 18142 48934 18194 48986
rect 18206 48934 18258 48986
rect 8392 48875 8444 48884
rect 8392 48841 8401 48875
rect 8401 48841 8435 48875
rect 8435 48841 8444 48875
rect 8392 48832 8444 48841
rect 9496 48628 9548 48680
rect 9128 48560 9180 48612
rect 9956 48492 10008 48544
rect 25136 48492 25188 48544
rect 2950 48390 3002 48442
rect 3014 48390 3066 48442
rect 3078 48390 3130 48442
rect 3142 48390 3194 48442
rect 3206 48390 3258 48442
rect 12950 48390 13002 48442
rect 13014 48390 13066 48442
rect 13078 48390 13130 48442
rect 13142 48390 13194 48442
rect 13206 48390 13258 48442
rect 22950 48390 23002 48442
rect 23014 48390 23066 48442
rect 23078 48390 23130 48442
rect 23142 48390 23194 48442
rect 23206 48390 23258 48442
rect 7748 48084 7800 48136
rect 25136 48127 25188 48136
rect 25136 48093 25145 48127
rect 25145 48093 25179 48127
rect 25179 48093 25188 48127
rect 25136 48084 25188 48093
rect 26332 48016 26384 48068
rect 12624 47948 12676 48000
rect 7950 47846 8002 47898
rect 8014 47846 8066 47898
rect 8078 47846 8130 47898
rect 8142 47846 8194 47898
rect 8206 47846 8258 47898
rect 17950 47846 18002 47898
rect 18014 47846 18066 47898
rect 18078 47846 18130 47898
rect 18142 47846 18194 47898
rect 18206 47846 18258 47898
rect 9220 47744 9272 47796
rect 9404 47744 9456 47796
rect 8300 47608 8352 47660
rect 10324 47608 10376 47660
rect 25320 47651 25372 47660
rect 25320 47617 25329 47651
rect 25329 47617 25363 47651
rect 25363 47617 25372 47651
rect 25320 47608 25372 47617
rect 9496 47447 9548 47456
rect 9496 47413 9505 47447
rect 9505 47413 9539 47447
rect 9539 47413 9548 47447
rect 9496 47404 9548 47413
rect 26424 47404 26476 47456
rect 2950 47302 3002 47354
rect 3014 47302 3066 47354
rect 3078 47302 3130 47354
rect 3142 47302 3194 47354
rect 3206 47302 3258 47354
rect 12950 47302 13002 47354
rect 13014 47302 13066 47354
rect 13078 47302 13130 47354
rect 13142 47302 13194 47354
rect 13206 47302 13258 47354
rect 22950 47302 23002 47354
rect 23014 47302 23066 47354
rect 23078 47302 23130 47354
rect 23142 47302 23194 47354
rect 23206 47302 23258 47354
rect 9220 46996 9272 47048
rect 13728 46928 13780 46980
rect 25320 46860 25372 46912
rect 7950 46758 8002 46810
rect 8014 46758 8066 46810
rect 8078 46758 8130 46810
rect 8142 46758 8194 46810
rect 8206 46758 8258 46810
rect 17950 46758 18002 46810
rect 18014 46758 18066 46810
rect 18078 46758 18130 46810
rect 18142 46758 18194 46810
rect 18206 46758 18258 46810
rect 9772 46656 9824 46708
rect 10784 46699 10836 46708
rect 10784 46665 10793 46699
rect 10793 46665 10827 46699
rect 10827 46665 10836 46699
rect 10784 46656 10836 46665
rect 10324 46563 10376 46572
rect 10324 46529 10333 46563
rect 10333 46529 10367 46563
rect 10367 46529 10376 46563
rect 10324 46520 10376 46529
rect 13728 46588 13780 46640
rect 13912 46563 13964 46572
rect 13912 46529 13921 46563
rect 13921 46529 13955 46563
rect 13955 46529 13964 46563
rect 13912 46520 13964 46529
rect 25320 46563 25372 46572
rect 25320 46529 25329 46563
rect 25329 46529 25363 46563
rect 25363 46529 25372 46563
rect 25320 46520 25372 46529
rect 15752 46495 15804 46504
rect 15752 46461 15761 46495
rect 15761 46461 15795 46495
rect 15795 46461 15804 46495
rect 15752 46452 15804 46461
rect 10416 46359 10468 46368
rect 10416 46325 10425 46359
rect 10425 46325 10459 46359
rect 10459 46325 10468 46359
rect 10416 46316 10468 46325
rect 15016 46316 15068 46368
rect 25412 46316 25464 46368
rect 2950 46214 3002 46266
rect 3014 46214 3066 46266
rect 3078 46214 3130 46266
rect 3142 46214 3194 46266
rect 3206 46214 3258 46266
rect 12950 46214 13002 46266
rect 13014 46214 13066 46266
rect 13078 46214 13130 46266
rect 13142 46214 13194 46266
rect 13206 46214 13258 46266
rect 22950 46214 23002 46266
rect 23014 46214 23066 46266
rect 23078 46214 23130 46266
rect 23142 46214 23194 46266
rect 23206 46214 23258 46266
rect 8484 46155 8536 46164
rect 8484 46121 8493 46155
rect 8493 46121 8527 46155
rect 8527 46121 8536 46155
rect 8484 46112 8536 46121
rect 7748 45976 7800 46028
rect 15660 46044 15712 46096
rect 15016 46019 15068 46028
rect 15016 45985 15025 46019
rect 15025 45985 15059 46019
rect 15059 45985 15068 46019
rect 15016 45976 15068 45985
rect 16488 46019 16540 46028
rect 16488 45985 16497 46019
rect 16497 45985 16531 46019
rect 16531 45985 16540 46019
rect 16488 45976 16540 45985
rect 7840 45908 7892 45960
rect 12532 45908 12584 45960
rect 25320 45951 25372 45960
rect 25320 45917 25329 45951
rect 25329 45917 25363 45951
rect 25363 45917 25372 45951
rect 25320 45908 25372 45917
rect 15108 45772 15160 45824
rect 24860 45772 24912 45824
rect 7950 45670 8002 45722
rect 8014 45670 8066 45722
rect 8078 45670 8130 45722
rect 8142 45670 8194 45722
rect 8206 45670 8258 45722
rect 17950 45670 18002 45722
rect 18014 45670 18066 45722
rect 18078 45670 18130 45722
rect 18142 45670 18194 45722
rect 18206 45670 18258 45722
rect 10508 45500 10560 45552
rect 12532 45500 12584 45552
rect 12624 45500 12676 45552
rect 12716 45475 12768 45484
rect 12716 45441 12725 45475
rect 12725 45441 12759 45475
rect 12759 45441 12768 45475
rect 12716 45432 12768 45441
rect 14556 45407 14608 45416
rect 14556 45373 14565 45407
rect 14565 45373 14599 45407
rect 14599 45373 14608 45407
rect 14556 45364 14608 45373
rect 25320 45228 25372 45280
rect 2950 45126 3002 45178
rect 3014 45126 3066 45178
rect 3078 45126 3130 45178
rect 3142 45126 3194 45178
rect 3206 45126 3258 45178
rect 12950 45126 13002 45178
rect 13014 45126 13066 45178
rect 13078 45126 13130 45178
rect 13142 45126 13194 45178
rect 13206 45126 13258 45178
rect 22950 45126 23002 45178
rect 23014 45126 23066 45178
rect 23078 45126 23130 45178
rect 23142 45126 23194 45178
rect 23206 45126 23258 45178
rect 9404 45024 9456 45076
rect 9128 44931 9180 44940
rect 9128 44897 9137 44931
rect 9137 44897 9171 44931
rect 9171 44897 9180 44931
rect 9128 44888 9180 44897
rect 9404 44888 9456 44940
rect 9956 44888 10008 44940
rect 9680 44752 9732 44804
rect 16120 44888 16172 44940
rect 25320 44863 25372 44872
rect 25320 44829 25329 44863
rect 25329 44829 25363 44863
rect 25363 44829 25372 44863
rect 25320 44820 25372 44829
rect 10416 44684 10468 44736
rect 15108 44752 15160 44804
rect 19984 44752 20036 44804
rect 11520 44684 11572 44736
rect 25044 44684 25096 44736
rect 7950 44582 8002 44634
rect 8014 44582 8066 44634
rect 8078 44582 8130 44634
rect 8142 44582 8194 44634
rect 8206 44582 8258 44634
rect 17950 44582 18002 44634
rect 18014 44582 18066 44634
rect 18078 44582 18130 44634
rect 18142 44582 18194 44634
rect 18206 44582 18258 44634
rect 9588 44523 9640 44532
rect 9588 44489 9597 44523
rect 9597 44489 9631 44523
rect 9631 44489 9640 44523
rect 9588 44480 9640 44489
rect 9220 44344 9272 44396
rect 10324 44344 10376 44396
rect 24768 44387 24820 44396
rect 24768 44353 24777 44387
rect 24777 44353 24811 44387
rect 24811 44353 24820 44387
rect 24768 44344 24820 44353
rect 9036 44276 9088 44328
rect 10508 44208 10560 44260
rect 25872 44208 25924 44260
rect 10692 44183 10744 44192
rect 10692 44149 10701 44183
rect 10701 44149 10735 44183
rect 10735 44149 10744 44183
rect 10692 44140 10744 44149
rect 10968 44140 11020 44192
rect 2950 44038 3002 44090
rect 3014 44038 3066 44090
rect 3078 44038 3130 44090
rect 3142 44038 3194 44090
rect 3206 44038 3258 44090
rect 12950 44038 13002 44090
rect 13014 44038 13066 44090
rect 13078 44038 13130 44090
rect 13142 44038 13194 44090
rect 13206 44038 13258 44090
rect 22950 44038 23002 44090
rect 23014 44038 23066 44090
rect 23078 44038 23130 44090
rect 23142 44038 23194 44090
rect 23206 44038 23258 44090
rect 24952 43936 25004 43988
rect 21088 43800 21140 43852
rect 19524 43732 19576 43784
rect 21088 43664 21140 43716
rect 22100 43639 22152 43648
rect 22100 43605 22109 43639
rect 22109 43605 22143 43639
rect 22143 43605 22152 43639
rect 22100 43596 22152 43605
rect 25504 43639 25556 43648
rect 25504 43605 25513 43639
rect 25513 43605 25547 43639
rect 25547 43605 25556 43639
rect 25504 43596 25556 43605
rect 7950 43494 8002 43546
rect 8014 43494 8066 43546
rect 8078 43494 8130 43546
rect 8142 43494 8194 43546
rect 8206 43494 8258 43546
rect 17950 43494 18002 43546
rect 18014 43494 18066 43546
rect 18078 43494 18130 43546
rect 18142 43494 18194 43546
rect 18206 43494 18258 43546
rect 25504 43324 25556 43376
rect 25964 43120 26016 43172
rect 2950 42950 3002 43002
rect 3014 42950 3066 43002
rect 3078 42950 3130 43002
rect 3142 42950 3194 43002
rect 3206 42950 3258 43002
rect 12950 42950 13002 43002
rect 13014 42950 13066 43002
rect 13078 42950 13130 43002
rect 13142 42950 13194 43002
rect 13206 42950 13258 43002
rect 22950 42950 23002 43002
rect 23014 42950 23066 43002
rect 23078 42950 23130 43002
rect 23142 42950 23194 43002
rect 23206 42950 23258 43002
rect 9772 42755 9824 42764
rect 9772 42721 9781 42755
rect 9781 42721 9815 42755
rect 9815 42721 9824 42755
rect 9772 42712 9824 42721
rect 10232 42755 10284 42764
rect 10232 42721 10241 42755
rect 10241 42721 10275 42755
rect 10275 42721 10284 42755
rect 10232 42712 10284 42721
rect 8944 42644 8996 42696
rect 25136 42619 25188 42628
rect 25136 42585 25145 42619
rect 25145 42585 25179 42619
rect 25179 42585 25188 42619
rect 25136 42576 25188 42585
rect 25688 42576 25740 42628
rect 7950 42406 8002 42458
rect 8014 42406 8066 42458
rect 8078 42406 8130 42458
rect 8142 42406 8194 42458
rect 8206 42406 8258 42458
rect 17950 42406 18002 42458
rect 18014 42406 18066 42458
rect 18078 42406 18130 42458
rect 18142 42406 18194 42458
rect 18206 42406 18258 42458
rect 9680 42304 9732 42356
rect 11520 42236 11572 42288
rect 9404 42143 9456 42152
rect 9404 42109 9413 42143
rect 9413 42109 9447 42143
rect 9447 42109 9456 42143
rect 9404 42100 9456 42109
rect 9772 42100 9824 42152
rect 10692 42100 10744 42152
rect 11520 42007 11572 42016
rect 11520 41973 11529 42007
rect 11529 41973 11563 42007
rect 11563 41973 11572 42007
rect 11520 41964 11572 41973
rect 25136 41964 25188 42016
rect 2950 41862 3002 41914
rect 3014 41862 3066 41914
rect 3078 41862 3130 41914
rect 3142 41862 3194 41914
rect 3206 41862 3258 41914
rect 12950 41862 13002 41914
rect 13014 41862 13066 41914
rect 13078 41862 13130 41914
rect 13142 41862 13194 41914
rect 13206 41862 13258 41914
rect 22950 41862 23002 41914
rect 23014 41862 23066 41914
rect 23078 41862 23130 41914
rect 23142 41862 23194 41914
rect 23206 41862 23258 41914
rect 10876 41803 10928 41812
rect 10876 41769 10885 41803
rect 10885 41769 10919 41803
rect 10919 41769 10928 41803
rect 10876 41760 10928 41769
rect 10968 41624 11020 41676
rect 9220 41556 9272 41608
rect 25136 41599 25188 41608
rect 25136 41565 25145 41599
rect 25145 41565 25179 41599
rect 25179 41565 25188 41599
rect 25136 41556 25188 41565
rect 26148 41488 26200 41540
rect 7950 41318 8002 41370
rect 8014 41318 8066 41370
rect 8078 41318 8130 41370
rect 8142 41318 8194 41370
rect 8206 41318 8258 41370
rect 17950 41318 18002 41370
rect 18014 41318 18066 41370
rect 18078 41318 18130 41370
rect 18142 41318 18194 41370
rect 18206 41318 18258 41370
rect 25320 41123 25372 41132
rect 25320 41089 25329 41123
rect 25329 41089 25363 41123
rect 25363 41089 25372 41123
rect 25320 41080 25372 41089
rect 25596 40876 25648 40928
rect 2950 40774 3002 40826
rect 3014 40774 3066 40826
rect 3078 40774 3130 40826
rect 3142 40774 3194 40826
rect 3206 40774 3258 40826
rect 12950 40774 13002 40826
rect 13014 40774 13066 40826
rect 13078 40774 13130 40826
rect 13142 40774 13194 40826
rect 13206 40774 13258 40826
rect 22950 40774 23002 40826
rect 23014 40774 23066 40826
rect 23078 40774 23130 40826
rect 23142 40774 23194 40826
rect 23206 40774 23258 40826
rect 25504 40375 25556 40384
rect 25504 40341 25513 40375
rect 25513 40341 25547 40375
rect 25547 40341 25556 40375
rect 25504 40332 25556 40341
rect 7950 40230 8002 40282
rect 8014 40230 8066 40282
rect 8078 40230 8130 40282
rect 8142 40230 8194 40282
rect 8206 40230 8258 40282
rect 17950 40230 18002 40282
rect 18014 40230 18066 40282
rect 18078 40230 18130 40282
rect 18142 40230 18194 40282
rect 18206 40230 18258 40282
rect 23388 40128 23440 40180
rect 25504 40060 25556 40112
rect 2950 39686 3002 39738
rect 3014 39686 3066 39738
rect 3078 39686 3130 39738
rect 3142 39686 3194 39738
rect 3206 39686 3258 39738
rect 12950 39686 13002 39738
rect 13014 39686 13066 39738
rect 13078 39686 13130 39738
rect 13142 39686 13194 39738
rect 13206 39686 13258 39738
rect 22950 39686 23002 39738
rect 23014 39686 23066 39738
rect 23078 39686 23130 39738
rect 23142 39686 23194 39738
rect 23206 39686 23258 39738
rect 25320 39423 25372 39432
rect 25320 39389 25329 39423
rect 25329 39389 25363 39423
rect 25363 39389 25372 39423
rect 25320 39380 25372 39389
rect 21916 39244 21968 39296
rect 7950 39142 8002 39194
rect 8014 39142 8066 39194
rect 8078 39142 8130 39194
rect 8142 39142 8194 39194
rect 8206 39142 8258 39194
rect 17950 39142 18002 39194
rect 18014 39142 18066 39194
rect 18078 39142 18130 39194
rect 18142 39142 18194 39194
rect 18206 39142 18258 39194
rect 25320 38700 25372 38752
rect 2950 38598 3002 38650
rect 3014 38598 3066 38650
rect 3078 38598 3130 38650
rect 3142 38598 3194 38650
rect 3206 38598 3258 38650
rect 12950 38598 13002 38650
rect 13014 38598 13066 38650
rect 13078 38598 13130 38650
rect 13142 38598 13194 38650
rect 13206 38598 13258 38650
rect 22950 38598 23002 38650
rect 23014 38598 23066 38650
rect 23078 38598 23130 38650
rect 23142 38598 23194 38650
rect 23206 38598 23258 38650
rect 25320 38335 25372 38344
rect 25320 38301 25329 38335
rect 25329 38301 25363 38335
rect 25363 38301 25372 38335
rect 25320 38292 25372 38301
rect 25044 38156 25096 38208
rect 7950 38054 8002 38106
rect 8014 38054 8066 38106
rect 8078 38054 8130 38106
rect 8142 38054 8194 38106
rect 8206 38054 8258 38106
rect 17950 38054 18002 38106
rect 18014 38054 18066 38106
rect 18078 38054 18130 38106
rect 18142 38054 18194 38106
rect 18206 38054 18258 38106
rect 7840 37952 7892 38004
rect 8852 37859 8904 37868
rect 8852 37825 8861 37859
rect 8861 37825 8895 37859
rect 8895 37825 8904 37859
rect 8852 37816 8904 37825
rect 25136 37859 25188 37868
rect 25136 37825 25145 37859
rect 25145 37825 25179 37859
rect 25179 37825 25188 37859
rect 25136 37816 25188 37825
rect 26056 37680 26108 37732
rect 2950 37510 3002 37562
rect 3014 37510 3066 37562
rect 3078 37510 3130 37562
rect 3142 37510 3194 37562
rect 3206 37510 3258 37562
rect 12950 37510 13002 37562
rect 13014 37510 13066 37562
rect 13078 37510 13130 37562
rect 13142 37510 13194 37562
rect 13206 37510 13258 37562
rect 22950 37510 23002 37562
rect 23014 37510 23066 37562
rect 23078 37510 23130 37562
rect 23142 37510 23194 37562
rect 23206 37510 23258 37562
rect 25504 37111 25556 37120
rect 25504 37077 25513 37111
rect 25513 37077 25547 37111
rect 25547 37077 25556 37111
rect 25504 37068 25556 37077
rect 7950 36966 8002 37018
rect 8014 36966 8066 37018
rect 8078 36966 8130 37018
rect 8142 36966 8194 37018
rect 8206 36966 8258 37018
rect 17950 36966 18002 37018
rect 18014 36966 18066 37018
rect 18078 36966 18130 37018
rect 18142 36966 18194 37018
rect 18206 36966 18258 37018
rect 25504 36796 25556 36848
rect 26700 36592 26752 36644
rect 2950 36422 3002 36474
rect 3014 36422 3066 36474
rect 3078 36422 3130 36474
rect 3142 36422 3194 36474
rect 3206 36422 3258 36474
rect 12950 36422 13002 36474
rect 13014 36422 13066 36474
rect 13078 36422 13130 36474
rect 13142 36422 13194 36474
rect 13206 36422 13258 36474
rect 22950 36422 23002 36474
rect 23014 36422 23066 36474
rect 23078 36422 23130 36474
rect 23142 36422 23194 36474
rect 23206 36422 23258 36474
rect 25320 36159 25372 36168
rect 25320 36125 25329 36159
rect 25329 36125 25363 36159
rect 25363 36125 25372 36159
rect 25320 36116 25372 36125
rect 26608 35980 26660 36032
rect 7950 35878 8002 35930
rect 8014 35878 8066 35930
rect 8078 35878 8130 35930
rect 8142 35878 8194 35930
rect 8206 35878 8258 35930
rect 17950 35878 18002 35930
rect 18014 35878 18066 35930
rect 18078 35878 18130 35930
rect 18142 35878 18194 35930
rect 18206 35878 18258 35930
rect 9772 35776 9824 35828
rect 11520 35819 11572 35828
rect 11520 35785 11529 35819
rect 11529 35785 11563 35819
rect 11563 35785 11572 35819
rect 11520 35776 11572 35785
rect 24860 35776 24912 35828
rect 12716 35708 12768 35760
rect 25412 35708 25464 35760
rect 9404 35615 9456 35624
rect 9404 35581 9413 35615
rect 9413 35581 9447 35615
rect 9447 35581 9456 35615
rect 9404 35572 9456 35581
rect 9680 35615 9732 35624
rect 9680 35581 9689 35615
rect 9689 35581 9723 35615
rect 9723 35581 9732 35615
rect 9680 35572 9732 35581
rect 19340 35504 19392 35556
rect 21824 35640 21876 35692
rect 21272 35615 21324 35624
rect 21272 35581 21281 35615
rect 21281 35581 21315 35615
rect 21315 35581 21324 35615
rect 21272 35572 21324 35581
rect 22468 35572 22520 35624
rect 15752 35436 15804 35488
rect 22376 35504 22428 35556
rect 22008 35479 22060 35488
rect 22008 35445 22017 35479
rect 22017 35445 22051 35479
rect 22051 35445 22060 35479
rect 22008 35436 22060 35445
rect 25320 35436 25372 35488
rect 2950 35334 3002 35386
rect 3014 35334 3066 35386
rect 3078 35334 3130 35386
rect 3142 35334 3194 35386
rect 3206 35334 3258 35386
rect 12950 35334 13002 35386
rect 13014 35334 13066 35386
rect 13078 35334 13130 35386
rect 13142 35334 13194 35386
rect 13206 35334 13258 35386
rect 22950 35334 23002 35386
rect 23014 35334 23066 35386
rect 23078 35334 23130 35386
rect 23142 35334 23194 35386
rect 23206 35334 23258 35386
rect 23296 35139 23348 35148
rect 23296 35105 23305 35139
rect 23305 35105 23339 35139
rect 23339 35105 23348 35139
rect 23296 35096 23348 35105
rect 24952 35028 25004 35080
rect 25320 35071 25372 35080
rect 25320 35037 25329 35071
rect 25329 35037 25363 35071
rect 25363 35037 25372 35071
rect 25320 35028 25372 35037
rect 19984 34960 20036 35012
rect 20628 34960 20680 35012
rect 16488 34892 16540 34944
rect 21824 34935 21876 34944
rect 21824 34901 21833 34935
rect 21833 34901 21867 34935
rect 21867 34901 21876 34935
rect 21824 34892 21876 34901
rect 22560 34892 22612 34944
rect 25780 34892 25832 34944
rect 7950 34790 8002 34842
rect 8014 34790 8066 34842
rect 8078 34790 8130 34842
rect 8142 34790 8194 34842
rect 8206 34790 8258 34842
rect 17950 34790 18002 34842
rect 18014 34790 18066 34842
rect 18078 34790 18130 34842
rect 18142 34790 18194 34842
rect 18206 34790 18258 34842
rect 20720 34688 20772 34740
rect 25320 34595 25372 34604
rect 25320 34561 25329 34595
rect 25329 34561 25363 34595
rect 25363 34561 25372 34595
rect 25320 34552 25372 34561
rect 20444 34416 20496 34468
rect 23940 34416 23992 34468
rect 21088 34348 21140 34400
rect 21364 34391 21416 34400
rect 21364 34357 21373 34391
rect 21373 34357 21407 34391
rect 21407 34357 21416 34391
rect 21364 34348 21416 34357
rect 2950 34246 3002 34298
rect 3014 34246 3066 34298
rect 3078 34246 3130 34298
rect 3142 34246 3194 34298
rect 3206 34246 3258 34298
rect 12950 34246 13002 34298
rect 13014 34246 13066 34298
rect 13078 34246 13130 34298
rect 13142 34246 13194 34298
rect 13206 34246 13258 34298
rect 22950 34246 23002 34298
rect 23014 34246 23066 34298
rect 23078 34246 23130 34298
rect 23142 34246 23194 34298
rect 23206 34246 23258 34298
rect 9036 34144 9088 34196
rect 21364 34144 21416 34196
rect 9404 34008 9456 34060
rect 19708 34008 19760 34060
rect 22284 34008 22336 34060
rect 9312 33983 9364 33992
rect 9312 33949 9321 33983
rect 9321 33949 9355 33983
rect 9355 33949 9364 33983
rect 9312 33940 9364 33949
rect 19432 33983 19484 33992
rect 19432 33949 19441 33983
rect 19441 33949 19475 33983
rect 19475 33949 19484 33983
rect 19432 33940 19484 33949
rect 23572 33940 23624 33992
rect 25320 33983 25372 33992
rect 25320 33949 25329 33983
rect 25329 33949 25363 33983
rect 25363 33949 25372 33983
rect 25320 33940 25372 33949
rect 15384 33872 15436 33924
rect 19800 33872 19852 33924
rect 21180 33847 21232 33856
rect 21180 33813 21189 33847
rect 21189 33813 21223 33847
rect 21223 33813 21232 33847
rect 21180 33804 21232 33813
rect 21272 33804 21324 33856
rect 22928 33804 22980 33856
rect 23204 33804 23256 33856
rect 26240 33804 26292 33856
rect 7950 33702 8002 33754
rect 8014 33702 8066 33754
rect 8078 33702 8130 33754
rect 8142 33702 8194 33754
rect 8206 33702 8258 33754
rect 17950 33702 18002 33754
rect 18014 33702 18066 33754
rect 18078 33702 18130 33754
rect 18142 33702 18194 33754
rect 18206 33702 18258 33754
rect 22468 33600 22520 33652
rect 23204 33600 23256 33652
rect 21272 33532 21324 33584
rect 19524 33507 19576 33516
rect 19524 33473 19533 33507
rect 19533 33473 19567 33507
rect 19567 33473 19576 33507
rect 19524 33464 19576 33473
rect 22284 33532 22336 33584
rect 23572 33532 23624 33584
rect 25504 33464 25556 33516
rect 19800 33396 19852 33448
rect 20536 33396 20588 33448
rect 22376 33396 22428 33448
rect 22744 33396 22796 33448
rect 22928 33396 22980 33448
rect 21272 33260 21324 33312
rect 24584 33303 24636 33312
rect 24584 33269 24593 33303
rect 24593 33269 24627 33303
rect 24627 33269 24636 33303
rect 24584 33260 24636 33269
rect 25412 33260 25464 33312
rect 2950 33158 3002 33210
rect 3014 33158 3066 33210
rect 3078 33158 3130 33210
rect 3142 33158 3194 33210
rect 3206 33158 3258 33210
rect 12950 33158 13002 33210
rect 13014 33158 13066 33210
rect 13078 33158 13130 33210
rect 13142 33158 13194 33210
rect 13206 33158 13258 33210
rect 22950 33158 23002 33210
rect 23014 33158 23066 33210
rect 23078 33158 23130 33210
rect 23142 33158 23194 33210
rect 23206 33158 23258 33210
rect 16580 33099 16632 33108
rect 16580 33065 16589 33099
rect 16589 33065 16623 33099
rect 16623 33065 16632 33099
rect 16580 33056 16632 33065
rect 17316 33056 17368 33108
rect 22376 33056 22428 33108
rect 23296 33056 23348 33108
rect 16856 33031 16908 33040
rect 16856 32997 16865 33031
rect 16865 32997 16899 33031
rect 16899 32997 16908 33031
rect 16856 32988 16908 32997
rect 17132 32988 17184 33040
rect 16120 32963 16172 32972
rect 16120 32929 16129 32963
rect 16129 32929 16163 32963
rect 16163 32929 16172 32963
rect 16120 32920 16172 32929
rect 22100 32920 22152 32972
rect 19432 32852 19484 32904
rect 12624 32716 12676 32768
rect 24952 32988 25004 33040
rect 22284 32963 22336 32972
rect 22284 32929 22293 32963
rect 22293 32929 22327 32963
rect 22327 32929 22336 32963
rect 22284 32920 22336 32929
rect 16856 32716 16908 32768
rect 19616 32759 19668 32768
rect 19616 32725 19625 32759
rect 19625 32725 19659 32759
rect 19659 32725 19668 32759
rect 19616 32716 19668 32725
rect 21824 32716 21876 32768
rect 22376 32716 22428 32768
rect 22836 32716 22888 32768
rect 23572 32784 23624 32836
rect 24584 32852 24636 32904
rect 24768 32852 24820 32904
rect 25596 32852 25648 32904
rect 24492 32716 24544 32768
rect 24584 32759 24636 32768
rect 24584 32725 24593 32759
rect 24593 32725 24627 32759
rect 24627 32725 24636 32759
rect 24584 32716 24636 32725
rect 25044 32716 25096 32768
rect 7950 32614 8002 32666
rect 8014 32614 8066 32666
rect 8078 32614 8130 32666
rect 8142 32614 8194 32666
rect 8206 32614 8258 32666
rect 17950 32614 18002 32666
rect 18014 32614 18066 32666
rect 18078 32614 18130 32666
rect 18142 32614 18194 32666
rect 18206 32614 18258 32666
rect 15384 32487 15436 32496
rect 15384 32453 15393 32487
rect 15393 32453 15427 32487
rect 15427 32453 15436 32487
rect 19616 32512 19668 32564
rect 21272 32512 21324 32564
rect 23572 32512 23624 32564
rect 25044 32512 25096 32564
rect 15384 32444 15436 32453
rect 19800 32444 19852 32496
rect 22284 32444 22336 32496
rect 21824 32376 21876 32428
rect 25504 32444 25556 32496
rect 25780 32444 25832 32496
rect 13360 32308 13412 32360
rect 16764 32308 16816 32360
rect 21180 32308 21232 32360
rect 24952 32308 25004 32360
rect 24860 32240 24912 32292
rect 25044 32240 25096 32292
rect 19432 32172 19484 32224
rect 20904 32172 20956 32224
rect 21824 32172 21876 32224
rect 22100 32172 22152 32224
rect 26792 32172 26844 32224
rect 2950 32070 3002 32122
rect 3014 32070 3066 32122
rect 3078 32070 3130 32122
rect 3142 32070 3194 32122
rect 3206 32070 3258 32122
rect 12950 32070 13002 32122
rect 13014 32070 13066 32122
rect 13078 32070 13130 32122
rect 13142 32070 13194 32122
rect 13206 32070 13258 32122
rect 22950 32070 23002 32122
rect 23014 32070 23066 32122
rect 23078 32070 23130 32122
rect 23142 32070 23194 32122
rect 23206 32070 23258 32122
rect 18512 31968 18564 32020
rect 12532 31900 12584 31952
rect 18052 31900 18104 31952
rect 22100 31968 22152 32020
rect 22468 31968 22520 32020
rect 23204 31968 23256 32020
rect 16120 31875 16172 31884
rect 16120 31841 16129 31875
rect 16129 31841 16163 31875
rect 16163 31841 16172 31875
rect 16120 31832 16172 31841
rect 17684 31832 17736 31884
rect 19708 31875 19760 31884
rect 19708 31841 19717 31875
rect 19717 31841 19751 31875
rect 19751 31841 19760 31875
rect 19708 31832 19760 31841
rect 21916 31832 21968 31884
rect 22744 31900 22796 31952
rect 23388 31900 23440 31952
rect 16764 31807 16816 31816
rect 16764 31773 16773 31807
rect 16773 31773 16807 31807
rect 16807 31773 16816 31807
rect 16764 31764 16816 31773
rect 19432 31807 19484 31816
rect 19432 31773 19441 31807
rect 19441 31773 19475 31807
rect 19475 31773 19484 31807
rect 19432 31764 19484 31773
rect 23020 31764 23072 31816
rect 25044 31900 25096 31952
rect 25320 31807 25372 31816
rect 25320 31773 25329 31807
rect 25329 31773 25363 31807
rect 25363 31773 25372 31807
rect 25320 31764 25372 31773
rect 16672 31696 16724 31748
rect 19800 31696 19852 31748
rect 23204 31696 23256 31748
rect 16488 31628 16540 31680
rect 20996 31628 21048 31680
rect 21640 31671 21692 31680
rect 21640 31637 21649 31671
rect 21649 31637 21683 31671
rect 21683 31637 21692 31671
rect 21640 31628 21692 31637
rect 21732 31628 21784 31680
rect 22008 31671 22060 31680
rect 22008 31637 22017 31671
rect 22017 31637 22051 31671
rect 22051 31637 22060 31671
rect 22008 31628 22060 31637
rect 22468 31628 22520 31680
rect 22652 31628 22704 31680
rect 24676 31671 24728 31680
rect 24676 31637 24685 31671
rect 24685 31637 24719 31671
rect 24719 31637 24728 31671
rect 24676 31628 24728 31637
rect 7950 31526 8002 31578
rect 8014 31526 8066 31578
rect 8078 31526 8130 31578
rect 8142 31526 8194 31578
rect 8206 31526 8258 31578
rect 17950 31526 18002 31578
rect 18014 31526 18066 31578
rect 18078 31526 18130 31578
rect 18142 31526 18194 31578
rect 18206 31526 18258 31578
rect 16488 31467 16540 31476
rect 16488 31433 16497 31467
rect 16497 31433 16531 31467
rect 16531 31433 16540 31467
rect 16488 31424 16540 31433
rect 17868 31424 17920 31476
rect 19708 31424 19760 31476
rect 21272 31467 21324 31476
rect 21272 31433 21281 31467
rect 21281 31433 21315 31467
rect 21315 31433 21324 31467
rect 21272 31424 21324 31433
rect 23572 31424 23624 31476
rect 14924 31356 14976 31408
rect 17776 31356 17828 31408
rect 20628 31356 20680 31408
rect 21364 31356 21416 31408
rect 22652 31356 22704 31408
rect 23020 31356 23072 31408
rect 24676 31356 24728 31408
rect 16764 31288 16816 31340
rect 19708 31288 19760 31340
rect 13360 31263 13412 31272
rect 13360 31229 13369 31263
rect 13369 31229 13403 31263
rect 13403 31229 13412 31263
rect 13360 31220 13412 31229
rect 16120 31220 16172 31272
rect 16672 31263 16724 31272
rect 16672 31229 16681 31263
rect 16681 31229 16715 31263
rect 16715 31229 16724 31263
rect 16672 31220 16724 31229
rect 17224 31220 17276 31272
rect 20444 31220 20496 31272
rect 20628 31263 20680 31272
rect 20628 31229 20637 31263
rect 20637 31229 20671 31263
rect 20671 31229 20680 31263
rect 20628 31220 20680 31229
rect 22008 31220 22060 31272
rect 22100 31220 22152 31272
rect 22284 31288 22336 31340
rect 25504 31288 25556 31340
rect 25136 31220 25188 31272
rect 12348 31084 12400 31136
rect 17500 31084 17552 31136
rect 23756 31152 23808 31204
rect 18788 31084 18840 31136
rect 20628 31084 20680 31136
rect 24676 31084 24728 31136
rect 25136 31127 25188 31136
rect 25136 31093 25145 31127
rect 25145 31093 25179 31127
rect 25179 31093 25188 31127
rect 25136 31084 25188 31093
rect 2950 30982 3002 31034
rect 3014 30982 3066 31034
rect 3078 30982 3130 31034
rect 3142 30982 3194 31034
rect 3206 30982 3258 31034
rect 12950 30982 13002 31034
rect 13014 30982 13066 31034
rect 13078 30982 13130 31034
rect 13142 30982 13194 31034
rect 13206 30982 13258 31034
rect 22950 30982 23002 31034
rect 23014 30982 23066 31034
rect 23078 30982 23130 31034
rect 23142 30982 23194 31034
rect 23206 30982 23258 31034
rect 9220 30880 9272 30932
rect 15384 30880 15436 30932
rect 18512 30923 18564 30932
rect 18512 30889 18521 30923
rect 18521 30889 18555 30923
rect 18555 30889 18564 30923
rect 18512 30880 18564 30889
rect 18788 30880 18840 30932
rect 18880 30880 18932 30932
rect 19708 30880 19760 30932
rect 22652 30880 22704 30932
rect 25504 30923 25556 30932
rect 25504 30889 25513 30923
rect 25513 30889 25547 30923
rect 25547 30889 25556 30923
rect 25504 30880 25556 30889
rect 19432 30744 19484 30796
rect 8760 30676 8812 30728
rect 14096 30676 14148 30728
rect 15384 30676 15436 30728
rect 15108 30651 15160 30660
rect 15108 30617 15117 30651
rect 15117 30617 15151 30651
rect 15151 30617 15160 30651
rect 15108 30608 15160 30617
rect 20996 30651 21048 30660
rect 20996 30617 21005 30651
rect 21005 30617 21039 30651
rect 21039 30617 21048 30651
rect 20996 30608 21048 30617
rect 21272 30608 21324 30660
rect 18696 30540 18748 30592
rect 18788 30583 18840 30592
rect 18788 30549 18797 30583
rect 18797 30549 18831 30583
rect 18831 30549 18840 30583
rect 18788 30540 18840 30549
rect 20076 30583 20128 30592
rect 20076 30549 20085 30583
rect 20085 30549 20119 30583
rect 20119 30549 20128 30583
rect 20076 30540 20128 30549
rect 22928 30540 22980 30592
rect 7950 30438 8002 30490
rect 8014 30438 8066 30490
rect 8078 30438 8130 30490
rect 8142 30438 8194 30490
rect 8206 30438 8258 30490
rect 17950 30438 18002 30490
rect 18014 30438 18066 30490
rect 18078 30438 18130 30490
rect 18142 30438 18194 30490
rect 18206 30438 18258 30490
rect 13360 30336 13412 30388
rect 8484 30200 8536 30252
rect 12716 30268 12768 30320
rect 14096 30311 14148 30320
rect 14096 30277 14105 30311
rect 14105 30277 14139 30311
rect 14139 30277 14148 30311
rect 14096 30268 14148 30277
rect 14556 30268 14608 30320
rect 20076 30336 20128 30388
rect 22652 30336 22704 30388
rect 23296 30336 23348 30388
rect 19984 30268 20036 30320
rect 21916 30268 21968 30320
rect 22560 30268 22612 30320
rect 16948 30243 17000 30252
rect 16948 30209 16957 30243
rect 16957 30209 16991 30243
rect 16991 30209 17000 30243
rect 16948 30200 17000 30209
rect 12072 30175 12124 30184
rect 12072 30141 12081 30175
rect 12081 30141 12115 30175
rect 12115 30141 12124 30175
rect 12072 30132 12124 30141
rect 13360 30132 13412 30184
rect 8944 30107 8996 30116
rect 8944 30073 8953 30107
rect 8953 30073 8987 30107
rect 8987 30073 8996 30107
rect 8944 30064 8996 30073
rect 16028 30175 16080 30184
rect 16028 30141 16037 30175
rect 16037 30141 16071 30175
rect 16071 30141 16080 30175
rect 16028 30132 16080 30141
rect 16764 30175 16816 30184
rect 16764 30141 16773 30175
rect 16773 30141 16807 30175
rect 16807 30141 16816 30175
rect 16764 30132 16816 30141
rect 20260 30132 20312 30184
rect 20536 30175 20588 30184
rect 20536 30141 20545 30175
rect 20545 30141 20579 30175
rect 20579 30141 20588 30175
rect 20536 30132 20588 30141
rect 24676 30200 24728 30252
rect 22284 30132 22336 30184
rect 22836 30132 22888 30184
rect 23296 30175 23348 30184
rect 23296 30141 23305 30175
rect 23305 30141 23339 30175
rect 23339 30141 23348 30175
rect 23296 30132 23348 30141
rect 23664 30132 23716 30184
rect 16488 30064 16540 30116
rect 22468 30064 22520 30116
rect 24952 30132 25004 30184
rect 11336 29996 11388 30048
rect 13636 29996 13688 30048
rect 15936 29996 15988 30048
rect 18788 29996 18840 30048
rect 19800 29996 19852 30048
rect 21916 29996 21968 30048
rect 2950 29894 3002 29946
rect 3014 29894 3066 29946
rect 3078 29894 3130 29946
rect 3142 29894 3194 29946
rect 3206 29894 3258 29946
rect 12950 29894 13002 29946
rect 13014 29894 13066 29946
rect 13078 29894 13130 29946
rect 13142 29894 13194 29946
rect 13206 29894 13258 29946
rect 22950 29894 23002 29946
rect 23014 29894 23066 29946
rect 23078 29894 23130 29946
rect 23142 29894 23194 29946
rect 23206 29894 23258 29946
rect 12072 29792 12124 29844
rect 16488 29835 16540 29844
rect 16488 29801 16497 29835
rect 16497 29801 16531 29835
rect 16531 29801 16540 29835
rect 16488 29792 16540 29801
rect 18696 29792 18748 29844
rect 11428 29656 11480 29708
rect 13360 29656 13412 29708
rect 18420 29724 18472 29776
rect 20260 29724 20312 29776
rect 26516 29792 26568 29844
rect 23204 29724 23256 29776
rect 16028 29656 16080 29708
rect 19340 29656 19392 29708
rect 16488 29588 16540 29640
rect 18880 29588 18932 29640
rect 11060 29520 11112 29572
rect 12716 29520 12768 29572
rect 13728 29520 13780 29572
rect 15568 29563 15620 29572
rect 15568 29529 15577 29563
rect 15577 29529 15611 29563
rect 15611 29529 15620 29563
rect 15568 29520 15620 29529
rect 15200 29495 15252 29504
rect 15200 29461 15209 29495
rect 15209 29461 15243 29495
rect 15243 29461 15252 29495
rect 15200 29452 15252 29461
rect 16304 29495 16356 29504
rect 16304 29461 16313 29495
rect 16313 29461 16347 29495
rect 16347 29461 16356 29495
rect 16304 29452 16356 29461
rect 18788 29520 18840 29572
rect 20720 29520 20772 29572
rect 24492 29588 24544 29640
rect 25320 29631 25372 29640
rect 25320 29597 25329 29631
rect 25329 29597 25363 29631
rect 25363 29597 25372 29631
rect 25320 29588 25372 29597
rect 24952 29520 25004 29572
rect 18880 29452 18932 29504
rect 19156 29452 19208 29504
rect 19984 29452 20036 29504
rect 22652 29452 22704 29504
rect 24308 29452 24360 29504
rect 24492 29495 24544 29504
rect 24492 29461 24501 29495
rect 24501 29461 24535 29495
rect 24535 29461 24544 29495
rect 24492 29452 24544 29461
rect 7950 29350 8002 29402
rect 8014 29350 8066 29402
rect 8078 29350 8130 29402
rect 8142 29350 8194 29402
rect 8206 29350 8258 29402
rect 17950 29350 18002 29402
rect 18014 29350 18066 29402
rect 18078 29350 18130 29402
rect 18142 29350 18194 29402
rect 18206 29350 18258 29402
rect 8852 29248 8904 29300
rect 12532 29291 12584 29300
rect 12532 29257 12541 29291
rect 12541 29257 12575 29291
rect 12575 29257 12584 29291
rect 12532 29248 12584 29257
rect 12624 29291 12676 29300
rect 12624 29257 12633 29291
rect 12633 29257 12667 29291
rect 12667 29257 12676 29291
rect 12624 29248 12676 29257
rect 13452 29248 13504 29300
rect 10324 29180 10376 29232
rect 14924 29180 14976 29232
rect 15200 29248 15252 29300
rect 16304 29248 16356 29300
rect 15844 29180 15896 29232
rect 15936 29223 15988 29232
rect 15936 29189 15945 29223
rect 15945 29189 15979 29223
rect 15979 29189 15988 29223
rect 15936 29180 15988 29189
rect 17132 29180 17184 29232
rect 17408 29248 17460 29300
rect 19156 29291 19208 29300
rect 19156 29257 19165 29291
rect 19165 29257 19199 29291
rect 19199 29257 19208 29291
rect 19156 29248 19208 29257
rect 19432 29248 19484 29300
rect 19984 29291 20036 29300
rect 19984 29257 19993 29291
rect 19993 29257 20027 29291
rect 20027 29257 20036 29291
rect 19984 29248 20036 29257
rect 20168 29248 20220 29300
rect 24124 29248 24176 29300
rect 24768 29248 24820 29300
rect 25320 29248 25372 29300
rect 10232 29112 10284 29164
rect 13360 29155 13412 29164
rect 13360 29121 13369 29155
rect 13369 29121 13403 29155
rect 13403 29121 13412 29155
rect 13360 29112 13412 29121
rect 9680 29044 9732 29096
rect 10876 29044 10928 29096
rect 11152 29044 11204 29096
rect 12348 29044 12400 29096
rect 13636 29044 13688 29096
rect 17316 29087 17368 29096
rect 17316 29053 17325 29087
rect 17325 29053 17359 29087
rect 17359 29053 17368 29087
rect 17316 29044 17368 29053
rect 17408 29087 17460 29096
rect 17408 29053 17417 29087
rect 17417 29053 17451 29087
rect 17451 29053 17460 29087
rect 17408 29044 17460 29053
rect 20904 29044 20956 29096
rect 12256 28976 12308 29028
rect 14096 28908 14148 28960
rect 14188 28908 14240 28960
rect 15752 28976 15804 29028
rect 17500 28976 17552 29028
rect 19064 28976 19116 29028
rect 21824 29019 21876 29028
rect 21824 28985 21833 29019
rect 21833 28985 21867 29019
rect 21867 28985 21876 29019
rect 23388 29044 23440 29096
rect 26424 29180 26476 29232
rect 26884 29112 26936 29164
rect 24216 29087 24268 29096
rect 24216 29053 24225 29087
rect 24225 29053 24259 29087
rect 24259 29053 24268 29087
rect 24216 29044 24268 29053
rect 24952 29044 25004 29096
rect 21824 28976 21876 28985
rect 24400 28976 24452 29028
rect 22100 28908 22152 28960
rect 22468 28908 22520 28960
rect 25228 28951 25280 28960
rect 25228 28917 25237 28951
rect 25237 28917 25271 28951
rect 25271 28917 25280 28951
rect 25228 28908 25280 28917
rect 2950 28806 3002 28858
rect 3014 28806 3066 28858
rect 3078 28806 3130 28858
rect 3142 28806 3194 28858
rect 3206 28806 3258 28858
rect 12950 28806 13002 28858
rect 13014 28806 13066 28858
rect 13078 28806 13130 28858
rect 13142 28806 13194 28858
rect 13206 28806 13258 28858
rect 22950 28806 23002 28858
rect 23014 28806 23066 28858
rect 23078 28806 23130 28858
rect 23142 28806 23194 28858
rect 23206 28806 23258 28858
rect 10876 28747 10928 28756
rect 10876 28713 10885 28747
rect 10885 28713 10919 28747
rect 10919 28713 10928 28747
rect 10876 28704 10928 28713
rect 13728 28704 13780 28756
rect 15016 28704 15068 28756
rect 18788 28704 18840 28756
rect 18880 28747 18932 28756
rect 18880 28713 18889 28747
rect 18889 28713 18923 28747
rect 18923 28713 18932 28747
rect 18880 28704 18932 28713
rect 21088 28704 21140 28756
rect 11428 28611 11480 28620
rect 11428 28577 11437 28611
rect 11437 28577 11471 28611
rect 11471 28577 11480 28611
rect 11428 28568 11480 28577
rect 14096 28568 14148 28620
rect 16212 28636 16264 28688
rect 22560 28636 22612 28688
rect 25504 28704 25556 28756
rect 15384 28611 15436 28620
rect 15384 28577 15393 28611
rect 15393 28577 15427 28611
rect 15427 28577 15436 28611
rect 15384 28568 15436 28577
rect 18972 28568 19024 28620
rect 20996 28568 21048 28620
rect 21456 28568 21508 28620
rect 25412 28636 25464 28688
rect 15108 28500 15160 28552
rect 19340 28500 19392 28552
rect 20628 28543 20680 28552
rect 20628 28509 20637 28543
rect 20637 28509 20671 28543
rect 20671 28509 20680 28543
rect 20628 28500 20680 28509
rect 23572 28568 23624 28620
rect 24860 28568 24912 28620
rect 23940 28500 23992 28552
rect 24584 28500 24636 28552
rect 24952 28543 25004 28552
rect 24952 28509 24961 28543
rect 24961 28509 24995 28543
rect 24995 28509 25004 28543
rect 24952 28500 25004 28509
rect 11336 28432 11388 28484
rect 9772 28364 9824 28416
rect 11244 28364 11296 28416
rect 12624 28364 12676 28416
rect 13728 28432 13780 28484
rect 18788 28432 18840 28484
rect 20904 28475 20956 28484
rect 20904 28441 20913 28475
rect 20913 28441 20947 28475
rect 20947 28441 20956 28475
rect 20904 28432 20956 28441
rect 21456 28432 21508 28484
rect 14832 28407 14884 28416
rect 14832 28373 14841 28407
rect 14841 28373 14875 28407
rect 14875 28373 14884 28407
rect 14832 28364 14884 28373
rect 16028 28407 16080 28416
rect 16028 28373 16037 28407
rect 16037 28373 16071 28407
rect 16071 28373 16080 28407
rect 16028 28364 16080 28373
rect 16212 28407 16264 28416
rect 16212 28373 16221 28407
rect 16221 28373 16255 28407
rect 16255 28373 16264 28407
rect 16212 28364 16264 28373
rect 19524 28364 19576 28416
rect 19708 28364 19760 28416
rect 21640 28364 21692 28416
rect 24216 28432 24268 28484
rect 22468 28364 22520 28416
rect 24492 28364 24544 28416
rect 7950 28262 8002 28314
rect 8014 28262 8066 28314
rect 8078 28262 8130 28314
rect 8142 28262 8194 28314
rect 8206 28262 8258 28314
rect 17950 28262 18002 28314
rect 18014 28262 18066 28314
rect 18078 28262 18130 28314
rect 18142 28262 18194 28314
rect 18206 28262 18258 28314
rect 3424 28160 3476 28212
rect 11244 28092 11296 28144
rect 13728 28135 13780 28144
rect 13728 28101 13737 28135
rect 13737 28101 13771 28135
rect 13771 28101 13780 28135
rect 13728 28092 13780 28101
rect 15936 28092 15988 28144
rect 16396 28135 16448 28144
rect 16396 28101 16405 28135
rect 16405 28101 16439 28135
rect 16439 28101 16448 28135
rect 16396 28092 16448 28101
rect 17224 28135 17276 28144
rect 17224 28101 17233 28135
rect 17233 28101 17267 28135
rect 17267 28101 17276 28135
rect 17224 28092 17276 28101
rect 18788 28160 18840 28212
rect 19708 28203 19760 28212
rect 19708 28169 19717 28203
rect 19717 28169 19751 28203
rect 19751 28169 19760 28203
rect 19708 28160 19760 28169
rect 20628 28092 20680 28144
rect 26240 28160 26292 28212
rect 22560 28092 22612 28144
rect 15660 28067 15712 28076
rect 15660 28033 15669 28067
rect 15669 28033 15703 28067
rect 15703 28033 15712 28067
rect 15660 28024 15712 28033
rect 16304 28024 16356 28076
rect 17868 28024 17920 28076
rect 11704 27999 11756 28008
rect 11704 27965 11713 27999
rect 11713 27965 11747 27999
rect 11747 27965 11756 27999
rect 11704 27956 11756 27965
rect 11980 27999 12032 28008
rect 11980 27965 11989 27999
rect 11989 27965 12023 27999
rect 12023 27965 12032 27999
rect 11980 27956 12032 27965
rect 10784 27888 10836 27940
rect 15384 27888 15436 27940
rect 17408 27999 17460 28008
rect 17408 27965 17417 27999
rect 17417 27965 17451 27999
rect 17451 27965 17460 27999
rect 17408 27956 17460 27965
rect 17960 27956 18012 28008
rect 18788 27956 18840 28008
rect 17684 27888 17736 27940
rect 21824 28024 21876 28076
rect 23388 28092 23440 28144
rect 23940 28092 23992 28144
rect 22560 27999 22612 28008
rect 22560 27965 22569 27999
rect 22569 27965 22603 27999
rect 22603 27965 22612 27999
rect 22560 27956 22612 27965
rect 23480 27999 23532 28008
rect 23480 27965 23489 27999
rect 23489 27965 23523 27999
rect 23523 27965 23532 27999
rect 23480 27956 23532 27965
rect 23940 27956 23992 28008
rect 25228 27999 25280 28008
rect 25228 27965 25237 27999
rect 25237 27965 25271 27999
rect 25271 27965 25280 27999
rect 25228 27956 25280 27965
rect 13820 27820 13872 27872
rect 16304 27863 16356 27872
rect 16304 27829 16313 27863
rect 16313 27829 16347 27863
rect 16347 27829 16356 27863
rect 16304 27820 16356 27829
rect 16856 27863 16908 27872
rect 16856 27829 16865 27863
rect 16865 27829 16899 27863
rect 16899 27829 16908 27863
rect 16856 27820 16908 27829
rect 17224 27820 17276 27872
rect 18512 27820 18564 27872
rect 20720 27820 20772 27872
rect 22376 27820 22428 27872
rect 25412 27863 25464 27872
rect 25412 27829 25421 27863
rect 25421 27829 25455 27863
rect 25455 27829 25464 27863
rect 25412 27820 25464 27829
rect 2950 27718 3002 27770
rect 3014 27718 3066 27770
rect 3078 27718 3130 27770
rect 3142 27718 3194 27770
rect 3206 27718 3258 27770
rect 12950 27718 13002 27770
rect 13014 27718 13066 27770
rect 13078 27718 13130 27770
rect 13142 27718 13194 27770
rect 13206 27718 13258 27770
rect 22950 27718 23002 27770
rect 23014 27718 23066 27770
rect 23078 27718 23130 27770
rect 23142 27718 23194 27770
rect 23206 27718 23258 27770
rect 11428 27616 11480 27668
rect 11796 27616 11848 27668
rect 10784 27523 10836 27532
rect 10784 27489 10793 27523
rect 10793 27489 10827 27523
rect 10827 27489 10836 27523
rect 10784 27480 10836 27489
rect 12440 27548 12492 27600
rect 12624 27591 12676 27600
rect 12624 27557 12633 27591
rect 12633 27557 12667 27591
rect 12667 27557 12676 27591
rect 12624 27548 12676 27557
rect 13084 27548 13136 27600
rect 15108 27616 15160 27668
rect 23572 27616 23624 27668
rect 23480 27548 23532 27600
rect 24768 27548 24820 27600
rect 9588 27276 9640 27328
rect 15108 27480 15160 27532
rect 17776 27480 17828 27532
rect 23388 27480 23440 27532
rect 24124 27523 24176 27532
rect 24124 27489 24133 27523
rect 24133 27489 24167 27523
rect 24167 27489 24176 27523
rect 24124 27480 24176 27489
rect 25044 27523 25096 27532
rect 25044 27489 25053 27523
rect 25053 27489 25087 27523
rect 25087 27489 25096 27523
rect 25044 27480 25096 27489
rect 14832 27412 14884 27464
rect 16212 27412 16264 27464
rect 17960 27412 18012 27464
rect 23940 27412 23992 27464
rect 25412 27412 25464 27464
rect 13820 27344 13872 27396
rect 21456 27344 21508 27396
rect 21824 27344 21876 27396
rect 22376 27387 22428 27396
rect 22376 27353 22385 27387
rect 22385 27353 22419 27387
rect 22419 27353 22428 27387
rect 22376 27344 22428 27353
rect 12624 27276 12676 27328
rect 13728 27276 13780 27328
rect 16028 27276 16080 27328
rect 16488 27276 16540 27328
rect 17592 27276 17644 27328
rect 21640 27319 21692 27328
rect 21640 27285 21649 27319
rect 21649 27285 21683 27319
rect 21683 27285 21692 27319
rect 21640 27276 21692 27285
rect 24584 27319 24636 27328
rect 24584 27285 24593 27319
rect 24593 27285 24627 27319
rect 24627 27285 24636 27319
rect 24584 27276 24636 27285
rect 24860 27276 24912 27328
rect 25320 27276 25372 27328
rect 7950 27174 8002 27226
rect 8014 27174 8066 27226
rect 8078 27174 8130 27226
rect 8142 27174 8194 27226
rect 8206 27174 8258 27226
rect 17950 27174 18002 27226
rect 18014 27174 18066 27226
rect 18078 27174 18130 27226
rect 18142 27174 18194 27226
rect 18206 27174 18258 27226
rect 11060 27115 11112 27124
rect 11060 27081 11069 27115
rect 11069 27081 11103 27115
rect 11103 27081 11112 27115
rect 11060 27072 11112 27081
rect 9588 27047 9640 27056
rect 9588 27013 9597 27047
rect 9597 27013 9631 27047
rect 9631 27013 9640 27047
rect 9588 27004 9640 27013
rect 11244 27004 11296 27056
rect 12440 27072 12492 27124
rect 13544 27072 13596 27124
rect 13452 27004 13504 27056
rect 16856 27072 16908 27124
rect 15752 27047 15804 27056
rect 15752 27013 15761 27047
rect 15761 27013 15795 27047
rect 15795 27013 15804 27047
rect 15752 27004 15804 27013
rect 19248 27072 19300 27124
rect 22744 27072 22796 27124
rect 12716 26936 12768 26988
rect 13084 26979 13136 26988
rect 13084 26945 13093 26979
rect 13093 26945 13127 26979
rect 13127 26945 13136 26979
rect 13084 26936 13136 26945
rect 14740 26936 14792 26988
rect 16764 26936 16816 26988
rect 20076 27004 20128 27056
rect 22928 26936 22980 26988
rect 22100 26868 22152 26920
rect 22560 26868 22612 26920
rect 23664 27072 23716 27124
rect 24768 27072 24820 27124
rect 23940 27004 23992 27056
rect 25228 27004 25280 27056
rect 25504 27004 25556 27056
rect 25780 26936 25832 26988
rect 26056 26936 26108 26988
rect 23388 26868 23440 26920
rect 25504 26868 25556 26920
rect 9680 26732 9732 26784
rect 12072 26732 12124 26784
rect 22468 26800 22520 26852
rect 22836 26800 22888 26852
rect 14924 26732 14976 26784
rect 18972 26732 19024 26784
rect 20076 26775 20128 26784
rect 20076 26741 20085 26775
rect 20085 26741 20119 26775
rect 20119 26741 20128 26775
rect 21824 26775 21876 26784
rect 20076 26732 20128 26741
rect 21824 26741 21833 26775
rect 21833 26741 21867 26775
rect 21867 26741 21876 26775
rect 21824 26732 21876 26741
rect 22192 26732 22244 26784
rect 2950 26630 3002 26682
rect 3014 26630 3066 26682
rect 3078 26630 3130 26682
rect 3142 26630 3194 26682
rect 3206 26630 3258 26682
rect 12950 26630 13002 26682
rect 13014 26630 13066 26682
rect 13078 26630 13130 26682
rect 13142 26630 13194 26682
rect 13206 26630 13258 26682
rect 22950 26630 23002 26682
rect 23014 26630 23066 26682
rect 23078 26630 23130 26682
rect 23142 26630 23194 26682
rect 23206 26630 23258 26682
rect 11980 26528 12032 26580
rect 12348 26528 12400 26580
rect 13544 26528 13596 26580
rect 16948 26571 17000 26580
rect 16948 26537 16957 26571
rect 16957 26537 16991 26571
rect 16991 26537 17000 26571
rect 16948 26528 17000 26537
rect 22100 26528 22152 26580
rect 24952 26528 25004 26580
rect 11244 26503 11296 26512
rect 11244 26469 11253 26503
rect 11253 26469 11287 26503
rect 11287 26469 11296 26503
rect 11244 26460 11296 26469
rect 13636 26460 13688 26512
rect 15936 26460 15988 26512
rect 17224 26503 17276 26512
rect 17224 26469 17233 26503
rect 17233 26469 17267 26503
rect 17267 26469 17276 26503
rect 17224 26460 17276 26469
rect 22468 26460 22520 26512
rect 25044 26460 25096 26512
rect 7748 26392 7800 26444
rect 11152 26392 11204 26444
rect 14464 26392 14516 26444
rect 14740 26435 14792 26444
rect 14740 26401 14749 26435
rect 14749 26401 14783 26435
rect 14783 26401 14792 26435
rect 14740 26392 14792 26401
rect 14832 26435 14884 26444
rect 14832 26401 14841 26435
rect 14841 26401 14875 26435
rect 14875 26401 14884 26435
rect 14832 26392 14884 26401
rect 15108 26392 15160 26444
rect 16764 26435 16816 26444
rect 16764 26401 16773 26435
rect 16773 26401 16807 26435
rect 16807 26401 16816 26435
rect 16764 26392 16816 26401
rect 19432 26435 19484 26444
rect 19432 26401 19441 26435
rect 19441 26401 19475 26435
rect 19475 26401 19484 26435
rect 19432 26392 19484 26401
rect 20996 26392 21048 26444
rect 21640 26392 21692 26444
rect 22376 26392 22428 26444
rect 10968 26324 11020 26376
rect 12716 26324 12768 26376
rect 9680 26256 9732 26308
rect 11244 26256 11296 26308
rect 11796 26256 11848 26308
rect 16948 26324 17000 26376
rect 23296 26324 23348 26376
rect 24032 26367 24084 26376
rect 24032 26333 24041 26367
rect 24041 26333 24075 26367
rect 24075 26333 24084 26367
rect 24032 26324 24084 26333
rect 25228 26528 25280 26580
rect 25596 26528 25648 26580
rect 25872 26528 25924 26580
rect 25228 26435 25280 26444
rect 25228 26401 25237 26435
rect 25237 26401 25271 26435
rect 25271 26401 25280 26435
rect 25228 26392 25280 26401
rect 25596 26324 25648 26376
rect 10876 26188 10928 26240
rect 15936 26256 15988 26308
rect 16304 26256 16356 26308
rect 17408 26256 17460 26308
rect 21088 26256 21140 26308
rect 21824 26256 21876 26308
rect 22836 26256 22888 26308
rect 23480 26256 23532 26308
rect 24584 26256 24636 26308
rect 25136 26256 25188 26308
rect 18328 26188 18380 26240
rect 7950 26086 8002 26138
rect 8014 26086 8066 26138
rect 8078 26086 8130 26138
rect 8142 26086 8194 26138
rect 8206 26086 8258 26138
rect 17950 26086 18002 26138
rect 18014 26086 18066 26138
rect 18078 26086 18130 26138
rect 18142 26086 18194 26138
rect 18206 26086 18258 26138
rect 12624 26027 12676 26036
rect 12624 25993 12633 26027
rect 12633 25993 12667 26027
rect 12667 25993 12676 26027
rect 12624 25984 12676 25993
rect 13820 25984 13872 26036
rect 9680 25916 9732 25968
rect 12532 25891 12584 25900
rect 12532 25857 12541 25891
rect 12541 25857 12575 25891
rect 12575 25857 12584 25891
rect 12532 25848 12584 25857
rect 14188 25848 14240 25900
rect 11060 25780 11112 25832
rect 14004 25823 14056 25832
rect 14004 25789 14013 25823
rect 14013 25789 14047 25823
rect 14047 25789 14056 25823
rect 14004 25780 14056 25789
rect 14096 25823 14148 25832
rect 14096 25789 14105 25823
rect 14105 25789 14139 25823
rect 14139 25789 14148 25823
rect 14096 25780 14148 25789
rect 16304 25984 16356 26036
rect 18328 25984 18380 26036
rect 19156 25984 19208 26036
rect 22284 25984 22336 26036
rect 22652 25984 22704 26036
rect 18420 25916 18472 25968
rect 16580 25848 16632 25900
rect 17592 25848 17644 25900
rect 18696 25780 18748 25832
rect 21456 25848 21508 25900
rect 25412 25984 25464 26036
rect 24860 25916 24912 25968
rect 23940 25891 23992 25900
rect 23940 25857 23949 25891
rect 23949 25857 23983 25891
rect 23983 25857 23992 25891
rect 23940 25848 23992 25857
rect 17592 25712 17644 25764
rect 19984 25712 20036 25764
rect 22560 25823 22612 25832
rect 22560 25789 22569 25823
rect 22569 25789 22603 25823
rect 22603 25789 22612 25823
rect 22560 25780 22612 25789
rect 25136 25823 25188 25832
rect 25136 25789 25145 25823
rect 25145 25789 25179 25823
rect 25179 25789 25188 25823
rect 25136 25780 25188 25789
rect 24768 25712 24820 25764
rect 16580 25644 16632 25696
rect 16856 25687 16908 25696
rect 16856 25653 16865 25687
rect 16865 25653 16899 25687
rect 16899 25653 16908 25687
rect 16856 25644 16908 25653
rect 18604 25644 18656 25696
rect 19156 25644 19208 25696
rect 21456 25644 21508 25696
rect 23296 25687 23348 25696
rect 23296 25653 23305 25687
rect 23305 25653 23339 25687
rect 23339 25653 23348 25687
rect 23296 25644 23348 25653
rect 2950 25542 3002 25594
rect 3014 25542 3066 25594
rect 3078 25542 3130 25594
rect 3142 25542 3194 25594
rect 3206 25542 3258 25594
rect 12950 25542 13002 25594
rect 13014 25542 13066 25594
rect 13078 25542 13130 25594
rect 13142 25542 13194 25594
rect 13206 25542 13258 25594
rect 22950 25542 23002 25594
rect 23014 25542 23066 25594
rect 23078 25542 23130 25594
rect 23142 25542 23194 25594
rect 23206 25542 23258 25594
rect 11704 25440 11756 25492
rect 15568 25440 15620 25492
rect 12992 25415 13044 25424
rect 12992 25381 13001 25415
rect 13001 25381 13035 25415
rect 13035 25381 13044 25415
rect 12992 25372 13044 25381
rect 13544 25372 13596 25424
rect 15108 25372 15160 25424
rect 10876 25347 10928 25356
rect 10876 25313 10885 25347
rect 10885 25313 10919 25347
rect 10919 25313 10928 25347
rect 10876 25304 10928 25313
rect 14740 25304 14792 25356
rect 14832 25347 14884 25356
rect 14832 25313 14841 25347
rect 14841 25313 14875 25347
rect 14875 25313 14884 25347
rect 14832 25304 14884 25313
rect 13360 25236 13412 25288
rect 12992 25168 13044 25220
rect 15568 25168 15620 25220
rect 18512 25440 18564 25492
rect 20076 25440 20128 25492
rect 23940 25440 23992 25492
rect 24860 25440 24912 25492
rect 16856 25304 16908 25356
rect 17132 25279 17184 25288
rect 17132 25245 17141 25279
rect 17141 25245 17175 25279
rect 17175 25245 17184 25279
rect 17132 25236 17184 25245
rect 17592 25236 17644 25288
rect 18604 25236 18656 25288
rect 24032 25372 24084 25424
rect 25320 25279 25372 25288
rect 25320 25245 25329 25279
rect 25329 25245 25363 25279
rect 25363 25245 25372 25279
rect 25320 25236 25372 25245
rect 12624 25143 12676 25152
rect 12624 25109 12633 25143
rect 12633 25109 12667 25143
rect 12667 25109 12676 25143
rect 12624 25100 12676 25109
rect 15384 25100 15436 25152
rect 15752 25143 15804 25152
rect 15752 25109 15761 25143
rect 15761 25109 15795 25143
rect 15795 25109 15804 25143
rect 15752 25100 15804 25109
rect 16212 25143 16264 25152
rect 16212 25109 16221 25143
rect 16221 25109 16255 25143
rect 16255 25109 16264 25143
rect 16212 25100 16264 25109
rect 19156 25168 19208 25220
rect 18512 25100 18564 25152
rect 19892 25143 19944 25152
rect 19892 25109 19901 25143
rect 19901 25109 19935 25143
rect 19935 25109 19944 25143
rect 19892 25100 19944 25109
rect 23848 25211 23900 25220
rect 23848 25177 23857 25211
rect 23857 25177 23891 25211
rect 23891 25177 23900 25211
rect 23848 25168 23900 25177
rect 25412 25168 25464 25220
rect 23756 25100 23808 25152
rect 25136 25143 25188 25152
rect 25136 25109 25145 25143
rect 25145 25109 25179 25143
rect 25179 25109 25188 25143
rect 25136 25100 25188 25109
rect 7950 24998 8002 25050
rect 8014 24998 8066 25050
rect 8078 24998 8130 25050
rect 8142 24998 8194 25050
rect 8206 24998 8258 25050
rect 17950 24998 18002 25050
rect 18014 24998 18066 25050
rect 18078 24998 18130 25050
rect 18142 24998 18194 25050
rect 18206 24998 18258 25050
rect 10140 24828 10192 24880
rect 11244 24828 11296 24880
rect 13544 24828 13596 24880
rect 12256 24760 12308 24812
rect 12716 24760 12768 24812
rect 17132 24896 17184 24948
rect 17224 24939 17276 24948
rect 17224 24905 17233 24939
rect 17233 24905 17267 24939
rect 17267 24905 17276 24939
rect 17224 24896 17276 24905
rect 18328 24896 18380 24948
rect 16212 24828 16264 24880
rect 18604 24828 18656 24880
rect 24124 24828 24176 24880
rect 25412 24828 25464 24880
rect 11152 24692 11204 24744
rect 12348 24735 12400 24744
rect 12348 24701 12357 24735
rect 12357 24701 12391 24735
rect 12391 24701 12400 24735
rect 12348 24692 12400 24701
rect 13912 24692 13964 24744
rect 10876 24624 10928 24676
rect 11060 24556 11112 24608
rect 15384 24803 15436 24812
rect 15384 24769 15393 24803
rect 15393 24769 15427 24803
rect 15427 24769 15436 24803
rect 15384 24760 15436 24769
rect 16396 24760 16448 24812
rect 14740 24735 14792 24744
rect 14740 24701 14749 24735
rect 14749 24701 14783 24735
rect 14783 24701 14792 24735
rect 14740 24692 14792 24701
rect 15016 24692 15068 24744
rect 18420 24803 18472 24812
rect 18420 24769 18429 24803
rect 18429 24769 18463 24803
rect 18463 24769 18472 24803
rect 18420 24760 18472 24769
rect 18696 24760 18748 24812
rect 19432 24760 19484 24812
rect 21088 24760 21140 24812
rect 23480 24760 23532 24812
rect 17040 24624 17092 24676
rect 20444 24692 20496 24744
rect 22376 24692 22428 24744
rect 22652 24735 22704 24744
rect 22652 24701 22661 24735
rect 22661 24701 22695 24735
rect 22695 24701 22704 24735
rect 22652 24692 22704 24701
rect 22192 24624 22244 24676
rect 23388 24624 23440 24676
rect 25228 24692 25280 24744
rect 25504 24692 25556 24744
rect 14740 24556 14792 24608
rect 15476 24556 15528 24608
rect 17868 24556 17920 24608
rect 22376 24556 22428 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 10876 24352 10928 24404
rect 14832 24352 14884 24404
rect 20444 24352 20496 24404
rect 25320 24395 25372 24404
rect 25320 24361 25329 24395
rect 25329 24361 25363 24395
rect 25363 24361 25372 24395
rect 25320 24352 25372 24361
rect 13544 24284 13596 24336
rect 14740 24284 14792 24336
rect 25596 24284 25648 24336
rect 10140 24216 10192 24268
rect 7840 24148 7892 24200
rect 11060 24216 11112 24268
rect 12348 24216 12400 24268
rect 18972 24216 19024 24268
rect 19432 24259 19484 24268
rect 19432 24225 19441 24259
rect 19441 24225 19475 24259
rect 19475 24225 19484 24259
rect 19432 24216 19484 24225
rect 22192 24216 22244 24268
rect 24124 24216 24176 24268
rect 17684 24191 17736 24200
rect 17684 24157 17693 24191
rect 17693 24157 17727 24191
rect 17727 24157 17736 24191
rect 17684 24148 17736 24157
rect 18512 24191 18564 24200
rect 18512 24157 18521 24191
rect 18521 24157 18555 24191
rect 18555 24157 18564 24191
rect 18512 24148 18564 24157
rect 9312 24080 9364 24132
rect 10140 24080 10192 24132
rect 11060 24012 11112 24064
rect 11980 24080 12032 24132
rect 18880 24080 18932 24132
rect 19708 24123 19760 24132
rect 19708 24089 19717 24123
rect 19717 24089 19751 24123
rect 19751 24089 19760 24123
rect 19708 24080 19760 24089
rect 21088 24080 21140 24132
rect 22284 24080 22336 24132
rect 12624 24012 12676 24064
rect 12900 24012 12952 24064
rect 13912 24012 13964 24064
rect 18420 24012 18472 24064
rect 20720 24012 20772 24064
rect 21548 24055 21600 24064
rect 21548 24021 21557 24055
rect 21557 24021 21591 24055
rect 21591 24021 21600 24055
rect 21548 24012 21600 24021
rect 23572 24012 23624 24064
rect 25320 24012 25372 24064
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 9772 23851 9824 23860
rect 9772 23817 9781 23851
rect 9781 23817 9815 23851
rect 9815 23817 9824 23851
rect 9772 23808 9824 23817
rect 10324 23808 10376 23860
rect 13820 23808 13872 23860
rect 7840 23672 7892 23724
rect 9680 23604 9732 23656
rect 13636 23783 13688 23792
rect 13636 23749 13645 23783
rect 13645 23749 13679 23783
rect 13679 23749 13688 23783
rect 13636 23740 13688 23749
rect 13728 23783 13780 23792
rect 13728 23749 13737 23783
rect 13737 23749 13771 23783
rect 13771 23749 13780 23783
rect 13728 23740 13780 23749
rect 14924 23851 14976 23860
rect 14924 23817 14933 23851
rect 14933 23817 14967 23851
rect 14967 23817 14976 23851
rect 14924 23808 14976 23817
rect 16764 23808 16816 23860
rect 18144 23808 18196 23860
rect 18236 23808 18288 23860
rect 18696 23808 18748 23860
rect 18880 23851 18932 23860
rect 18880 23817 18889 23851
rect 18889 23817 18923 23851
rect 18923 23817 18932 23851
rect 18880 23808 18932 23817
rect 19156 23808 19208 23860
rect 14004 23672 14056 23724
rect 17316 23715 17368 23724
rect 17316 23681 17325 23715
rect 17325 23681 17359 23715
rect 17359 23681 17368 23715
rect 19708 23740 19760 23792
rect 17316 23672 17368 23681
rect 10048 23604 10100 23656
rect 10968 23647 11020 23656
rect 10968 23613 10977 23647
rect 10977 23613 11011 23647
rect 11011 23613 11020 23647
rect 10968 23604 11020 23613
rect 12900 23536 12952 23588
rect 13912 23604 13964 23656
rect 15660 23647 15712 23656
rect 15660 23613 15669 23647
rect 15669 23613 15703 23647
rect 15703 23613 15712 23647
rect 15660 23604 15712 23613
rect 16580 23604 16632 23656
rect 19616 23715 19668 23724
rect 19616 23681 19625 23715
rect 19625 23681 19659 23715
rect 19659 23681 19668 23715
rect 19616 23672 19668 23681
rect 20168 23672 20220 23724
rect 14556 23536 14608 23588
rect 19340 23604 19392 23656
rect 19708 23647 19760 23656
rect 19708 23613 19717 23647
rect 19717 23613 19751 23647
rect 19751 23613 19760 23647
rect 19708 23604 19760 23613
rect 20812 23715 20864 23724
rect 20812 23681 20821 23715
rect 20821 23681 20855 23715
rect 20855 23681 20864 23715
rect 20812 23672 20864 23681
rect 22560 23740 22612 23792
rect 22284 23672 22336 23724
rect 25228 23808 25280 23860
rect 25596 23808 25648 23860
rect 25228 23672 25280 23724
rect 20904 23647 20956 23656
rect 20904 23613 20913 23647
rect 20913 23613 20947 23647
rect 20947 23613 20956 23647
rect 20904 23604 20956 23613
rect 20996 23647 21048 23656
rect 20996 23613 21005 23647
rect 21005 23613 21039 23647
rect 21039 23613 21048 23647
rect 20996 23604 21048 23613
rect 22192 23604 22244 23656
rect 23572 23604 23624 23656
rect 10140 23511 10192 23520
rect 10140 23477 10149 23511
rect 10149 23477 10183 23511
rect 10183 23477 10192 23511
rect 10140 23468 10192 23477
rect 12440 23468 12492 23520
rect 17316 23468 17368 23520
rect 18144 23468 18196 23520
rect 19156 23468 19208 23520
rect 19248 23511 19300 23520
rect 19248 23477 19257 23511
rect 19257 23477 19291 23511
rect 19291 23477 19300 23511
rect 19248 23468 19300 23477
rect 19340 23468 19392 23520
rect 20260 23468 20312 23520
rect 20628 23468 20680 23520
rect 21548 23511 21600 23520
rect 21548 23477 21557 23511
rect 21557 23477 21591 23511
rect 21591 23477 21600 23511
rect 21548 23468 21600 23477
rect 22836 23468 22888 23520
rect 23940 23468 23992 23520
rect 25228 23511 25280 23520
rect 25228 23477 25237 23511
rect 25237 23477 25271 23511
rect 25271 23477 25280 23511
rect 25228 23468 25280 23477
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 9220 23264 9272 23316
rect 14464 23264 14516 23316
rect 9404 23196 9456 23248
rect 8668 23128 8720 23180
rect 11704 23171 11756 23180
rect 11704 23137 11713 23171
rect 11713 23137 11747 23171
rect 11747 23137 11756 23171
rect 11704 23128 11756 23137
rect 12624 23196 12676 23248
rect 9864 23060 9916 23112
rect 13636 23128 13688 23180
rect 14464 23060 14516 23112
rect 15660 23060 15712 23112
rect 10416 22992 10468 23044
rect 11796 22992 11848 23044
rect 9772 22924 9824 22976
rect 10508 22924 10560 22976
rect 12164 22924 12216 22976
rect 16764 23264 16816 23316
rect 26332 23264 26384 23316
rect 18696 23196 18748 23248
rect 19708 23196 19760 23248
rect 18512 23171 18564 23180
rect 18512 23137 18521 23171
rect 18521 23137 18555 23171
rect 18555 23137 18564 23171
rect 18512 23128 18564 23137
rect 18604 23128 18656 23180
rect 18788 23128 18840 23180
rect 19984 23171 20036 23180
rect 19984 23137 19993 23171
rect 19993 23137 20027 23171
rect 20027 23137 20036 23171
rect 19984 23128 20036 23137
rect 20444 23128 20496 23180
rect 20812 23128 20864 23180
rect 24308 23128 24360 23180
rect 25320 23128 25372 23180
rect 18328 23060 18380 23112
rect 19248 23060 19300 23112
rect 16856 22992 16908 23044
rect 23756 23060 23808 23112
rect 25596 23060 25648 23112
rect 24860 22992 24912 23044
rect 16580 22924 16632 22976
rect 18236 22924 18288 22976
rect 18604 22924 18656 22976
rect 19248 22924 19300 22976
rect 22100 22924 22152 22976
rect 22560 22924 22612 22976
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 9312 22720 9364 22772
rect 10140 22763 10192 22772
rect 10140 22729 10149 22763
rect 10149 22729 10183 22763
rect 10183 22729 10192 22763
rect 10140 22720 10192 22729
rect 8944 22652 8996 22704
rect 14740 22720 14792 22772
rect 16856 22763 16908 22772
rect 16856 22729 16865 22763
rect 16865 22729 16899 22763
rect 16899 22729 16908 22763
rect 16856 22720 16908 22729
rect 18328 22720 18380 22772
rect 18972 22720 19024 22772
rect 19616 22720 19668 22772
rect 25136 22720 25188 22772
rect 18604 22652 18656 22704
rect 20904 22652 20956 22704
rect 7840 22584 7892 22636
rect 12348 22627 12400 22636
rect 12348 22593 12357 22627
rect 12357 22593 12391 22627
rect 12391 22593 12400 22627
rect 12348 22584 12400 22593
rect 10876 22516 10928 22568
rect 13360 22516 13412 22568
rect 20444 22584 20496 22636
rect 21456 22584 21508 22636
rect 22100 22627 22152 22636
rect 22100 22593 22109 22627
rect 22109 22593 22143 22627
rect 22143 22593 22152 22627
rect 22100 22584 22152 22593
rect 22836 22584 22888 22636
rect 18604 22516 18656 22568
rect 19156 22516 19208 22568
rect 19524 22516 19576 22568
rect 19800 22516 19852 22568
rect 20168 22516 20220 22568
rect 23388 22516 23440 22568
rect 24768 22559 24820 22568
rect 24768 22525 24777 22559
rect 24777 22525 24811 22559
rect 24811 22525 24820 22559
rect 24768 22516 24820 22525
rect 6920 22380 6972 22432
rect 9864 22423 9916 22432
rect 9864 22389 9873 22423
rect 9873 22389 9907 22423
rect 9907 22389 9916 22423
rect 9864 22380 9916 22389
rect 12072 22380 12124 22432
rect 22284 22448 22336 22500
rect 22836 22448 22888 22500
rect 14096 22423 14148 22432
rect 14096 22389 14105 22423
rect 14105 22389 14139 22423
rect 14139 22389 14148 22423
rect 14096 22380 14148 22389
rect 20444 22423 20496 22432
rect 20444 22389 20453 22423
rect 20453 22389 20487 22423
rect 20487 22389 20496 22423
rect 20444 22380 20496 22389
rect 20720 22423 20772 22432
rect 20720 22389 20729 22423
rect 20729 22389 20763 22423
rect 20763 22389 20772 22423
rect 20720 22380 20772 22389
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 11060 22176 11112 22228
rect 12072 22108 12124 22160
rect 23296 22176 23348 22228
rect 23756 22219 23808 22228
rect 23756 22185 23765 22219
rect 23765 22185 23799 22219
rect 23799 22185 23808 22219
rect 23756 22176 23808 22185
rect 8944 22083 8996 22092
rect 8944 22049 8953 22083
rect 8953 22049 8987 22083
rect 8987 22049 8996 22083
rect 8944 22040 8996 22049
rect 11336 22083 11388 22092
rect 11336 22049 11345 22083
rect 11345 22049 11379 22083
rect 11379 22049 11388 22083
rect 11336 22040 11388 22049
rect 12440 22083 12492 22092
rect 12440 22049 12449 22083
rect 12449 22049 12483 22083
rect 12483 22049 12492 22083
rect 12440 22040 12492 22049
rect 15752 22108 15804 22160
rect 9496 21972 9548 22024
rect 10324 21879 10376 21888
rect 10324 21845 10333 21879
rect 10333 21845 10367 21879
rect 10367 21845 10376 21879
rect 10324 21836 10376 21845
rect 10692 21879 10744 21888
rect 10692 21845 10701 21879
rect 10701 21845 10735 21879
rect 10735 21845 10744 21879
rect 10692 21836 10744 21845
rect 11060 21879 11112 21888
rect 11060 21845 11069 21879
rect 11069 21845 11103 21879
rect 11103 21845 11112 21879
rect 11060 21836 11112 21845
rect 14096 21972 14148 22024
rect 18788 22040 18840 22092
rect 20352 22083 20404 22092
rect 20352 22049 20361 22083
rect 20361 22049 20395 22083
rect 20395 22049 20404 22083
rect 20352 22040 20404 22049
rect 22192 22040 22244 22092
rect 22836 22040 22888 22092
rect 25044 22083 25096 22092
rect 25044 22049 25053 22083
rect 25053 22049 25087 22083
rect 25087 22049 25096 22083
rect 25044 22040 25096 22049
rect 25504 22108 25556 22160
rect 14832 21879 14884 21888
rect 14832 21845 14841 21879
rect 14841 21845 14875 21879
rect 14875 21845 14884 21879
rect 14832 21836 14884 21845
rect 15200 21879 15252 21888
rect 15200 21845 15209 21879
rect 15209 21845 15243 21879
rect 15243 21845 15252 21879
rect 15200 21836 15252 21845
rect 21364 21972 21416 22024
rect 23940 22015 23992 22024
rect 23940 21981 23949 22015
rect 23949 21981 23983 22015
rect 23983 21981 23992 22015
rect 23940 21972 23992 21981
rect 16396 21947 16448 21956
rect 16396 21913 16405 21947
rect 16405 21913 16439 21947
rect 16439 21913 16448 21947
rect 16396 21904 16448 21913
rect 16580 21836 16632 21888
rect 17776 21904 17828 21956
rect 21548 21904 21600 21956
rect 17040 21836 17092 21888
rect 17132 21836 17184 21888
rect 19892 21836 19944 21888
rect 20076 21879 20128 21888
rect 20076 21845 20085 21879
rect 20085 21845 20119 21879
rect 20119 21845 20128 21879
rect 20076 21836 20128 21845
rect 24032 21836 24084 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 8944 21564 8996 21616
rect 10232 21632 10284 21684
rect 11060 21632 11112 21684
rect 9956 21496 10008 21548
rect 8852 21428 8904 21480
rect 8944 21428 8996 21480
rect 7748 21292 7800 21344
rect 8300 21292 8352 21344
rect 8668 21335 8720 21344
rect 8668 21301 8677 21335
rect 8677 21301 8711 21335
rect 8711 21301 8720 21335
rect 8668 21292 8720 21301
rect 9588 21292 9640 21344
rect 10692 21564 10744 21616
rect 14096 21632 14148 21684
rect 15108 21632 15160 21684
rect 20076 21632 20128 21684
rect 21364 21675 21416 21684
rect 21364 21641 21373 21675
rect 21373 21641 21407 21675
rect 21407 21641 21416 21675
rect 21364 21632 21416 21641
rect 22468 21675 22520 21684
rect 22468 21641 22477 21675
rect 22477 21641 22511 21675
rect 22511 21641 22520 21675
rect 22468 21632 22520 21641
rect 22652 21632 22704 21684
rect 22836 21632 22888 21684
rect 23296 21632 23348 21684
rect 11520 21496 11572 21548
rect 10876 21471 10928 21480
rect 10876 21437 10885 21471
rect 10885 21437 10919 21471
rect 10919 21437 10928 21471
rect 10876 21428 10928 21437
rect 10968 21471 11020 21480
rect 10968 21437 10977 21471
rect 10977 21437 11011 21471
rect 11011 21437 11020 21471
rect 10968 21428 11020 21437
rect 14832 21564 14884 21616
rect 22192 21564 22244 21616
rect 12348 21428 12400 21480
rect 12716 21428 12768 21480
rect 22008 21496 22060 21548
rect 24124 21564 24176 21616
rect 19064 21428 19116 21480
rect 19156 21428 19208 21480
rect 20168 21471 20220 21480
rect 20168 21437 20177 21471
rect 20177 21437 20211 21471
rect 20211 21437 20220 21471
rect 20168 21428 20220 21437
rect 12532 21292 12584 21344
rect 14648 21360 14700 21412
rect 15292 21360 15344 21412
rect 14096 21292 14148 21344
rect 14372 21292 14424 21344
rect 15016 21292 15068 21344
rect 21088 21360 21140 21412
rect 19156 21335 19208 21344
rect 19156 21301 19165 21335
rect 19165 21301 19199 21335
rect 19199 21301 19208 21335
rect 19156 21292 19208 21301
rect 20444 21292 20496 21344
rect 21548 21335 21600 21344
rect 21548 21301 21557 21335
rect 21557 21301 21591 21335
rect 21591 21301 21600 21335
rect 21548 21292 21600 21301
rect 21732 21292 21784 21344
rect 25320 21428 25372 21480
rect 23572 21292 23624 21344
rect 24124 21292 24176 21344
rect 25136 21292 25188 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 3516 21088 3568 21140
rect 15292 21088 15344 21140
rect 15568 21088 15620 21140
rect 13360 21020 13412 21072
rect 16580 21020 16632 21072
rect 20076 21020 20128 21072
rect 9956 20995 10008 21004
rect 9956 20961 9965 20995
rect 9965 20961 9999 20995
rect 9999 20961 10008 20995
rect 9956 20952 10008 20961
rect 19708 20952 19760 21004
rect 20904 21088 20956 21140
rect 10692 20927 10744 20936
rect 10692 20893 10701 20927
rect 10701 20893 10735 20927
rect 10735 20893 10744 20927
rect 10692 20884 10744 20893
rect 18604 20884 18656 20936
rect 22008 20995 22060 21004
rect 22008 20961 22017 20995
rect 22017 20961 22051 20995
rect 22051 20961 22060 20995
rect 22008 20952 22060 20961
rect 24860 20952 24912 21004
rect 24952 20952 25004 21004
rect 23940 20884 23992 20936
rect 10876 20816 10928 20868
rect 8944 20748 8996 20800
rect 15752 20816 15804 20868
rect 14648 20791 14700 20800
rect 14648 20757 14657 20791
rect 14657 20757 14691 20791
rect 14691 20757 14700 20791
rect 14648 20748 14700 20757
rect 16396 20748 16448 20800
rect 20260 20816 20312 20868
rect 17776 20748 17828 20800
rect 18788 20748 18840 20800
rect 18972 20748 19024 20800
rect 24584 20791 24636 20800
rect 24584 20757 24593 20791
rect 24593 20757 24627 20791
rect 24627 20757 24636 20791
rect 24584 20748 24636 20757
rect 24860 20748 24912 20800
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 8852 20544 8904 20596
rect 8300 20476 8352 20528
rect 9036 20476 9088 20528
rect 9312 20476 9364 20528
rect 9588 20476 9640 20528
rect 10416 20587 10468 20596
rect 10416 20553 10425 20587
rect 10425 20553 10459 20587
rect 10459 20553 10468 20587
rect 10416 20544 10468 20553
rect 12624 20544 12676 20596
rect 13636 20544 13688 20596
rect 15476 20587 15528 20596
rect 15476 20553 15485 20587
rect 15485 20553 15519 20587
rect 15519 20553 15528 20587
rect 15476 20544 15528 20553
rect 14648 20476 14700 20528
rect 19432 20544 19484 20596
rect 20904 20587 20956 20596
rect 20904 20553 20913 20587
rect 20913 20553 20947 20587
rect 20947 20553 20956 20587
rect 20904 20544 20956 20553
rect 17132 20519 17184 20528
rect 17132 20485 17141 20519
rect 17141 20485 17175 20519
rect 17175 20485 17184 20519
rect 17132 20476 17184 20485
rect 17776 20476 17828 20528
rect 18788 20476 18840 20528
rect 25320 20587 25372 20596
rect 25320 20553 25329 20587
rect 25329 20553 25363 20587
rect 25363 20553 25372 20587
rect 25320 20544 25372 20553
rect 21088 20476 21140 20528
rect 7748 20383 7800 20392
rect 7748 20349 7757 20383
rect 7757 20349 7791 20383
rect 7791 20349 7800 20383
rect 7748 20340 7800 20349
rect 9772 20383 9824 20392
rect 9772 20349 9781 20383
rect 9781 20349 9815 20383
rect 9815 20349 9824 20383
rect 9772 20340 9824 20349
rect 10232 20340 10284 20392
rect 19524 20408 19576 20460
rect 12716 20383 12768 20392
rect 12716 20349 12725 20383
rect 12725 20349 12759 20383
rect 12759 20349 12768 20383
rect 12716 20340 12768 20349
rect 13452 20340 13504 20392
rect 14372 20340 14424 20392
rect 17224 20340 17276 20392
rect 18512 20340 18564 20392
rect 21824 20408 21876 20460
rect 22192 20451 22244 20460
rect 22192 20417 22201 20451
rect 22201 20417 22235 20451
rect 22235 20417 22244 20451
rect 22192 20408 22244 20417
rect 24124 20476 24176 20528
rect 23388 20340 23440 20392
rect 23572 20383 23624 20392
rect 23572 20349 23581 20383
rect 23581 20349 23615 20383
rect 23615 20349 23624 20383
rect 23572 20340 23624 20349
rect 25136 20340 25188 20392
rect 14464 20247 14516 20256
rect 14464 20213 14473 20247
rect 14473 20213 14507 20247
rect 14507 20213 14516 20247
rect 14464 20204 14516 20213
rect 19156 20272 19208 20324
rect 19064 20247 19116 20256
rect 19064 20213 19073 20247
rect 19073 20213 19107 20247
rect 19107 20213 19116 20247
rect 19064 20204 19116 20213
rect 19524 20204 19576 20256
rect 21272 20204 21324 20256
rect 22744 20247 22796 20256
rect 22744 20213 22753 20247
rect 22753 20213 22787 20247
rect 22787 20213 22796 20247
rect 22744 20204 22796 20213
rect 23664 20204 23716 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 8392 20000 8444 20052
rect 9036 20000 9088 20052
rect 14004 20000 14056 20052
rect 15752 20000 15804 20052
rect 22192 20000 22244 20052
rect 23940 20000 23992 20052
rect 17132 19932 17184 19984
rect 7748 19796 7800 19848
rect 9036 19796 9088 19848
rect 10692 19864 10744 19916
rect 11980 19907 12032 19916
rect 11980 19873 11989 19907
rect 11989 19873 12023 19907
rect 12023 19873 12032 19907
rect 11980 19864 12032 19873
rect 14556 19907 14608 19916
rect 14556 19873 14565 19907
rect 14565 19873 14599 19907
rect 14599 19873 14608 19907
rect 14556 19864 14608 19873
rect 14648 19864 14700 19916
rect 17776 19864 17828 19916
rect 17960 19907 18012 19916
rect 17960 19873 17969 19907
rect 17969 19873 18003 19907
rect 18003 19873 18012 19907
rect 17960 19864 18012 19873
rect 20260 19864 20312 19916
rect 22836 19864 22888 19916
rect 23112 19864 23164 19916
rect 24860 19864 24912 19916
rect 12716 19796 12768 19848
rect 15844 19796 15896 19848
rect 8300 19728 8352 19780
rect 9404 19771 9456 19780
rect 9404 19737 9413 19771
rect 9413 19737 9447 19771
rect 9447 19737 9456 19771
rect 9404 19728 9456 19737
rect 11244 19728 11296 19780
rect 14648 19728 14700 19780
rect 15936 19728 15988 19780
rect 19616 19796 19668 19848
rect 21548 19796 21600 19848
rect 21824 19796 21876 19848
rect 9588 19660 9640 19712
rect 10876 19703 10928 19712
rect 10876 19669 10885 19703
rect 10885 19669 10919 19703
rect 10919 19669 10928 19703
rect 10876 19660 10928 19669
rect 11704 19703 11756 19712
rect 11704 19669 11713 19703
rect 11713 19669 11747 19703
rect 11747 19669 11756 19703
rect 11704 19660 11756 19669
rect 14556 19660 14608 19712
rect 15384 19660 15436 19712
rect 19800 19728 19852 19780
rect 20168 19771 20220 19780
rect 20168 19737 20177 19771
rect 20177 19737 20211 19771
rect 20211 19737 20220 19771
rect 20168 19728 20220 19737
rect 18512 19660 18564 19712
rect 21640 19703 21692 19712
rect 21640 19669 21649 19703
rect 21649 19669 21683 19703
rect 21683 19669 21692 19703
rect 21640 19660 21692 19669
rect 21824 19660 21876 19712
rect 24124 19703 24176 19712
rect 24124 19669 24133 19703
rect 24133 19669 24167 19703
rect 24167 19669 24176 19703
rect 25412 19703 25464 19712
rect 24124 19660 24176 19669
rect 25412 19669 25421 19703
rect 25421 19669 25455 19703
rect 25455 19669 25464 19703
rect 25412 19660 25464 19669
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 8760 19499 8812 19508
rect 8760 19465 8769 19499
rect 8769 19465 8803 19499
rect 8803 19465 8812 19499
rect 8760 19456 8812 19465
rect 9588 19456 9640 19508
rect 8392 19388 8444 19440
rect 8668 19388 8720 19440
rect 9220 19388 9272 19440
rect 6552 19295 6604 19304
rect 6552 19261 6561 19295
rect 6561 19261 6595 19295
rect 6595 19261 6604 19295
rect 6552 19252 6604 19261
rect 6920 19252 6972 19304
rect 10140 19320 10192 19372
rect 11704 19499 11756 19508
rect 11704 19465 11713 19499
rect 11713 19465 11747 19499
rect 11747 19465 11756 19499
rect 11704 19456 11756 19465
rect 11796 19456 11848 19508
rect 14648 19388 14700 19440
rect 15292 19456 15344 19508
rect 17316 19499 17368 19508
rect 17316 19465 17325 19499
rect 17325 19465 17359 19499
rect 17359 19465 17368 19499
rect 17316 19456 17368 19465
rect 19248 19456 19300 19508
rect 20444 19499 20496 19508
rect 20444 19465 20453 19499
rect 20453 19465 20487 19499
rect 20487 19465 20496 19499
rect 20444 19456 20496 19465
rect 20720 19456 20772 19508
rect 22468 19456 22520 19508
rect 22560 19456 22612 19508
rect 25136 19499 25188 19508
rect 25136 19465 25145 19499
rect 25145 19465 25179 19499
rect 25179 19465 25188 19499
rect 25136 19456 25188 19465
rect 25412 19499 25464 19508
rect 25412 19465 25421 19499
rect 25421 19465 25455 19499
rect 25455 19465 25464 19499
rect 25412 19456 25464 19465
rect 8576 19184 8628 19236
rect 11428 19252 11480 19304
rect 8392 19116 8444 19168
rect 11244 19159 11296 19168
rect 11244 19125 11253 19159
rect 11253 19125 11287 19159
rect 11287 19125 11296 19159
rect 11244 19116 11296 19125
rect 14464 19252 14516 19304
rect 15568 19320 15620 19372
rect 16488 19320 16540 19372
rect 16672 19320 16724 19372
rect 21548 19388 21600 19440
rect 15752 19252 15804 19304
rect 19156 19363 19208 19372
rect 19156 19329 19165 19363
rect 19165 19329 19199 19363
rect 19199 19329 19208 19363
rect 19156 19320 19208 19329
rect 23572 19388 23624 19440
rect 23940 19388 23992 19440
rect 24124 19388 24176 19440
rect 19340 19252 19392 19304
rect 21640 19252 21692 19304
rect 23296 19252 23348 19304
rect 12808 19116 12860 19168
rect 14372 19116 14424 19168
rect 14648 19159 14700 19168
rect 14648 19125 14657 19159
rect 14657 19125 14691 19159
rect 14691 19125 14700 19159
rect 14648 19116 14700 19125
rect 20996 19116 21048 19168
rect 21824 19159 21876 19168
rect 21824 19125 21833 19159
rect 21833 19125 21867 19159
rect 21867 19125 21876 19159
rect 21824 19116 21876 19125
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 8668 18955 8720 18964
rect 8668 18921 8677 18955
rect 8677 18921 8711 18955
rect 8711 18921 8720 18955
rect 8668 18912 8720 18921
rect 10048 18955 10100 18964
rect 10048 18921 10057 18955
rect 10057 18921 10091 18955
rect 10091 18921 10100 18955
rect 10048 18912 10100 18921
rect 15844 18912 15896 18964
rect 16856 18912 16908 18964
rect 25964 18912 26016 18964
rect 9956 18844 10008 18896
rect 8392 18776 8444 18828
rect 9680 18776 9732 18828
rect 10600 18819 10652 18828
rect 10600 18785 10609 18819
rect 10609 18785 10643 18819
rect 10643 18785 10652 18819
rect 10600 18776 10652 18785
rect 10876 18776 10928 18828
rect 6644 18751 6696 18760
rect 6644 18717 6653 18751
rect 6653 18717 6687 18751
rect 6687 18717 6696 18751
rect 6644 18708 6696 18717
rect 8668 18708 8720 18760
rect 8852 18708 8904 18760
rect 9404 18708 9456 18760
rect 7012 18572 7064 18624
rect 9588 18640 9640 18692
rect 10600 18640 10652 18692
rect 11704 18640 11756 18692
rect 12164 18708 12216 18760
rect 16948 18776 17000 18828
rect 12532 18708 12584 18760
rect 17776 18776 17828 18828
rect 17316 18708 17368 18760
rect 24492 18844 24544 18896
rect 23848 18819 23900 18828
rect 23848 18785 23857 18819
rect 23857 18785 23891 18819
rect 23891 18785 23900 18819
rect 23848 18776 23900 18785
rect 21548 18708 21600 18760
rect 22744 18751 22796 18760
rect 22744 18717 22753 18751
rect 22753 18717 22787 18751
rect 22787 18717 22796 18751
rect 22744 18708 22796 18717
rect 26608 18708 26660 18760
rect 12440 18640 12492 18692
rect 16948 18640 17000 18692
rect 17684 18640 17736 18692
rect 25412 18640 25464 18692
rect 8300 18572 8352 18624
rect 8944 18572 8996 18624
rect 10508 18615 10560 18624
rect 10508 18581 10517 18615
rect 10517 18581 10551 18615
rect 10551 18581 10560 18615
rect 10508 18572 10560 18581
rect 11336 18572 11388 18624
rect 12624 18572 12676 18624
rect 14280 18615 14332 18624
rect 14280 18581 14289 18615
rect 14289 18581 14323 18615
rect 14323 18581 14332 18615
rect 14280 18572 14332 18581
rect 16764 18572 16816 18624
rect 17592 18572 17644 18624
rect 21364 18572 21416 18624
rect 22100 18572 22152 18624
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 10048 18368 10100 18420
rect 10416 18411 10468 18420
rect 10416 18377 10425 18411
rect 10425 18377 10459 18411
rect 10459 18377 10468 18411
rect 10416 18368 10468 18377
rect 10508 18368 10560 18420
rect 16856 18368 16908 18420
rect 8668 18300 8720 18352
rect 9588 18232 9640 18284
rect 6644 18164 6696 18216
rect 8392 18164 8444 18216
rect 11428 18300 11480 18352
rect 11612 18300 11664 18352
rect 12440 18343 12492 18352
rect 12440 18309 12449 18343
rect 12449 18309 12483 18343
rect 12483 18309 12492 18343
rect 12440 18300 12492 18309
rect 17040 18300 17092 18352
rect 17224 18300 17276 18352
rect 13544 18232 13596 18284
rect 16304 18275 16356 18284
rect 16304 18241 16313 18275
rect 16313 18241 16347 18275
rect 16347 18241 16356 18275
rect 16304 18232 16356 18241
rect 16580 18232 16632 18284
rect 22192 18300 22244 18352
rect 24860 18300 24912 18352
rect 12808 18164 12860 18216
rect 14096 18164 14148 18216
rect 14464 18207 14516 18216
rect 14464 18173 14473 18207
rect 14473 18173 14507 18207
rect 14507 18173 14516 18207
rect 14464 18164 14516 18173
rect 9036 18096 9088 18148
rect 9588 18096 9640 18148
rect 11796 18096 11848 18148
rect 9404 18028 9456 18080
rect 17592 18028 17644 18080
rect 18328 18028 18380 18080
rect 22100 18275 22152 18284
rect 22100 18241 22109 18275
rect 22109 18241 22143 18275
rect 22143 18241 22152 18275
rect 22100 18232 22152 18241
rect 23664 18232 23716 18284
rect 24676 18207 24728 18216
rect 24676 18173 24685 18207
rect 24685 18173 24719 18207
rect 24719 18173 24728 18207
rect 24676 18164 24728 18173
rect 19156 18028 19208 18080
rect 21548 18028 21600 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 8484 17824 8536 17876
rect 15200 17824 15252 17876
rect 21824 17824 21876 17876
rect 21916 17824 21968 17876
rect 26056 17824 26108 17876
rect 9772 17756 9824 17808
rect 7840 17688 7892 17740
rect 24308 17756 24360 17808
rect 24584 17756 24636 17808
rect 11704 17688 11756 17740
rect 13360 17688 13412 17740
rect 13912 17688 13964 17740
rect 14648 17688 14700 17740
rect 16212 17688 16264 17740
rect 17408 17731 17460 17740
rect 17408 17697 17417 17731
rect 17417 17697 17451 17731
rect 17451 17697 17460 17731
rect 17408 17688 17460 17697
rect 17500 17731 17552 17740
rect 17500 17697 17509 17731
rect 17509 17697 17543 17731
rect 17543 17697 17552 17731
rect 17500 17688 17552 17697
rect 18328 17688 18380 17740
rect 19800 17688 19852 17740
rect 9588 17620 9640 17672
rect 14280 17620 14332 17672
rect 17316 17663 17368 17672
rect 17316 17629 17325 17663
rect 17325 17629 17359 17663
rect 17359 17629 17368 17663
rect 17316 17620 17368 17629
rect 8852 17552 8904 17604
rect 11428 17552 11480 17604
rect 14096 17552 14148 17604
rect 15568 17552 15620 17604
rect 18696 17552 18748 17604
rect 19340 17620 19392 17672
rect 24952 17688 25004 17740
rect 25136 17731 25188 17740
rect 25136 17697 25145 17731
rect 25145 17697 25179 17731
rect 25179 17697 25188 17731
rect 25136 17688 25188 17697
rect 22192 17595 22244 17604
rect 22192 17561 22201 17595
rect 22201 17561 22235 17595
rect 22235 17561 22244 17595
rect 22192 17552 22244 17561
rect 24584 17620 24636 17672
rect 25872 17552 25924 17604
rect 7196 17527 7248 17536
rect 7196 17493 7205 17527
rect 7205 17493 7239 17527
rect 7239 17493 7248 17527
rect 7196 17484 7248 17493
rect 7748 17484 7800 17536
rect 9404 17484 9456 17536
rect 12716 17527 12768 17536
rect 12716 17493 12725 17527
rect 12725 17493 12759 17527
rect 12759 17493 12768 17527
rect 12716 17484 12768 17493
rect 13176 17484 13228 17536
rect 15752 17527 15804 17536
rect 15752 17493 15761 17527
rect 15761 17493 15795 17527
rect 15795 17493 15804 17527
rect 15752 17484 15804 17493
rect 16212 17484 16264 17536
rect 17224 17484 17276 17536
rect 20904 17484 20956 17536
rect 23572 17484 23624 17536
rect 24676 17484 24728 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 7196 17280 7248 17332
rect 9404 17323 9456 17332
rect 9404 17289 9413 17323
rect 9413 17289 9447 17323
rect 9447 17289 9456 17323
rect 9404 17280 9456 17289
rect 11612 17323 11664 17332
rect 9496 17212 9548 17264
rect 9588 17212 9640 17264
rect 11612 17289 11621 17323
rect 11621 17289 11655 17323
rect 11655 17289 11664 17323
rect 11612 17280 11664 17289
rect 13176 17323 13228 17332
rect 13176 17289 13185 17323
rect 13185 17289 13219 17323
rect 13219 17289 13228 17323
rect 13176 17280 13228 17289
rect 13360 17280 13412 17332
rect 14464 17280 14516 17332
rect 11428 17212 11480 17264
rect 11888 17255 11940 17264
rect 11888 17221 11897 17255
rect 11897 17221 11931 17255
rect 11931 17221 11940 17255
rect 11888 17212 11940 17221
rect 16396 17280 16448 17332
rect 16580 17280 16632 17332
rect 17408 17323 17460 17332
rect 17408 17289 17417 17323
rect 17417 17289 17451 17323
rect 17451 17289 17460 17323
rect 17408 17280 17460 17289
rect 7656 17144 7708 17196
rect 3332 17076 3384 17128
rect 13728 17144 13780 17196
rect 16212 17212 16264 17264
rect 18972 17280 19024 17332
rect 20168 17280 20220 17332
rect 24400 17280 24452 17332
rect 18604 17212 18656 17264
rect 20996 17212 21048 17264
rect 9496 17119 9548 17128
rect 9496 17085 9505 17119
rect 9505 17085 9539 17119
rect 9539 17085 9548 17119
rect 9496 17076 9548 17085
rect 9312 17008 9364 17060
rect 9772 17076 9824 17128
rect 13360 17076 13412 17128
rect 13452 17119 13504 17128
rect 13452 17085 13461 17119
rect 13461 17085 13495 17119
rect 13495 17085 13504 17119
rect 13452 17076 13504 17085
rect 14832 17119 14884 17128
rect 14832 17085 14841 17119
rect 14841 17085 14875 17119
rect 14875 17085 14884 17119
rect 14832 17076 14884 17085
rect 14924 17076 14976 17128
rect 23480 17187 23532 17196
rect 23480 17153 23489 17187
rect 23489 17153 23523 17187
rect 23523 17153 23532 17187
rect 23480 17144 23532 17153
rect 24860 17144 24912 17196
rect 17868 17076 17920 17128
rect 18972 17076 19024 17128
rect 21916 17076 21968 17128
rect 22836 17076 22888 17128
rect 13636 17008 13688 17060
rect 17132 17051 17184 17060
rect 17132 17017 17141 17051
rect 17141 17017 17175 17051
rect 17175 17017 17184 17051
rect 17132 17008 17184 17017
rect 11152 16940 11204 16992
rect 11888 16940 11940 16992
rect 13912 16940 13964 16992
rect 15384 16940 15436 16992
rect 22560 16940 22612 16992
rect 24216 17076 24268 17128
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 10048 16600 10100 16652
rect 10968 16600 11020 16652
rect 10416 16532 10468 16584
rect 11428 16600 11480 16652
rect 12808 16736 12860 16788
rect 13912 16779 13964 16788
rect 13912 16745 13921 16779
rect 13921 16745 13955 16779
rect 13955 16745 13964 16779
rect 13912 16736 13964 16745
rect 14280 16779 14332 16788
rect 14280 16745 14289 16779
rect 14289 16745 14323 16779
rect 14323 16745 14332 16779
rect 14280 16736 14332 16745
rect 18972 16736 19024 16788
rect 20996 16736 21048 16788
rect 22284 16736 22336 16788
rect 24584 16779 24636 16788
rect 24584 16745 24593 16779
rect 24593 16745 24627 16779
rect 24627 16745 24636 16779
rect 24584 16736 24636 16745
rect 14372 16668 14424 16720
rect 13636 16600 13688 16652
rect 15844 16600 15896 16652
rect 16304 16643 16356 16652
rect 16304 16609 16313 16643
rect 16313 16609 16347 16643
rect 16347 16609 16356 16643
rect 16304 16600 16356 16609
rect 16396 16600 16448 16652
rect 17868 16600 17920 16652
rect 19340 16643 19392 16652
rect 10324 16464 10376 16516
rect 13912 16464 13964 16516
rect 9864 16439 9916 16448
rect 9864 16405 9873 16439
rect 9873 16405 9907 16439
rect 9907 16405 9916 16439
rect 9864 16396 9916 16405
rect 10232 16439 10284 16448
rect 10232 16405 10241 16439
rect 10241 16405 10275 16439
rect 10275 16405 10284 16439
rect 10232 16396 10284 16405
rect 12256 16396 12308 16448
rect 13636 16396 13688 16448
rect 15476 16464 15528 16516
rect 15752 16532 15804 16584
rect 16948 16575 17000 16584
rect 16948 16541 16957 16575
rect 16957 16541 16991 16575
rect 16991 16541 17000 16575
rect 16948 16532 17000 16541
rect 19340 16609 19349 16643
rect 19349 16609 19383 16643
rect 19383 16609 19392 16643
rect 19340 16600 19392 16609
rect 20260 16643 20312 16652
rect 20260 16609 20269 16643
rect 20269 16609 20303 16643
rect 20303 16609 20312 16643
rect 20260 16600 20312 16609
rect 19800 16575 19852 16584
rect 19800 16541 19809 16575
rect 19809 16541 19843 16575
rect 19843 16541 19852 16575
rect 19800 16532 19852 16541
rect 22376 16532 22428 16584
rect 23848 16575 23900 16584
rect 23848 16541 23857 16575
rect 23857 16541 23891 16575
rect 23891 16541 23900 16575
rect 23848 16532 23900 16541
rect 15016 16439 15068 16448
rect 15016 16405 15025 16439
rect 15025 16405 15059 16439
rect 15059 16405 15068 16439
rect 15016 16396 15068 16405
rect 15936 16396 15988 16448
rect 19616 16439 19668 16448
rect 19616 16405 19625 16439
rect 19625 16405 19659 16439
rect 19659 16405 19668 16439
rect 19616 16396 19668 16405
rect 20536 16507 20588 16516
rect 20536 16473 20545 16507
rect 20545 16473 20579 16507
rect 20579 16473 20588 16507
rect 20536 16464 20588 16473
rect 20996 16464 21048 16516
rect 21916 16396 21968 16448
rect 22284 16396 22336 16448
rect 23664 16396 23716 16448
rect 24860 16396 24912 16448
rect 25136 16396 25188 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 8576 16192 8628 16244
rect 8668 16235 8720 16244
rect 8668 16201 8677 16235
rect 8677 16201 8711 16235
rect 8711 16201 8720 16235
rect 8668 16192 8720 16201
rect 11060 16192 11112 16244
rect 14188 16192 14240 16244
rect 15016 16192 15068 16244
rect 15476 16192 15528 16244
rect 16856 16235 16908 16244
rect 16856 16201 16865 16235
rect 16865 16201 16899 16235
rect 16899 16201 16908 16235
rect 16856 16192 16908 16201
rect 14280 16124 14332 16176
rect 20260 16192 20312 16244
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 11704 16056 11756 16108
rect 12164 16056 12216 16108
rect 8484 15988 8536 16040
rect 9588 15988 9640 16040
rect 14740 16056 14792 16108
rect 13820 16031 13872 16040
rect 13820 15997 13829 16031
rect 13829 15997 13863 16031
rect 13863 15997 13872 16031
rect 13820 15988 13872 15997
rect 11704 15920 11756 15972
rect 14280 15988 14332 16040
rect 14372 15920 14424 15972
rect 18420 16056 18472 16108
rect 19340 16056 19392 16108
rect 20352 16124 20404 16176
rect 20628 16124 20680 16176
rect 21916 16124 21968 16176
rect 20444 16056 20496 16108
rect 20812 16056 20864 16108
rect 22284 16192 22336 16244
rect 23296 16192 23348 16244
rect 23664 16124 23716 16176
rect 24860 16192 24912 16244
rect 23296 16056 23348 16108
rect 23848 16056 23900 16108
rect 19892 15988 19944 16040
rect 17684 15920 17736 15972
rect 18236 15920 18288 15972
rect 19800 15920 19852 15972
rect 22008 15920 22060 15972
rect 12256 15852 12308 15904
rect 17316 15895 17368 15904
rect 17316 15861 17325 15895
rect 17325 15861 17359 15895
rect 17359 15861 17368 15895
rect 17316 15852 17368 15861
rect 17776 15852 17828 15904
rect 18512 15895 18564 15904
rect 18512 15861 18521 15895
rect 18521 15861 18555 15895
rect 18555 15861 18564 15895
rect 18512 15852 18564 15861
rect 21456 15852 21508 15904
rect 22744 15988 22796 16040
rect 22836 15988 22888 16040
rect 24584 15988 24636 16040
rect 23756 15895 23808 15904
rect 23756 15861 23765 15895
rect 23765 15861 23799 15895
rect 23799 15861 23808 15895
rect 23756 15852 23808 15861
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 9220 15648 9272 15700
rect 10416 15648 10468 15700
rect 11520 15648 11572 15700
rect 17684 15648 17736 15700
rect 17868 15648 17920 15700
rect 9588 15512 9640 15564
rect 12164 15555 12216 15564
rect 12164 15521 12173 15555
rect 12173 15521 12207 15555
rect 12207 15521 12216 15555
rect 12164 15512 12216 15521
rect 16396 15555 16448 15564
rect 16396 15521 16405 15555
rect 16405 15521 16439 15555
rect 16439 15521 16448 15555
rect 16396 15512 16448 15521
rect 18328 15512 18380 15564
rect 19156 15648 19208 15700
rect 21456 15648 21508 15700
rect 22744 15648 22796 15700
rect 22928 15648 22980 15700
rect 25136 15691 25188 15700
rect 25136 15657 25145 15691
rect 25145 15657 25179 15691
rect 25179 15657 25188 15691
rect 25136 15648 25188 15657
rect 20260 15512 20312 15564
rect 9220 15376 9272 15428
rect 12532 15376 12584 15428
rect 10048 15308 10100 15360
rect 12072 15351 12124 15360
rect 12072 15317 12081 15351
rect 12081 15317 12115 15351
rect 12115 15317 12124 15351
rect 12072 15308 12124 15317
rect 14280 15351 14332 15360
rect 14280 15317 14289 15351
rect 14289 15317 14323 15351
rect 14323 15317 14332 15351
rect 14280 15308 14332 15317
rect 15752 15351 15804 15360
rect 15752 15317 15761 15351
rect 15761 15317 15795 15351
rect 15795 15317 15804 15351
rect 15752 15308 15804 15317
rect 16396 15308 16448 15360
rect 19708 15419 19760 15428
rect 19708 15385 19717 15419
rect 19717 15385 19751 15419
rect 19751 15385 19760 15419
rect 19708 15376 19760 15385
rect 22284 15555 22336 15564
rect 22284 15521 22293 15555
rect 22293 15521 22327 15555
rect 22327 15521 22336 15555
rect 22284 15512 22336 15521
rect 23756 15512 23808 15564
rect 24676 15512 24728 15564
rect 21824 15487 21876 15496
rect 21824 15453 21833 15487
rect 21833 15453 21867 15487
rect 21867 15453 21876 15487
rect 21824 15444 21876 15453
rect 23664 15444 23716 15496
rect 21088 15376 21140 15428
rect 20536 15308 20588 15360
rect 25228 15376 25280 15428
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 10140 15147 10192 15156
rect 10140 15113 10149 15147
rect 10149 15113 10183 15147
rect 10183 15113 10192 15147
rect 10140 15104 10192 15113
rect 10416 15104 10468 15156
rect 10876 15104 10928 15156
rect 14280 15104 14332 15156
rect 15568 15147 15620 15156
rect 15568 15113 15577 15147
rect 15577 15113 15611 15147
rect 15611 15113 15620 15147
rect 15568 15104 15620 15113
rect 15752 15104 15804 15156
rect 20076 15147 20128 15156
rect 20076 15113 20085 15147
rect 20085 15113 20119 15147
rect 20119 15113 20128 15147
rect 20076 15104 20128 15113
rect 20168 15104 20220 15156
rect 25688 15104 25740 15156
rect 8668 15036 8720 15088
rect 11520 15036 11572 15088
rect 19248 15036 19300 15088
rect 21088 15036 21140 15088
rect 23296 15079 23348 15088
rect 23296 15045 23305 15079
rect 23305 15045 23339 15079
rect 23339 15045 23348 15079
rect 23296 15036 23348 15045
rect 9588 14968 9640 15020
rect 8576 14900 8628 14952
rect 9312 14900 9364 14952
rect 11428 14968 11480 15020
rect 19432 14968 19484 15020
rect 11888 14900 11940 14952
rect 15384 14900 15436 14952
rect 15476 14900 15528 14952
rect 17040 14900 17092 14952
rect 20536 14900 20588 14952
rect 22100 15011 22152 15020
rect 22100 14977 22109 15011
rect 22109 14977 22143 15011
rect 22143 14977 22152 15011
rect 22100 14968 22152 14977
rect 24124 15011 24176 15020
rect 24124 14977 24133 15011
rect 24133 14977 24167 15011
rect 24167 14977 24176 15011
rect 24124 14968 24176 14977
rect 24032 14900 24084 14952
rect 24768 14943 24820 14952
rect 24768 14909 24777 14943
rect 24777 14909 24811 14943
rect 24811 14909 24820 14943
rect 24768 14900 24820 14909
rect 16672 14832 16724 14884
rect 18880 14875 18932 14884
rect 18880 14841 18889 14875
rect 18889 14841 18923 14875
rect 18923 14841 18932 14875
rect 18880 14832 18932 14841
rect 8300 14764 8352 14816
rect 20720 14764 20772 14816
rect 24032 14764 24084 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 7840 14560 7892 14612
rect 8668 14560 8720 14612
rect 9312 14560 9364 14612
rect 6460 14467 6512 14476
rect 6460 14433 6469 14467
rect 6469 14433 6503 14467
rect 6503 14433 6512 14467
rect 6460 14424 6512 14433
rect 8300 14424 8352 14476
rect 12624 14560 12676 14612
rect 25044 14560 25096 14612
rect 9772 14424 9824 14476
rect 11704 14424 11756 14476
rect 9588 14356 9640 14408
rect 9404 14288 9456 14340
rect 10876 14288 10928 14340
rect 13452 14424 13504 14476
rect 15752 14492 15804 14544
rect 20352 14492 20404 14544
rect 24308 14492 24360 14544
rect 14924 14424 14976 14476
rect 21272 14424 21324 14476
rect 23204 14424 23256 14476
rect 23388 14424 23440 14476
rect 24860 14424 24912 14476
rect 20168 14356 20220 14408
rect 21732 14356 21784 14408
rect 24492 14356 24544 14408
rect 10968 14220 11020 14272
rect 20904 14288 20956 14340
rect 24400 14288 24452 14340
rect 12808 14263 12860 14272
rect 12808 14229 12817 14263
rect 12817 14229 12851 14263
rect 12851 14229 12860 14263
rect 12808 14220 12860 14229
rect 13360 14220 13412 14272
rect 13544 14263 13596 14272
rect 13544 14229 13553 14263
rect 13553 14229 13587 14263
rect 13587 14229 13596 14263
rect 13544 14220 13596 14229
rect 14464 14220 14516 14272
rect 14740 14263 14792 14272
rect 14740 14229 14749 14263
rect 14749 14229 14783 14263
rect 14783 14229 14792 14263
rect 14740 14220 14792 14229
rect 16580 14220 16632 14272
rect 20260 14263 20312 14272
rect 20260 14229 20269 14263
rect 20269 14229 20303 14263
rect 20303 14229 20312 14263
rect 20260 14220 20312 14229
rect 21824 14263 21876 14272
rect 21824 14229 21833 14263
rect 21833 14229 21867 14263
rect 21867 14229 21876 14263
rect 21824 14220 21876 14229
rect 22008 14220 22060 14272
rect 22468 14220 22520 14272
rect 24860 14263 24912 14272
rect 24860 14229 24869 14263
rect 24869 14229 24903 14263
rect 24903 14229 24912 14263
rect 24860 14220 24912 14229
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 8300 14016 8352 14068
rect 9588 14016 9640 14068
rect 7932 13948 7984 14000
rect 8668 13948 8720 14000
rect 9772 13991 9824 14000
rect 9772 13957 9781 13991
rect 9781 13957 9815 13991
rect 9815 13957 9824 13991
rect 9772 13948 9824 13957
rect 11612 14016 11664 14068
rect 12348 14016 12400 14068
rect 13544 14016 13596 14068
rect 14832 14016 14884 14068
rect 13268 13948 13320 14000
rect 16396 14016 16448 14068
rect 18604 14059 18656 14068
rect 18604 14025 18613 14059
rect 18613 14025 18647 14059
rect 18647 14025 18656 14059
rect 18604 14016 18656 14025
rect 18788 14016 18840 14068
rect 18972 14016 19024 14068
rect 19156 14016 19208 14068
rect 21088 14016 21140 14068
rect 23480 14016 23532 14068
rect 19248 13948 19300 14000
rect 9588 13880 9640 13932
rect 13544 13880 13596 13932
rect 20352 13923 20404 13932
rect 20352 13889 20361 13923
rect 20361 13889 20395 13923
rect 20395 13889 20404 13923
rect 20352 13880 20404 13889
rect 21916 13880 21968 13932
rect 22652 13948 22704 14000
rect 23664 13948 23716 14000
rect 22284 13880 22336 13932
rect 24400 13880 24452 13932
rect 11060 13812 11112 13864
rect 12716 13812 12768 13864
rect 11152 13676 11204 13728
rect 12256 13676 12308 13728
rect 12624 13719 12676 13728
rect 12624 13685 12633 13719
rect 12633 13685 12667 13719
rect 12667 13685 12676 13719
rect 12624 13676 12676 13685
rect 13820 13855 13872 13864
rect 13820 13821 13829 13855
rect 13829 13821 13863 13855
rect 13863 13821 13872 13855
rect 13820 13812 13872 13821
rect 16856 13855 16908 13864
rect 16856 13821 16865 13855
rect 16865 13821 16899 13855
rect 16899 13821 16908 13855
rect 16856 13812 16908 13821
rect 19892 13812 19944 13864
rect 15108 13744 15160 13796
rect 15660 13744 15712 13796
rect 21916 13744 21968 13796
rect 22376 13812 22428 13864
rect 22652 13812 22704 13864
rect 23204 13812 23256 13864
rect 13912 13676 13964 13728
rect 14096 13719 14148 13728
rect 14096 13685 14126 13719
rect 14126 13685 14148 13719
rect 14096 13676 14148 13685
rect 17132 13719 17184 13728
rect 17132 13685 17162 13719
rect 17162 13685 17184 13719
rect 17132 13676 17184 13685
rect 17500 13676 17552 13728
rect 22468 13676 22520 13728
rect 22836 13676 22888 13728
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 8484 13472 8536 13524
rect 8668 13515 8720 13524
rect 8668 13481 8677 13515
rect 8677 13481 8711 13515
rect 8711 13481 8720 13515
rect 8668 13472 8720 13481
rect 8852 13472 8904 13524
rect 13636 13472 13688 13524
rect 14280 13472 14332 13524
rect 17316 13472 17368 13524
rect 17408 13515 17460 13524
rect 17408 13481 17417 13515
rect 17417 13481 17451 13515
rect 17451 13481 17460 13515
rect 17408 13472 17460 13481
rect 18328 13472 18380 13524
rect 21180 13472 21232 13524
rect 24492 13472 24544 13524
rect 9404 13404 9456 13456
rect 9588 13404 9640 13456
rect 6460 13336 6512 13388
rect 9680 13336 9732 13388
rect 13176 13404 13228 13456
rect 15108 13404 15160 13456
rect 16488 13404 16540 13456
rect 19800 13404 19852 13456
rect 20904 13404 20956 13456
rect 22100 13404 22152 13456
rect 22836 13404 22888 13456
rect 23664 13404 23716 13456
rect 11704 13336 11756 13388
rect 13820 13336 13872 13388
rect 15752 13379 15804 13388
rect 15752 13345 15761 13379
rect 15761 13345 15795 13379
rect 15795 13345 15804 13379
rect 15752 13336 15804 13345
rect 16212 13336 16264 13388
rect 17316 13336 17368 13388
rect 17868 13336 17920 13388
rect 18604 13336 18656 13388
rect 13912 13268 13964 13320
rect 15108 13268 15160 13320
rect 8668 13200 8720 13252
rect 9680 13175 9732 13184
rect 9680 13141 9689 13175
rect 9689 13141 9723 13175
rect 9723 13141 9732 13175
rect 9680 13132 9732 13141
rect 11152 13200 11204 13252
rect 12348 13200 12400 13252
rect 11980 13132 12032 13184
rect 12164 13175 12216 13184
rect 12164 13141 12173 13175
rect 12173 13141 12207 13175
rect 12207 13141 12216 13175
rect 12164 13132 12216 13141
rect 12900 13200 12952 13252
rect 15844 13268 15896 13320
rect 16120 13268 16172 13320
rect 20996 13336 21048 13388
rect 21088 13336 21140 13388
rect 19340 13268 19392 13320
rect 17408 13200 17460 13252
rect 13912 13175 13964 13184
rect 13912 13141 13921 13175
rect 13921 13141 13955 13175
rect 13955 13141 13964 13175
rect 13912 13132 13964 13141
rect 15200 13175 15252 13184
rect 15200 13141 15209 13175
rect 15209 13141 15243 13175
rect 15243 13141 15252 13175
rect 15200 13132 15252 13141
rect 16304 13175 16356 13184
rect 16304 13141 16313 13175
rect 16313 13141 16347 13175
rect 16347 13141 16356 13175
rect 16304 13132 16356 13141
rect 18972 13200 19024 13252
rect 20444 13200 20496 13252
rect 23480 13268 23532 13320
rect 23848 13379 23900 13388
rect 23848 13345 23857 13379
rect 23857 13345 23891 13379
rect 23891 13345 23900 13379
rect 23848 13336 23900 13345
rect 25136 13200 25188 13252
rect 19156 13132 19208 13184
rect 20168 13132 20220 13184
rect 22560 13132 22612 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 7012 12928 7064 12980
rect 9220 12928 9272 12980
rect 9404 12971 9456 12980
rect 9404 12937 9413 12971
rect 9413 12937 9447 12971
rect 9447 12937 9456 12971
rect 9404 12928 9456 12937
rect 10048 12928 10100 12980
rect 11060 12928 11112 12980
rect 12256 12971 12308 12980
rect 12256 12937 12265 12971
rect 12265 12937 12299 12971
rect 12299 12937 12308 12971
rect 12256 12928 12308 12937
rect 13084 12928 13136 12980
rect 15476 12971 15528 12980
rect 15476 12937 15485 12971
rect 15485 12937 15519 12971
rect 15519 12937 15528 12971
rect 15476 12928 15528 12937
rect 16120 12971 16172 12980
rect 6920 12860 6972 12912
rect 7012 12835 7064 12844
rect 7012 12801 7021 12835
rect 7021 12801 7055 12835
rect 7055 12801 7064 12835
rect 7012 12792 7064 12801
rect 6920 12724 6972 12776
rect 8208 12835 8260 12844
rect 8208 12801 8217 12835
rect 8217 12801 8251 12835
rect 8251 12801 8260 12835
rect 8208 12792 8260 12801
rect 12624 12860 12676 12912
rect 14004 12860 14056 12912
rect 14280 12903 14332 12912
rect 14280 12869 14289 12903
rect 14289 12869 14323 12903
rect 14323 12869 14332 12903
rect 14280 12860 14332 12869
rect 16120 12937 16129 12971
rect 16129 12937 16163 12971
rect 16163 12937 16172 12971
rect 16120 12928 16172 12937
rect 17224 12928 17276 12980
rect 15936 12860 15988 12912
rect 19800 12928 19852 12980
rect 21180 12971 21232 12980
rect 21180 12937 21189 12971
rect 21189 12937 21223 12971
rect 21223 12937 21232 12971
rect 21180 12928 21232 12937
rect 18052 12860 18104 12912
rect 22284 12860 22336 12912
rect 22376 12860 22428 12912
rect 23664 12928 23716 12980
rect 23388 12903 23440 12912
rect 23388 12869 23397 12903
rect 23397 12869 23431 12903
rect 23431 12869 23440 12903
rect 23388 12860 23440 12869
rect 7656 12724 7708 12776
rect 8392 12767 8444 12776
rect 8392 12733 8401 12767
rect 8401 12733 8435 12767
rect 8435 12733 8444 12767
rect 8392 12724 8444 12733
rect 9772 12724 9824 12776
rect 9956 12724 10008 12776
rect 10968 12767 11020 12776
rect 10968 12733 10977 12767
rect 10977 12733 11011 12767
rect 11011 12733 11020 12767
rect 10968 12724 11020 12733
rect 11796 12792 11848 12844
rect 12900 12792 12952 12844
rect 13544 12792 13596 12844
rect 13728 12792 13780 12844
rect 14924 12792 14976 12844
rect 16488 12792 16540 12844
rect 17224 12835 17276 12844
rect 17224 12801 17233 12835
rect 17233 12801 17267 12835
rect 17267 12801 17276 12835
rect 17224 12792 17276 12801
rect 13176 12724 13228 12776
rect 13452 12724 13504 12776
rect 14280 12724 14332 12776
rect 14832 12724 14884 12776
rect 15108 12724 15160 12776
rect 15660 12724 15712 12776
rect 19156 12835 19208 12844
rect 19156 12801 19165 12835
rect 19165 12801 19199 12835
rect 19199 12801 19208 12835
rect 19156 12792 19208 12801
rect 20168 12835 20220 12844
rect 20168 12801 20177 12835
rect 20177 12801 20211 12835
rect 20211 12801 20220 12835
rect 20168 12792 20220 12801
rect 20352 12792 20404 12844
rect 18788 12724 18840 12776
rect 20628 12724 20680 12776
rect 11336 12656 11388 12708
rect 12348 12656 12400 12708
rect 11244 12588 11296 12640
rect 11796 12588 11848 12640
rect 12440 12588 12492 12640
rect 16580 12588 16632 12640
rect 17408 12588 17460 12640
rect 18052 12631 18104 12640
rect 18052 12597 18061 12631
rect 18061 12597 18095 12631
rect 18095 12597 18104 12631
rect 18052 12588 18104 12597
rect 20812 12656 20864 12708
rect 22652 12724 22704 12776
rect 21916 12588 21968 12640
rect 22836 12588 22888 12640
rect 23388 12588 23440 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 7748 12384 7800 12436
rect 11428 12427 11480 12436
rect 11428 12393 11437 12427
rect 11437 12393 11471 12427
rect 11471 12393 11480 12427
rect 11428 12384 11480 12393
rect 12532 12384 12584 12436
rect 13912 12384 13964 12436
rect 17316 12384 17368 12436
rect 12072 12316 12124 12368
rect 13084 12316 13136 12368
rect 14188 12316 14240 12368
rect 14648 12316 14700 12368
rect 18880 12384 18932 12436
rect 19248 12384 19300 12436
rect 20076 12427 20128 12436
rect 20076 12393 20085 12427
rect 20085 12393 20119 12427
rect 20119 12393 20128 12427
rect 20076 12384 20128 12393
rect 17592 12316 17644 12368
rect 19524 12316 19576 12368
rect 19708 12316 19760 12368
rect 24124 12384 24176 12436
rect 7012 12248 7064 12300
rect 8208 12291 8260 12300
rect 8208 12257 8217 12291
rect 8217 12257 8251 12291
rect 8251 12257 8260 12291
rect 8208 12248 8260 12257
rect 9588 12248 9640 12300
rect 10968 12248 11020 12300
rect 12164 12248 12216 12300
rect 13636 12248 13688 12300
rect 13912 12248 13964 12300
rect 14556 12248 14608 12300
rect 15108 12248 15160 12300
rect 16396 12248 16448 12300
rect 18420 12248 18472 12300
rect 19156 12248 19208 12300
rect 20444 12291 20496 12300
rect 20444 12257 20453 12291
rect 20453 12257 20487 12291
rect 20487 12257 20496 12291
rect 20444 12248 20496 12257
rect 21272 12248 21324 12300
rect 12440 12180 12492 12232
rect 12532 12180 12584 12232
rect 13728 12180 13780 12232
rect 17316 12223 17368 12232
rect 17316 12189 17325 12223
rect 17325 12189 17359 12223
rect 17359 12189 17368 12223
rect 17316 12180 17368 12189
rect 20076 12180 20128 12232
rect 21824 12180 21876 12232
rect 22376 12180 22428 12232
rect 22836 12223 22888 12232
rect 22836 12189 22845 12223
rect 22845 12189 22879 12223
rect 22879 12189 22888 12223
rect 22836 12180 22888 12189
rect 12624 12112 12676 12164
rect 10600 12087 10652 12096
rect 10600 12053 10609 12087
rect 10609 12053 10643 12087
rect 10643 12053 10652 12087
rect 10600 12044 10652 12053
rect 13452 12112 13504 12164
rect 16396 12112 16448 12164
rect 16948 12112 17000 12164
rect 15016 12044 15068 12096
rect 15292 12044 15344 12096
rect 15844 12044 15896 12096
rect 18420 12044 18472 12096
rect 18972 12044 19024 12096
rect 20996 12044 21048 12096
rect 24952 12112 25004 12164
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 5264 11840 5316 11892
rect 9588 11840 9640 11892
rect 9680 11840 9732 11892
rect 11152 11840 11204 11892
rect 12808 11840 12860 11892
rect 13084 11883 13136 11892
rect 13084 11849 13093 11883
rect 13093 11849 13127 11883
rect 13127 11849 13136 11883
rect 13084 11840 13136 11849
rect 13452 11840 13504 11892
rect 14188 11840 14240 11892
rect 14372 11840 14424 11892
rect 16764 11840 16816 11892
rect 8668 11704 8720 11756
rect 11796 11772 11848 11824
rect 12348 11772 12400 11824
rect 14464 11772 14516 11824
rect 12072 11704 12124 11756
rect 17500 11772 17552 11824
rect 18420 11883 18472 11892
rect 18420 11849 18429 11883
rect 18429 11849 18463 11883
rect 18463 11849 18472 11883
rect 18420 11840 18472 11849
rect 19432 11772 19484 11824
rect 19984 11772 20036 11824
rect 25780 11840 25832 11892
rect 24860 11772 24912 11824
rect 14648 11747 14700 11756
rect 14648 11713 14657 11747
rect 14657 11713 14691 11747
rect 14691 11713 14700 11747
rect 14648 11704 14700 11713
rect 16120 11704 16172 11756
rect 19340 11747 19392 11756
rect 19340 11713 19349 11747
rect 19349 11713 19383 11747
rect 19383 11713 19392 11747
rect 19340 11704 19392 11713
rect 11060 11636 11112 11688
rect 10508 11568 10560 11620
rect 11888 11568 11940 11620
rect 8300 11500 8352 11552
rect 11612 11500 11664 11552
rect 12348 11500 12400 11552
rect 13452 11568 13504 11620
rect 13636 11636 13688 11688
rect 14372 11636 14424 11688
rect 15108 11636 15160 11688
rect 16672 11636 16724 11688
rect 18236 11636 18288 11688
rect 19708 11636 19760 11688
rect 19984 11636 20036 11688
rect 15476 11568 15528 11620
rect 16488 11568 16540 11620
rect 16764 11568 16816 11620
rect 21732 11568 21784 11620
rect 23940 11704 23992 11756
rect 24952 11704 25004 11756
rect 24768 11679 24820 11688
rect 24768 11645 24777 11679
rect 24777 11645 24811 11679
rect 24811 11645 24820 11679
rect 24768 11636 24820 11645
rect 26148 11568 26200 11620
rect 14832 11500 14884 11552
rect 15016 11500 15068 11552
rect 15384 11500 15436 11552
rect 17684 11500 17736 11552
rect 19708 11500 19760 11552
rect 20720 11500 20772 11552
rect 23756 11500 23808 11552
rect 24124 11500 24176 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 7196 11296 7248 11348
rect 10508 11296 10560 11348
rect 10600 11296 10652 11348
rect 13268 11296 13320 11348
rect 13452 11296 13504 11348
rect 12808 11228 12860 11280
rect 13176 11228 13228 11280
rect 13820 11228 13872 11280
rect 9128 11135 9180 11144
rect 9128 11101 9137 11135
rect 9137 11101 9171 11135
rect 9171 11101 9180 11135
rect 9128 11092 9180 11101
rect 11888 11203 11940 11212
rect 11888 11169 11897 11203
rect 11897 11169 11931 11203
rect 11931 11169 11940 11203
rect 11888 11160 11940 11169
rect 12256 11160 12308 11212
rect 12072 11092 12124 11144
rect 12716 11092 12768 11144
rect 8668 11024 8720 11076
rect 9864 11024 9916 11076
rect 11060 11024 11112 11076
rect 13544 11160 13596 11212
rect 15200 11296 15252 11348
rect 16304 11296 16356 11348
rect 19432 11296 19484 11348
rect 21640 11296 21692 11348
rect 22836 11296 22888 11348
rect 14464 11228 14516 11280
rect 14832 11228 14884 11280
rect 16672 11271 16724 11280
rect 16672 11237 16681 11271
rect 16681 11237 16715 11271
rect 16715 11237 16724 11271
rect 16672 11228 16724 11237
rect 16764 11228 16816 11280
rect 21364 11228 21416 11280
rect 23756 11228 23808 11280
rect 14372 11160 14424 11212
rect 14740 11160 14792 11212
rect 16948 11160 17000 11212
rect 17316 11160 17368 11212
rect 17500 11160 17552 11212
rect 17960 11160 18012 11212
rect 14188 11092 14240 11144
rect 14556 11092 14608 11144
rect 19984 11135 20036 11144
rect 19984 11101 19993 11135
rect 19993 11101 20027 11135
rect 20027 11101 20036 11135
rect 19984 11092 20036 11101
rect 22468 11160 22520 11212
rect 20812 11092 20864 11144
rect 21088 11092 21140 11144
rect 21732 11135 21784 11144
rect 21732 11101 21741 11135
rect 21741 11101 21775 11135
rect 21775 11101 21784 11135
rect 21732 11092 21784 11101
rect 23480 11092 23532 11144
rect 15108 11024 15160 11076
rect 15200 11067 15252 11076
rect 15200 11033 15209 11067
rect 15209 11033 15243 11067
rect 15243 11033 15252 11067
rect 15200 11024 15252 11033
rect 9680 10956 9732 11008
rect 10876 10999 10928 11008
rect 10876 10965 10885 10999
rect 10885 10965 10919 10999
rect 10919 10965 10928 10999
rect 10876 10956 10928 10965
rect 11888 10956 11940 11008
rect 12072 10956 12124 11008
rect 12440 10956 12492 11008
rect 13452 10956 13504 11008
rect 14280 10999 14332 11008
rect 14280 10965 14289 10999
rect 14289 10965 14323 10999
rect 14323 10965 14332 10999
rect 14280 10956 14332 10965
rect 14832 10956 14884 11008
rect 15476 11024 15528 11076
rect 15384 10956 15436 11008
rect 17684 11024 17736 11076
rect 18236 10956 18288 11008
rect 18512 11067 18564 11076
rect 18512 11033 18521 11067
rect 18521 11033 18555 11067
rect 18555 11033 18564 11067
rect 18512 11024 18564 11033
rect 19616 11024 19668 11076
rect 26700 11160 26752 11212
rect 25228 11135 25280 11144
rect 25228 11101 25237 11135
rect 25237 11101 25271 11135
rect 25271 11101 25280 11135
rect 25228 11092 25280 11101
rect 23848 11067 23900 11076
rect 23848 11033 23857 11067
rect 23857 11033 23891 11067
rect 23891 11033 23900 11067
rect 23848 11024 23900 11033
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 8668 10752 8720 10804
rect 9956 10795 10008 10804
rect 9956 10761 9965 10795
rect 9965 10761 9999 10795
rect 9999 10761 10008 10795
rect 9956 10752 10008 10761
rect 14280 10752 14332 10804
rect 14372 10752 14424 10804
rect 7104 10684 7156 10736
rect 9864 10684 9916 10736
rect 12348 10684 12400 10736
rect 10876 10616 10928 10668
rect 12808 10727 12860 10736
rect 12808 10693 12817 10727
rect 12817 10693 12851 10727
rect 12851 10693 12860 10727
rect 12808 10684 12860 10693
rect 15292 10684 15344 10736
rect 12072 10548 12124 10600
rect 13360 10616 13412 10668
rect 14188 10659 14240 10668
rect 14188 10625 14197 10659
rect 14197 10625 14231 10659
rect 14231 10625 14240 10659
rect 14188 10616 14240 10625
rect 14280 10659 14332 10668
rect 14280 10625 14289 10659
rect 14289 10625 14323 10659
rect 14323 10625 14332 10659
rect 14280 10616 14332 10625
rect 15292 10548 15344 10600
rect 14004 10480 14056 10532
rect 16028 10591 16080 10600
rect 16028 10557 16037 10591
rect 16037 10557 16071 10591
rect 16071 10557 16080 10591
rect 16028 10548 16080 10557
rect 17592 10727 17644 10736
rect 17592 10693 17601 10727
rect 17601 10693 17635 10727
rect 17635 10693 17644 10727
rect 17592 10684 17644 10693
rect 16488 10548 16540 10600
rect 20628 10752 20680 10804
rect 18420 10659 18472 10668
rect 18420 10625 18429 10659
rect 18429 10625 18463 10659
rect 18463 10625 18472 10659
rect 18420 10616 18472 10625
rect 21364 10684 21416 10736
rect 19248 10616 19300 10668
rect 21088 10659 21140 10668
rect 21088 10625 21097 10659
rect 21097 10625 21131 10659
rect 21131 10625 21140 10659
rect 21088 10616 21140 10625
rect 23572 10752 23624 10804
rect 23388 10727 23440 10736
rect 23388 10693 23397 10727
rect 23397 10693 23431 10727
rect 23431 10693 23440 10727
rect 23388 10684 23440 10693
rect 22652 10616 22704 10668
rect 19432 10548 19484 10600
rect 19984 10591 20036 10600
rect 19984 10557 19993 10591
rect 19993 10557 20027 10591
rect 20027 10557 20036 10591
rect 19984 10548 20036 10557
rect 20168 10591 20220 10600
rect 20168 10557 20177 10591
rect 20177 10557 20211 10591
rect 20211 10557 20220 10591
rect 20168 10548 20220 10557
rect 21272 10591 21324 10600
rect 21272 10557 21281 10591
rect 21281 10557 21315 10591
rect 21315 10557 21324 10591
rect 21272 10548 21324 10557
rect 21916 10548 21968 10600
rect 24400 10548 24452 10600
rect 20352 10480 20404 10532
rect 8300 10412 8352 10464
rect 9128 10412 9180 10464
rect 9588 10412 9640 10464
rect 15660 10412 15712 10464
rect 16856 10455 16908 10464
rect 16856 10421 16865 10455
rect 16865 10421 16899 10455
rect 16899 10421 16908 10455
rect 16856 10412 16908 10421
rect 17040 10412 17092 10464
rect 18880 10455 18932 10464
rect 18880 10421 18889 10455
rect 18889 10421 18923 10455
rect 18923 10421 18932 10455
rect 18880 10412 18932 10421
rect 21364 10412 21416 10464
rect 21824 10412 21876 10464
rect 23388 10412 23440 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 11060 10251 11112 10260
rect 11060 10217 11069 10251
rect 11069 10217 11103 10251
rect 11103 10217 11112 10251
rect 11060 10208 11112 10217
rect 11520 10208 11572 10260
rect 11980 10208 12032 10260
rect 14556 10251 14608 10260
rect 14556 10217 14565 10251
rect 14565 10217 14599 10251
rect 14599 10217 14608 10251
rect 14556 10208 14608 10217
rect 14740 10208 14792 10260
rect 12716 10140 12768 10192
rect 13728 10140 13780 10192
rect 16028 10140 16080 10192
rect 16304 10140 16356 10192
rect 9588 10072 9640 10124
rect 12164 10115 12216 10124
rect 12164 10081 12173 10115
rect 12173 10081 12207 10115
rect 12207 10081 12216 10115
rect 12164 10072 12216 10081
rect 13544 10072 13596 10124
rect 14924 10072 14976 10124
rect 16856 10208 16908 10260
rect 20996 10208 21048 10260
rect 24584 10251 24636 10260
rect 24584 10217 24593 10251
rect 24593 10217 24627 10251
rect 24627 10217 24636 10251
rect 24584 10208 24636 10217
rect 18328 10140 18380 10192
rect 17684 10072 17736 10124
rect 17776 10072 17828 10124
rect 19800 10140 19852 10192
rect 19984 10140 20036 10192
rect 22284 10183 22336 10192
rect 22284 10149 22293 10183
rect 22293 10149 22327 10183
rect 22327 10149 22336 10183
rect 22284 10140 22336 10149
rect 18880 10072 18932 10124
rect 19524 10072 19576 10124
rect 20812 10115 20864 10124
rect 20812 10081 20821 10115
rect 20821 10081 20855 10115
rect 20855 10081 20864 10115
rect 20812 10072 20864 10081
rect 22008 10072 22060 10124
rect 23388 10115 23440 10124
rect 23388 10081 23397 10115
rect 23397 10081 23431 10115
rect 23431 10081 23440 10115
rect 23388 10072 23440 10081
rect 12072 10004 12124 10056
rect 9312 9936 9364 9988
rect 9864 9936 9916 9988
rect 13728 9936 13780 9988
rect 15016 10004 15068 10056
rect 16948 10004 17000 10056
rect 21916 10004 21968 10056
rect 24032 10004 24084 10056
rect 19064 9936 19116 9988
rect 12808 9868 12860 9920
rect 13452 9868 13504 9920
rect 13912 9911 13964 9920
rect 13912 9877 13921 9911
rect 13921 9877 13955 9911
rect 13955 9877 13964 9911
rect 13912 9868 13964 9877
rect 14832 9868 14884 9920
rect 15384 9868 15436 9920
rect 16120 9911 16172 9920
rect 16120 9877 16129 9911
rect 16129 9877 16163 9911
rect 16163 9877 16172 9911
rect 16120 9868 16172 9877
rect 16764 9868 16816 9920
rect 17684 9868 17736 9920
rect 18696 9868 18748 9920
rect 21180 9868 21232 9920
rect 23296 9936 23348 9988
rect 24216 9868 24268 9920
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 7104 9664 7156 9716
rect 9864 9596 9916 9648
rect 11152 9596 11204 9648
rect 11704 9571 11756 9580
rect 11704 9537 11713 9571
rect 11713 9537 11747 9571
rect 11747 9537 11756 9571
rect 11704 9528 11756 9537
rect 12532 9460 12584 9512
rect 11152 9324 11204 9376
rect 13912 9596 13964 9648
rect 14004 9596 14056 9648
rect 14464 9528 14516 9580
rect 14096 9460 14148 9512
rect 16120 9664 16172 9716
rect 20996 9664 21048 9716
rect 21088 9664 21140 9716
rect 22376 9664 22428 9716
rect 17868 9596 17920 9648
rect 19432 9596 19484 9648
rect 19340 9528 19392 9580
rect 22468 9528 22520 9580
rect 24032 9528 24084 9580
rect 14924 9460 14976 9512
rect 15660 9460 15712 9512
rect 16212 9460 16264 9512
rect 16948 9460 17000 9512
rect 17592 9503 17644 9512
rect 17592 9469 17601 9503
rect 17601 9469 17635 9503
rect 17635 9469 17644 9503
rect 17592 9460 17644 9469
rect 17960 9460 18012 9512
rect 19064 9460 19116 9512
rect 13728 9392 13780 9444
rect 15108 9435 15160 9444
rect 15108 9401 15117 9435
rect 15117 9401 15151 9435
rect 15151 9401 15160 9435
rect 15108 9392 15160 9401
rect 22008 9460 22060 9512
rect 22652 9503 22704 9512
rect 22652 9469 22661 9503
rect 22661 9469 22695 9503
rect 22695 9469 22704 9503
rect 22652 9460 22704 9469
rect 23388 9460 23440 9512
rect 17408 9324 17460 9376
rect 20444 9392 20496 9444
rect 21732 9392 21784 9444
rect 19156 9324 19208 9376
rect 19432 9367 19484 9376
rect 19432 9333 19441 9367
rect 19441 9333 19475 9367
rect 19475 9333 19484 9367
rect 19432 9324 19484 9333
rect 20352 9324 20404 9376
rect 21640 9324 21692 9376
rect 22744 9324 22796 9376
rect 24032 9392 24084 9444
rect 24400 9392 24452 9444
rect 24860 9367 24912 9376
rect 24860 9333 24869 9367
rect 24869 9333 24903 9367
rect 24903 9333 24912 9367
rect 24860 9324 24912 9333
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 11152 9163 11204 9172
rect 11152 9129 11161 9163
rect 11161 9129 11195 9163
rect 11195 9129 11204 9163
rect 11152 9120 11204 9129
rect 12808 9120 12860 9172
rect 15660 9120 15712 9172
rect 18512 9120 18564 9172
rect 18696 9120 18748 9172
rect 21548 9120 21600 9172
rect 21640 9120 21692 9172
rect 22744 9120 22796 9172
rect 23940 9120 23992 9172
rect 12624 9052 12676 9104
rect 13636 9052 13688 9104
rect 17868 9052 17920 9104
rect 19156 9052 19208 9104
rect 11060 8984 11112 9036
rect 11704 8984 11756 9036
rect 13544 9027 13596 9036
rect 13544 8993 13553 9027
rect 13553 8993 13587 9027
rect 13587 8993 13596 9027
rect 13544 8984 13596 8993
rect 14924 9027 14976 9036
rect 14924 8993 14933 9027
rect 14933 8993 14967 9027
rect 14967 8993 14976 9027
rect 14924 8984 14976 8993
rect 16488 9027 16540 9036
rect 16488 8993 16497 9027
rect 16497 8993 16531 9027
rect 16531 8993 16540 9027
rect 16488 8984 16540 8993
rect 14648 8959 14700 8968
rect 14648 8925 14657 8959
rect 14657 8925 14691 8959
rect 14691 8925 14700 8959
rect 14648 8916 14700 8925
rect 17408 8984 17460 9036
rect 18512 8984 18564 9036
rect 20444 8984 20496 9036
rect 9680 8848 9732 8900
rect 9864 8848 9916 8900
rect 10968 8780 11020 8832
rect 14188 8780 14240 8832
rect 14648 8780 14700 8832
rect 15936 8780 15988 8832
rect 16856 8780 16908 8832
rect 18696 8891 18748 8900
rect 18696 8857 18705 8891
rect 18705 8857 18739 8891
rect 18739 8857 18748 8891
rect 18696 8848 18748 8857
rect 19432 8848 19484 8900
rect 17500 8823 17552 8832
rect 17500 8789 17509 8823
rect 17509 8789 17543 8823
rect 17543 8789 17552 8823
rect 17500 8780 17552 8789
rect 17684 8780 17736 8832
rect 21640 8916 21692 8968
rect 22008 8959 22060 8968
rect 22008 8925 22017 8959
rect 22017 8925 22051 8959
rect 22051 8925 22060 8959
rect 22008 8916 22060 8925
rect 22652 8959 22704 8968
rect 22652 8925 22661 8959
rect 22661 8925 22695 8959
rect 22695 8925 22704 8959
rect 22652 8916 22704 8925
rect 23756 8916 23808 8968
rect 19984 8848 20036 8900
rect 20628 8780 20680 8832
rect 20812 8780 20864 8832
rect 23572 8848 23624 8900
rect 24952 8848 25004 8900
rect 22744 8780 22796 8832
rect 23940 8780 23992 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 15752 8576 15804 8628
rect 16856 8576 16908 8628
rect 17500 8576 17552 8628
rect 20260 8576 20312 8628
rect 21272 8576 21324 8628
rect 22468 8576 22520 8628
rect 24400 8576 24452 8628
rect 14280 8440 14332 8492
rect 11704 8415 11756 8424
rect 11704 8381 11713 8415
rect 11713 8381 11747 8415
rect 11747 8381 11756 8415
rect 11704 8372 11756 8381
rect 13360 8372 13412 8424
rect 10508 8304 10560 8356
rect 14096 8347 14148 8356
rect 14096 8313 14105 8347
rect 14105 8313 14139 8347
rect 14139 8313 14148 8347
rect 14096 8304 14148 8313
rect 14832 8415 14884 8424
rect 14832 8381 14841 8415
rect 14841 8381 14875 8415
rect 14875 8381 14884 8415
rect 14832 8372 14884 8381
rect 16120 8415 16172 8424
rect 16120 8381 16129 8415
rect 16129 8381 16163 8415
rect 16163 8381 16172 8415
rect 16120 8372 16172 8381
rect 17408 8415 17460 8424
rect 17408 8381 17417 8415
rect 17417 8381 17451 8415
rect 17451 8381 17460 8415
rect 17408 8372 17460 8381
rect 17776 8440 17828 8492
rect 18236 8483 18288 8492
rect 18236 8449 18245 8483
rect 18245 8449 18279 8483
rect 18279 8449 18288 8483
rect 18236 8440 18288 8449
rect 20076 8483 20128 8492
rect 20076 8449 20085 8483
rect 20085 8449 20119 8483
rect 20119 8449 20128 8483
rect 20076 8440 20128 8449
rect 17684 8372 17736 8424
rect 20536 8372 20588 8424
rect 21640 8372 21692 8424
rect 22284 8483 22336 8492
rect 22284 8449 22293 8483
rect 22293 8449 22327 8483
rect 22327 8449 22336 8483
rect 22284 8440 22336 8449
rect 22468 8372 22520 8424
rect 24768 8415 24820 8424
rect 24768 8381 24777 8415
rect 24777 8381 24811 8415
rect 24811 8381 24820 8415
rect 24768 8372 24820 8381
rect 19248 8304 19300 8356
rect 11152 8236 11204 8288
rect 17224 8236 17276 8288
rect 17960 8236 18012 8288
rect 22836 8236 22888 8288
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 11152 8032 11204 8084
rect 13544 8032 13596 8084
rect 14188 8032 14240 8084
rect 16488 8032 16540 8084
rect 21824 8032 21876 8084
rect 12532 7964 12584 8016
rect 11612 7939 11664 7948
rect 11612 7905 11621 7939
rect 11621 7905 11655 7939
rect 11655 7905 11664 7939
rect 11612 7896 11664 7905
rect 14556 7896 14608 7948
rect 15016 7964 15068 8016
rect 18420 7964 18472 8016
rect 20352 7964 20404 8016
rect 23480 8032 23532 8084
rect 16212 7896 16264 7948
rect 17500 7896 17552 7948
rect 20260 7896 20312 7948
rect 11704 7828 11756 7880
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 16120 7828 16172 7880
rect 2228 7692 2280 7744
rect 11152 7692 11204 7744
rect 12624 7692 12676 7744
rect 13360 7692 13412 7744
rect 15752 7760 15804 7812
rect 17960 7828 18012 7880
rect 19800 7828 19852 7880
rect 19892 7828 19944 7880
rect 20168 7828 20220 7880
rect 24032 7964 24084 8016
rect 22376 7939 22428 7948
rect 22376 7905 22385 7939
rect 22385 7905 22419 7939
rect 22419 7905 22428 7939
rect 22376 7896 22428 7905
rect 21732 7828 21784 7880
rect 23940 7828 23992 7880
rect 17776 7760 17828 7812
rect 18328 7760 18380 7812
rect 15016 7692 15068 7744
rect 16488 7692 16540 7744
rect 16856 7692 16908 7744
rect 17132 7692 17184 7744
rect 17868 7692 17920 7744
rect 21088 7760 21140 7812
rect 21456 7803 21508 7812
rect 21456 7769 21465 7803
rect 21465 7769 21499 7803
rect 21499 7769 21508 7803
rect 21456 7760 21508 7769
rect 20812 7692 20864 7744
rect 23848 7735 23900 7744
rect 23848 7701 23857 7735
rect 23857 7701 23891 7735
rect 23891 7701 23900 7735
rect 23848 7692 23900 7701
rect 23940 7692 23992 7744
rect 24768 7692 24820 7744
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 9588 7420 9640 7472
rect 11520 7420 11572 7472
rect 12624 7531 12676 7540
rect 12624 7497 12633 7531
rect 12633 7497 12667 7531
rect 12667 7497 12676 7531
rect 12624 7488 12676 7497
rect 13636 7488 13688 7540
rect 17776 7531 17828 7540
rect 17776 7497 17785 7531
rect 17785 7497 17819 7531
rect 17819 7497 17828 7531
rect 17776 7488 17828 7497
rect 19156 7488 19208 7540
rect 14280 7420 14332 7472
rect 15016 7420 15068 7472
rect 18788 7420 18840 7472
rect 20260 7488 20312 7540
rect 25320 7488 25372 7540
rect 20352 7420 20404 7472
rect 20996 7420 21048 7472
rect 21180 7420 21232 7472
rect 16396 7352 16448 7404
rect 17684 7395 17736 7404
rect 17684 7361 17693 7395
rect 17693 7361 17727 7395
rect 17727 7361 17736 7395
rect 17684 7352 17736 7361
rect 18512 7395 18564 7404
rect 18512 7361 18521 7395
rect 18521 7361 18555 7395
rect 18555 7361 18564 7395
rect 18512 7352 18564 7361
rect 25136 7463 25188 7472
rect 25136 7429 25145 7463
rect 25145 7429 25179 7463
rect 25179 7429 25188 7463
rect 25136 7420 25188 7429
rect 10968 7284 11020 7336
rect 11428 7284 11480 7336
rect 10784 7191 10836 7200
rect 10784 7157 10793 7191
rect 10793 7157 10827 7191
rect 10827 7157 10836 7191
rect 10784 7148 10836 7157
rect 11520 7148 11572 7200
rect 16672 7284 16724 7336
rect 17592 7284 17644 7336
rect 18880 7284 18932 7336
rect 19248 7284 19300 7336
rect 15108 7148 15160 7200
rect 15476 7148 15528 7200
rect 18328 7216 18380 7268
rect 19892 7216 19944 7268
rect 24860 7284 24912 7336
rect 24124 7216 24176 7268
rect 17224 7148 17276 7200
rect 17776 7148 17828 7200
rect 19248 7148 19300 7200
rect 22560 7148 22612 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 11612 6944 11664 6996
rect 16856 6944 16908 6996
rect 17132 6944 17184 6996
rect 19248 6944 19300 6996
rect 23940 6944 23992 6996
rect 11060 6808 11112 6860
rect 11520 6808 11572 6860
rect 12532 6851 12584 6860
rect 12532 6817 12541 6851
rect 12541 6817 12575 6851
rect 12575 6817 12584 6851
rect 12532 6808 12584 6817
rect 13728 6783 13780 6792
rect 13728 6749 13737 6783
rect 13737 6749 13771 6783
rect 13771 6749 13780 6783
rect 13728 6740 13780 6749
rect 14740 6740 14792 6792
rect 15016 6740 15068 6792
rect 21180 6876 21232 6928
rect 23848 6876 23900 6928
rect 15384 6808 15436 6860
rect 15752 6808 15804 6860
rect 16396 6740 16448 6792
rect 16948 6740 17000 6792
rect 19892 6808 19944 6860
rect 19984 6808 20036 6860
rect 23756 6808 23808 6860
rect 20352 6740 20404 6792
rect 20904 6783 20956 6792
rect 20904 6749 20913 6783
rect 20913 6749 20947 6783
rect 20947 6749 20956 6783
rect 20904 6740 20956 6749
rect 22652 6783 22704 6792
rect 22652 6749 22661 6783
rect 22661 6749 22695 6783
rect 22695 6749 22704 6783
rect 22652 6740 22704 6749
rect 24952 6740 25004 6792
rect 11336 6672 11388 6724
rect 11520 6672 11572 6724
rect 12808 6672 12860 6724
rect 15476 6715 15528 6724
rect 15476 6681 15485 6715
rect 15485 6681 15519 6715
rect 15519 6681 15528 6715
rect 15476 6672 15528 6681
rect 15844 6672 15896 6724
rect 16580 6672 16632 6724
rect 17408 6715 17460 6724
rect 17408 6681 17417 6715
rect 17417 6681 17451 6715
rect 17451 6681 17460 6715
rect 17408 6672 17460 6681
rect 13544 6647 13596 6656
rect 13544 6613 13553 6647
rect 13553 6613 13587 6647
rect 13587 6613 13596 6647
rect 13544 6604 13596 6613
rect 14372 6647 14424 6656
rect 14372 6613 14381 6647
rect 14381 6613 14415 6647
rect 14415 6613 14424 6647
rect 14372 6604 14424 6613
rect 15016 6604 15068 6656
rect 17224 6604 17276 6656
rect 19156 6672 19208 6724
rect 20996 6672 21048 6724
rect 22836 6672 22888 6724
rect 19892 6647 19944 6656
rect 19892 6613 19901 6647
rect 19901 6613 19935 6647
rect 19935 6613 19944 6647
rect 19892 6604 19944 6613
rect 21180 6604 21232 6656
rect 21364 6604 21416 6656
rect 24584 6647 24636 6656
rect 24584 6613 24593 6647
rect 24593 6613 24627 6647
rect 24627 6613 24636 6647
rect 24584 6604 24636 6613
rect 24676 6604 24728 6656
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 11428 6400 11480 6452
rect 13360 6400 13412 6452
rect 13820 6443 13872 6452
rect 13820 6409 13829 6443
rect 13829 6409 13863 6443
rect 13863 6409 13872 6443
rect 13820 6400 13872 6409
rect 14372 6400 14424 6452
rect 20812 6400 20864 6452
rect 6368 6264 6420 6316
rect 12072 6307 12124 6316
rect 12072 6273 12081 6307
rect 12081 6273 12115 6307
rect 12115 6273 12124 6307
rect 12072 6264 12124 6273
rect 13268 6332 13320 6384
rect 13544 6332 13596 6384
rect 10876 6239 10928 6248
rect 10876 6205 10885 6239
rect 10885 6205 10919 6239
rect 10919 6205 10928 6239
rect 10876 6196 10928 6205
rect 10968 6239 11020 6248
rect 10968 6205 10977 6239
rect 10977 6205 11011 6239
rect 11011 6205 11020 6239
rect 10968 6196 11020 6205
rect 12348 6239 12400 6248
rect 12348 6205 12357 6239
rect 12357 6205 12391 6239
rect 12391 6205 12400 6239
rect 12348 6196 12400 6205
rect 8300 6060 8352 6112
rect 13820 6264 13872 6316
rect 12900 6239 12952 6248
rect 12900 6205 12909 6239
rect 12909 6205 12943 6239
rect 12943 6205 12952 6239
rect 12900 6196 12952 6205
rect 13636 6128 13688 6180
rect 16120 6239 16172 6248
rect 16120 6205 16129 6239
rect 16129 6205 16163 6239
rect 16163 6205 16172 6239
rect 16120 6196 16172 6205
rect 17316 6264 17368 6316
rect 19248 6332 19300 6384
rect 22192 6400 22244 6452
rect 22376 6400 22428 6452
rect 24584 6400 24636 6452
rect 25228 6400 25280 6452
rect 18328 6264 18380 6316
rect 19892 6264 19944 6316
rect 20260 6307 20312 6316
rect 20260 6273 20269 6307
rect 20269 6273 20303 6307
rect 20303 6273 20312 6307
rect 20260 6264 20312 6273
rect 21824 6264 21876 6316
rect 16856 6239 16908 6248
rect 16856 6205 16865 6239
rect 16865 6205 16899 6239
rect 16899 6205 16908 6239
rect 16856 6196 16908 6205
rect 20628 6128 20680 6180
rect 21732 6196 21784 6248
rect 23848 6264 23900 6316
rect 24216 6375 24268 6384
rect 24216 6341 24225 6375
rect 24225 6341 24259 6375
rect 24259 6341 24268 6375
rect 24216 6332 24268 6341
rect 24768 6264 24820 6316
rect 25044 6307 25096 6316
rect 25044 6273 25053 6307
rect 25053 6273 25087 6307
rect 25087 6273 25096 6307
rect 25044 6264 25096 6273
rect 23756 6239 23808 6248
rect 23756 6205 23765 6239
rect 23765 6205 23799 6239
rect 23799 6205 23808 6239
rect 23756 6196 23808 6205
rect 22008 6128 22060 6180
rect 13360 6103 13412 6112
rect 13360 6069 13369 6103
rect 13369 6069 13403 6103
rect 13403 6069 13412 6103
rect 13360 6060 13412 6069
rect 16396 6060 16448 6112
rect 17592 6060 17644 6112
rect 22100 6060 22152 6112
rect 24768 6060 24820 6112
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 11336 5856 11388 5908
rect 12348 5856 12400 5908
rect 14740 5899 14792 5908
rect 14740 5865 14749 5899
rect 14749 5865 14783 5899
rect 14783 5865 14792 5899
rect 14740 5856 14792 5865
rect 14924 5788 14976 5840
rect 10784 5720 10836 5772
rect 13360 5720 13412 5772
rect 17408 5856 17460 5908
rect 20260 5856 20312 5908
rect 9588 5652 9640 5704
rect 11428 5652 11480 5704
rect 13452 5652 13504 5704
rect 15016 5652 15068 5704
rect 15108 5652 15160 5704
rect 16948 5720 17000 5772
rect 17224 5720 17276 5772
rect 19340 5720 19392 5772
rect 17316 5652 17368 5704
rect 17592 5652 17644 5704
rect 19616 5695 19668 5704
rect 19616 5661 19625 5695
rect 19625 5661 19659 5695
rect 19659 5661 19668 5695
rect 19616 5652 19668 5661
rect 11704 5584 11756 5636
rect 15752 5584 15804 5636
rect 20628 5788 20680 5840
rect 20720 5720 20772 5772
rect 23572 5720 23624 5772
rect 21088 5652 21140 5704
rect 22744 5652 22796 5704
rect 23664 5652 23716 5704
rect 13544 5559 13596 5568
rect 13544 5525 13553 5559
rect 13553 5525 13587 5559
rect 13587 5525 13596 5559
rect 13544 5516 13596 5525
rect 16856 5516 16908 5568
rect 18328 5516 18380 5568
rect 23756 5584 23808 5636
rect 25136 5516 25188 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 7840 5312 7892 5364
rect 11244 5312 11296 5364
rect 13636 5312 13688 5364
rect 18880 5312 18932 5364
rect 21180 5312 21232 5364
rect 15016 5244 15068 5296
rect 15476 5244 15528 5296
rect 19156 5244 19208 5296
rect 20352 5244 20404 5296
rect 20444 5244 20496 5296
rect 11060 5108 11112 5160
rect 18144 5151 18196 5160
rect 18144 5117 18153 5151
rect 18153 5117 18187 5151
rect 18187 5117 18196 5151
rect 18144 5108 18196 5117
rect 17960 5040 18012 5092
rect 13912 4972 13964 5024
rect 14188 4972 14240 5024
rect 14924 5015 14976 5024
rect 14924 4981 14933 5015
rect 14933 4981 14967 5015
rect 14967 4981 14976 5015
rect 14924 4972 14976 4981
rect 18512 5176 18564 5228
rect 21088 5219 21140 5228
rect 21088 5185 21097 5219
rect 21097 5185 21131 5219
rect 21131 5185 21140 5219
rect 21088 5176 21140 5185
rect 22100 5219 22152 5228
rect 22100 5185 22109 5219
rect 22109 5185 22143 5219
rect 22143 5185 22152 5219
rect 22100 5176 22152 5185
rect 23756 5176 23808 5228
rect 21180 5108 21232 5160
rect 21364 5108 21416 5160
rect 20444 4972 20496 5024
rect 23848 4972 23900 5024
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 12256 4743 12308 4752
rect 12256 4709 12265 4743
rect 12265 4709 12299 4743
rect 12299 4709 12308 4743
rect 12256 4700 12308 4709
rect 9588 4632 9640 4684
rect 11428 4564 11480 4616
rect 12624 4700 12676 4752
rect 17224 4768 17276 4820
rect 19064 4768 19116 4820
rect 21088 4768 21140 4820
rect 21180 4768 21232 4820
rect 24032 4768 24084 4820
rect 13820 4632 13872 4684
rect 15108 4675 15160 4684
rect 15108 4641 15117 4675
rect 15117 4641 15151 4675
rect 15151 4641 15160 4675
rect 15108 4632 15160 4641
rect 17316 4700 17368 4752
rect 17408 4632 17460 4684
rect 17500 4632 17552 4684
rect 18512 4632 18564 4684
rect 19800 4675 19852 4684
rect 19800 4641 19809 4675
rect 19809 4641 19843 4675
rect 19843 4641 19852 4675
rect 19800 4632 19852 4641
rect 19892 4632 19944 4684
rect 22376 4632 22428 4684
rect 5356 4539 5408 4548
rect 5356 4505 5365 4539
rect 5365 4505 5399 4539
rect 5399 4505 5408 4539
rect 5356 4496 5408 4505
rect 7104 4539 7156 4548
rect 7104 4505 7113 4539
rect 7113 4505 7147 4539
rect 7147 4505 7156 4539
rect 7104 4496 7156 4505
rect 15108 4496 15160 4548
rect 15384 4539 15436 4548
rect 15384 4505 15393 4539
rect 15393 4505 15427 4539
rect 15427 4505 15436 4539
rect 15384 4496 15436 4505
rect 15476 4496 15528 4548
rect 15844 4496 15896 4548
rect 24308 4564 24360 4616
rect 24492 4564 24544 4616
rect 19524 4496 19576 4548
rect 20352 4496 20404 4548
rect 1492 4471 1544 4480
rect 1492 4437 1501 4471
rect 1501 4437 1535 4471
rect 1535 4437 1544 4471
rect 1492 4428 1544 4437
rect 11152 4428 11204 4480
rect 14924 4428 14976 4480
rect 18144 4428 18196 4480
rect 22284 4428 22336 4480
rect 23756 4471 23808 4480
rect 23756 4437 23765 4471
rect 23765 4437 23799 4471
rect 23799 4437 23808 4471
rect 23756 4428 23808 4437
rect 24768 4428 24820 4480
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 14188 4199 14240 4208
rect 14188 4165 14197 4199
rect 14197 4165 14231 4199
rect 14231 4165 14240 4199
rect 14188 4156 14240 4165
rect 14924 4156 14976 4208
rect 18328 4224 18380 4276
rect 20352 4224 20404 4276
rect 21824 4224 21876 4276
rect 17132 4156 17184 4208
rect 17408 4156 17460 4208
rect 19616 4156 19668 4208
rect 1492 4088 1544 4140
rect 1860 4088 1912 4140
rect 4068 4088 4120 4140
rect 9220 4088 9272 4140
rect 10968 4131 11020 4140
rect 10968 4097 10977 4131
rect 10977 4097 11011 4131
rect 11011 4097 11020 4131
rect 10968 4088 11020 4097
rect 12256 4131 12308 4140
rect 12256 4097 12265 4131
rect 12265 4097 12299 4131
rect 12299 4097 12308 4131
rect 12256 4088 12308 4097
rect 13912 4131 13964 4140
rect 13912 4097 13921 4131
rect 13921 4097 13955 4131
rect 13955 4097 13964 4131
rect 13912 4088 13964 4097
rect 18696 4088 18748 4140
rect 18788 4131 18840 4140
rect 18788 4097 18797 4131
rect 18797 4097 18831 4131
rect 18831 4097 18840 4131
rect 18788 4088 18840 4097
rect 19524 4088 19576 4140
rect 20904 4131 20956 4140
rect 20904 4097 20913 4131
rect 20913 4097 20947 4131
rect 20947 4097 20956 4131
rect 20904 4088 20956 4097
rect 20996 4131 21048 4140
rect 20996 4097 21005 4131
rect 21005 4097 21039 4131
rect 21039 4097 21048 4131
rect 20996 4088 21048 4097
rect 5356 4020 5408 4072
rect 2228 3995 2280 4004
rect 2228 3961 2237 3995
rect 2237 3961 2271 3995
rect 2271 3961 2280 3995
rect 2228 3952 2280 3961
rect 6920 3952 6972 4004
rect 12808 4020 12860 4072
rect 16028 4020 16080 4072
rect 16212 4020 16264 4072
rect 18328 4020 18380 4072
rect 20536 4020 20588 4072
rect 21548 4088 21600 4140
rect 22100 4088 22152 4140
rect 22376 4088 22428 4140
rect 21180 4063 21232 4072
rect 21180 4029 21189 4063
rect 21189 4029 21223 4063
rect 21223 4029 21232 4063
rect 21180 4020 21232 4029
rect 23848 4131 23900 4140
rect 23848 4097 23857 4131
rect 23857 4097 23891 4131
rect 23891 4097 23900 4131
rect 23848 4088 23900 4097
rect 25412 4088 25464 4140
rect 9404 3952 9456 4004
rect 12440 3952 12492 4004
rect 15476 3952 15528 4004
rect 20996 3952 21048 4004
rect 2872 3927 2924 3936
rect 2872 3893 2881 3927
rect 2881 3893 2915 3927
rect 2915 3893 2924 3927
rect 2872 3884 2924 3893
rect 10600 3927 10652 3936
rect 10600 3893 10609 3927
rect 10609 3893 10643 3927
rect 10643 3893 10652 3927
rect 10600 3884 10652 3893
rect 11612 3927 11664 3936
rect 11612 3893 11621 3927
rect 11621 3893 11655 3927
rect 11655 3893 11664 3927
rect 11612 3884 11664 3893
rect 12532 3884 12584 3936
rect 13360 3884 13412 3936
rect 20168 3884 20220 3936
rect 20536 3927 20588 3936
rect 20536 3893 20545 3927
rect 20545 3893 20579 3927
rect 20579 3893 20588 3927
rect 20536 3884 20588 3893
rect 21548 3884 21600 3936
rect 22376 3884 22428 3936
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 3332 3680 3384 3732
rect 7656 3680 7708 3732
rect 10876 3680 10928 3732
rect 10968 3680 11020 3732
rect 15936 3680 15988 3732
rect 17960 3723 18012 3732
rect 17960 3689 17969 3723
rect 17969 3689 18003 3723
rect 18003 3689 18012 3723
rect 17960 3680 18012 3689
rect 22100 3680 22152 3732
rect 22744 3680 22796 3732
rect 6368 3655 6420 3664
rect 6368 3621 6377 3655
rect 6377 3621 6411 3655
rect 6411 3621 6420 3655
rect 6368 3612 6420 3621
rect 9404 3612 9456 3664
rect 2872 3544 2924 3596
rect 3700 3544 3752 3596
rect 5172 3587 5224 3596
rect 5172 3553 5181 3587
rect 5181 3553 5215 3587
rect 5215 3553 5224 3587
rect 5172 3544 5224 3553
rect 5448 3544 5500 3596
rect 12716 3612 12768 3664
rect 16028 3612 16080 3664
rect 23480 3612 23532 3664
rect 24952 3655 25004 3664
rect 24952 3621 24961 3655
rect 24961 3621 24995 3655
rect 24995 3621 25004 3655
rect 24952 3612 25004 3621
rect 12532 3544 12584 3596
rect 12808 3587 12860 3596
rect 12808 3553 12817 3587
rect 12817 3553 12851 3587
rect 12851 3553 12860 3587
rect 12808 3544 12860 3553
rect 14004 3544 14056 3596
rect 15476 3544 15528 3596
rect 17684 3544 17736 3596
rect 2228 3476 2280 3528
rect 4436 3519 4488 3528
rect 4436 3485 4445 3519
rect 4445 3485 4479 3519
rect 4479 3485 4488 3519
rect 4436 3476 4488 3485
rect 4896 3519 4948 3528
rect 4896 3485 4905 3519
rect 4905 3485 4939 3519
rect 4939 3485 4948 3519
rect 4896 3476 4948 3485
rect 6276 3476 6328 3528
rect 7012 3476 7064 3528
rect 8484 3476 8536 3528
rect 9588 3476 9640 3528
rect 10600 3519 10652 3528
rect 10600 3485 10609 3519
rect 10609 3485 10643 3519
rect 10643 3485 10652 3519
rect 10600 3476 10652 3485
rect 9312 3408 9364 3460
rect 13360 3476 13412 3528
rect 14464 3519 14516 3528
rect 14464 3485 14473 3519
rect 14473 3485 14507 3519
rect 14507 3485 14516 3519
rect 14464 3476 14516 3485
rect 17040 3476 17092 3528
rect 19248 3476 19300 3528
rect 19432 3519 19484 3528
rect 19432 3485 19441 3519
rect 19441 3485 19475 3519
rect 19475 3485 19484 3519
rect 19432 3476 19484 3485
rect 20812 3476 20864 3528
rect 3424 3383 3476 3392
rect 3424 3349 3433 3383
rect 3433 3349 3467 3383
rect 3467 3349 3476 3383
rect 3424 3340 3476 3349
rect 7380 3340 7432 3392
rect 10416 3383 10468 3392
rect 10416 3349 10425 3383
rect 10425 3349 10459 3383
rect 10459 3349 10468 3383
rect 10416 3340 10468 3349
rect 14280 3340 14332 3392
rect 14556 3408 14608 3460
rect 18880 3408 18932 3460
rect 23940 3544 23992 3596
rect 22560 3476 22612 3528
rect 25136 3519 25188 3528
rect 25136 3485 25145 3519
rect 25145 3485 25179 3519
rect 25179 3485 25188 3519
rect 25136 3476 25188 3485
rect 21824 3408 21876 3460
rect 24768 3408 24820 3460
rect 14648 3340 14700 3392
rect 20812 3340 20864 3392
rect 21272 3340 21324 3392
rect 21456 3340 21508 3392
rect 22836 3340 22888 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 4436 3136 4488 3188
rect 4896 3136 4948 3188
rect 7840 3068 7892 3120
rect 10968 3179 11020 3188
rect 10968 3145 10977 3179
rect 10977 3145 11011 3179
rect 11011 3145 11020 3179
rect 10968 3136 11020 3145
rect 12072 3136 12124 3188
rect 20444 3136 20496 3188
rect 20904 3136 20956 3188
rect 24676 3136 24728 3188
rect 24768 3136 24820 3188
rect 2596 3000 2648 3052
rect 3424 3043 3476 3052
rect 3424 3009 3433 3043
rect 3433 3009 3467 3043
rect 3467 3009 3476 3043
rect 3424 3000 3476 3009
rect 5264 3000 5316 3052
rect 5448 3043 5500 3052
rect 5448 3009 5457 3043
rect 5457 3009 5491 3043
rect 5491 3009 5500 3043
rect 5448 3000 5500 3009
rect 6644 3000 6696 3052
rect 7380 3043 7432 3052
rect 7380 3009 7389 3043
rect 7389 3009 7423 3043
rect 7423 3009 7432 3043
rect 7380 3000 7432 3009
rect 10324 3000 10376 3052
rect 11796 3068 11848 3120
rect 11060 3000 11112 3052
rect 11152 3043 11204 3052
rect 11152 3009 11161 3043
rect 11161 3009 11195 3043
rect 11195 3009 11204 3043
rect 11152 3000 11204 3009
rect 11612 3000 11664 3052
rect 13912 3068 13964 3120
rect 16580 3068 16632 3120
rect 13176 3043 13228 3052
rect 13176 3009 13185 3043
rect 13185 3009 13219 3043
rect 13219 3009 13228 3043
rect 13176 3000 13228 3009
rect 14096 3000 14148 3052
rect 15016 3000 15068 3052
rect 15384 3000 15436 3052
rect 18604 3000 18656 3052
rect 18972 3000 19024 3052
rect 5172 2975 5224 2984
rect 5172 2941 5181 2975
rect 5181 2941 5215 2975
rect 5215 2941 5224 2975
rect 5172 2932 5224 2941
rect 7748 2932 7800 2984
rect 10416 2932 10468 2984
rect 8944 2864 8996 2916
rect 13636 2975 13688 2984
rect 13636 2941 13645 2975
rect 13645 2941 13679 2975
rect 13679 2941 13688 2975
rect 13636 2932 13688 2941
rect 14740 2932 14792 2984
rect 15844 2932 15896 2984
rect 22192 3068 22244 3120
rect 20812 3043 20864 3052
rect 20812 3009 20821 3043
rect 20821 3009 20855 3043
rect 20855 3009 20864 3043
rect 20812 3000 20864 3009
rect 23572 3043 23624 3052
rect 23572 3009 23581 3043
rect 23581 3009 23615 3043
rect 23615 3009 23624 3043
rect 23572 3000 23624 3009
rect 20076 2932 20128 2984
rect 7196 2839 7248 2848
rect 7196 2805 7205 2839
rect 7205 2805 7239 2839
rect 7239 2805 7248 2839
rect 7196 2796 7248 2805
rect 9036 2839 9088 2848
rect 9036 2805 9045 2839
rect 9045 2805 9079 2839
rect 9079 2805 9088 2839
rect 9036 2796 9088 2805
rect 10508 2796 10560 2848
rect 16304 2864 16356 2916
rect 16948 2864 17000 2916
rect 20352 2864 20404 2916
rect 22100 2864 22152 2916
rect 15016 2796 15068 2848
rect 15108 2796 15160 2848
rect 17316 2796 17368 2848
rect 18420 2796 18472 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 11888 2592 11940 2644
rect 15200 2592 15252 2644
rect 19616 2592 19668 2644
rect 23572 2592 23624 2644
rect 24308 2592 24360 2644
rect 9680 2524 9732 2576
rect 5448 2499 5500 2508
rect 5448 2465 5457 2499
rect 5457 2465 5491 2499
rect 5491 2465 5500 2499
rect 5448 2456 5500 2465
rect 2964 2388 3016 2440
rect 5540 2388 5592 2440
rect 5908 2320 5960 2372
rect 2596 2252 2648 2304
rect 5172 2252 5224 2304
rect 6644 2252 6696 2304
rect 8300 2456 8352 2508
rect 7840 2388 7892 2440
rect 9036 2388 9088 2440
rect 12624 2524 12676 2576
rect 13544 2524 13596 2576
rect 12164 2456 12216 2508
rect 14372 2456 14424 2508
rect 8852 2320 8904 2372
rect 9956 2320 10008 2372
rect 10968 2363 11020 2372
rect 10968 2329 10977 2363
rect 10977 2329 11011 2363
rect 11011 2329 11020 2363
rect 10968 2320 11020 2329
rect 7748 2295 7800 2304
rect 7748 2261 7757 2295
rect 7757 2261 7791 2295
rect 7791 2261 7800 2295
rect 7748 2252 7800 2261
rect 8392 2295 8444 2304
rect 8392 2261 8401 2295
rect 8401 2261 8435 2295
rect 8435 2261 8444 2295
rect 8392 2252 8444 2261
rect 11704 2295 11756 2304
rect 11704 2261 11713 2295
rect 11713 2261 11747 2295
rect 11747 2261 11756 2295
rect 11704 2252 11756 2261
rect 13268 2363 13320 2372
rect 13268 2329 13277 2363
rect 13277 2329 13311 2363
rect 13311 2329 13320 2363
rect 13268 2320 13320 2329
rect 16120 2524 16172 2576
rect 22284 2524 22336 2576
rect 22652 2524 22704 2576
rect 17316 2499 17368 2508
rect 17316 2465 17325 2499
rect 17325 2465 17359 2499
rect 17359 2465 17368 2499
rect 17316 2456 17368 2465
rect 16028 2388 16080 2440
rect 16764 2388 16816 2440
rect 20536 2456 20588 2508
rect 19708 2388 19760 2440
rect 20352 2431 20404 2440
rect 20352 2397 20361 2431
rect 20361 2397 20395 2431
rect 20395 2397 20404 2431
rect 20352 2388 20404 2397
rect 16304 2363 16356 2372
rect 16304 2329 16313 2363
rect 16313 2329 16347 2363
rect 16347 2329 16356 2363
rect 16304 2320 16356 2329
rect 16672 2320 16724 2372
rect 22192 2456 22244 2508
rect 15660 2252 15712 2304
rect 17776 2252 17828 2304
rect 23388 2388 23440 2440
rect 24952 2388 25004 2440
rect 23848 2295 23900 2304
rect 23848 2261 23857 2295
rect 23857 2261 23891 2295
rect 23891 2261 23900 2295
rect 23848 2252 23900 2261
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 13728 1980 13780 2032
rect 23848 1980 23900 2032
rect 8392 1912 8444 1964
rect 15568 1912 15620 1964
rect 10968 1776 11020 1828
rect 22100 1776 22152 1828
rect 21640 1232 21692 1284
rect 23204 1232 23256 1284
<< metal2 >>
rect 1030 56200 1086 57000
rect 2410 56200 2466 57000
rect 3790 56200 3846 57000
rect 5170 56200 5226 57000
rect 6550 56200 6606 57000
rect 7930 56200 7986 57000
rect 9310 56200 9366 57000
rect 10690 56200 10746 57000
rect 12070 56200 12126 57000
rect 12176 56222 12388 56250
rect 1044 53650 1072 56200
rect 2424 54126 2452 56200
rect 2412 54120 2464 54126
rect 2412 54062 2464 54068
rect 2950 53884 3258 53893
rect 2950 53882 2956 53884
rect 3012 53882 3036 53884
rect 3092 53882 3116 53884
rect 3172 53882 3196 53884
rect 3252 53882 3258 53884
rect 3012 53830 3014 53882
rect 3194 53830 3196 53882
rect 2950 53828 2956 53830
rect 3012 53828 3036 53830
rect 3092 53828 3116 53830
rect 3172 53828 3196 53830
rect 3252 53828 3258 53830
rect 2950 53819 3258 53828
rect 3804 53650 3832 56200
rect 4068 54188 4120 54194
rect 4068 54130 4120 54136
rect 4804 54188 4856 54194
rect 4804 54130 4856 54136
rect 1032 53644 1084 53650
rect 1032 53586 1084 53592
rect 3792 53644 3844 53650
rect 3792 53586 3844 53592
rect 4080 53242 4108 54130
rect 4160 53576 4212 53582
rect 4160 53518 4212 53524
rect 4068 53236 4120 53242
rect 4068 53178 4120 53184
rect 2950 52796 3258 52805
rect 2950 52794 2956 52796
rect 3012 52794 3036 52796
rect 3092 52794 3116 52796
rect 3172 52794 3196 52796
rect 3252 52794 3258 52796
rect 3012 52742 3014 52794
rect 3194 52742 3196 52794
rect 2950 52740 2956 52742
rect 3012 52740 3036 52742
rect 3092 52740 3116 52742
rect 3172 52740 3196 52742
rect 3252 52740 3258 52742
rect 2950 52731 3258 52740
rect 4172 52698 4200 53518
rect 4160 52692 4212 52698
rect 4160 52634 4212 52640
rect 2950 51708 3258 51717
rect 2950 51706 2956 51708
rect 3012 51706 3036 51708
rect 3092 51706 3116 51708
rect 3172 51706 3196 51708
rect 3252 51706 3258 51708
rect 3012 51654 3014 51706
rect 3194 51654 3196 51706
rect 2950 51652 2956 51654
rect 3012 51652 3036 51654
rect 3092 51652 3116 51654
rect 3172 51652 3196 51654
rect 3252 51652 3258 51654
rect 2950 51643 3258 51652
rect 4816 51406 4844 54130
rect 5184 54126 5212 56200
rect 5172 54120 5224 54126
rect 5172 54062 5224 54068
rect 6564 53650 6592 56200
rect 7944 55214 7972 56200
rect 7852 55186 7972 55214
rect 7380 54188 7432 54194
rect 7380 54130 7432 54136
rect 6552 53644 6604 53650
rect 6552 53586 6604 53592
rect 5540 53508 5592 53514
rect 5540 53450 5592 53456
rect 4804 51400 4856 51406
rect 4804 51342 4856 51348
rect 2950 50620 3258 50629
rect 2950 50618 2956 50620
rect 3012 50618 3036 50620
rect 3092 50618 3116 50620
rect 3172 50618 3196 50620
rect 3252 50618 3258 50620
rect 3012 50566 3014 50618
rect 3194 50566 3196 50618
rect 2950 50564 2956 50566
rect 3012 50564 3036 50566
rect 3092 50564 3116 50566
rect 3172 50564 3196 50566
rect 3252 50564 3258 50566
rect 2950 50555 3258 50564
rect 5552 50522 5580 53450
rect 7392 51610 7420 54130
rect 7852 54126 7880 55186
rect 7950 54428 8258 54437
rect 7950 54426 7956 54428
rect 8012 54426 8036 54428
rect 8092 54426 8116 54428
rect 8172 54426 8196 54428
rect 8252 54426 8258 54428
rect 8012 54374 8014 54426
rect 8194 54374 8196 54426
rect 7950 54372 7956 54374
rect 8012 54372 8036 54374
rect 8092 54372 8116 54374
rect 8172 54372 8196 54374
rect 8252 54372 8258 54374
rect 7950 54363 8258 54372
rect 9324 54126 9352 56200
rect 9588 54188 9640 54194
rect 9588 54130 9640 54136
rect 7840 54120 7892 54126
rect 7840 54062 7892 54068
rect 9312 54120 9364 54126
rect 9312 54062 9364 54068
rect 8300 54052 8352 54058
rect 8300 53994 8352 54000
rect 7840 53576 7892 53582
rect 7840 53518 7892 53524
rect 7748 53100 7800 53106
rect 7748 53042 7800 53048
rect 7380 51604 7432 51610
rect 7380 51546 7432 51552
rect 5540 50516 5592 50522
rect 5540 50458 5592 50464
rect 7760 50454 7788 53042
rect 7852 51542 7880 53518
rect 7950 53340 8258 53349
rect 7950 53338 7956 53340
rect 8012 53338 8036 53340
rect 8092 53338 8116 53340
rect 8172 53338 8196 53340
rect 8252 53338 8258 53340
rect 8012 53286 8014 53338
rect 8194 53286 8196 53338
rect 7950 53284 7956 53286
rect 8012 53284 8036 53286
rect 8092 53284 8116 53286
rect 8172 53284 8196 53286
rect 8252 53284 8258 53286
rect 7950 53275 8258 53284
rect 7950 52252 8258 52261
rect 7950 52250 7956 52252
rect 8012 52250 8036 52252
rect 8092 52250 8116 52252
rect 8172 52250 8196 52252
rect 8252 52250 8258 52252
rect 8012 52198 8014 52250
rect 8194 52198 8196 52250
rect 7950 52196 7956 52198
rect 8012 52196 8036 52198
rect 8092 52196 8116 52198
rect 8172 52196 8196 52198
rect 8252 52196 8258 52198
rect 7950 52187 8258 52196
rect 7840 51536 7892 51542
rect 7840 51478 7892 51484
rect 7950 51164 8258 51173
rect 7950 51162 7956 51164
rect 8012 51162 8036 51164
rect 8092 51162 8116 51164
rect 8172 51162 8196 51164
rect 8252 51162 8258 51164
rect 8012 51110 8014 51162
rect 8194 51110 8196 51162
rect 7950 51108 7956 51110
rect 8012 51108 8036 51110
rect 8092 51108 8116 51110
rect 8172 51108 8196 51110
rect 8252 51108 8258 51110
rect 7950 51099 8258 51108
rect 7748 50448 7800 50454
rect 7748 50390 7800 50396
rect 2950 49532 3258 49541
rect 2950 49530 2956 49532
rect 3012 49530 3036 49532
rect 3092 49530 3116 49532
rect 3172 49530 3196 49532
rect 3252 49530 3258 49532
rect 3012 49478 3014 49530
rect 3194 49478 3196 49530
rect 2950 49476 2956 49478
rect 3012 49476 3036 49478
rect 3092 49476 3116 49478
rect 3172 49476 3196 49478
rect 3252 49476 3258 49478
rect 2950 49467 3258 49476
rect 2950 48444 3258 48453
rect 2950 48442 2956 48444
rect 3012 48442 3036 48444
rect 3092 48442 3116 48444
rect 3172 48442 3196 48444
rect 3252 48442 3258 48444
rect 3012 48390 3014 48442
rect 3194 48390 3196 48442
rect 2950 48388 2956 48390
rect 3012 48388 3036 48390
rect 3092 48388 3116 48390
rect 3172 48388 3196 48390
rect 3252 48388 3258 48390
rect 2950 48379 3258 48388
rect 7760 48142 7788 50390
rect 8312 50318 8340 53994
rect 9404 52488 9456 52494
rect 9404 52430 9456 52436
rect 8484 51400 8536 51406
rect 8484 51342 8536 51348
rect 8392 50516 8444 50522
rect 8392 50458 8444 50464
rect 8300 50312 8352 50318
rect 8300 50254 8352 50260
rect 7950 50076 8258 50085
rect 7950 50074 7956 50076
rect 8012 50074 8036 50076
rect 8092 50074 8116 50076
rect 8172 50074 8196 50076
rect 8252 50074 8258 50076
rect 8012 50022 8014 50074
rect 8194 50022 8196 50074
rect 7950 50020 7956 50022
rect 8012 50020 8036 50022
rect 8092 50020 8116 50022
rect 8172 50020 8196 50022
rect 8252 50020 8258 50022
rect 7950 50011 8258 50020
rect 7950 48988 8258 48997
rect 7950 48986 7956 48988
rect 8012 48986 8036 48988
rect 8092 48986 8116 48988
rect 8172 48986 8196 48988
rect 8252 48986 8258 48988
rect 8012 48934 8014 48986
rect 8194 48934 8196 48986
rect 7950 48932 7956 48934
rect 8012 48932 8036 48934
rect 8092 48932 8116 48934
rect 8172 48932 8196 48934
rect 8252 48932 8258 48934
rect 7950 48923 8258 48932
rect 7748 48136 7800 48142
rect 7748 48078 7800 48084
rect 2950 47356 3258 47365
rect 2950 47354 2956 47356
rect 3012 47354 3036 47356
rect 3092 47354 3116 47356
rect 3172 47354 3196 47356
rect 3252 47354 3258 47356
rect 3012 47302 3014 47354
rect 3194 47302 3196 47354
rect 2950 47300 2956 47302
rect 3012 47300 3036 47302
rect 3092 47300 3116 47302
rect 3172 47300 3196 47302
rect 3252 47300 3258 47302
rect 2950 47291 3258 47300
rect 2950 46268 3258 46277
rect 2950 46266 2956 46268
rect 3012 46266 3036 46268
rect 3092 46266 3116 46268
rect 3172 46266 3196 46268
rect 3252 46266 3258 46268
rect 3012 46214 3014 46266
rect 3194 46214 3196 46266
rect 2950 46212 2956 46214
rect 3012 46212 3036 46214
rect 3092 46212 3116 46214
rect 3172 46212 3196 46214
rect 3252 46212 3258 46214
rect 2950 46203 3258 46212
rect 7760 46034 7788 48078
rect 7950 47900 8258 47909
rect 7950 47898 7956 47900
rect 8012 47898 8036 47900
rect 8092 47898 8116 47900
rect 8172 47898 8196 47900
rect 8252 47898 8258 47900
rect 8012 47846 8014 47898
rect 8194 47846 8196 47898
rect 7950 47844 7956 47846
rect 8012 47844 8036 47846
rect 8092 47844 8116 47846
rect 8172 47844 8196 47846
rect 8252 47844 8258 47846
rect 7950 47835 8258 47844
rect 8312 47666 8340 50254
rect 8404 48890 8432 50458
rect 8392 48884 8444 48890
rect 8392 48826 8444 48832
rect 8300 47660 8352 47666
rect 8300 47602 8352 47608
rect 7950 46812 8258 46821
rect 7950 46810 7956 46812
rect 8012 46810 8036 46812
rect 8092 46810 8116 46812
rect 8172 46810 8196 46812
rect 8252 46810 8258 46812
rect 8012 46758 8014 46810
rect 8194 46758 8196 46810
rect 7950 46756 7956 46758
rect 8012 46756 8036 46758
rect 8092 46756 8116 46758
rect 8172 46756 8196 46758
rect 8252 46756 8258 46758
rect 7950 46747 8258 46756
rect 8496 46170 8524 51342
rect 9128 48612 9180 48618
rect 9128 48554 9180 48560
rect 8484 46164 8536 46170
rect 8484 46106 8536 46112
rect 7748 46028 7800 46034
rect 7748 45970 7800 45976
rect 7840 45960 7892 45966
rect 7840 45902 7892 45908
rect 2950 45180 3258 45189
rect 2950 45178 2956 45180
rect 3012 45178 3036 45180
rect 3092 45178 3116 45180
rect 3172 45178 3196 45180
rect 3252 45178 3258 45180
rect 3012 45126 3014 45178
rect 3194 45126 3196 45178
rect 2950 45124 2956 45126
rect 3012 45124 3036 45126
rect 3092 45124 3116 45126
rect 3172 45124 3196 45126
rect 3252 45124 3258 45126
rect 2950 45115 3258 45124
rect 2950 44092 3258 44101
rect 2950 44090 2956 44092
rect 3012 44090 3036 44092
rect 3092 44090 3116 44092
rect 3172 44090 3196 44092
rect 3252 44090 3258 44092
rect 3012 44038 3014 44090
rect 3194 44038 3196 44090
rect 2950 44036 2956 44038
rect 3012 44036 3036 44038
rect 3092 44036 3116 44038
rect 3172 44036 3196 44038
rect 3252 44036 3258 44038
rect 2950 44027 3258 44036
rect 2950 43004 3258 43013
rect 2950 43002 2956 43004
rect 3012 43002 3036 43004
rect 3092 43002 3116 43004
rect 3172 43002 3196 43004
rect 3252 43002 3258 43004
rect 3012 42950 3014 43002
rect 3194 42950 3196 43002
rect 2950 42948 2956 42950
rect 3012 42948 3036 42950
rect 3092 42948 3116 42950
rect 3172 42948 3196 42950
rect 3252 42948 3258 42950
rect 2950 42939 3258 42948
rect 2950 41916 3258 41925
rect 2950 41914 2956 41916
rect 3012 41914 3036 41916
rect 3092 41914 3116 41916
rect 3172 41914 3196 41916
rect 3252 41914 3258 41916
rect 3012 41862 3014 41914
rect 3194 41862 3196 41914
rect 2950 41860 2956 41862
rect 3012 41860 3036 41862
rect 3092 41860 3116 41862
rect 3172 41860 3196 41862
rect 3252 41860 3258 41862
rect 2950 41851 3258 41860
rect 2950 40828 3258 40837
rect 2950 40826 2956 40828
rect 3012 40826 3036 40828
rect 3092 40826 3116 40828
rect 3172 40826 3196 40828
rect 3252 40826 3258 40828
rect 3012 40774 3014 40826
rect 3194 40774 3196 40826
rect 2950 40772 2956 40774
rect 3012 40772 3036 40774
rect 3092 40772 3116 40774
rect 3172 40772 3196 40774
rect 3252 40772 3258 40774
rect 2950 40763 3258 40772
rect 2950 39740 3258 39749
rect 2950 39738 2956 39740
rect 3012 39738 3036 39740
rect 3092 39738 3116 39740
rect 3172 39738 3196 39740
rect 3252 39738 3258 39740
rect 3012 39686 3014 39738
rect 3194 39686 3196 39738
rect 2950 39684 2956 39686
rect 3012 39684 3036 39686
rect 3092 39684 3116 39686
rect 3172 39684 3196 39686
rect 3252 39684 3258 39686
rect 2950 39675 3258 39684
rect 2950 38652 3258 38661
rect 2950 38650 2956 38652
rect 3012 38650 3036 38652
rect 3092 38650 3116 38652
rect 3172 38650 3196 38652
rect 3252 38650 3258 38652
rect 3012 38598 3014 38650
rect 3194 38598 3196 38650
rect 2950 38596 2956 38598
rect 3012 38596 3036 38598
rect 3092 38596 3116 38598
rect 3172 38596 3196 38598
rect 3252 38596 3258 38598
rect 2950 38587 3258 38596
rect 7852 38010 7880 45902
rect 7950 45724 8258 45733
rect 7950 45722 7956 45724
rect 8012 45722 8036 45724
rect 8092 45722 8116 45724
rect 8172 45722 8196 45724
rect 8252 45722 8258 45724
rect 8012 45670 8014 45722
rect 8194 45670 8196 45722
rect 7950 45668 7956 45670
rect 8012 45668 8036 45670
rect 8092 45668 8116 45670
rect 8172 45668 8196 45670
rect 8252 45668 8258 45670
rect 7950 45659 8258 45668
rect 9140 44946 9168 48554
rect 9416 47802 9444 52430
rect 9600 50522 9628 54130
rect 10704 53718 10732 56200
rect 12084 56114 12112 56200
rect 12176 56114 12204 56222
rect 12084 56086 12204 56114
rect 11704 54188 11756 54194
rect 11704 54130 11756 54136
rect 10692 53712 10744 53718
rect 10692 53654 10744 53660
rect 10692 53576 10744 53582
rect 10692 53518 10744 53524
rect 10508 51400 10560 51406
rect 10508 51342 10560 51348
rect 9588 50516 9640 50522
rect 9588 50458 9640 50464
rect 9588 50312 9640 50318
rect 9588 50254 9640 50260
rect 9496 48680 9548 48686
rect 9496 48622 9548 48628
rect 9220 47796 9272 47802
rect 9220 47738 9272 47744
rect 9404 47796 9456 47802
rect 9404 47738 9456 47744
rect 9232 47054 9260 47738
rect 9508 47462 9536 48622
rect 9496 47456 9548 47462
rect 9496 47398 9548 47404
rect 9220 47048 9272 47054
rect 9220 46990 9272 46996
rect 9128 44940 9180 44946
rect 9128 44882 9180 44888
rect 7950 44636 8258 44645
rect 7950 44634 7956 44636
rect 8012 44634 8036 44636
rect 8092 44634 8116 44636
rect 8172 44634 8196 44636
rect 8252 44634 8258 44636
rect 8012 44582 8014 44634
rect 8194 44582 8196 44634
rect 7950 44580 7956 44582
rect 8012 44580 8036 44582
rect 8092 44580 8116 44582
rect 8172 44580 8196 44582
rect 8252 44580 8258 44582
rect 7950 44571 8258 44580
rect 9232 44402 9260 46990
rect 9508 45554 9536 47398
rect 9416 45526 9536 45554
rect 9416 45082 9444 45526
rect 9404 45076 9456 45082
rect 9404 45018 9456 45024
rect 9404 44940 9456 44946
rect 9404 44882 9456 44888
rect 9220 44396 9272 44402
rect 9220 44338 9272 44344
rect 9036 44328 9088 44334
rect 9036 44270 9088 44276
rect 7950 43548 8258 43557
rect 7950 43546 7956 43548
rect 8012 43546 8036 43548
rect 8092 43546 8116 43548
rect 8172 43546 8196 43548
rect 8252 43546 8258 43548
rect 8012 43494 8014 43546
rect 8194 43494 8196 43546
rect 7950 43492 7956 43494
rect 8012 43492 8036 43494
rect 8092 43492 8116 43494
rect 8172 43492 8196 43494
rect 8252 43492 8258 43494
rect 7950 43483 8258 43492
rect 8944 42696 8996 42702
rect 8944 42638 8996 42644
rect 7950 42460 8258 42469
rect 7950 42458 7956 42460
rect 8012 42458 8036 42460
rect 8092 42458 8116 42460
rect 8172 42458 8196 42460
rect 8252 42458 8258 42460
rect 8012 42406 8014 42458
rect 8194 42406 8196 42458
rect 7950 42404 7956 42406
rect 8012 42404 8036 42406
rect 8092 42404 8116 42406
rect 8172 42404 8196 42406
rect 8252 42404 8258 42406
rect 7950 42395 8258 42404
rect 7950 41372 8258 41381
rect 7950 41370 7956 41372
rect 8012 41370 8036 41372
rect 8092 41370 8116 41372
rect 8172 41370 8196 41372
rect 8252 41370 8258 41372
rect 8012 41318 8014 41370
rect 8194 41318 8196 41370
rect 7950 41316 7956 41318
rect 8012 41316 8036 41318
rect 8092 41316 8116 41318
rect 8172 41316 8196 41318
rect 8252 41316 8258 41318
rect 7950 41307 8258 41316
rect 7950 40284 8258 40293
rect 7950 40282 7956 40284
rect 8012 40282 8036 40284
rect 8092 40282 8116 40284
rect 8172 40282 8196 40284
rect 8252 40282 8258 40284
rect 8012 40230 8014 40282
rect 8194 40230 8196 40282
rect 7950 40228 7956 40230
rect 8012 40228 8036 40230
rect 8092 40228 8116 40230
rect 8172 40228 8196 40230
rect 8252 40228 8258 40230
rect 7950 40219 8258 40228
rect 7950 39196 8258 39205
rect 7950 39194 7956 39196
rect 8012 39194 8036 39196
rect 8092 39194 8116 39196
rect 8172 39194 8196 39196
rect 8252 39194 8258 39196
rect 8012 39142 8014 39194
rect 8194 39142 8196 39194
rect 7950 39140 7956 39142
rect 8012 39140 8036 39142
rect 8092 39140 8116 39142
rect 8172 39140 8196 39142
rect 8252 39140 8258 39142
rect 7950 39131 8258 39140
rect 7950 38108 8258 38117
rect 7950 38106 7956 38108
rect 8012 38106 8036 38108
rect 8092 38106 8116 38108
rect 8172 38106 8196 38108
rect 8252 38106 8258 38108
rect 8012 38054 8014 38106
rect 8194 38054 8196 38106
rect 7950 38052 7956 38054
rect 8012 38052 8036 38054
rect 8092 38052 8116 38054
rect 8172 38052 8196 38054
rect 8252 38052 8258 38054
rect 7950 38043 8258 38052
rect 7840 38004 7892 38010
rect 7840 37946 7892 37952
rect 8852 37868 8904 37874
rect 8852 37810 8904 37816
rect 2950 37564 3258 37573
rect 2950 37562 2956 37564
rect 3012 37562 3036 37564
rect 3092 37562 3116 37564
rect 3172 37562 3196 37564
rect 3252 37562 3258 37564
rect 3012 37510 3014 37562
rect 3194 37510 3196 37562
rect 2950 37508 2956 37510
rect 3012 37508 3036 37510
rect 3092 37508 3116 37510
rect 3172 37508 3196 37510
rect 3252 37508 3258 37510
rect 2950 37499 3258 37508
rect 7950 37020 8258 37029
rect 7950 37018 7956 37020
rect 8012 37018 8036 37020
rect 8092 37018 8116 37020
rect 8172 37018 8196 37020
rect 8252 37018 8258 37020
rect 8012 36966 8014 37018
rect 8194 36966 8196 37018
rect 7950 36964 7956 36966
rect 8012 36964 8036 36966
rect 8092 36964 8116 36966
rect 8172 36964 8196 36966
rect 8252 36964 8258 36966
rect 7950 36955 8258 36964
rect 2950 36476 3258 36485
rect 2950 36474 2956 36476
rect 3012 36474 3036 36476
rect 3092 36474 3116 36476
rect 3172 36474 3196 36476
rect 3252 36474 3258 36476
rect 3012 36422 3014 36474
rect 3194 36422 3196 36474
rect 2950 36420 2956 36422
rect 3012 36420 3036 36422
rect 3092 36420 3116 36422
rect 3172 36420 3196 36422
rect 3252 36420 3258 36422
rect 2950 36411 3258 36420
rect 7950 35932 8258 35941
rect 7950 35930 7956 35932
rect 8012 35930 8036 35932
rect 8092 35930 8116 35932
rect 8172 35930 8196 35932
rect 8252 35930 8258 35932
rect 8012 35878 8014 35930
rect 8194 35878 8196 35930
rect 7950 35876 7956 35878
rect 8012 35876 8036 35878
rect 8092 35876 8116 35878
rect 8172 35876 8196 35878
rect 8252 35876 8258 35878
rect 7950 35867 8258 35876
rect 2950 35388 3258 35397
rect 2950 35386 2956 35388
rect 3012 35386 3036 35388
rect 3092 35386 3116 35388
rect 3172 35386 3196 35388
rect 3252 35386 3258 35388
rect 3012 35334 3014 35386
rect 3194 35334 3196 35386
rect 2950 35332 2956 35334
rect 3012 35332 3036 35334
rect 3092 35332 3116 35334
rect 3172 35332 3196 35334
rect 3252 35332 3258 35334
rect 2950 35323 3258 35332
rect 7950 34844 8258 34853
rect 7950 34842 7956 34844
rect 8012 34842 8036 34844
rect 8092 34842 8116 34844
rect 8172 34842 8196 34844
rect 8252 34842 8258 34844
rect 8012 34790 8014 34842
rect 8194 34790 8196 34842
rect 7950 34788 7956 34790
rect 8012 34788 8036 34790
rect 8092 34788 8116 34790
rect 8172 34788 8196 34790
rect 8252 34788 8258 34790
rect 7950 34779 8258 34788
rect 2950 34300 3258 34309
rect 2950 34298 2956 34300
rect 3012 34298 3036 34300
rect 3092 34298 3116 34300
rect 3172 34298 3196 34300
rect 3252 34298 3258 34300
rect 3012 34246 3014 34298
rect 3194 34246 3196 34298
rect 2950 34244 2956 34246
rect 3012 34244 3036 34246
rect 3092 34244 3116 34246
rect 3172 34244 3196 34246
rect 3252 34244 3258 34246
rect 2950 34235 3258 34244
rect 7950 33756 8258 33765
rect 7950 33754 7956 33756
rect 8012 33754 8036 33756
rect 8092 33754 8116 33756
rect 8172 33754 8196 33756
rect 8252 33754 8258 33756
rect 8012 33702 8014 33754
rect 8194 33702 8196 33754
rect 7950 33700 7956 33702
rect 8012 33700 8036 33702
rect 8092 33700 8116 33702
rect 8172 33700 8196 33702
rect 8252 33700 8258 33702
rect 7950 33691 8258 33700
rect 2950 33212 3258 33221
rect 2950 33210 2956 33212
rect 3012 33210 3036 33212
rect 3092 33210 3116 33212
rect 3172 33210 3196 33212
rect 3252 33210 3258 33212
rect 3012 33158 3014 33210
rect 3194 33158 3196 33210
rect 2950 33156 2956 33158
rect 3012 33156 3036 33158
rect 3092 33156 3116 33158
rect 3172 33156 3196 33158
rect 3252 33156 3258 33158
rect 2950 33147 3258 33156
rect 7950 32668 8258 32677
rect 7950 32666 7956 32668
rect 8012 32666 8036 32668
rect 8092 32666 8116 32668
rect 8172 32666 8196 32668
rect 8252 32666 8258 32668
rect 8012 32614 8014 32666
rect 8194 32614 8196 32666
rect 7950 32612 7956 32614
rect 8012 32612 8036 32614
rect 8092 32612 8116 32614
rect 8172 32612 8196 32614
rect 8252 32612 8258 32614
rect 7950 32603 8258 32612
rect 2950 32124 3258 32133
rect 2950 32122 2956 32124
rect 3012 32122 3036 32124
rect 3092 32122 3116 32124
rect 3172 32122 3196 32124
rect 3252 32122 3258 32124
rect 3012 32070 3014 32122
rect 3194 32070 3196 32122
rect 2950 32068 2956 32070
rect 3012 32068 3036 32070
rect 3092 32068 3116 32070
rect 3172 32068 3196 32070
rect 3252 32068 3258 32070
rect 2950 32059 3258 32068
rect 7950 31580 8258 31589
rect 7950 31578 7956 31580
rect 8012 31578 8036 31580
rect 8092 31578 8116 31580
rect 8172 31578 8196 31580
rect 8252 31578 8258 31580
rect 8012 31526 8014 31578
rect 8194 31526 8196 31578
rect 7950 31524 7956 31526
rect 8012 31524 8036 31526
rect 8092 31524 8116 31526
rect 8172 31524 8196 31526
rect 8252 31524 8258 31526
rect 7950 31515 8258 31524
rect 2950 31036 3258 31045
rect 2950 31034 2956 31036
rect 3012 31034 3036 31036
rect 3092 31034 3116 31036
rect 3172 31034 3196 31036
rect 3252 31034 3258 31036
rect 3012 30982 3014 31034
rect 3194 30982 3196 31034
rect 2950 30980 2956 30982
rect 3012 30980 3036 30982
rect 3092 30980 3116 30982
rect 3172 30980 3196 30982
rect 3252 30980 3258 30982
rect 2950 30971 3258 30980
rect 8760 30728 8812 30734
rect 8760 30670 8812 30676
rect 7950 30492 8258 30501
rect 7950 30490 7956 30492
rect 8012 30490 8036 30492
rect 8092 30490 8116 30492
rect 8172 30490 8196 30492
rect 8252 30490 8258 30492
rect 8012 30438 8014 30490
rect 8194 30438 8196 30490
rect 7950 30436 7956 30438
rect 8012 30436 8036 30438
rect 8092 30436 8116 30438
rect 8172 30436 8196 30438
rect 8252 30436 8258 30438
rect 7950 30427 8258 30436
rect 8484 30252 8536 30258
rect 8484 30194 8536 30200
rect 2950 29948 3258 29957
rect 2950 29946 2956 29948
rect 3012 29946 3036 29948
rect 3092 29946 3116 29948
rect 3172 29946 3196 29948
rect 3252 29946 3258 29948
rect 3012 29894 3014 29946
rect 3194 29894 3196 29946
rect 2950 29892 2956 29894
rect 3012 29892 3036 29894
rect 3092 29892 3116 29894
rect 3172 29892 3196 29894
rect 3252 29892 3258 29894
rect 2950 29883 3258 29892
rect 7950 29404 8258 29413
rect 7950 29402 7956 29404
rect 8012 29402 8036 29404
rect 8092 29402 8116 29404
rect 8172 29402 8196 29404
rect 8252 29402 8258 29404
rect 8012 29350 8014 29402
rect 8194 29350 8196 29402
rect 7950 29348 7956 29350
rect 8012 29348 8036 29350
rect 8092 29348 8116 29350
rect 8172 29348 8196 29350
rect 8252 29348 8258 29350
rect 7950 29339 8258 29348
rect 2950 28860 3258 28869
rect 2950 28858 2956 28860
rect 3012 28858 3036 28860
rect 3092 28858 3116 28860
rect 3172 28858 3196 28860
rect 3252 28858 3258 28860
rect 3012 28806 3014 28858
rect 3194 28806 3196 28858
rect 2950 28804 2956 28806
rect 3012 28804 3036 28806
rect 3092 28804 3116 28806
rect 3172 28804 3196 28806
rect 3252 28804 3258 28806
rect 2950 28795 3258 28804
rect 7950 28316 8258 28325
rect 7950 28314 7956 28316
rect 8012 28314 8036 28316
rect 8092 28314 8116 28316
rect 8172 28314 8196 28316
rect 8252 28314 8258 28316
rect 8012 28262 8014 28314
rect 8194 28262 8196 28314
rect 7950 28260 7956 28262
rect 8012 28260 8036 28262
rect 8092 28260 8116 28262
rect 8172 28260 8196 28262
rect 8252 28260 8258 28262
rect 7950 28251 8258 28260
rect 3424 28212 3476 28218
rect 3424 28154 3476 28160
rect 2950 27772 3258 27781
rect 2950 27770 2956 27772
rect 3012 27770 3036 27772
rect 3092 27770 3116 27772
rect 3172 27770 3196 27772
rect 3252 27770 3258 27772
rect 3012 27718 3014 27770
rect 3194 27718 3196 27770
rect 2950 27716 2956 27718
rect 3012 27716 3036 27718
rect 3092 27716 3116 27718
rect 3172 27716 3196 27718
rect 3252 27716 3258 27718
rect 2950 27707 3258 27716
rect 2950 26684 3258 26693
rect 2950 26682 2956 26684
rect 3012 26682 3036 26684
rect 3092 26682 3116 26684
rect 3172 26682 3196 26684
rect 3252 26682 3258 26684
rect 3012 26630 3014 26682
rect 3194 26630 3196 26682
rect 2950 26628 2956 26630
rect 3012 26628 3036 26630
rect 3092 26628 3116 26630
rect 3172 26628 3196 26630
rect 3252 26628 3258 26630
rect 2950 26619 3258 26628
rect 2950 25596 3258 25605
rect 2950 25594 2956 25596
rect 3012 25594 3036 25596
rect 3092 25594 3116 25596
rect 3172 25594 3196 25596
rect 3252 25594 3258 25596
rect 3012 25542 3014 25594
rect 3194 25542 3196 25594
rect 2950 25540 2956 25542
rect 3012 25540 3036 25542
rect 3092 25540 3116 25542
rect 3172 25540 3196 25542
rect 3252 25540 3258 25542
rect 2950 25531 3258 25540
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 3332 17128 3384 17134
rect 3332 17070 3384 17076
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 2228 7744 2280 7750
rect 2228 7686 2280 7692
rect 1492 4480 1544 4486
rect 1492 4422 1544 4428
rect 1504 4146 1532 4422
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 1504 800 1532 4082
rect 1872 800 1900 4082
rect 2240 4010 2268 7686
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 2228 4004 2280 4010
rect 2228 3946 2280 3952
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2884 3602 2912 3878
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 3344 3738 3372 17070
rect 3436 6497 3464 28154
rect 7950 27228 8258 27237
rect 7950 27226 7956 27228
rect 8012 27226 8036 27228
rect 8092 27226 8116 27228
rect 8172 27226 8196 27228
rect 8252 27226 8258 27228
rect 8012 27174 8014 27226
rect 8194 27174 8196 27226
rect 7950 27172 7956 27174
rect 8012 27172 8036 27174
rect 8092 27172 8116 27174
rect 8172 27172 8196 27174
rect 8252 27172 8258 27174
rect 7950 27163 8258 27172
rect 7748 26444 7800 26450
rect 7748 26386 7800 26392
rect 6920 22432 6972 22438
rect 6920 22374 6972 22380
rect 3516 21140 3568 21146
rect 3516 21082 3568 21088
rect 3528 8809 3556 21082
rect 6932 19310 6960 22374
rect 7760 22094 7788 26386
rect 7950 26140 8258 26149
rect 7950 26138 7956 26140
rect 8012 26138 8036 26140
rect 8092 26138 8116 26140
rect 8172 26138 8196 26140
rect 8252 26138 8258 26140
rect 8012 26086 8014 26138
rect 8194 26086 8196 26138
rect 7950 26084 7956 26086
rect 8012 26084 8036 26086
rect 8092 26084 8116 26086
rect 8172 26084 8196 26086
rect 8252 26084 8258 26086
rect 7950 26075 8258 26084
rect 7950 25052 8258 25061
rect 7950 25050 7956 25052
rect 8012 25050 8036 25052
rect 8092 25050 8116 25052
rect 8172 25050 8196 25052
rect 8252 25050 8258 25052
rect 8012 24998 8014 25050
rect 8194 24998 8196 25050
rect 7950 24996 7956 24998
rect 8012 24996 8036 24998
rect 8092 24996 8116 24998
rect 8172 24996 8196 24998
rect 8252 24996 8258 24998
rect 7950 24987 8258 24996
rect 7840 24200 7892 24206
rect 7840 24142 7892 24148
rect 7852 23730 7880 24142
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 7840 23724 7892 23730
rect 7840 23666 7892 23672
rect 7852 22642 7880 23666
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 7668 22066 7788 22094
rect 6552 19304 6604 19310
rect 6552 19246 6604 19252
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 6564 18748 6592 19246
rect 6644 18760 6696 18766
rect 6564 18720 6644 18748
rect 6644 18702 6696 18708
rect 6656 18222 6684 18702
rect 6644 18216 6696 18222
rect 6564 18176 6644 18204
rect 6564 16114 6592 18176
rect 6644 18158 6696 18164
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6472 13394 6500 14418
rect 6460 13388 6512 13394
rect 6460 13330 6512 13336
rect 6932 12918 6960 19246
rect 7012 18624 7064 18630
rect 7012 18566 7064 18572
rect 7024 12986 7052 18566
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7208 17338 7236 17478
rect 7196 17332 7248 17338
rect 7196 17274 7248 17280
rect 7668 17202 7696 22066
rect 7748 21344 7800 21350
rect 7852 21332 7880 22578
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 7800 21304 7880 21332
rect 8300 21344 8352 21350
rect 7748 21286 7800 21292
rect 8300 21286 8352 21292
rect 7760 20398 7788 21286
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8312 20534 8340 21286
rect 8300 20528 8352 20534
rect 8300 20470 8352 20476
rect 7748 20392 7800 20398
rect 7748 20334 7800 20340
rect 7760 19854 7788 20334
rect 8392 20052 8444 20058
rect 8392 19994 8444 20000
rect 7748 19848 7800 19854
rect 7748 19790 7800 19796
rect 8300 19780 8352 19786
rect 8300 19722 8352 19728
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 8312 18630 8340 19722
rect 8404 19446 8432 19994
rect 8392 19440 8444 19446
rect 8392 19382 8444 19388
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8404 18834 8432 19110
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 8312 18034 8340 18566
rect 8404 18222 8432 18770
rect 8392 18216 8444 18222
rect 8392 18158 8444 18164
rect 8312 18006 8432 18034
rect 7840 17740 7892 17746
rect 7840 17682 7892 17688
rect 7748 17536 7800 17542
rect 7748 17478 7800 17484
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 3514 8800 3570 8809
rect 3514 8735 3570 8744
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 3700 3596 3752 3602
rect 3700 3538 3752 3544
rect 2228 3528 2280 3534
rect 2228 3470 2280 3476
rect 2240 800 2268 3470
rect 3424 3392 3476 3398
rect 3424 3334 3476 3340
rect 3436 3058 3464 3334
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 3424 3052 3476 3058
rect 3424 2994 3476 3000
rect 2608 2310 2636 2994
rect 3436 2774 3464 2994
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 3344 2746 3464 2774
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 2596 2304 2648 2310
rect 2596 2246 2648 2252
rect 2608 800 2636 2246
rect 2976 800 3004 2382
rect 3344 800 3372 2746
rect 3712 800 3740 3538
rect 4080 800 4108 4082
rect 5170 3632 5226 3641
rect 5170 3567 5172 3576
rect 5224 3567 5226 3576
rect 5172 3538 5224 3544
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 4448 3194 4476 3470
rect 4908 3194 4936 3470
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 4448 800 4476 3130
rect 4908 2774 4936 3130
rect 5276 3058 5304 11834
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 5368 4078 5396 4490
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 6380 3670 6408 6258
rect 6932 4010 6960 12718
rect 7024 12306 7052 12786
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7104 10736 7156 10742
rect 7104 10678 7156 10684
rect 7116 9722 7144 10678
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7116 4554 7144 9658
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 6920 4004 6972 4010
rect 6920 3946 6972 3952
rect 6368 3664 6420 3670
rect 6368 3606 6420 3612
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5460 3058 5488 3538
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 7012 3528 7064 3534
rect 7012 3470 7064 3476
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 4816 2746 4936 2774
rect 4816 800 4844 2746
rect 5184 2310 5212 2926
rect 5446 2544 5502 2553
rect 5446 2479 5448 2488
rect 5500 2479 5502 2488
rect 5448 2450 5500 2456
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 5184 800 5212 2246
rect 5552 800 5580 2382
rect 5908 2372 5960 2378
rect 5908 2314 5960 2320
rect 5920 800 5948 2314
rect 6288 800 6316 3470
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6656 2310 6684 2994
rect 6644 2304 6696 2310
rect 6644 2246 6696 2252
rect 6656 800 6684 2246
rect 7024 800 7052 3470
rect 7208 2854 7236 11290
rect 7668 3738 7696 12718
rect 7760 12442 7788 17478
rect 7852 14618 7880 17682
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7852 13954 7880 14554
rect 8312 14482 8340 14758
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 8312 14074 8340 14418
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 7932 14000 7984 14006
rect 7852 13948 7932 13954
rect 7852 13942 7984 13948
rect 7852 13926 7972 13942
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 8220 12306 8248 12786
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 8312 11558 8340 14010
rect 8404 12782 8432 18006
rect 8496 17882 8524 30194
rect 8668 23180 8720 23186
rect 8668 23122 8720 23128
rect 8680 21350 8708 23122
rect 8668 21344 8720 21350
rect 8668 21286 8720 21292
rect 8772 19514 8800 30670
rect 8864 29306 8892 37810
rect 8956 30122 8984 42638
rect 9048 34202 9076 44270
rect 9416 42158 9444 44882
rect 9600 44538 9628 50254
rect 10232 49156 10284 49162
rect 10232 49098 10284 49104
rect 9956 48544 10008 48550
rect 9956 48486 10008 48492
rect 9772 46708 9824 46714
rect 9772 46650 9824 46656
rect 9680 44804 9732 44810
rect 9680 44746 9732 44752
rect 9588 44532 9640 44538
rect 9588 44474 9640 44480
rect 9692 42362 9720 44746
rect 9784 42770 9812 46650
rect 9968 44946 9996 48486
rect 9956 44940 10008 44946
rect 9956 44882 10008 44888
rect 10244 42770 10272 49098
rect 10324 47660 10376 47666
rect 10324 47602 10376 47608
rect 10336 46578 10364 47602
rect 10324 46572 10376 46578
rect 10324 46514 10376 46520
rect 10336 44402 10364 46514
rect 10416 46368 10468 46374
rect 10416 46310 10468 46316
rect 10428 44742 10456 46310
rect 10520 45558 10548 51342
rect 10704 49366 10732 53518
rect 10784 51332 10836 51338
rect 10784 51274 10836 51280
rect 10692 49360 10744 49366
rect 10692 49302 10744 49308
rect 10796 46714 10824 51274
rect 11716 49366 11744 54130
rect 12360 54126 12388 56222
rect 13450 56200 13506 57000
rect 13556 56222 13768 56250
rect 13464 56114 13492 56200
rect 13556 56114 13584 56222
rect 13464 56086 13584 56114
rect 13740 55214 13768 56222
rect 14830 56200 14886 57000
rect 16210 56200 16266 57000
rect 16316 56222 16528 56250
rect 13740 55186 13860 55214
rect 13832 54330 13860 55186
rect 13820 54324 13872 54330
rect 13820 54266 13872 54272
rect 14844 54194 14872 56200
rect 16224 56114 16252 56200
rect 16316 56114 16344 56222
rect 16224 56086 16344 56114
rect 14832 54188 14884 54194
rect 16500 54176 16528 56222
rect 17590 56200 17646 57000
rect 18970 56200 19026 57000
rect 20350 56200 20406 57000
rect 20456 56222 20668 56250
rect 17604 54194 17632 56200
rect 17950 54428 18258 54437
rect 17950 54426 17956 54428
rect 18012 54426 18036 54428
rect 18092 54426 18116 54428
rect 18172 54426 18196 54428
rect 18252 54426 18258 54428
rect 18012 54374 18014 54426
rect 18194 54374 18196 54426
rect 17950 54372 17956 54374
rect 18012 54372 18036 54374
rect 18092 54372 18116 54374
rect 18172 54372 18196 54374
rect 18252 54372 18258 54374
rect 17950 54363 18258 54372
rect 18984 54330 19012 56200
rect 20364 56114 20392 56200
rect 20456 56114 20484 56222
rect 20364 56086 20484 56114
rect 18972 54324 19024 54330
rect 18972 54266 19024 54272
rect 16580 54188 16632 54194
rect 16500 54148 16580 54176
rect 14832 54130 14884 54136
rect 16580 54130 16632 54136
rect 17592 54188 17644 54194
rect 20640 54176 20668 56222
rect 21730 56200 21786 57000
rect 23110 56200 23166 57000
rect 24490 56200 24546 57000
rect 25870 56200 25926 57000
rect 21744 54194 21772 56200
rect 23124 54194 23152 56200
rect 23386 56128 23442 56137
rect 23386 56063 23442 56072
rect 20720 54188 20772 54194
rect 20640 54148 20720 54176
rect 17592 54130 17644 54136
rect 20720 54130 20772 54136
rect 21732 54188 21784 54194
rect 21732 54130 21784 54136
rect 23112 54188 23164 54194
rect 23112 54130 23164 54136
rect 12348 54120 12400 54126
rect 12348 54062 12400 54068
rect 16672 54120 16724 54126
rect 16672 54062 16724 54068
rect 13912 54052 13964 54058
rect 13912 53994 13964 54000
rect 16120 54052 16172 54058
rect 16120 53994 16172 54000
rect 12716 53984 12768 53990
rect 12716 53926 12768 53932
rect 11704 49360 11756 49366
rect 11704 49302 11756 49308
rect 10876 49156 10928 49162
rect 10876 49098 10928 49104
rect 10784 46708 10836 46714
rect 10784 46650 10836 46656
rect 10508 45552 10560 45558
rect 10508 45494 10560 45500
rect 10416 44736 10468 44742
rect 10416 44678 10468 44684
rect 10324 44396 10376 44402
rect 10324 44338 10376 44344
rect 10520 44266 10548 45494
rect 10508 44260 10560 44266
rect 10508 44202 10560 44208
rect 10692 44192 10744 44198
rect 10692 44134 10744 44140
rect 9772 42764 9824 42770
rect 9772 42706 9824 42712
rect 10232 42764 10284 42770
rect 10232 42706 10284 42712
rect 9680 42356 9732 42362
rect 9680 42298 9732 42304
rect 10704 42158 10732 44134
rect 9404 42152 9456 42158
rect 9404 42094 9456 42100
rect 9772 42152 9824 42158
rect 9772 42094 9824 42100
rect 10692 42152 10744 42158
rect 10692 42094 10744 42100
rect 9220 41608 9272 41614
rect 9220 41550 9272 41556
rect 9036 34196 9088 34202
rect 9036 34138 9088 34144
rect 9232 30938 9260 41550
rect 9416 35630 9444 42094
rect 9784 35834 9812 42094
rect 10888 41818 10916 49098
rect 12624 48000 12676 48006
rect 12624 47942 12676 47948
rect 12532 45960 12584 45966
rect 12532 45902 12584 45908
rect 12544 45558 12572 45902
rect 12636 45558 12664 47942
rect 12532 45552 12584 45558
rect 12532 45494 12584 45500
rect 12624 45552 12676 45558
rect 12624 45494 12676 45500
rect 12728 45490 12756 53926
rect 12950 53884 13258 53893
rect 12950 53882 12956 53884
rect 13012 53882 13036 53884
rect 13092 53882 13116 53884
rect 13172 53882 13196 53884
rect 13252 53882 13258 53884
rect 13012 53830 13014 53882
rect 13194 53830 13196 53882
rect 12950 53828 12956 53830
rect 13012 53828 13036 53830
rect 13092 53828 13116 53830
rect 13172 53828 13196 53830
rect 13252 53828 13258 53830
rect 12950 53819 13258 53828
rect 12950 52796 13258 52805
rect 12950 52794 12956 52796
rect 13012 52794 13036 52796
rect 13092 52794 13116 52796
rect 13172 52794 13196 52796
rect 13252 52794 13258 52796
rect 13012 52742 13014 52794
rect 13194 52742 13196 52794
rect 12950 52740 12956 52742
rect 13012 52740 13036 52742
rect 13092 52740 13116 52742
rect 13172 52740 13196 52742
rect 13252 52740 13258 52742
rect 12950 52731 13258 52740
rect 12950 51708 13258 51717
rect 12950 51706 12956 51708
rect 13012 51706 13036 51708
rect 13092 51706 13116 51708
rect 13172 51706 13196 51708
rect 13252 51706 13258 51708
rect 13012 51654 13014 51706
rect 13194 51654 13196 51706
rect 12950 51652 12956 51654
rect 13012 51652 13036 51654
rect 13092 51652 13116 51654
rect 13172 51652 13196 51654
rect 13252 51652 13258 51654
rect 12950 51643 13258 51652
rect 12950 50620 13258 50629
rect 12950 50618 12956 50620
rect 13012 50618 13036 50620
rect 13092 50618 13116 50620
rect 13172 50618 13196 50620
rect 13252 50618 13258 50620
rect 13012 50566 13014 50618
rect 13194 50566 13196 50618
rect 12950 50564 12956 50566
rect 13012 50564 13036 50566
rect 13092 50564 13116 50566
rect 13172 50564 13196 50566
rect 13252 50564 13258 50566
rect 12950 50555 13258 50564
rect 12950 49532 13258 49541
rect 12950 49530 12956 49532
rect 13012 49530 13036 49532
rect 13092 49530 13116 49532
rect 13172 49530 13196 49532
rect 13252 49530 13258 49532
rect 13012 49478 13014 49530
rect 13194 49478 13196 49530
rect 12950 49476 12956 49478
rect 13012 49476 13036 49478
rect 13092 49476 13116 49478
rect 13172 49476 13196 49478
rect 13252 49476 13258 49478
rect 12950 49467 13258 49476
rect 12950 48444 13258 48453
rect 12950 48442 12956 48444
rect 13012 48442 13036 48444
rect 13092 48442 13116 48444
rect 13172 48442 13196 48444
rect 13252 48442 13258 48444
rect 13012 48390 13014 48442
rect 13194 48390 13196 48442
rect 12950 48388 12956 48390
rect 13012 48388 13036 48390
rect 13092 48388 13116 48390
rect 13172 48388 13196 48390
rect 13252 48388 13258 48390
rect 12950 48379 13258 48388
rect 12950 47356 13258 47365
rect 12950 47354 12956 47356
rect 13012 47354 13036 47356
rect 13092 47354 13116 47356
rect 13172 47354 13196 47356
rect 13252 47354 13258 47356
rect 13012 47302 13014 47354
rect 13194 47302 13196 47354
rect 12950 47300 12956 47302
rect 13012 47300 13036 47302
rect 13092 47300 13116 47302
rect 13172 47300 13196 47302
rect 13252 47300 13258 47302
rect 12950 47291 13258 47300
rect 13728 46980 13780 46986
rect 13728 46922 13780 46928
rect 13740 46646 13768 46922
rect 13728 46640 13780 46646
rect 13728 46582 13780 46588
rect 13924 46578 13952 53994
rect 15660 53984 15712 53990
rect 15660 53926 15712 53932
rect 15568 52964 15620 52970
rect 15568 52906 15620 52912
rect 13912 46572 13964 46578
rect 13912 46514 13964 46520
rect 15016 46368 15068 46374
rect 15016 46310 15068 46316
rect 12950 46268 13258 46277
rect 12950 46266 12956 46268
rect 13012 46266 13036 46268
rect 13092 46266 13116 46268
rect 13172 46266 13196 46268
rect 13252 46266 13258 46268
rect 13012 46214 13014 46266
rect 13194 46214 13196 46266
rect 12950 46212 12956 46214
rect 13012 46212 13036 46214
rect 13092 46212 13116 46214
rect 13172 46212 13196 46214
rect 13252 46212 13258 46214
rect 12950 46203 13258 46212
rect 15028 46034 15056 46310
rect 15016 46028 15068 46034
rect 15016 45970 15068 45976
rect 15108 45824 15160 45830
rect 15108 45766 15160 45772
rect 12716 45484 12768 45490
rect 12716 45426 12768 45432
rect 14556 45416 14608 45422
rect 14556 45358 14608 45364
rect 12950 45180 13258 45189
rect 12950 45178 12956 45180
rect 13012 45178 13036 45180
rect 13092 45178 13116 45180
rect 13172 45178 13196 45180
rect 13252 45178 13258 45180
rect 13012 45126 13014 45178
rect 13194 45126 13196 45178
rect 12950 45124 12956 45126
rect 13012 45124 13036 45126
rect 13092 45124 13116 45126
rect 13172 45124 13196 45126
rect 13252 45124 13258 45126
rect 12950 45115 13258 45124
rect 11520 44736 11572 44742
rect 11520 44678 11572 44684
rect 10968 44192 11020 44198
rect 10968 44134 11020 44140
rect 10876 41812 10928 41818
rect 10876 41754 10928 41760
rect 10980 41682 11008 44134
rect 11532 42294 11560 44678
rect 12950 44092 13258 44101
rect 12950 44090 12956 44092
rect 13012 44090 13036 44092
rect 13092 44090 13116 44092
rect 13172 44090 13196 44092
rect 13252 44090 13258 44092
rect 13012 44038 13014 44090
rect 13194 44038 13196 44090
rect 12950 44036 12956 44038
rect 13012 44036 13036 44038
rect 13092 44036 13116 44038
rect 13172 44036 13196 44038
rect 13252 44036 13258 44038
rect 12950 44027 13258 44036
rect 12950 43004 13258 43013
rect 12950 43002 12956 43004
rect 13012 43002 13036 43004
rect 13092 43002 13116 43004
rect 13172 43002 13196 43004
rect 13252 43002 13258 43004
rect 13012 42950 13014 43002
rect 13194 42950 13196 43002
rect 12950 42948 12956 42950
rect 13012 42948 13036 42950
rect 13092 42948 13116 42950
rect 13172 42948 13196 42950
rect 13252 42948 13258 42950
rect 12950 42939 13258 42948
rect 11520 42288 11572 42294
rect 11520 42230 11572 42236
rect 11532 42022 11560 42230
rect 11520 42016 11572 42022
rect 11520 41958 11572 41964
rect 10968 41676 11020 41682
rect 10968 41618 11020 41624
rect 11532 35834 11560 41958
rect 12950 41916 13258 41925
rect 12950 41914 12956 41916
rect 13012 41914 13036 41916
rect 13092 41914 13116 41916
rect 13172 41914 13196 41916
rect 13252 41914 13258 41916
rect 13012 41862 13014 41914
rect 13194 41862 13196 41914
rect 12950 41860 12956 41862
rect 13012 41860 13036 41862
rect 13092 41860 13116 41862
rect 13172 41860 13196 41862
rect 13252 41860 13258 41862
rect 12950 41851 13258 41860
rect 12950 40828 13258 40837
rect 12950 40826 12956 40828
rect 13012 40826 13036 40828
rect 13092 40826 13116 40828
rect 13172 40826 13196 40828
rect 13252 40826 13258 40828
rect 13012 40774 13014 40826
rect 13194 40774 13196 40826
rect 12950 40772 12956 40774
rect 13012 40772 13036 40774
rect 13092 40772 13116 40774
rect 13172 40772 13196 40774
rect 13252 40772 13258 40774
rect 12950 40763 13258 40772
rect 12950 39740 13258 39749
rect 12950 39738 12956 39740
rect 13012 39738 13036 39740
rect 13092 39738 13116 39740
rect 13172 39738 13196 39740
rect 13252 39738 13258 39740
rect 13012 39686 13014 39738
rect 13194 39686 13196 39738
rect 12950 39684 12956 39686
rect 13012 39684 13036 39686
rect 13092 39684 13116 39686
rect 13172 39684 13196 39686
rect 13252 39684 13258 39686
rect 12950 39675 13258 39684
rect 12950 38652 13258 38661
rect 12950 38650 12956 38652
rect 13012 38650 13036 38652
rect 13092 38650 13116 38652
rect 13172 38650 13196 38652
rect 13252 38650 13258 38652
rect 13012 38598 13014 38650
rect 13194 38598 13196 38650
rect 12950 38596 12956 38598
rect 13012 38596 13036 38598
rect 13092 38596 13116 38598
rect 13172 38596 13196 38598
rect 13252 38596 13258 38598
rect 12950 38587 13258 38596
rect 12950 37564 13258 37573
rect 12950 37562 12956 37564
rect 13012 37562 13036 37564
rect 13092 37562 13116 37564
rect 13172 37562 13196 37564
rect 13252 37562 13258 37564
rect 13012 37510 13014 37562
rect 13194 37510 13196 37562
rect 12950 37508 12956 37510
rect 13012 37508 13036 37510
rect 13092 37508 13116 37510
rect 13172 37508 13196 37510
rect 13252 37508 13258 37510
rect 12950 37499 13258 37508
rect 12950 36476 13258 36485
rect 12950 36474 12956 36476
rect 13012 36474 13036 36476
rect 13092 36474 13116 36476
rect 13172 36474 13196 36476
rect 13252 36474 13258 36476
rect 13012 36422 13014 36474
rect 13194 36422 13196 36474
rect 12950 36420 12956 36422
rect 13012 36420 13036 36422
rect 13092 36420 13116 36422
rect 13172 36420 13196 36422
rect 13252 36420 13258 36422
rect 12950 36411 13258 36420
rect 9772 35828 9824 35834
rect 9772 35770 9824 35776
rect 11520 35828 11572 35834
rect 11520 35770 11572 35776
rect 12716 35760 12768 35766
rect 12716 35702 12768 35708
rect 9404 35624 9456 35630
rect 9404 35566 9456 35572
rect 9680 35624 9732 35630
rect 9680 35566 9732 35572
rect 9416 34066 9444 35566
rect 9404 34060 9456 34066
rect 9404 34002 9456 34008
rect 9312 33992 9364 33998
rect 9312 33934 9364 33940
rect 9220 30932 9272 30938
rect 9220 30874 9272 30880
rect 8944 30116 8996 30122
rect 8944 30058 8996 30064
rect 8852 29300 8904 29306
rect 8852 29242 8904 29248
rect 9324 26234 9352 33934
rect 9692 29102 9720 35566
rect 12624 32768 12676 32774
rect 12624 32710 12676 32716
rect 12532 31952 12584 31958
rect 12532 31894 12584 31900
rect 12348 31136 12400 31142
rect 12348 31078 12400 31084
rect 12072 30184 12124 30190
rect 12072 30126 12124 30132
rect 11336 30048 11388 30054
rect 11336 29990 11388 29996
rect 11060 29572 11112 29578
rect 11060 29514 11112 29520
rect 10324 29232 10376 29238
rect 10324 29174 10376 29180
rect 10232 29164 10284 29170
rect 10232 29106 10284 29112
rect 9680 29096 9732 29102
rect 9680 29038 9732 29044
rect 9772 28416 9824 28422
rect 9772 28358 9824 28364
rect 9588 27328 9640 27334
rect 9588 27270 9640 27276
rect 9600 27062 9628 27270
rect 9588 27056 9640 27062
rect 9588 26998 9640 27004
rect 9232 26206 9352 26234
rect 9232 23322 9260 26206
rect 9312 24132 9364 24138
rect 9312 24074 9364 24080
rect 9220 23316 9272 23322
rect 9220 23258 9272 23264
rect 9324 23202 9352 24074
rect 9232 23174 9352 23202
rect 9404 23248 9456 23254
rect 9404 23190 9456 23196
rect 8944 22704 8996 22710
rect 8944 22646 8996 22652
rect 8956 22098 8984 22646
rect 8944 22092 8996 22098
rect 8944 22034 8996 22040
rect 8956 21622 8984 22034
rect 8944 21616 8996 21622
rect 8996 21564 9076 21570
rect 8944 21558 9076 21564
rect 8956 21542 9076 21558
rect 8852 21480 8904 21486
rect 8852 21422 8904 21428
rect 8944 21480 8996 21486
rect 8944 21422 8996 21428
rect 8864 20602 8892 21422
rect 8956 20806 8984 21422
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 8852 20596 8904 20602
rect 8852 20538 8904 20544
rect 8760 19508 8812 19514
rect 8760 19450 8812 19456
rect 8668 19440 8720 19446
rect 8668 19382 8720 19388
rect 8576 19236 8628 19242
rect 8576 19178 8628 19184
rect 8484 17876 8536 17882
rect 8484 17818 8536 17824
rect 8588 16250 8616 19178
rect 8680 18970 8708 19382
rect 8668 18964 8720 18970
rect 8668 18906 8720 18912
rect 8680 18766 8708 18906
rect 8864 18766 8892 20538
rect 8668 18760 8720 18766
rect 8668 18702 8720 18708
rect 8852 18760 8904 18766
rect 8852 18702 8904 18708
rect 8680 18358 8708 18702
rect 8956 18630 8984 20742
rect 9048 20534 9076 21542
rect 9036 20528 9088 20534
rect 9036 20470 9088 20476
rect 9048 20058 9076 20470
rect 9232 20346 9260 23174
rect 9312 22772 9364 22778
rect 9312 22714 9364 22720
rect 9324 20534 9352 22714
rect 9312 20528 9364 20534
rect 9312 20470 9364 20476
rect 9232 20318 9352 20346
rect 9036 20052 9088 20058
rect 9036 19994 9088 20000
rect 9036 19848 9088 19854
rect 9036 19790 9088 19796
rect 8944 18624 8996 18630
rect 8944 18566 8996 18572
rect 8668 18352 8720 18358
rect 8668 18294 8720 18300
rect 8680 16250 8708 18294
rect 8852 17604 8904 17610
rect 8852 17546 8904 17552
rect 8576 16244 8628 16250
rect 8576 16186 8628 16192
rect 8668 16244 8720 16250
rect 8668 16186 8720 16192
rect 8484 16040 8536 16046
rect 8484 15982 8536 15988
rect 8496 13530 8524 15982
rect 8588 14958 8616 16186
rect 8680 15094 8708 16186
rect 8668 15088 8720 15094
rect 8668 15030 8720 15036
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 8680 14618 8708 15030
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8680 14006 8708 14554
rect 8668 14000 8720 14006
rect 8668 13942 8720 13948
rect 8680 13530 8708 13942
rect 8864 13530 8892 17546
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 8680 13258 8708 13466
rect 8668 13252 8720 13258
rect 8668 13194 8720 13200
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8680 11762 8708 13194
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 8312 10470 8340 11494
rect 8680 11082 8708 11698
rect 8668 11076 8720 11082
rect 8668 11018 8720 11024
rect 8680 10810 8708 11018
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7656 3732 7708 3738
rect 7656 3674 7708 3680
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7392 3058 7420 3334
rect 7852 3126 7880 5306
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 7840 3120 7892 3126
rect 7840 3062 7892 3068
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 7196 2848 7248 2854
rect 7196 2790 7248 2796
rect 7392 800 7420 2994
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7760 2310 7788 2926
rect 8312 2514 8340 6054
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8300 2508 8352 2514
rect 8300 2450 8352 2456
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 7760 800 7788 2246
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 7852 762 7880 2382
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 8404 1970 8432 2246
rect 8392 1964 8444 1970
rect 8392 1906 8444 1912
rect 8036 870 8156 898
rect 8036 762 8064 870
rect 8128 800 8156 870
rect 8496 800 8524 3470
rect 8956 2922 8984 18566
rect 9048 18154 9076 19790
rect 9220 19440 9272 19446
rect 9220 19382 9272 19388
rect 9036 18148 9088 18154
rect 9036 18090 9088 18096
rect 9232 15706 9260 19382
rect 9324 17066 9352 20318
rect 9416 19786 9444 23190
rect 9496 22024 9548 22030
rect 9496 21966 9548 21972
rect 9404 19780 9456 19786
rect 9404 19722 9456 19728
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 9416 18086 9444 18702
rect 9404 18080 9456 18086
rect 9404 18022 9456 18028
rect 9404 17536 9456 17542
rect 9404 17478 9456 17484
rect 9416 17338 9444 17478
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9508 17270 9536 21966
rect 9600 21350 9628 26998
rect 9680 26784 9732 26790
rect 9680 26726 9732 26732
rect 9692 26314 9720 26726
rect 9680 26308 9732 26314
rect 9680 26250 9732 26256
rect 9680 25968 9732 25974
rect 9680 25910 9732 25916
rect 9692 23662 9720 25910
rect 9784 23866 9812 28358
rect 10140 24880 10192 24886
rect 10140 24822 10192 24828
rect 10152 24274 10180 24822
rect 10140 24268 10192 24274
rect 10140 24210 10192 24216
rect 10152 24138 10180 24210
rect 10140 24132 10192 24138
rect 10140 24074 10192 24080
rect 9772 23860 9824 23866
rect 9772 23802 9824 23808
rect 9680 23656 9732 23662
rect 9680 23598 9732 23604
rect 10048 23656 10100 23662
rect 10048 23598 10100 23604
rect 9588 21344 9640 21350
rect 9588 21286 9640 21292
rect 9588 20528 9640 20534
rect 9588 20470 9640 20476
rect 9600 19718 9628 20470
rect 9588 19712 9640 19718
rect 9588 19654 9640 19660
rect 9600 19514 9628 19654
rect 9588 19508 9640 19514
rect 9588 19450 9640 19456
rect 9692 18834 9720 23598
rect 9864 23112 9916 23118
rect 9864 23054 9916 23060
rect 9772 22976 9824 22982
rect 9772 22918 9824 22924
rect 9784 22094 9812 22918
rect 9876 22438 9904 23054
rect 9864 22432 9916 22438
rect 9864 22374 9916 22380
rect 9784 22066 9904 22094
rect 9876 20890 9904 22066
rect 9956 21548 10008 21554
rect 9956 21490 10008 21496
rect 9968 21010 9996 21490
rect 9956 21004 10008 21010
rect 9956 20946 10008 20952
rect 9876 20862 9996 20890
rect 9772 20392 9824 20398
rect 9772 20334 9824 20340
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9588 18692 9640 18698
rect 9588 18634 9640 18640
rect 9600 18290 9628 18634
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 9588 18148 9640 18154
rect 9588 18090 9640 18096
rect 9600 17678 9628 18090
rect 9784 17814 9812 20334
rect 9968 18902 9996 20862
rect 10060 18970 10088 23598
rect 10152 23526 10180 24074
rect 10140 23520 10192 23526
rect 10140 23462 10192 23468
rect 10152 22778 10180 23462
rect 10140 22772 10192 22778
rect 10140 22714 10192 22720
rect 10244 21690 10272 29106
rect 10336 23866 10364 29174
rect 10876 29096 10928 29102
rect 10876 29038 10928 29044
rect 10888 28762 10916 29038
rect 10876 28756 10928 28762
rect 10876 28698 10928 28704
rect 10784 27940 10836 27946
rect 10784 27882 10836 27888
rect 10796 27538 10824 27882
rect 10784 27532 10836 27538
rect 10784 27474 10836 27480
rect 11072 27130 11100 29514
rect 11152 29096 11204 29102
rect 11152 29038 11204 29044
rect 11060 27124 11112 27130
rect 11060 27066 11112 27072
rect 10968 26376 11020 26382
rect 10968 26318 11020 26324
rect 10876 26240 10928 26246
rect 10980 26234 11008 26318
rect 10928 26206 11008 26234
rect 10876 26182 10928 26188
rect 10888 25362 10916 26182
rect 11072 25838 11100 27066
rect 11164 26450 11192 29038
rect 11348 28490 11376 29990
rect 12084 29850 12112 30126
rect 12072 29844 12124 29850
rect 12072 29786 12124 29792
rect 11428 29708 11480 29714
rect 11428 29650 11480 29656
rect 11440 28626 11468 29650
rect 12360 29102 12388 31078
rect 12544 29306 12572 31894
rect 12636 29306 12664 32710
rect 12728 30326 12756 35702
rect 12950 35388 13258 35397
rect 12950 35386 12956 35388
rect 13012 35386 13036 35388
rect 13092 35386 13116 35388
rect 13172 35386 13196 35388
rect 13252 35386 13258 35388
rect 13012 35334 13014 35386
rect 13194 35334 13196 35386
rect 12950 35332 12956 35334
rect 13012 35332 13036 35334
rect 13092 35332 13116 35334
rect 13172 35332 13196 35334
rect 13252 35332 13258 35334
rect 12950 35323 13258 35332
rect 12950 34300 13258 34309
rect 12950 34298 12956 34300
rect 13012 34298 13036 34300
rect 13092 34298 13116 34300
rect 13172 34298 13196 34300
rect 13252 34298 13258 34300
rect 13012 34246 13014 34298
rect 13194 34246 13196 34298
rect 12950 34244 12956 34246
rect 13012 34244 13036 34246
rect 13092 34244 13116 34246
rect 13172 34244 13196 34246
rect 13252 34244 13258 34246
rect 12950 34235 13258 34244
rect 12950 33212 13258 33221
rect 12950 33210 12956 33212
rect 13012 33210 13036 33212
rect 13092 33210 13116 33212
rect 13172 33210 13196 33212
rect 13252 33210 13258 33212
rect 13012 33158 13014 33210
rect 13194 33158 13196 33210
rect 12950 33156 12956 33158
rect 13012 33156 13036 33158
rect 13092 33156 13116 33158
rect 13172 33156 13196 33158
rect 13252 33156 13258 33158
rect 12950 33147 13258 33156
rect 13360 32360 13412 32366
rect 13360 32302 13412 32308
rect 12950 32124 13258 32133
rect 12950 32122 12956 32124
rect 13012 32122 13036 32124
rect 13092 32122 13116 32124
rect 13172 32122 13196 32124
rect 13252 32122 13258 32124
rect 13012 32070 13014 32122
rect 13194 32070 13196 32122
rect 12950 32068 12956 32070
rect 13012 32068 13036 32070
rect 13092 32068 13116 32070
rect 13172 32068 13196 32070
rect 13252 32068 13258 32070
rect 12950 32059 13258 32068
rect 13372 31278 13400 32302
rect 13360 31272 13412 31278
rect 13360 31214 13412 31220
rect 12950 31036 13258 31045
rect 12950 31034 12956 31036
rect 13012 31034 13036 31036
rect 13092 31034 13116 31036
rect 13172 31034 13196 31036
rect 13252 31034 13258 31036
rect 13012 30982 13014 31034
rect 13194 30982 13196 31034
rect 12950 30980 12956 30982
rect 13012 30980 13036 30982
rect 13092 30980 13116 30982
rect 13172 30980 13196 30982
rect 13252 30980 13258 30982
rect 12950 30971 13258 30980
rect 13372 30394 13400 31214
rect 14096 30728 14148 30734
rect 14096 30670 14148 30676
rect 13360 30388 13412 30394
rect 13360 30330 13412 30336
rect 14108 30326 14136 30670
rect 14568 30326 14596 45358
rect 15120 44810 15148 45766
rect 15580 45554 15608 52906
rect 15672 46102 15700 53926
rect 16028 50516 16080 50522
rect 16028 50458 16080 50464
rect 15752 46504 15804 46510
rect 15752 46446 15804 46452
rect 15660 46096 15712 46102
rect 15660 46038 15712 46044
rect 15580 45526 15700 45554
rect 15108 44804 15160 44810
rect 15108 44746 15160 44752
rect 15384 33924 15436 33930
rect 15384 33866 15436 33872
rect 15396 32502 15424 33866
rect 15384 32496 15436 32502
rect 15384 32438 15436 32444
rect 14924 31408 14976 31414
rect 14924 31350 14976 31356
rect 12716 30320 12768 30326
rect 12716 30262 12768 30268
rect 14096 30320 14148 30326
rect 14096 30262 14148 30268
rect 14556 30320 14608 30326
rect 14556 30262 14608 30268
rect 12728 29578 12756 30262
rect 13360 30184 13412 30190
rect 13360 30126 13412 30132
rect 12950 29948 13258 29957
rect 12950 29946 12956 29948
rect 13012 29946 13036 29948
rect 13092 29946 13116 29948
rect 13172 29946 13196 29948
rect 13252 29946 13258 29948
rect 13012 29894 13014 29946
rect 13194 29894 13196 29946
rect 12950 29892 12956 29894
rect 13012 29892 13036 29894
rect 13092 29892 13116 29894
rect 13172 29892 13196 29894
rect 13252 29892 13258 29894
rect 12950 29883 13258 29892
rect 13372 29714 13400 30126
rect 13636 30048 13688 30054
rect 13636 29990 13688 29996
rect 13360 29708 13412 29714
rect 13360 29650 13412 29656
rect 12716 29572 12768 29578
rect 12716 29514 12768 29520
rect 12532 29300 12584 29306
rect 12532 29242 12584 29248
rect 12624 29300 12676 29306
rect 12624 29242 12676 29248
rect 13372 29170 13400 29650
rect 13452 29300 13504 29306
rect 13452 29242 13504 29248
rect 13360 29164 13412 29170
rect 13360 29106 13412 29112
rect 12348 29096 12400 29102
rect 12348 29038 12400 29044
rect 12256 29028 12308 29034
rect 12256 28970 12308 28976
rect 11428 28620 11480 28626
rect 11428 28562 11480 28568
rect 11336 28484 11388 28490
rect 11336 28426 11388 28432
rect 11244 28416 11296 28422
rect 11244 28358 11296 28364
rect 11256 28150 11284 28358
rect 11244 28144 11296 28150
rect 11244 28086 11296 28092
rect 11244 27056 11296 27062
rect 11244 26998 11296 27004
rect 11256 26518 11284 26998
rect 11244 26512 11296 26518
rect 11244 26454 11296 26460
rect 11152 26444 11204 26450
rect 11152 26386 11204 26392
rect 11256 26314 11284 26454
rect 11244 26308 11296 26314
rect 11244 26250 11296 26256
rect 11060 25832 11112 25838
rect 11060 25774 11112 25780
rect 10876 25356 10928 25362
rect 10876 25298 10928 25304
rect 11244 24880 11296 24886
rect 11244 24822 11296 24828
rect 11152 24744 11204 24750
rect 11152 24686 11204 24692
rect 10876 24676 10928 24682
rect 10876 24618 10928 24624
rect 10888 24410 10916 24618
rect 11060 24608 11112 24614
rect 11060 24550 11112 24556
rect 10876 24404 10928 24410
rect 10876 24346 10928 24352
rect 10324 23860 10376 23866
rect 10324 23802 10376 23808
rect 10416 23044 10468 23050
rect 10416 22986 10468 22992
rect 10324 21888 10376 21894
rect 10324 21830 10376 21836
rect 10232 21684 10284 21690
rect 10232 21626 10284 21632
rect 10232 20392 10284 20398
rect 10232 20334 10284 20340
rect 10140 19372 10192 19378
rect 10140 19314 10192 19320
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 9956 18896 10008 18902
rect 9956 18838 10008 18844
rect 10048 18420 10100 18426
rect 10048 18362 10100 18368
rect 9772 17808 9824 17814
rect 9772 17750 9824 17756
rect 9588 17672 9640 17678
rect 9588 17614 9640 17620
rect 9600 17270 9628 17614
rect 9496 17264 9548 17270
rect 9496 17206 9548 17212
rect 9588 17264 9640 17270
rect 9588 17206 9640 17212
rect 9784 17134 9812 17750
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9312 17060 9364 17066
rect 9312 17002 9364 17008
rect 9220 15700 9272 15706
rect 9220 15642 9272 15648
rect 9220 15428 9272 15434
rect 9220 15370 9272 15376
rect 9232 12986 9260 15370
rect 9312 14952 9364 14958
rect 9312 14894 9364 14900
rect 9324 14618 9352 14894
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9140 10470 9168 11086
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 9324 9994 9352 14554
rect 9404 14340 9456 14346
rect 9404 14282 9456 14288
rect 9416 13462 9444 14282
rect 9404 13456 9456 13462
rect 9404 13398 9456 13404
rect 9508 13274 9536 17070
rect 10060 16658 10088 18362
rect 10048 16652 10100 16658
rect 10048 16594 10100 16600
rect 9864 16448 9916 16454
rect 9864 16390 9916 16396
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9600 15570 9628 15982
rect 9588 15564 9640 15570
rect 9588 15506 9640 15512
rect 9600 15026 9628 15506
rect 9588 15020 9640 15026
rect 9588 14962 9640 14968
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9588 14408 9640 14414
rect 9588 14350 9640 14356
rect 9600 14074 9628 14350
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 9600 13938 9628 14010
rect 9784 14006 9812 14418
rect 9772 14000 9824 14006
rect 9772 13942 9824 13948
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9416 13246 9536 13274
rect 9416 12986 9444 13246
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9312 9988 9364 9994
rect 9312 9930 9364 9936
rect 9416 4162 9444 12922
rect 9600 12306 9628 13398
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9692 13274 9720 13330
rect 9692 13246 9812 13274
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 9600 11898 9628 12242
rect 9692 11898 9720 13126
rect 9784 12782 9812 13246
rect 9772 12776 9824 12782
rect 9772 12718 9824 12724
rect 9876 12628 9904 16390
rect 10048 15360 10100 15366
rect 10048 15302 10100 15308
rect 10060 12986 10088 15302
rect 10152 15162 10180 19314
rect 10244 16454 10272 20334
rect 10336 16522 10364 21830
rect 10428 20602 10456 22986
rect 10508 22976 10560 22982
rect 10508 22918 10560 22924
rect 10416 20596 10468 20602
rect 10416 20538 10468 20544
rect 10520 20210 10548 22918
rect 10888 22574 10916 24346
rect 11072 24274 11100 24550
rect 11060 24268 11112 24274
rect 11060 24210 11112 24216
rect 11164 24154 11192 24686
rect 11072 24126 11192 24154
rect 11072 24070 11100 24126
rect 11060 24064 11112 24070
rect 11060 24006 11112 24012
rect 10968 23656 11020 23662
rect 10968 23598 11020 23604
rect 10876 22568 10928 22574
rect 10876 22510 10928 22516
rect 10692 21888 10744 21894
rect 10692 21830 10744 21836
rect 10704 21622 10732 21830
rect 10692 21616 10744 21622
rect 10692 21558 10744 21564
rect 10980 21486 11008 23598
rect 11072 22234 11100 24006
rect 11060 22228 11112 22234
rect 11060 22170 11112 22176
rect 11256 22094 11284 24822
rect 11348 22098 11376 28426
rect 11440 27674 11468 28562
rect 11704 28008 11756 28014
rect 11704 27950 11756 27956
rect 11980 28008 12032 28014
rect 11980 27950 12032 27956
rect 11716 27826 11744 27950
rect 11716 27798 11836 27826
rect 11808 27674 11836 27798
rect 11428 27668 11480 27674
rect 11428 27610 11480 27616
rect 11796 27668 11848 27674
rect 11796 27610 11848 27616
rect 11992 26586 12020 27950
rect 12072 26784 12124 26790
rect 12072 26726 12124 26732
rect 11980 26580 12032 26586
rect 11980 26522 12032 26528
rect 11796 26308 11848 26314
rect 11796 26250 11848 26256
rect 11704 25492 11756 25498
rect 11704 25434 11756 25440
rect 11716 23186 11744 25434
rect 11704 23180 11756 23186
rect 11704 23122 11756 23128
rect 11808 23050 11836 26250
rect 12084 26234 12112 26726
rect 11992 26206 12112 26234
rect 11992 24138 12020 26206
rect 12268 24818 12296 28970
rect 12950 28860 13258 28869
rect 12950 28858 12956 28860
rect 13012 28858 13036 28860
rect 13092 28858 13116 28860
rect 13172 28858 13196 28860
rect 13252 28858 13258 28860
rect 13012 28806 13014 28858
rect 13194 28806 13196 28858
rect 12950 28804 12956 28806
rect 13012 28804 13036 28806
rect 13092 28804 13116 28806
rect 13172 28804 13196 28806
rect 13252 28804 13258 28806
rect 12950 28795 13258 28804
rect 12624 28416 12676 28422
rect 12624 28358 12676 28364
rect 12636 27606 12664 28358
rect 12950 27772 13258 27781
rect 12950 27770 12956 27772
rect 13012 27770 13036 27772
rect 13092 27770 13116 27772
rect 13172 27770 13196 27772
rect 13252 27770 13258 27772
rect 13012 27718 13014 27770
rect 13194 27718 13196 27770
rect 12950 27716 12956 27718
rect 13012 27716 13036 27718
rect 13092 27716 13116 27718
rect 13172 27716 13196 27718
rect 13252 27716 13258 27718
rect 12950 27707 13258 27716
rect 12440 27600 12492 27606
rect 12440 27542 12492 27548
rect 12624 27600 12676 27606
rect 12624 27542 12676 27548
rect 13084 27600 13136 27606
rect 13084 27542 13136 27548
rect 12452 27130 12480 27542
rect 12624 27328 12676 27334
rect 12624 27270 12676 27276
rect 12440 27124 12492 27130
rect 12440 27066 12492 27072
rect 12348 26580 12400 26586
rect 12348 26522 12400 26528
rect 12256 24812 12308 24818
rect 12256 24754 12308 24760
rect 12360 24750 12388 26522
rect 12636 26042 12664 27270
rect 13096 26994 13124 27542
rect 13464 27062 13492 29242
rect 13648 29102 13676 29990
rect 13728 29572 13780 29578
rect 13728 29514 13780 29520
rect 13636 29096 13688 29102
rect 13636 29038 13688 29044
rect 13740 28762 13768 29514
rect 14936 29238 14964 31350
rect 15396 30938 15424 32438
rect 15384 30932 15436 30938
rect 15384 30874 15436 30880
rect 15396 30734 15424 30874
rect 15384 30728 15436 30734
rect 15384 30670 15436 30676
rect 15108 30660 15160 30666
rect 15108 30602 15160 30608
rect 14924 29232 14976 29238
rect 14924 29174 14976 29180
rect 14016 29022 14228 29050
rect 13728 28756 13780 28762
rect 13728 28698 13780 28704
rect 13740 28490 13768 28698
rect 13728 28484 13780 28490
rect 13728 28426 13780 28432
rect 13740 28150 13768 28426
rect 13728 28144 13780 28150
rect 13728 28086 13780 28092
rect 13820 27872 13872 27878
rect 13820 27814 13872 27820
rect 13832 27402 13860 27814
rect 13820 27396 13872 27402
rect 13820 27338 13872 27344
rect 13728 27328 13780 27334
rect 13728 27270 13780 27276
rect 13544 27124 13596 27130
rect 13544 27066 13596 27072
rect 13452 27056 13504 27062
rect 13452 26998 13504 27004
rect 12716 26988 12768 26994
rect 12716 26930 12768 26936
rect 13084 26988 13136 26994
rect 13084 26930 13136 26936
rect 12728 26382 12756 26930
rect 12950 26684 13258 26693
rect 12950 26682 12956 26684
rect 13012 26682 13036 26684
rect 13092 26682 13116 26684
rect 13172 26682 13196 26684
rect 13252 26682 13258 26684
rect 13012 26630 13014 26682
rect 13194 26630 13196 26682
rect 12950 26628 12956 26630
rect 13012 26628 13036 26630
rect 13092 26628 13116 26630
rect 13172 26628 13196 26630
rect 13252 26628 13258 26630
rect 12950 26619 13258 26628
rect 13556 26586 13584 27066
rect 13544 26580 13596 26586
rect 13544 26522 13596 26528
rect 12716 26376 12768 26382
rect 12716 26318 12768 26324
rect 12624 26036 12676 26042
rect 12624 25978 12676 25984
rect 12532 25900 12584 25906
rect 12532 25842 12584 25848
rect 12348 24744 12400 24750
rect 12348 24686 12400 24692
rect 12348 24268 12400 24274
rect 12348 24210 12400 24216
rect 11980 24132 12032 24138
rect 11980 24074 12032 24080
rect 11796 23044 11848 23050
rect 11796 22986 11848 22992
rect 11164 22066 11284 22094
rect 11336 22092 11388 22098
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 11072 21690 11100 21830
rect 11060 21684 11112 21690
rect 11060 21626 11112 21632
rect 10876 21480 10928 21486
rect 10876 21422 10928 21428
rect 10968 21480 11020 21486
rect 10968 21422 11020 21428
rect 10888 21332 10916 21422
rect 10888 21304 11100 21332
rect 10692 20936 10744 20942
rect 10692 20878 10744 20884
rect 10428 20182 10548 20210
rect 10428 18426 10456 20182
rect 10704 19922 10732 20878
rect 10876 20868 10928 20874
rect 10876 20810 10928 20816
rect 10692 19916 10744 19922
rect 10692 19858 10744 19864
rect 10888 19718 10916 20810
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 10888 18834 10916 19654
rect 10600 18828 10652 18834
rect 10600 18770 10652 18776
rect 10876 18828 10928 18834
rect 10876 18770 10928 18776
rect 10612 18698 10640 18770
rect 10600 18692 10652 18698
rect 10600 18634 10652 18640
rect 10508 18624 10560 18630
rect 10508 18566 10560 18572
rect 10520 18426 10548 18566
rect 10416 18420 10468 18426
rect 10416 18362 10468 18368
rect 10508 18420 10560 18426
rect 10508 18362 10560 18368
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10324 16516 10376 16522
rect 10324 16458 10376 16464
rect 10232 16448 10284 16454
rect 10232 16390 10284 16396
rect 10428 15706 10456 16526
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10428 15162 10456 15642
rect 10140 15156 10192 15162
rect 10140 15098 10192 15104
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 10888 14346 10916 15098
rect 10876 14340 10928 14346
rect 10876 14282 10928 14288
rect 10888 14090 10916 14282
rect 10980 14278 11008 16594
rect 11072 16250 11100 21304
rect 11164 16998 11192 22066
rect 11336 22034 11388 22040
rect 11520 21548 11572 21554
rect 11520 21490 11572 21496
rect 11244 19780 11296 19786
rect 11244 19722 11296 19728
rect 11256 19174 11284 19722
rect 11428 19304 11480 19310
rect 11428 19246 11480 19252
rect 11244 19168 11296 19174
rect 11244 19110 11296 19116
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 10888 14062 11192 14090
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11072 12986 11100 13806
rect 11164 13734 11192 14062
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 11164 13258 11192 13670
rect 11152 13252 11204 13258
rect 11152 13194 11204 13200
rect 11256 13138 11284 19110
rect 11336 18624 11388 18630
rect 11336 18566 11388 18572
rect 11164 13110 11284 13138
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 9956 12776 10008 12782
rect 9956 12718 10008 12724
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 9784 12600 9904 12628
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9600 10130 9628 10406
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9600 7478 9628 10066
rect 9692 8906 9720 10950
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 9600 5710 9628 7414
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9600 4690 9628 5646
rect 9588 4684 9640 4690
rect 9588 4626 9640 4632
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9324 4134 9444 4162
rect 8944 2916 8996 2922
rect 8944 2858 8996 2864
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 9048 2446 9076 2790
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 8852 2372 8904 2378
rect 8852 2314 8904 2320
rect 8864 800 8892 2314
rect 9232 800 9260 4082
rect 9324 3466 9352 4134
rect 9404 4004 9456 4010
rect 9404 3946 9456 3952
rect 9416 3670 9444 3946
rect 9404 3664 9456 3670
rect 9404 3606 9456 3612
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9312 3460 9364 3466
rect 9312 3402 9364 3408
rect 9600 800 9628 3470
rect 9784 2774 9812 12600
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 9876 10742 9904 11018
rect 9968 10810 9996 12718
rect 10980 12306 11008 12718
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10508 11620 10560 11626
rect 10508 11562 10560 11568
rect 10520 11354 10548 11562
rect 10612 11354 10640 12038
rect 11164 11898 11192 13110
rect 11348 12714 11376 18566
rect 11440 18358 11468 19246
rect 11428 18352 11480 18358
rect 11428 18294 11480 18300
rect 11440 17610 11468 18294
rect 11428 17604 11480 17610
rect 11428 17546 11480 17552
rect 11440 17270 11468 17546
rect 11428 17264 11480 17270
rect 11428 17206 11480 17212
rect 11440 16658 11468 17206
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 11532 15706 11560 21490
rect 11992 19922 12020 24074
rect 12164 22976 12216 22982
rect 12164 22918 12216 22924
rect 12072 22432 12124 22438
rect 12072 22374 12124 22380
rect 12084 22166 12112 22374
rect 12072 22160 12124 22166
rect 12072 22102 12124 22108
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 11704 19712 11756 19718
rect 11704 19654 11756 19660
rect 11716 19514 11744 19654
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 11796 19508 11848 19514
rect 11796 19450 11848 19456
rect 11704 18692 11756 18698
rect 11704 18634 11756 18640
rect 11612 18352 11664 18358
rect 11612 18294 11664 18300
rect 11624 17338 11652 18294
rect 11716 17746 11744 18634
rect 11808 18154 11836 19450
rect 12176 18766 12204 22918
rect 12360 22642 12388 24210
rect 12440 23520 12492 23526
rect 12440 23462 12492 23468
rect 12348 22636 12400 22642
rect 12348 22578 12400 22584
rect 12360 21486 12388 22578
rect 12452 22098 12480 23462
rect 12440 22092 12492 22098
rect 12440 22034 12492 22040
rect 12348 21480 12400 21486
rect 12348 21422 12400 21428
rect 12544 21350 12572 25842
rect 12624 25152 12676 25158
rect 12624 25094 12676 25100
rect 12636 24070 12664 25094
rect 12728 24818 12756 26318
rect 12950 25596 13258 25605
rect 12950 25594 12956 25596
rect 13012 25594 13036 25596
rect 13092 25594 13116 25596
rect 13172 25594 13196 25596
rect 13252 25594 13258 25596
rect 13012 25542 13014 25594
rect 13194 25542 13196 25594
rect 12950 25540 12956 25542
rect 13012 25540 13036 25542
rect 13092 25540 13116 25542
rect 13172 25540 13196 25542
rect 13252 25540 13258 25542
rect 12950 25531 13258 25540
rect 13556 25430 13584 26522
rect 13636 26512 13688 26518
rect 13636 26454 13688 26460
rect 12992 25424 13044 25430
rect 12992 25366 13044 25372
rect 13544 25424 13596 25430
rect 13544 25366 13596 25372
rect 13004 25226 13032 25366
rect 13360 25288 13412 25294
rect 13360 25230 13412 25236
rect 12992 25220 13044 25226
rect 12992 25162 13044 25168
rect 12716 24812 12768 24818
rect 12716 24754 12768 24760
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12624 24064 12676 24070
rect 12624 24006 12676 24012
rect 12900 24064 12952 24070
rect 12900 24006 12952 24012
rect 12912 23594 12940 24006
rect 12900 23588 12952 23594
rect 12900 23530 12952 23536
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 12624 23248 12676 23254
rect 12624 23190 12676 23196
rect 12532 21344 12584 21350
rect 12532 21286 12584 21292
rect 12636 20602 12664 23190
rect 13372 22574 13400 25230
rect 13556 24886 13584 25366
rect 13544 24880 13596 24886
rect 13544 24822 13596 24828
rect 13556 24342 13584 24822
rect 13544 24336 13596 24342
rect 13544 24278 13596 24284
rect 13648 23798 13676 26454
rect 13740 23798 13768 27270
rect 13820 26036 13872 26042
rect 13820 25978 13872 25984
rect 13832 23866 13860 25978
rect 14016 25838 14044 29022
rect 14200 28966 14228 29022
rect 14936 28994 14964 29174
rect 14936 28966 15056 28994
rect 14096 28960 14148 28966
rect 14096 28902 14148 28908
rect 14188 28960 14240 28966
rect 14188 28902 14240 28908
rect 14108 28626 14136 28902
rect 15028 28762 15056 28966
rect 15016 28756 15068 28762
rect 15016 28698 15068 28704
rect 14096 28620 14148 28626
rect 14096 28562 14148 28568
rect 14108 25838 14136 28562
rect 15120 28558 15148 30602
rect 15568 29572 15620 29578
rect 15568 29514 15620 29520
rect 15200 29504 15252 29510
rect 15200 29446 15252 29452
rect 15212 29306 15240 29446
rect 15200 29300 15252 29306
rect 15200 29242 15252 29248
rect 15384 28620 15436 28626
rect 15384 28562 15436 28568
rect 15108 28552 15160 28558
rect 15108 28494 15160 28500
rect 14832 28416 14884 28422
rect 14832 28358 14884 28364
rect 14844 27470 14872 28358
rect 15120 27674 15148 28494
rect 15396 27946 15424 28562
rect 15384 27940 15436 27946
rect 15384 27882 15436 27888
rect 15108 27668 15160 27674
rect 15108 27610 15160 27616
rect 15108 27532 15160 27538
rect 15108 27474 15160 27480
rect 14832 27464 14884 27470
rect 14832 27406 14884 27412
rect 14740 26988 14792 26994
rect 14740 26930 14792 26936
rect 14752 26450 14780 26930
rect 14924 26784 14976 26790
rect 14924 26726 14976 26732
rect 14464 26444 14516 26450
rect 14464 26386 14516 26392
rect 14740 26444 14792 26450
rect 14740 26386 14792 26392
rect 14832 26444 14884 26450
rect 14832 26386 14884 26392
rect 14188 25900 14240 25906
rect 14188 25842 14240 25848
rect 14004 25832 14056 25838
rect 14004 25774 14056 25780
rect 14096 25832 14148 25838
rect 14096 25774 14148 25780
rect 13912 24744 13964 24750
rect 13912 24686 13964 24692
rect 13924 24070 13952 24686
rect 13912 24064 13964 24070
rect 13912 24006 13964 24012
rect 13820 23860 13872 23866
rect 13820 23802 13872 23808
rect 13636 23792 13688 23798
rect 13636 23734 13688 23740
rect 13728 23792 13780 23798
rect 13728 23734 13780 23740
rect 13924 23662 13952 24006
rect 14004 23724 14056 23730
rect 14004 23666 14056 23672
rect 13912 23656 13964 23662
rect 13912 23598 13964 23604
rect 13636 23180 13688 23186
rect 13636 23122 13688 23128
rect 13360 22568 13412 22574
rect 13360 22510 13412 22516
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 12716 21480 12768 21486
rect 12716 21422 12768 21428
rect 12624 20596 12676 20602
rect 12624 20538 12676 20544
rect 12728 20398 12756 21422
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 13372 21078 13400 22510
rect 13648 22094 13676 23122
rect 13556 22066 13676 22094
rect 13360 21072 13412 21078
rect 13360 21014 13412 21020
rect 12716 20392 12768 20398
rect 12716 20334 12768 20340
rect 12728 19854 12756 20334
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 12716 19848 12768 19854
rect 12716 19790 12768 19796
rect 12728 19666 12756 19790
rect 12728 19638 12848 19666
rect 12820 19174 12848 19638
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12440 18692 12492 18698
rect 12440 18634 12492 18640
rect 12452 18358 12480 18634
rect 12440 18352 12492 18358
rect 12440 18294 12492 18300
rect 11796 18148 11848 18154
rect 11796 18090 11848 18096
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11612 17332 11664 17338
rect 11612 17274 11664 17280
rect 11520 15700 11572 15706
rect 11520 15642 11572 15648
rect 11520 15088 11572 15094
rect 11520 15030 11572 15036
rect 11428 15020 11480 15026
rect 11428 14962 11480 14968
rect 11336 12708 11388 12714
rect 11336 12650 11388 12656
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 10508 11348 10560 11354
rect 10508 11290 10560 11296
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 11072 11082 11100 11630
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 10876 11008 10928 11014
rect 10876 10950 10928 10956
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 9864 10736 9916 10742
rect 9864 10678 9916 10684
rect 9876 9994 9904 10678
rect 10888 10674 10916 10950
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 11072 10266 11100 11018
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 9864 9988 9916 9994
rect 9864 9930 9916 9936
rect 9876 9654 9904 9930
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 11152 9648 11204 9654
rect 11152 9590 11204 9596
rect 9876 8906 9904 9590
rect 11164 9382 11192 9590
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 11164 9178 11192 9318
rect 11152 9172 11204 9178
rect 11152 9114 11204 9120
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 9692 2746 9812 2774
rect 9692 2582 9720 2746
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 9956 2372 10008 2378
rect 9956 2314 10008 2320
rect 9968 800 9996 2314
rect 10336 800 10364 2994
rect 10428 2990 10456 3334
rect 10416 2984 10468 2990
rect 10416 2926 10468 2932
rect 10520 2854 10548 8298
rect 10980 7342 11008 8774
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10796 5778 10824 7142
rect 10980 6254 11008 7278
rect 11072 6866 11100 8978
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11164 8090 11192 8230
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 11152 7744 11204 7750
rect 11152 7686 11204 7692
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 10876 6248 10928 6254
rect 10874 6216 10876 6225
rect 10968 6248 11020 6254
rect 10928 6216 10930 6225
rect 10968 6190 11020 6196
rect 10874 6151 10930 6160
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 11072 5166 11100 6802
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 11164 4570 11192 7686
rect 11256 5370 11284 12582
rect 11440 12442 11468 14962
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11532 10266 11560 15030
rect 11624 14074 11652 17274
rect 11716 16114 11744 17682
rect 11888 17264 11940 17270
rect 11888 17206 11940 17212
rect 11900 16998 11928 17206
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 12544 16674 12572 18702
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12452 16646 12572 16674
rect 12256 16448 12308 16454
rect 12256 16390 12308 16396
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 12164 16108 12216 16114
rect 12164 16050 12216 16056
rect 11704 15972 11756 15978
rect 11704 15914 11756 15920
rect 11716 14482 11744 15914
rect 12176 15570 12204 16050
rect 12268 15910 12296 16390
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 12164 15564 12216 15570
rect 12164 15506 12216 15512
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 11888 14952 11940 14958
rect 11888 14894 11940 14900
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11716 13954 11744 14418
rect 11624 13926 11744 13954
rect 11624 11558 11652 13926
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11716 9586 11744 13330
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11808 12646 11836 12786
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11794 11928 11850 11937
rect 11794 11863 11850 11872
rect 11808 11830 11836 11863
rect 11796 11824 11848 11830
rect 11796 11766 11848 11772
rect 11900 11626 11928 14894
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11888 11620 11940 11626
rect 11888 11562 11940 11568
rect 11886 11248 11942 11257
rect 11886 11183 11888 11192
rect 11940 11183 11942 11192
rect 11888 11154 11940 11160
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11716 9042 11744 9522
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11520 7472 11572 7478
rect 11520 7414 11572 7420
rect 11428 7336 11480 7342
rect 11428 7278 11480 7284
rect 11336 6724 11388 6730
rect 11336 6666 11388 6672
rect 11348 5914 11376 6666
rect 11440 6458 11468 7278
rect 11532 7206 11560 7414
rect 11520 7200 11572 7206
rect 11520 7142 11572 7148
rect 11532 6866 11560 7142
rect 11624 7002 11652 7890
rect 11716 7886 11744 8366
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 11520 6860 11572 6866
rect 11520 6802 11572 6808
rect 11532 6730 11560 6802
rect 11520 6724 11572 6730
rect 11520 6666 11572 6672
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 11532 6066 11560 6666
rect 11440 6038 11560 6066
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11440 5710 11468 6038
rect 11428 5704 11480 5710
rect 11428 5646 11480 5652
rect 11244 5364 11296 5370
rect 11244 5306 11296 5312
rect 11440 4622 11468 5646
rect 11704 5636 11756 5642
rect 11704 5578 11756 5584
rect 11072 4542 11192 4570
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 10980 4049 11008 4082
rect 10966 4040 11022 4049
rect 10966 3975 11022 3984
rect 10600 3936 10652 3942
rect 11072 3890 11100 4542
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 10600 3878 10652 3884
rect 10612 3534 10640 3878
rect 10888 3862 11100 3890
rect 10888 3738 10916 3862
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 10508 2848 10560 2854
rect 10508 2790 10560 2796
rect 10612 2774 10640 3470
rect 10980 3194 11008 3674
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 11164 3058 11192 4422
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 11624 3058 11652 3878
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 10612 2746 10732 2774
rect 10704 800 10732 2746
rect 10968 2372 11020 2378
rect 10968 2314 11020 2320
rect 10980 1834 11008 2314
rect 10968 1828 11020 1834
rect 10968 1770 11020 1776
rect 11072 800 11100 2994
rect 11624 2774 11652 2994
rect 11440 2746 11652 2774
rect 11440 800 11468 2746
rect 11716 2310 11744 5578
rect 11796 3120 11848 3126
rect 11796 3062 11848 3068
rect 11704 2304 11756 2310
rect 11704 2246 11756 2252
rect 11808 800 11836 3062
rect 11900 2650 11928 10950
rect 11992 10266 12020 13126
rect 12084 12374 12112 15302
rect 12348 14068 12400 14074
rect 12348 14010 12400 14016
rect 12256 13728 12308 13734
rect 12256 13670 12308 13676
rect 12164 13184 12216 13190
rect 12164 13126 12216 13132
rect 12176 12434 12204 13126
rect 12268 12986 12296 13670
rect 12360 13258 12388 14010
rect 12348 13252 12400 13258
rect 12348 13194 12400 13200
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12348 12708 12400 12714
rect 12348 12650 12400 12656
rect 12176 12406 12296 12434
rect 12072 12368 12124 12374
rect 12072 12310 12124 12316
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12070 11792 12126 11801
rect 12070 11727 12072 11736
rect 12124 11727 12126 11736
rect 12072 11698 12124 11704
rect 12072 11144 12124 11150
rect 12072 11086 12124 11092
rect 12084 11014 12112 11086
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 12072 10600 12124 10606
rect 12072 10542 12124 10548
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 12084 10062 12112 10542
rect 12176 10130 12204 12242
rect 12268 11218 12296 12406
rect 12360 12050 12388 12650
rect 12452 12646 12480 16646
rect 12532 15428 12584 15434
rect 12532 15370 12584 15376
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12438 12472 12494 12481
rect 12544 12442 12572 15370
rect 12636 14618 12664 18566
rect 12820 18222 12848 19110
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 12808 18216 12860 18222
rect 12808 18158 12860 18164
rect 12716 17536 12768 17542
rect 12714 17504 12716 17513
rect 12768 17504 12770 17513
rect 12714 17439 12770 17448
rect 12820 16794 12848 18158
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 13372 17746 13400 21014
rect 13452 20392 13504 20398
rect 13452 20334 13504 20340
rect 13360 17740 13412 17746
rect 13360 17682 13412 17688
rect 13176 17536 13228 17542
rect 13176 17478 13228 17484
rect 13188 17338 13216 17478
rect 13176 17332 13228 17338
rect 13176 17274 13228 17280
rect 13360 17332 13412 17338
rect 13360 17274 13412 17280
rect 13372 17134 13400 17274
rect 13464 17134 13492 20334
rect 13556 18290 13584 22066
rect 13636 20596 13688 20602
rect 13636 20538 13688 20544
rect 13544 18284 13596 18290
rect 13544 18226 13596 18232
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 13452 17128 13504 17134
rect 13452 17070 13504 17076
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 13372 14498 13400 17070
rect 13648 17066 13676 20538
rect 14016 20058 14044 23666
rect 14096 22432 14148 22438
rect 14096 22374 14148 22380
rect 14108 22030 14136 22374
rect 14096 22024 14148 22030
rect 14096 21966 14148 21972
rect 14108 21690 14136 21966
rect 14096 21684 14148 21690
rect 14096 21626 14148 21632
rect 14200 21434 14228 25842
rect 14476 23322 14504 26386
rect 14844 25362 14872 26386
rect 14740 25356 14792 25362
rect 14740 25298 14792 25304
rect 14832 25356 14884 25362
rect 14832 25298 14884 25304
rect 14752 24750 14780 25298
rect 14740 24744 14792 24750
rect 14740 24686 14792 24692
rect 14740 24608 14792 24614
rect 14740 24550 14792 24556
rect 14752 24342 14780 24550
rect 14844 24410 14872 25298
rect 14832 24404 14884 24410
rect 14832 24346 14884 24352
rect 14740 24336 14792 24342
rect 14740 24278 14792 24284
rect 14556 23588 14608 23594
rect 14556 23530 14608 23536
rect 14464 23316 14516 23322
rect 14464 23258 14516 23264
rect 14476 23118 14504 23258
rect 14464 23112 14516 23118
rect 14464 23054 14516 23060
rect 14108 21406 14228 21434
rect 14108 21350 14136 21406
rect 14096 21344 14148 21350
rect 14096 21286 14148 21292
rect 14372 21344 14424 21350
rect 14372 21286 14424 21292
rect 14384 20398 14412 21286
rect 14372 20392 14424 20398
rect 14372 20334 14424 20340
rect 14464 20256 14516 20262
rect 14464 20198 14516 20204
rect 14004 20052 14056 20058
rect 14004 19994 14056 20000
rect 14476 19310 14504 20198
rect 14568 19922 14596 23530
rect 14752 22778 14780 24278
rect 14936 23866 14964 26726
rect 15120 26450 15148 27474
rect 15108 26444 15160 26450
rect 15108 26386 15160 26392
rect 15120 25430 15148 26386
rect 15580 25498 15608 29514
rect 15672 28082 15700 45526
rect 15764 35494 15792 46446
rect 15752 35488 15804 35494
rect 15752 35430 15804 35436
rect 16040 30274 16068 50458
rect 16132 44946 16160 53994
rect 16396 52692 16448 52698
rect 16396 52634 16448 52640
rect 16120 44940 16172 44946
rect 16120 44882 16172 44888
rect 16120 32972 16172 32978
rect 16120 32914 16172 32920
rect 16132 31890 16160 32914
rect 16120 31884 16172 31890
rect 16120 31826 16172 31832
rect 16132 31278 16160 31826
rect 16408 31770 16436 52634
rect 16488 46028 16540 46034
rect 16488 45970 16540 45976
rect 16500 34950 16528 45970
rect 16684 45554 16712 54062
rect 22192 53984 22244 53990
rect 22192 53926 22244 53932
rect 22652 53984 22704 53990
rect 22652 53926 22704 53932
rect 17950 53340 18258 53349
rect 17950 53338 17956 53340
rect 18012 53338 18036 53340
rect 18092 53338 18116 53340
rect 18172 53338 18196 53340
rect 18252 53338 18258 53340
rect 18012 53286 18014 53338
rect 18194 53286 18196 53338
rect 17950 53284 17956 53286
rect 18012 53284 18036 53286
rect 18092 53284 18116 53286
rect 18172 53284 18196 53286
rect 18252 53284 18258 53286
rect 17950 53275 18258 53284
rect 17950 52252 18258 52261
rect 17950 52250 17956 52252
rect 18012 52250 18036 52252
rect 18092 52250 18116 52252
rect 18172 52250 18196 52252
rect 18252 52250 18258 52252
rect 18012 52198 18014 52250
rect 18194 52198 18196 52250
rect 17950 52196 17956 52198
rect 18012 52196 18036 52198
rect 18092 52196 18116 52198
rect 18172 52196 18196 52198
rect 18252 52196 18258 52198
rect 17950 52187 18258 52196
rect 17950 51164 18258 51173
rect 17950 51162 17956 51164
rect 18012 51162 18036 51164
rect 18092 51162 18116 51164
rect 18172 51162 18196 51164
rect 18252 51162 18258 51164
rect 18012 51110 18014 51162
rect 18194 51110 18196 51162
rect 17950 51108 17956 51110
rect 18012 51108 18036 51110
rect 18092 51108 18116 51110
rect 18172 51108 18196 51110
rect 18252 51108 18258 51110
rect 17950 51099 18258 51108
rect 17950 50076 18258 50085
rect 17950 50074 17956 50076
rect 18012 50074 18036 50076
rect 18092 50074 18116 50076
rect 18172 50074 18196 50076
rect 18252 50074 18258 50076
rect 18012 50022 18014 50074
rect 18194 50022 18196 50074
rect 17950 50020 17956 50022
rect 18012 50020 18036 50022
rect 18092 50020 18116 50022
rect 18172 50020 18196 50022
rect 18252 50020 18258 50022
rect 17950 50011 18258 50020
rect 17950 48988 18258 48997
rect 17950 48986 17956 48988
rect 18012 48986 18036 48988
rect 18092 48986 18116 48988
rect 18172 48986 18196 48988
rect 18252 48986 18258 48988
rect 18012 48934 18014 48986
rect 18194 48934 18196 48986
rect 17950 48932 17956 48934
rect 18012 48932 18036 48934
rect 18092 48932 18116 48934
rect 18172 48932 18196 48934
rect 18252 48932 18258 48934
rect 17950 48923 18258 48932
rect 17950 47900 18258 47909
rect 17950 47898 17956 47900
rect 18012 47898 18036 47900
rect 18092 47898 18116 47900
rect 18172 47898 18196 47900
rect 18252 47898 18258 47900
rect 18012 47846 18014 47898
rect 18194 47846 18196 47898
rect 17950 47844 17956 47846
rect 18012 47844 18036 47846
rect 18092 47844 18116 47846
rect 18172 47844 18196 47846
rect 18252 47844 18258 47846
rect 17950 47835 18258 47844
rect 17950 46812 18258 46821
rect 17950 46810 17956 46812
rect 18012 46810 18036 46812
rect 18092 46810 18116 46812
rect 18172 46810 18196 46812
rect 18252 46810 18258 46812
rect 18012 46758 18014 46810
rect 18194 46758 18196 46810
rect 17950 46756 17956 46758
rect 18012 46756 18036 46758
rect 18092 46756 18116 46758
rect 18172 46756 18196 46758
rect 18252 46756 18258 46758
rect 17950 46747 18258 46756
rect 17950 45724 18258 45733
rect 17950 45722 17956 45724
rect 18012 45722 18036 45724
rect 18092 45722 18116 45724
rect 18172 45722 18196 45724
rect 18252 45722 18258 45724
rect 18012 45670 18014 45722
rect 18194 45670 18196 45722
rect 17950 45668 17956 45670
rect 18012 45668 18036 45670
rect 18092 45668 18116 45670
rect 18172 45668 18196 45670
rect 18252 45668 18258 45670
rect 17950 45659 18258 45668
rect 16592 45526 16712 45554
rect 16488 34944 16540 34950
rect 16488 34886 16540 34892
rect 16592 33114 16620 45526
rect 19984 44804 20036 44810
rect 19984 44746 20036 44752
rect 17950 44636 18258 44645
rect 17950 44634 17956 44636
rect 18012 44634 18036 44636
rect 18092 44634 18116 44636
rect 18172 44634 18196 44636
rect 18252 44634 18258 44636
rect 18012 44582 18014 44634
rect 18194 44582 18196 44634
rect 17950 44580 17956 44582
rect 18012 44580 18036 44582
rect 18092 44580 18116 44582
rect 18172 44580 18196 44582
rect 18252 44580 18258 44582
rect 17950 44571 18258 44580
rect 19524 43784 19576 43790
rect 19524 43726 19576 43732
rect 17950 43548 18258 43557
rect 17950 43546 17956 43548
rect 18012 43546 18036 43548
rect 18092 43546 18116 43548
rect 18172 43546 18196 43548
rect 18252 43546 18258 43548
rect 18012 43494 18014 43546
rect 18194 43494 18196 43546
rect 17950 43492 17956 43494
rect 18012 43492 18036 43494
rect 18092 43492 18116 43494
rect 18172 43492 18196 43494
rect 18252 43492 18258 43494
rect 17950 43483 18258 43492
rect 17950 42460 18258 42469
rect 17950 42458 17956 42460
rect 18012 42458 18036 42460
rect 18092 42458 18116 42460
rect 18172 42458 18196 42460
rect 18252 42458 18258 42460
rect 18012 42406 18014 42458
rect 18194 42406 18196 42458
rect 17950 42404 17956 42406
rect 18012 42404 18036 42406
rect 18092 42404 18116 42406
rect 18172 42404 18196 42406
rect 18252 42404 18258 42406
rect 17950 42395 18258 42404
rect 17950 41372 18258 41381
rect 17950 41370 17956 41372
rect 18012 41370 18036 41372
rect 18092 41370 18116 41372
rect 18172 41370 18196 41372
rect 18252 41370 18258 41372
rect 18012 41318 18014 41370
rect 18194 41318 18196 41370
rect 17950 41316 17956 41318
rect 18012 41316 18036 41318
rect 18092 41316 18116 41318
rect 18172 41316 18196 41318
rect 18252 41316 18258 41318
rect 17950 41307 18258 41316
rect 17950 40284 18258 40293
rect 17950 40282 17956 40284
rect 18012 40282 18036 40284
rect 18092 40282 18116 40284
rect 18172 40282 18196 40284
rect 18252 40282 18258 40284
rect 18012 40230 18014 40282
rect 18194 40230 18196 40282
rect 17950 40228 17956 40230
rect 18012 40228 18036 40230
rect 18092 40228 18116 40230
rect 18172 40228 18196 40230
rect 18252 40228 18258 40230
rect 17950 40219 18258 40228
rect 17950 39196 18258 39205
rect 17950 39194 17956 39196
rect 18012 39194 18036 39196
rect 18092 39194 18116 39196
rect 18172 39194 18196 39196
rect 18252 39194 18258 39196
rect 18012 39142 18014 39194
rect 18194 39142 18196 39194
rect 17950 39140 17956 39142
rect 18012 39140 18036 39142
rect 18092 39140 18116 39142
rect 18172 39140 18196 39142
rect 18252 39140 18258 39142
rect 17950 39131 18258 39140
rect 17950 38108 18258 38117
rect 17950 38106 17956 38108
rect 18012 38106 18036 38108
rect 18092 38106 18116 38108
rect 18172 38106 18196 38108
rect 18252 38106 18258 38108
rect 18012 38054 18014 38106
rect 18194 38054 18196 38106
rect 17950 38052 17956 38054
rect 18012 38052 18036 38054
rect 18092 38052 18116 38054
rect 18172 38052 18196 38054
rect 18252 38052 18258 38054
rect 17950 38043 18258 38052
rect 17950 37020 18258 37029
rect 17950 37018 17956 37020
rect 18012 37018 18036 37020
rect 18092 37018 18116 37020
rect 18172 37018 18196 37020
rect 18252 37018 18258 37020
rect 18012 36966 18014 37018
rect 18194 36966 18196 37018
rect 17950 36964 17956 36966
rect 18012 36964 18036 36966
rect 18092 36964 18116 36966
rect 18172 36964 18196 36966
rect 18252 36964 18258 36966
rect 17950 36955 18258 36964
rect 17950 35932 18258 35941
rect 17950 35930 17956 35932
rect 18012 35930 18036 35932
rect 18092 35930 18116 35932
rect 18172 35930 18196 35932
rect 18252 35930 18258 35932
rect 18012 35878 18014 35930
rect 18194 35878 18196 35930
rect 17950 35876 17956 35878
rect 18012 35876 18036 35878
rect 18092 35876 18116 35878
rect 18172 35876 18196 35878
rect 18252 35876 18258 35878
rect 17950 35867 18258 35876
rect 19340 35556 19392 35562
rect 19340 35498 19392 35504
rect 17950 34844 18258 34853
rect 17950 34842 17956 34844
rect 18012 34842 18036 34844
rect 18092 34842 18116 34844
rect 18172 34842 18196 34844
rect 18252 34842 18258 34844
rect 18012 34790 18014 34842
rect 18194 34790 18196 34842
rect 17950 34788 17956 34790
rect 18012 34788 18036 34790
rect 18092 34788 18116 34790
rect 18172 34788 18196 34790
rect 18252 34788 18258 34790
rect 17950 34779 18258 34788
rect 17950 33756 18258 33765
rect 17950 33754 17956 33756
rect 18012 33754 18036 33756
rect 18092 33754 18116 33756
rect 18172 33754 18196 33756
rect 18252 33754 18258 33756
rect 18012 33702 18014 33754
rect 18194 33702 18196 33754
rect 17950 33700 17956 33702
rect 18012 33700 18036 33702
rect 18092 33700 18116 33702
rect 18172 33700 18196 33702
rect 18252 33700 18258 33702
rect 17950 33691 18258 33700
rect 16580 33108 16632 33114
rect 16580 33050 16632 33056
rect 17316 33108 17368 33114
rect 17316 33050 17368 33056
rect 16856 33040 16908 33046
rect 16856 32982 16908 32988
rect 17132 33040 17184 33046
rect 17132 32982 17184 32988
rect 16868 32774 16896 32982
rect 16856 32768 16908 32774
rect 16856 32710 16908 32716
rect 16764 32360 16816 32366
rect 16764 32302 16816 32308
rect 16776 31822 16804 32302
rect 16764 31816 16816 31822
rect 16408 31726 16528 31770
rect 16764 31758 16816 31764
rect 16672 31748 16724 31754
rect 16120 31272 16172 31278
rect 16120 31214 16172 31220
rect 16040 30246 16160 30274
rect 16028 30184 16080 30190
rect 16028 30126 16080 30132
rect 15936 30048 15988 30054
rect 15936 29990 15988 29996
rect 15948 29238 15976 29990
rect 16040 29714 16068 30126
rect 16028 29708 16080 29714
rect 16028 29650 16080 29656
rect 16132 29560 16160 30246
rect 16040 29532 16160 29560
rect 15844 29232 15896 29238
rect 15844 29174 15896 29180
rect 15936 29232 15988 29238
rect 15936 29174 15988 29180
rect 15856 29073 15884 29174
rect 15842 29064 15898 29073
rect 15752 29028 15804 29034
rect 15842 28999 15898 29008
rect 15752 28970 15804 28976
rect 15660 28076 15712 28082
rect 15660 28018 15712 28024
rect 15764 27062 15792 28970
rect 16040 28422 16068 29532
rect 16304 29504 16356 29510
rect 16304 29446 16356 29452
rect 16316 29306 16344 29446
rect 16304 29300 16356 29306
rect 16304 29242 16356 29248
rect 16212 28688 16264 28694
rect 16212 28630 16264 28636
rect 16224 28422 16252 28630
rect 16028 28416 16080 28422
rect 16028 28358 16080 28364
rect 16212 28416 16264 28422
rect 16212 28358 16264 28364
rect 15936 28144 15988 28150
rect 15936 28086 15988 28092
rect 15752 27056 15804 27062
rect 15752 26998 15804 27004
rect 15948 26518 15976 28086
rect 16040 27334 16068 28358
rect 16224 27470 16252 28358
rect 16408 28150 16436 31726
rect 16672 31690 16724 31696
rect 16488 31680 16540 31686
rect 16488 31622 16540 31628
rect 16500 31482 16528 31622
rect 16488 31476 16540 31482
rect 16488 31418 16540 31424
rect 16684 31278 16712 31690
rect 16776 31346 16804 31758
rect 16764 31340 16816 31346
rect 16764 31282 16816 31288
rect 16672 31272 16724 31278
rect 16672 31214 16724 31220
rect 16948 30252 17000 30258
rect 16948 30194 17000 30200
rect 16764 30184 16816 30190
rect 16764 30126 16816 30132
rect 16488 30116 16540 30122
rect 16488 30058 16540 30064
rect 16500 29850 16528 30058
rect 16488 29844 16540 29850
rect 16488 29786 16540 29792
rect 16500 29646 16528 29786
rect 16488 29640 16540 29646
rect 16488 29582 16540 29588
rect 16396 28144 16448 28150
rect 16396 28086 16448 28092
rect 16304 28076 16356 28082
rect 16304 28018 16356 28024
rect 16316 27878 16344 28018
rect 16304 27872 16356 27878
rect 16304 27814 16356 27820
rect 16212 27464 16264 27470
rect 16212 27406 16264 27412
rect 16028 27328 16080 27334
rect 16028 27270 16080 27276
rect 15936 26512 15988 26518
rect 15936 26454 15988 26460
rect 15948 26314 15976 26454
rect 15936 26308 15988 26314
rect 15936 26250 15988 26256
rect 15568 25492 15620 25498
rect 15568 25434 15620 25440
rect 15108 25424 15160 25430
rect 15108 25366 15160 25372
rect 15580 25226 15608 25434
rect 15568 25220 15620 25226
rect 15568 25162 15620 25168
rect 15384 25152 15436 25158
rect 15580 25129 15608 25162
rect 15752 25152 15804 25158
rect 15384 25094 15436 25100
rect 15566 25120 15622 25129
rect 15396 24818 15424 25094
rect 15752 25094 15804 25100
rect 15566 25055 15622 25064
rect 15384 24812 15436 24818
rect 15384 24754 15436 24760
rect 15016 24744 15068 24750
rect 15016 24686 15068 24692
rect 14924 23860 14976 23866
rect 14924 23802 14976 23808
rect 14740 22772 14792 22778
rect 14740 22714 14792 22720
rect 14752 22094 14780 22714
rect 14660 22066 14780 22094
rect 14660 21418 14688 22066
rect 14832 21888 14884 21894
rect 14832 21830 14884 21836
rect 14844 21622 14872 21830
rect 14832 21616 14884 21622
rect 14832 21558 14884 21564
rect 14648 21412 14700 21418
rect 14648 21354 14700 21360
rect 14660 20806 14688 21354
rect 15028 21350 15056 24686
rect 15476 24608 15528 24614
rect 15476 24550 15528 24556
rect 15200 21888 15252 21894
rect 15200 21830 15252 21836
rect 15108 21684 15160 21690
rect 15108 21626 15160 21632
rect 15016 21344 15068 21350
rect 15016 21286 15068 21292
rect 14648 20800 14700 20806
rect 14648 20742 14700 20748
rect 14660 20534 14688 20742
rect 14648 20528 14700 20534
rect 14648 20470 14700 20476
rect 14660 19922 14688 20470
rect 14556 19916 14608 19922
rect 14556 19858 14608 19864
rect 14648 19916 14700 19922
rect 14648 19858 14700 19864
rect 14568 19718 14596 19858
rect 14660 19786 14688 19858
rect 14648 19780 14700 19786
rect 14648 19722 14700 19728
rect 14556 19712 14608 19718
rect 14556 19654 14608 19660
rect 14660 19446 14688 19722
rect 14648 19440 14700 19446
rect 14648 19382 14700 19388
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 14660 19174 14688 19382
rect 14372 19168 14424 19174
rect 14372 19110 14424 19116
rect 14648 19168 14700 19174
rect 14648 19110 14700 19116
rect 14280 18624 14332 18630
rect 14280 18566 14332 18572
rect 14096 18216 14148 18222
rect 14096 18158 14148 18164
rect 13912 17740 13964 17746
rect 13912 17682 13964 17688
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 13636 17060 13688 17066
rect 13636 17002 13688 17008
rect 13636 16652 13688 16658
rect 13636 16594 13688 16600
rect 13648 16454 13676 16594
rect 13636 16448 13688 16454
rect 13636 16390 13688 16396
rect 13280 14470 13400 14498
rect 13452 14476 13504 14482
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12636 12918 12664 13670
rect 12624 12912 12676 12918
rect 12624 12854 12676 12860
rect 12438 12407 12494 12416
rect 12532 12436 12584 12442
rect 12452 12238 12480 12407
rect 12532 12378 12584 12384
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 12360 12022 12480 12050
rect 12348 11824 12400 11830
rect 12346 11792 12348 11801
rect 12400 11792 12402 11801
rect 12346 11727 12402 11736
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12256 11212 12308 11218
rect 12256 11154 12308 11160
rect 12360 10742 12388 11494
rect 12452 11014 12480 12022
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12544 10826 12572 12174
rect 12624 12164 12676 12170
rect 12624 12106 12676 12112
rect 12452 10798 12572 10826
rect 12348 10736 12400 10742
rect 12348 10678 12400 10684
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 12072 6316 12124 6322
rect 12072 6258 12124 6264
rect 12084 3194 12112 6258
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 12360 5914 12388 6190
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12256 4752 12308 4758
rect 12254 4720 12256 4729
rect 12308 4720 12310 4729
rect 12254 4655 12310 4664
rect 12254 4584 12310 4593
rect 12254 4519 12310 4528
rect 12268 4146 12296 4519
rect 12256 4140 12308 4146
rect 12256 4082 12308 4088
rect 12452 4010 12480 10798
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12544 8022 12572 9454
rect 12636 9110 12664 12106
rect 12728 11150 12756 13806
rect 12820 11898 12848 14214
rect 13280 14006 13308 14470
rect 13452 14418 13504 14424
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 13268 14000 13320 14006
rect 13268 13942 13320 13948
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 13176 13456 13228 13462
rect 13176 13398 13228 13404
rect 12900 13252 12952 13258
rect 12900 13194 12952 13200
rect 12912 12850 12940 13194
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 13096 12753 13124 12922
rect 13188 12782 13216 13398
rect 13176 12776 13228 12782
rect 13082 12744 13138 12753
rect 13176 12718 13228 12724
rect 13082 12679 13138 12688
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 13084 12368 13136 12374
rect 13084 12310 13136 12316
rect 13096 11898 13124 12310
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 12808 11280 12860 11286
rect 13176 11280 13228 11286
rect 12808 11222 12860 11228
rect 13174 11248 13176 11257
rect 13228 11248 13230 11257
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12820 10742 12848 11222
rect 13174 11183 13230 11192
rect 12808 10736 12860 10742
rect 12808 10678 12860 10684
rect 13280 10520 13308 11290
rect 13372 10674 13400 14214
rect 13464 12782 13492 14418
rect 13544 14272 13596 14278
rect 13542 14240 13544 14249
rect 13596 14240 13598 14249
rect 13542 14175 13598 14184
rect 13556 14074 13584 14175
rect 13544 14068 13596 14074
rect 13544 14010 13596 14016
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13556 13410 13584 13874
rect 13648 13530 13676 16390
rect 13740 15994 13768 17138
rect 13924 16998 13952 17682
rect 14108 17610 14136 18158
rect 14292 17678 14320 18566
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14096 17604 14148 17610
rect 14096 17546 14148 17552
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 13924 16794 13952 16934
rect 13912 16788 13964 16794
rect 13912 16730 13964 16736
rect 14280 16788 14332 16794
rect 14280 16730 14332 16736
rect 13924 16522 13952 16730
rect 13912 16516 13964 16522
rect 13912 16458 13964 16464
rect 14188 16244 14240 16250
rect 14188 16186 14240 16192
rect 13820 16040 13872 16046
rect 13740 15988 13820 15994
rect 13740 15982 13872 15988
rect 13740 15966 13860 15982
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13556 13382 13676 13410
rect 13544 12844 13596 12850
rect 13544 12786 13596 12792
rect 13452 12776 13504 12782
rect 13452 12718 13504 12724
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 13464 11898 13492 12106
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 13452 11620 13504 11626
rect 13452 11562 13504 11568
rect 13464 11354 13492 11562
rect 13556 11370 13584 12786
rect 13648 12306 13676 13382
rect 13740 12968 13768 15966
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13832 13394 13860 13806
rect 13912 13728 13964 13734
rect 13912 13670 13964 13676
rect 14096 13728 14148 13734
rect 14096 13670 14148 13676
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 13924 13326 13952 13670
rect 13912 13320 13964 13326
rect 13912 13262 13964 13268
rect 13912 13184 13964 13190
rect 13912 13126 13964 13132
rect 13740 12940 13860 12968
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13636 12300 13688 12306
rect 13636 12242 13688 12248
rect 13648 11694 13676 12242
rect 13740 12238 13768 12786
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13832 12050 13860 12940
rect 13924 12442 13952 13126
rect 14004 12912 14056 12918
rect 14004 12854 14056 12860
rect 13912 12436 13964 12442
rect 13912 12378 13964 12384
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13740 12022 13860 12050
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 13452 11348 13504 11354
rect 13556 11342 13676 11370
rect 13452 11290 13504 11296
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13452 11008 13504 11014
rect 13452 10950 13504 10956
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13280 10492 13400 10520
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12716 10192 12768 10198
rect 12716 10134 12768 10140
rect 12624 9104 12676 9110
rect 12624 9046 12676 9052
rect 12532 8016 12584 8022
rect 12532 7958 12584 7964
rect 12544 6866 12572 7958
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12636 7546 12664 7686
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12624 4752 12676 4758
rect 12624 4694 12676 4700
rect 12440 4004 12492 4010
rect 12440 3946 12492 3952
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12544 3602 12572 3878
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 12164 2508 12216 2514
rect 12164 2450 12216 2456
rect 12176 800 12204 2450
rect 12544 800 12572 3538
rect 12636 2582 12664 4694
rect 12728 3670 12756 10134
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12820 9178 12848 9862
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 13372 9058 13400 10492
rect 13464 9926 13492 10950
rect 13556 10130 13584 11154
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13452 9920 13504 9926
rect 13452 9862 13504 9868
rect 12820 9030 13400 9058
rect 12820 6730 12848 9030
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 13372 7886 13400 8366
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 13266 6896 13322 6905
rect 13266 6831 13322 6840
rect 12808 6724 12860 6730
rect 12808 6666 12860 6672
rect 12820 4078 12848 6666
rect 13280 6390 13308 6831
rect 13372 6458 13400 7686
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 12900 6248 12952 6254
rect 12898 6216 12900 6225
rect 12952 6216 12954 6225
rect 12898 6151 12954 6160
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 13372 5778 13400 6054
rect 13360 5772 13412 5778
rect 13360 5714 13412 5720
rect 13464 5710 13492 9862
rect 13556 9042 13584 10066
rect 13648 9110 13676 11342
rect 13740 10198 13768 12022
rect 13820 11280 13872 11286
rect 13820 11222 13872 11228
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 13740 9450 13768 9930
rect 13728 9444 13780 9450
rect 13728 9386 13780 9392
rect 13832 9330 13860 11222
rect 13924 10418 13952 12242
rect 14016 10538 14044 12854
rect 14108 12220 14136 13670
rect 14200 12374 14228 16186
rect 14292 16182 14320 16730
rect 14384 16726 14412 19110
rect 14464 18216 14516 18222
rect 14464 18158 14516 18164
rect 14476 17338 14504 18158
rect 14660 17746 14688 19110
rect 14648 17740 14700 17746
rect 14648 17682 14700 17688
rect 14464 17332 14516 17338
rect 14464 17274 14516 17280
rect 14832 17128 14884 17134
rect 14832 17070 14884 17076
rect 14924 17128 14976 17134
rect 14924 17070 14976 17076
rect 14372 16720 14424 16726
rect 14372 16662 14424 16668
rect 14280 16176 14332 16182
rect 14280 16118 14332 16124
rect 14280 16040 14332 16046
rect 14280 15982 14332 15988
rect 14292 15450 14320 15982
rect 14384 15978 14412 16662
rect 14740 16108 14792 16114
rect 14740 16050 14792 16056
rect 14372 15972 14424 15978
rect 14372 15914 14424 15920
rect 14292 15422 14412 15450
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 14292 15162 14320 15302
rect 14280 15156 14332 15162
rect 14280 15098 14332 15104
rect 14280 13524 14332 13530
rect 14280 13466 14332 13472
rect 14292 12918 14320 13466
rect 14280 12912 14332 12918
rect 14280 12854 14332 12860
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14188 12368 14240 12374
rect 14188 12310 14240 12316
rect 14292 12220 14320 12718
rect 14108 12192 14320 12220
rect 14004 10532 14056 10538
rect 14004 10474 14056 10480
rect 13924 10390 14044 10418
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13924 9654 13952 9862
rect 14016 9654 14044 10390
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 14004 9648 14056 9654
rect 14004 9590 14056 9596
rect 13740 9302 13860 9330
rect 13636 9104 13688 9110
rect 13636 9046 13688 9052
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13542 8936 13598 8945
rect 13542 8871 13598 8880
rect 13556 8090 13584 8871
rect 13544 8084 13596 8090
rect 13544 8026 13596 8032
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 13556 6390 13584 6598
rect 13544 6384 13596 6390
rect 13544 6326 13596 6332
rect 13648 6186 13676 7482
rect 13740 6882 13768 9302
rect 13910 7848 13966 7857
rect 13910 7783 13966 7792
rect 13740 6854 13860 6882
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13636 6180 13688 6186
rect 13636 6122 13688 6128
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 13360 3936 13412 3942
rect 13360 3878 13412 3884
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 12716 3664 12768 3670
rect 12716 3606 12768 3612
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12624 2576 12676 2582
rect 12624 2518 12676 2524
rect 12820 1714 12848 3538
rect 13372 3534 13400 3878
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13174 3088 13230 3097
rect 13174 3023 13176 3032
rect 13228 3023 13230 3032
rect 13176 2994 13228 3000
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 13556 2582 13584 5510
rect 13648 5370 13676 6122
rect 13636 5364 13688 5370
rect 13636 5306 13688 5312
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 13544 2576 13596 2582
rect 13544 2518 13596 2524
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 12820 1686 12940 1714
rect 12912 800 12940 1686
rect 13280 800 13308 2314
rect 13648 800 13676 2926
rect 13740 2038 13768 6734
rect 13832 6458 13860 6854
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13832 6322 13860 6394
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 13924 5114 13952 7783
rect 13832 5086 13952 5114
rect 13832 4690 13860 5086
rect 13912 5024 13964 5030
rect 13912 4966 13964 4972
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 13924 4146 13952 4966
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 14016 4026 14044 9590
rect 14108 9518 14136 12192
rect 14384 11898 14412 15422
rect 14752 14278 14780 16050
rect 14844 14498 14872 17070
rect 14936 14770 14964 17070
rect 15016 16448 15068 16454
rect 15016 16390 15068 16396
rect 15028 16250 15056 16390
rect 15016 16244 15068 16250
rect 15016 16186 15068 16192
rect 14936 14742 15056 14770
rect 14844 14482 14964 14498
rect 14844 14476 14976 14482
rect 14844 14470 14924 14476
rect 14464 14272 14516 14278
rect 14740 14272 14792 14278
rect 14464 14214 14516 14220
rect 14738 14240 14740 14249
rect 14792 14240 14794 14249
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14372 11892 14424 11898
rect 14372 11834 14424 11840
rect 14200 11150 14228 11834
rect 14476 11830 14504 14214
rect 14738 14175 14794 14184
rect 14844 14074 14872 14470
rect 14924 14418 14976 14424
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 14554 12472 14610 12481
rect 14554 12407 14610 12416
rect 14568 12306 14596 12407
rect 14648 12368 14700 12374
rect 14844 12356 14872 12718
rect 14936 12481 14964 12786
rect 14922 12472 14978 12481
rect 14922 12407 14978 12416
rect 14844 12328 14964 12356
rect 14648 12310 14700 12316
rect 14556 12300 14608 12306
rect 14556 12242 14608 12248
rect 14464 11824 14516 11830
rect 14464 11766 14516 11772
rect 14660 11762 14688 12310
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14372 11688 14424 11694
rect 14372 11630 14424 11636
rect 14384 11218 14412 11630
rect 14464 11280 14516 11286
rect 14464 11222 14516 11228
rect 14372 11212 14424 11218
rect 14372 11154 14424 11160
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14292 10810 14320 10950
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14188 10668 14240 10674
rect 14188 10610 14240 10616
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14200 10577 14228 10610
rect 14186 10568 14242 10577
rect 14186 10503 14242 10512
rect 14096 9512 14148 9518
rect 14096 9454 14148 9460
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 14096 8356 14148 8362
rect 14096 8298 14148 8304
rect 13924 3998 14044 4026
rect 13924 3126 13952 3998
rect 14004 3596 14056 3602
rect 14004 3538 14056 3544
rect 13912 3120 13964 3126
rect 13912 3062 13964 3068
rect 13728 2032 13780 2038
rect 13728 1974 13780 1980
rect 14016 800 14044 3538
rect 14108 3058 14136 8298
rect 14200 8090 14228 8774
rect 14292 8498 14320 10610
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14292 7562 14320 8434
rect 14200 7534 14320 7562
rect 14200 7290 14228 7534
rect 14280 7472 14332 7478
rect 14384 7460 14412 10746
rect 14476 9586 14504 11222
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 14568 10266 14596 11086
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 14332 7432 14412 7460
rect 14280 7414 14332 7420
rect 14200 7262 14320 7290
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14200 4214 14228 4966
rect 14188 4208 14240 4214
rect 14188 4150 14240 4156
rect 14292 3398 14320 7262
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 14384 6458 14412 6598
rect 14372 6452 14424 6458
rect 14372 6394 14424 6400
rect 14476 5114 14504 9522
rect 14660 8974 14688 11698
rect 14832 11552 14884 11558
rect 14832 11494 14884 11500
rect 14844 11286 14872 11494
rect 14832 11280 14884 11286
rect 14832 11222 14884 11228
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 14752 10266 14780 11154
rect 14832 11008 14884 11014
rect 14832 10950 14884 10956
rect 14740 10260 14792 10266
rect 14740 10202 14792 10208
rect 14648 8968 14700 8974
rect 14648 8910 14700 8916
rect 14648 8832 14700 8838
rect 14752 8786 14780 10202
rect 14844 9926 14872 10950
rect 14936 10130 14964 12328
rect 15028 12102 15056 14742
rect 15120 13802 15148 21626
rect 15212 17882 15240 21830
rect 15292 21412 15344 21418
rect 15292 21354 15344 21360
rect 15304 21146 15332 21354
rect 15292 21140 15344 21146
rect 15292 21082 15344 21088
rect 15488 20602 15516 24550
rect 15660 23656 15712 23662
rect 15660 23598 15712 23604
rect 15672 23118 15700 23598
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 15764 22166 15792 25094
rect 15752 22160 15804 22166
rect 15752 22102 15804 22108
rect 15568 21140 15620 21146
rect 15568 21082 15620 21088
rect 15476 20596 15528 20602
rect 15476 20538 15528 20544
rect 15384 19712 15436 19718
rect 15384 19654 15436 19660
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 15108 13796 15160 13802
rect 15108 13738 15160 13744
rect 15120 13462 15148 13738
rect 15108 13456 15160 13462
rect 15108 13398 15160 13404
rect 15108 13320 15160 13326
rect 15108 13262 15160 13268
rect 15120 12782 15148 13262
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 15108 12300 15160 12306
rect 15108 12242 15160 12248
rect 15016 12096 15068 12102
rect 15016 12038 15068 12044
rect 15028 11558 15056 12038
rect 15120 11694 15148 12242
rect 15108 11688 15160 11694
rect 15108 11630 15160 11636
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 15212 11354 15240 13126
rect 15304 12102 15332 19450
rect 15396 16998 15424 19654
rect 15580 19378 15608 21082
rect 15752 20868 15804 20874
rect 15752 20810 15804 20816
rect 15764 20058 15792 20810
rect 15752 20052 15804 20058
rect 15752 19994 15804 20000
rect 15568 19372 15620 19378
rect 15568 19314 15620 19320
rect 15764 19310 15792 19994
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 15752 19304 15804 19310
rect 15752 19246 15804 19252
rect 15856 18970 15884 19790
rect 15936 19780 15988 19786
rect 15936 19722 15988 19728
rect 15844 18964 15896 18970
rect 15844 18906 15896 18912
rect 15568 17604 15620 17610
rect 15568 17546 15620 17552
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 15396 14958 15424 16934
rect 15476 16516 15528 16522
rect 15476 16458 15528 16464
rect 15488 16250 15516 16458
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15580 15162 15608 17546
rect 15752 17536 15804 17542
rect 15752 17478 15804 17484
rect 15764 16590 15792 17478
rect 15844 16652 15896 16658
rect 15844 16594 15896 16600
rect 15752 16584 15804 16590
rect 15752 16526 15804 16532
rect 15752 15360 15804 15366
rect 15752 15302 15804 15308
rect 15764 15162 15792 15302
rect 15568 15156 15620 15162
rect 15568 15098 15620 15104
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 15384 14952 15436 14958
rect 15384 14894 15436 14900
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15488 12986 15516 14894
rect 15752 14544 15804 14550
rect 15752 14486 15804 14492
rect 15660 13796 15712 13802
rect 15660 13738 15712 13744
rect 15672 13274 15700 13738
rect 15764 13394 15792 14486
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15856 13326 15884 16594
rect 15948 16454 15976 19722
rect 15936 16448 15988 16454
rect 15936 16390 15988 16396
rect 15844 13320 15896 13326
rect 15672 13246 15792 13274
rect 15844 13262 15896 13268
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15488 12434 15516 12922
rect 15660 12776 15712 12782
rect 15660 12718 15712 12724
rect 15488 12406 15608 12434
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15304 11937 15332 12038
rect 15290 11928 15346 11937
rect 15290 11863 15346 11872
rect 15476 11620 15528 11626
rect 15476 11562 15528 11568
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 15396 11234 15424 11494
rect 15212 11206 15424 11234
rect 15212 11082 15240 11206
rect 15488 11082 15516 11562
rect 15108 11076 15160 11082
rect 15108 11018 15160 11024
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 15476 11076 15528 11082
rect 15476 11018 15528 11024
rect 15014 10704 15070 10713
rect 15014 10639 15070 10648
rect 14924 10124 14976 10130
rect 14924 10066 14976 10072
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 14844 8922 14872 9862
rect 14936 9518 14964 10066
rect 15028 10062 15056 10639
rect 15016 10056 15068 10062
rect 15016 9998 15068 10004
rect 14924 9512 14976 9518
rect 14924 9454 14976 9460
rect 14936 9042 14964 9454
rect 15120 9450 15148 11018
rect 15108 9444 15160 9450
rect 15108 9386 15160 9392
rect 14924 9036 14976 9042
rect 14924 8978 14976 8984
rect 14844 8894 14964 8922
rect 14700 8780 14780 8786
rect 14648 8774 14780 8780
rect 14660 8758 14780 8774
rect 14554 7984 14610 7993
rect 14554 7919 14556 7928
rect 14608 7919 14610 7928
rect 14556 7890 14608 7896
rect 14476 5086 14596 5114
rect 14462 3632 14518 3641
rect 14462 3567 14518 3576
rect 14476 3534 14504 3567
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14568 3466 14596 5086
rect 14556 3460 14608 3466
rect 14556 3402 14608 3408
rect 14660 3398 14688 8758
rect 14832 8424 14884 8430
rect 14832 8366 14884 8372
rect 14740 6792 14792 6798
rect 14740 6734 14792 6740
rect 14752 5914 14780 6734
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 14844 3777 14872 8366
rect 14936 7460 14964 8894
rect 15016 8016 15068 8022
rect 15212 7993 15240 11018
rect 15384 11008 15436 11014
rect 15384 10950 15436 10956
rect 15292 10736 15344 10742
rect 15292 10678 15344 10684
rect 15304 10606 15332 10678
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15396 9926 15424 10950
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15396 8514 15424 9862
rect 15304 8486 15424 8514
rect 15016 7958 15068 7964
rect 15198 7984 15254 7993
rect 15028 7750 15056 7958
rect 15198 7919 15254 7928
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 15016 7472 15068 7478
rect 14936 7432 15016 7460
rect 15016 7414 15068 7420
rect 15028 6798 15056 7414
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 15028 6662 15056 6734
rect 15016 6656 15068 6662
rect 15016 6598 15068 6604
rect 14924 5840 14976 5846
rect 14924 5782 14976 5788
rect 14936 5030 14964 5782
rect 15028 5710 15056 6598
rect 15120 5710 15148 7142
rect 15016 5704 15068 5710
rect 15016 5646 15068 5652
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 15028 5302 15056 5646
rect 15016 5296 15068 5302
rect 15016 5238 15068 5244
rect 14924 5024 14976 5030
rect 14924 4966 14976 4972
rect 15120 4690 15148 5646
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 15108 4548 15160 4554
rect 15108 4490 15160 4496
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 15120 4434 15148 4490
rect 14936 4214 14964 4422
rect 15120 4406 15240 4434
rect 14924 4208 14976 4214
rect 14924 4150 14976 4156
rect 14830 3768 14886 3777
rect 14830 3703 14886 3712
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 14648 3392 14700 3398
rect 14648 3334 14700 3340
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 15016 3052 15068 3058
rect 15016 2994 15068 3000
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14372 2508 14424 2514
rect 14372 2450 14424 2456
rect 14384 800 14412 2450
rect 14752 800 14780 2926
rect 15028 2854 15056 2994
rect 15016 2848 15068 2854
rect 15016 2790 15068 2796
rect 15108 2848 15160 2854
rect 15108 2790 15160 2796
rect 15120 800 15148 2790
rect 15212 2650 15240 4406
rect 15304 4162 15332 8486
rect 15474 7304 15530 7313
rect 15474 7239 15530 7248
rect 15488 7206 15516 7239
rect 15476 7200 15528 7206
rect 15476 7142 15528 7148
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 15396 4554 15424 6802
rect 15488 6730 15516 7142
rect 15476 6724 15528 6730
rect 15476 6666 15528 6672
rect 15488 6225 15516 6666
rect 15474 6216 15530 6225
rect 15474 6151 15530 6160
rect 15476 5296 15528 5302
rect 15476 5238 15528 5244
rect 15488 4554 15516 5238
rect 15384 4548 15436 4554
rect 15384 4490 15436 4496
rect 15476 4548 15528 4554
rect 15476 4490 15528 4496
rect 15396 4298 15424 4490
rect 15396 4270 15516 4298
rect 15304 4134 15424 4162
rect 15396 3058 15424 4134
rect 15488 4010 15516 4270
rect 15476 4004 15528 4010
rect 15476 3946 15528 3952
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15488 800 15516 3538
rect 15580 1970 15608 12406
rect 15672 10470 15700 12718
rect 15660 10464 15712 10470
rect 15660 10406 15712 10412
rect 15660 9512 15712 9518
rect 15660 9454 15712 9460
rect 15672 9178 15700 9454
rect 15660 9172 15712 9178
rect 15660 9114 15712 9120
rect 15672 2310 15700 9114
rect 15764 8634 15792 13246
rect 15936 12912 15988 12918
rect 15936 12854 15988 12860
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15752 7812 15804 7818
rect 15752 7754 15804 7760
rect 15764 6866 15792 7754
rect 15752 6860 15804 6866
rect 15752 6802 15804 6808
rect 15764 5642 15792 6802
rect 15856 6730 15884 12038
rect 15948 10588 15976 12854
rect 16040 11257 16068 27270
rect 16224 25158 16252 27406
rect 16316 26314 16344 27814
rect 16500 27418 16528 29582
rect 16408 27390 16528 27418
rect 16304 26308 16356 26314
rect 16304 26250 16356 26256
rect 16304 26036 16356 26042
rect 16304 25978 16356 25984
rect 16212 25152 16264 25158
rect 16212 25094 16264 25100
rect 16224 24886 16252 25094
rect 16212 24880 16264 24886
rect 16212 24822 16264 24828
rect 16316 18290 16344 25978
rect 16408 24818 16436 27390
rect 16488 27328 16540 27334
rect 16488 27270 16540 27276
rect 16396 24812 16448 24818
rect 16396 24754 16448 24760
rect 16396 21956 16448 21962
rect 16396 21898 16448 21904
rect 16408 20806 16436 21898
rect 16396 20800 16448 20806
rect 16396 20742 16448 20748
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 16408 18170 16436 20742
rect 16500 19378 16528 27270
rect 16776 26994 16804 30126
rect 16856 27872 16908 27878
rect 16856 27814 16908 27820
rect 16868 27130 16896 27814
rect 16856 27124 16908 27130
rect 16856 27066 16908 27072
rect 16764 26988 16816 26994
rect 16764 26930 16816 26936
rect 16776 26450 16804 26930
rect 16960 26586 16988 30194
rect 17144 29238 17172 32982
rect 17224 31272 17276 31278
rect 17224 31214 17276 31220
rect 17132 29232 17184 29238
rect 17132 29174 17184 29180
rect 17236 28150 17264 31214
rect 17328 29186 17356 33050
rect 17950 32668 18258 32677
rect 17950 32666 17956 32668
rect 18012 32666 18036 32668
rect 18092 32666 18116 32668
rect 18172 32666 18196 32668
rect 18252 32666 18258 32668
rect 18012 32614 18014 32666
rect 18194 32614 18196 32666
rect 17950 32612 17956 32614
rect 18012 32612 18036 32614
rect 18092 32612 18116 32614
rect 18172 32612 18196 32614
rect 18252 32612 18258 32614
rect 17950 32603 18258 32612
rect 18512 32020 18564 32026
rect 18512 31962 18564 31968
rect 18052 31952 18104 31958
rect 18052 31894 18104 31900
rect 17684 31884 17736 31890
rect 17684 31826 17736 31832
rect 17696 31754 17724 31826
rect 18064 31770 18092 31894
rect 17696 31726 17816 31754
rect 17788 31414 17816 31726
rect 17880 31742 18092 31770
rect 17880 31482 17908 31742
rect 17950 31580 18258 31589
rect 17950 31578 17956 31580
rect 18012 31578 18036 31580
rect 18092 31578 18116 31580
rect 18172 31578 18196 31580
rect 18252 31578 18258 31580
rect 18012 31526 18014 31578
rect 18194 31526 18196 31578
rect 17950 31524 17956 31526
rect 18012 31524 18036 31526
rect 18092 31524 18116 31526
rect 18172 31524 18196 31526
rect 18252 31524 18258 31526
rect 17950 31515 18258 31524
rect 17868 31476 17920 31482
rect 17868 31418 17920 31424
rect 17776 31408 17828 31414
rect 17776 31350 17828 31356
rect 17500 31136 17552 31142
rect 17552 31096 17632 31124
rect 17500 31078 17552 31084
rect 17408 29300 17460 29306
rect 17408 29242 17460 29248
rect 17420 29186 17448 29242
rect 17328 29158 17448 29186
rect 17328 29102 17356 29158
rect 17316 29096 17368 29102
rect 17408 29096 17460 29102
rect 17316 29038 17368 29044
rect 17406 29064 17408 29073
rect 17460 29064 17462 29073
rect 17224 28144 17276 28150
rect 17224 28086 17276 28092
rect 17236 27878 17264 28086
rect 17224 27872 17276 27878
rect 17224 27814 17276 27820
rect 16948 26580 17000 26586
rect 16948 26522 17000 26528
rect 16764 26444 16816 26450
rect 16764 26386 16816 26392
rect 16580 25900 16632 25906
rect 16580 25842 16632 25848
rect 16592 25702 16620 25842
rect 16580 25696 16632 25702
rect 16580 25638 16632 25644
rect 16776 23866 16804 26386
rect 16960 26382 16988 26522
rect 17224 26512 17276 26518
rect 17224 26454 17276 26460
rect 16948 26376 17000 26382
rect 16948 26318 17000 26324
rect 16856 25696 16908 25702
rect 16856 25638 16908 25644
rect 16868 25362 16896 25638
rect 16856 25356 16908 25362
rect 16856 25298 16908 25304
rect 16764 23860 16816 23866
rect 16764 23802 16816 23808
rect 16580 23656 16632 23662
rect 16580 23598 16632 23604
rect 16592 22982 16620 23598
rect 16764 23316 16816 23322
rect 16764 23258 16816 23264
rect 16580 22976 16632 22982
rect 16580 22918 16632 22924
rect 16776 22817 16804 23258
rect 16856 23044 16908 23050
rect 16856 22986 16908 22992
rect 16762 22808 16818 22817
rect 16868 22778 16896 22986
rect 16762 22743 16818 22752
rect 16856 22772 16908 22778
rect 16856 22714 16908 22720
rect 16580 21888 16632 21894
rect 16580 21830 16632 21836
rect 16592 21078 16620 21830
rect 16580 21072 16632 21078
rect 16580 21014 16632 21020
rect 16488 19372 16540 19378
rect 16488 19314 16540 19320
rect 16592 18290 16620 21014
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16580 18284 16632 18290
rect 16580 18226 16632 18232
rect 16316 18142 16436 18170
rect 16212 17740 16264 17746
rect 16212 17682 16264 17688
rect 16224 17542 16252 17682
rect 16212 17536 16264 17542
rect 16212 17478 16264 17484
rect 16224 17270 16252 17478
rect 16212 17264 16264 17270
rect 16212 17206 16264 17212
rect 16224 15348 16252 17206
rect 16316 16658 16344 18142
rect 16592 17338 16620 18226
rect 16396 17332 16448 17338
rect 16396 17274 16448 17280
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16408 16658 16436 17274
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16396 16652 16448 16658
rect 16396 16594 16448 16600
rect 16408 15570 16436 16594
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16396 15360 16448 15366
rect 16224 15320 16396 15348
rect 16396 15302 16448 15308
rect 16408 14074 16436 15302
rect 16684 14890 16712 19314
rect 16856 18964 16908 18970
rect 16856 18906 16908 18912
rect 16764 18624 16816 18630
rect 16764 18566 16816 18572
rect 16672 14884 16724 14890
rect 16672 14826 16724 14832
rect 16580 14272 16632 14278
rect 16580 14214 16632 14220
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16212 13388 16264 13394
rect 16212 13330 16264 13336
rect 16120 13320 16172 13326
rect 16120 13262 16172 13268
rect 16132 12986 16160 13262
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16026 11248 16082 11257
rect 16026 11183 16082 11192
rect 16028 10600 16080 10606
rect 15948 10560 16028 10588
rect 16028 10542 16080 10548
rect 16040 10198 16068 10542
rect 16028 10192 16080 10198
rect 16028 10134 16080 10140
rect 16132 10010 16160 11698
rect 15948 9982 16160 10010
rect 15948 8945 15976 9982
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 16132 9722 16160 9862
rect 16120 9716 16172 9722
rect 16120 9658 16172 9664
rect 16224 9518 16252 13330
rect 16304 13184 16356 13190
rect 16304 13126 16356 13132
rect 16316 12481 16344 13126
rect 16302 12472 16358 12481
rect 16302 12407 16358 12416
rect 16408 12434 16436 14010
rect 16488 13456 16540 13462
rect 16488 13398 16540 13404
rect 16500 12850 16528 13398
rect 16488 12844 16540 12850
rect 16488 12786 16540 12792
rect 16592 12646 16620 14214
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16408 12406 16528 12434
rect 16396 12300 16448 12306
rect 16396 12242 16448 12248
rect 16408 12170 16436 12242
rect 16396 12164 16448 12170
rect 16396 12106 16448 12112
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16316 11257 16344 11290
rect 16302 11248 16358 11257
rect 16302 11183 16358 11192
rect 16304 10192 16356 10198
rect 16304 10134 16356 10140
rect 16212 9512 16264 9518
rect 16212 9454 16264 9460
rect 15934 8936 15990 8945
rect 15934 8871 15990 8880
rect 15936 8832 15988 8838
rect 15936 8774 15988 8780
rect 15844 6724 15896 6730
rect 15844 6666 15896 6672
rect 15752 5636 15804 5642
rect 15752 5578 15804 5584
rect 15844 4548 15896 4554
rect 15844 4490 15896 4496
rect 15856 3482 15884 4490
rect 15948 3738 15976 8774
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 16132 7886 16160 8366
rect 16224 7954 16252 9454
rect 16212 7948 16264 7954
rect 16212 7890 16264 7896
rect 16120 7880 16172 7886
rect 16316 7834 16344 10134
rect 16120 7822 16172 7828
rect 16224 7806 16344 7834
rect 16224 6746 16252 7806
rect 16408 7410 16436 12106
rect 16500 11626 16528 12406
rect 16776 11898 16804 18566
rect 16868 18426 16896 18906
rect 16960 18834 16988 26318
rect 17132 25288 17184 25294
rect 17132 25230 17184 25236
rect 17144 24954 17172 25230
rect 17236 24954 17264 26454
rect 17132 24948 17184 24954
rect 17132 24890 17184 24896
rect 17224 24948 17276 24954
rect 17224 24890 17276 24896
rect 17040 24676 17092 24682
rect 17040 24618 17092 24624
rect 17052 21894 17080 24618
rect 17328 23730 17356 29038
rect 17406 28999 17462 29008
rect 17500 29028 17552 29034
rect 17420 28014 17448 28999
rect 17500 28970 17552 28976
rect 17408 28008 17460 28014
rect 17408 27950 17460 27956
rect 17408 26308 17460 26314
rect 17408 26250 17460 26256
rect 17316 23724 17368 23730
rect 17316 23666 17368 23672
rect 17316 23520 17368 23526
rect 17316 23462 17368 23468
rect 17040 21888 17092 21894
rect 17040 21830 17092 21836
rect 17132 21888 17184 21894
rect 17132 21830 17184 21836
rect 17144 20534 17172 21830
rect 17132 20528 17184 20534
rect 17132 20470 17184 20476
rect 17144 19990 17172 20470
rect 17224 20392 17276 20398
rect 17224 20334 17276 20340
rect 17132 19984 17184 19990
rect 17132 19926 17184 19932
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 16948 18692 17000 18698
rect 16948 18634 17000 18640
rect 16856 18420 16908 18426
rect 16856 18362 16908 18368
rect 16868 18057 16896 18362
rect 16854 18048 16910 18057
rect 16854 17983 16910 17992
rect 16960 16590 16988 18634
rect 17236 18358 17264 20334
rect 17328 19514 17356 23462
rect 17316 19508 17368 19514
rect 17316 19450 17368 19456
rect 17316 18760 17368 18766
rect 17316 18702 17368 18708
rect 17040 18352 17092 18358
rect 17040 18294 17092 18300
rect 17224 18352 17276 18358
rect 17224 18294 17276 18300
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 16854 16280 16910 16289
rect 16854 16215 16856 16224
rect 16908 16215 16910 16224
rect 16856 16186 16908 16192
rect 17052 14958 17080 18294
rect 17328 17678 17356 18702
rect 17420 17746 17448 26250
rect 17512 22094 17540 28970
rect 17604 27334 17632 31096
rect 17684 27940 17736 27946
rect 17684 27882 17736 27888
rect 17592 27328 17644 27334
rect 17592 27270 17644 27276
rect 17590 25936 17646 25945
rect 17590 25871 17592 25880
rect 17644 25871 17646 25880
rect 17592 25842 17644 25848
rect 17592 25764 17644 25770
rect 17592 25706 17644 25712
rect 17604 25294 17632 25706
rect 17592 25288 17644 25294
rect 17592 25230 17644 25236
rect 17696 24206 17724 27882
rect 17788 27538 17816 31350
rect 17880 28082 17908 31418
rect 18524 30938 18552 31962
rect 18788 31136 18840 31142
rect 18788 31078 18840 31084
rect 18800 30938 18828 31078
rect 18512 30932 18564 30938
rect 18512 30874 18564 30880
rect 18788 30932 18840 30938
rect 18788 30874 18840 30880
rect 18880 30932 18932 30938
rect 18880 30874 18932 30880
rect 18696 30592 18748 30598
rect 18696 30534 18748 30540
rect 18788 30592 18840 30598
rect 18892 30580 18920 30874
rect 18840 30552 18920 30580
rect 18788 30534 18840 30540
rect 17950 30492 18258 30501
rect 17950 30490 17956 30492
rect 18012 30490 18036 30492
rect 18092 30490 18116 30492
rect 18172 30490 18196 30492
rect 18252 30490 18258 30492
rect 18012 30438 18014 30490
rect 18194 30438 18196 30490
rect 17950 30436 17956 30438
rect 18012 30436 18036 30438
rect 18092 30436 18116 30438
rect 18172 30436 18196 30438
rect 18252 30436 18258 30438
rect 17950 30427 18258 30436
rect 18708 29850 18736 30534
rect 18800 30054 18828 30534
rect 18788 30048 18840 30054
rect 18788 29990 18840 29996
rect 18696 29844 18748 29850
rect 18696 29786 18748 29792
rect 18420 29776 18472 29782
rect 18420 29718 18472 29724
rect 17950 29404 18258 29413
rect 17950 29402 17956 29404
rect 18012 29402 18036 29404
rect 18092 29402 18116 29404
rect 18172 29402 18196 29404
rect 18252 29402 18258 29404
rect 18012 29350 18014 29402
rect 18194 29350 18196 29402
rect 17950 29348 17956 29350
rect 18012 29348 18036 29350
rect 18092 29348 18116 29350
rect 18172 29348 18196 29350
rect 18252 29348 18258 29350
rect 17950 29339 18258 29348
rect 17950 28316 18258 28325
rect 17950 28314 17956 28316
rect 18012 28314 18036 28316
rect 18092 28314 18116 28316
rect 18172 28314 18196 28316
rect 18252 28314 18258 28316
rect 18012 28262 18014 28314
rect 18194 28262 18196 28314
rect 17950 28260 17956 28262
rect 18012 28260 18036 28262
rect 18092 28260 18116 28262
rect 18172 28260 18196 28262
rect 18252 28260 18258 28262
rect 17950 28251 18258 28260
rect 17868 28076 17920 28082
rect 17868 28018 17920 28024
rect 17960 28008 18012 28014
rect 17960 27950 18012 27956
rect 17776 27532 17828 27538
rect 17776 27474 17828 27480
rect 17972 27470 18000 27950
rect 17960 27464 18012 27470
rect 17960 27406 18012 27412
rect 17950 27228 18258 27237
rect 17950 27226 17956 27228
rect 18012 27226 18036 27228
rect 18092 27226 18116 27228
rect 18172 27226 18196 27228
rect 18252 27226 18258 27228
rect 18012 27174 18014 27226
rect 18194 27174 18196 27226
rect 17950 27172 17956 27174
rect 18012 27172 18036 27174
rect 18092 27172 18116 27174
rect 18172 27172 18196 27174
rect 18252 27172 18258 27174
rect 17950 27163 18258 27172
rect 18328 26240 18380 26246
rect 18328 26182 18380 26188
rect 17950 26140 18258 26149
rect 17950 26138 17956 26140
rect 18012 26138 18036 26140
rect 18092 26138 18116 26140
rect 18172 26138 18196 26140
rect 18252 26138 18258 26140
rect 18012 26086 18014 26138
rect 18194 26086 18196 26138
rect 17950 26084 17956 26086
rect 18012 26084 18036 26086
rect 18092 26084 18116 26086
rect 18172 26084 18196 26086
rect 18252 26084 18258 26086
rect 17950 26075 18258 26084
rect 18340 26042 18368 26182
rect 18328 26036 18380 26042
rect 18328 25978 18380 25984
rect 18432 25974 18460 29718
rect 18512 27872 18564 27878
rect 18512 27814 18564 27820
rect 18420 25968 18472 25974
rect 18420 25910 18472 25916
rect 18524 25498 18552 27814
rect 18708 25838 18736 29786
rect 18800 29578 18828 29990
rect 19352 29866 19380 35498
rect 19536 34082 19564 43726
rect 19996 35018 20024 44746
rect 21088 43852 21140 43858
rect 21088 43794 21140 43800
rect 21100 43722 21128 43794
rect 21088 43716 21140 43722
rect 21088 43658 21140 43664
rect 19984 35012 20036 35018
rect 19984 34954 20036 34960
rect 20628 35012 20680 35018
rect 20628 34954 20680 34960
rect 20444 34468 20496 34474
rect 20444 34410 20496 34416
rect 19536 34066 19748 34082
rect 19536 34060 19760 34066
rect 19536 34054 19708 34060
rect 19432 33992 19484 33998
rect 19432 33934 19484 33940
rect 19444 32910 19472 33934
rect 19536 33522 19564 34054
rect 19708 34002 19760 34008
rect 19800 33924 19852 33930
rect 19800 33866 19852 33872
rect 19524 33516 19576 33522
rect 19524 33458 19576 33464
rect 19812 33454 19840 33866
rect 19800 33448 19852 33454
rect 19800 33390 19852 33396
rect 19432 32904 19484 32910
rect 19432 32846 19484 32852
rect 19444 32230 19472 32846
rect 19616 32768 19668 32774
rect 19616 32710 19668 32716
rect 19628 32570 19656 32710
rect 19616 32564 19668 32570
rect 19616 32506 19668 32512
rect 19800 32496 19852 32502
rect 19800 32438 19852 32444
rect 19432 32224 19484 32230
rect 19432 32166 19484 32172
rect 19444 31822 19472 32166
rect 19708 31884 19760 31890
rect 19708 31826 19760 31832
rect 19432 31816 19484 31822
rect 19432 31758 19484 31764
rect 19444 30802 19472 31758
rect 19720 31482 19748 31826
rect 19812 31754 19840 32438
rect 19800 31748 19852 31754
rect 19800 31690 19852 31696
rect 19708 31476 19760 31482
rect 19708 31418 19760 31424
rect 19708 31340 19760 31346
rect 19812 31328 19840 31690
rect 19760 31300 19840 31328
rect 19708 31282 19760 31288
rect 19720 30938 19748 31282
rect 20456 31278 20484 34410
rect 20536 33448 20588 33454
rect 20536 33390 20588 33396
rect 20444 31272 20496 31278
rect 20444 31214 20496 31220
rect 19708 30932 19760 30938
rect 19708 30874 19760 30880
rect 19432 30796 19484 30802
rect 19432 30738 19484 30744
rect 20076 30592 20128 30598
rect 20076 30534 20128 30540
rect 20088 30394 20116 30534
rect 20076 30388 20128 30394
rect 20076 30330 20128 30336
rect 19984 30320 20036 30326
rect 19984 30262 20036 30268
rect 19800 30048 19852 30054
rect 19800 29990 19852 29996
rect 19352 29838 19472 29866
rect 19340 29708 19392 29714
rect 19340 29650 19392 29656
rect 18880 29640 18932 29646
rect 18880 29582 18932 29588
rect 18788 29572 18840 29578
rect 18788 29514 18840 29520
rect 18800 28762 18828 29514
rect 18892 29510 18920 29582
rect 18880 29504 18932 29510
rect 18880 29446 18932 29452
rect 19156 29504 19208 29510
rect 19156 29446 19208 29452
rect 18892 28762 18920 29446
rect 19168 29306 19196 29446
rect 19156 29300 19208 29306
rect 19156 29242 19208 29248
rect 19064 29028 19116 29034
rect 19064 28970 19116 28976
rect 18788 28756 18840 28762
rect 18788 28698 18840 28704
rect 18880 28756 18932 28762
rect 18880 28698 18932 28704
rect 18800 28490 18828 28698
rect 18972 28620 19024 28626
rect 18972 28562 19024 28568
rect 18788 28484 18840 28490
rect 18788 28426 18840 28432
rect 18800 28218 18828 28426
rect 18788 28212 18840 28218
rect 18788 28154 18840 28160
rect 18788 28008 18840 28014
rect 18788 27950 18840 27956
rect 18696 25832 18748 25838
rect 18696 25774 18748 25780
rect 18604 25696 18656 25702
rect 18604 25638 18656 25644
rect 18512 25492 18564 25498
rect 18512 25434 18564 25440
rect 18524 25378 18552 25434
rect 18432 25350 18552 25378
rect 17950 25052 18258 25061
rect 17950 25050 17956 25052
rect 18012 25050 18036 25052
rect 18092 25050 18116 25052
rect 18172 25050 18196 25052
rect 18252 25050 18258 25052
rect 18012 24998 18014 25050
rect 18194 24998 18196 25050
rect 17950 24996 17956 24998
rect 18012 24996 18036 24998
rect 18092 24996 18116 24998
rect 18172 24996 18196 24998
rect 18252 24996 18258 24998
rect 17950 24987 18258 24996
rect 18328 24948 18380 24954
rect 18328 24890 18380 24896
rect 17868 24608 17920 24614
rect 17868 24550 17920 24556
rect 17684 24200 17736 24206
rect 17684 24142 17736 24148
rect 17512 22066 17632 22094
rect 17604 18630 17632 22066
rect 17696 18698 17724 24142
rect 17776 21956 17828 21962
rect 17776 21898 17828 21904
rect 17788 20806 17816 21898
rect 17776 20800 17828 20806
rect 17776 20742 17828 20748
rect 17788 20534 17816 20742
rect 17776 20528 17828 20534
rect 17776 20470 17828 20476
rect 17788 19922 17816 20470
rect 17776 19916 17828 19922
rect 17880 19904 17908 24550
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 18144 23860 18196 23866
rect 18144 23802 18196 23808
rect 18236 23860 18288 23866
rect 18236 23802 18288 23808
rect 18156 23526 18184 23802
rect 18144 23520 18196 23526
rect 18144 23462 18196 23468
rect 18248 22982 18276 23802
rect 18340 23118 18368 24890
rect 18432 24818 18460 25350
rect 18616 25294 18644 25638
rect 18604 25288 18656 25294
rect 18604 25230 18656 25236
rect 18512 25152 18564 25158
rect 18512 25094 18564 25100
rect 18420 24812 18472 24818
rect 18420 24754 18472 24760
rect 18524 24206 18552 25094
rect 18616 24886 18644 25230
rect 18604 24880 18656 24886
rect 18604 24822 18656 24828
rect 18512 24200 18564 24206
rect 18512 24142 18564 24148
rect 18420 24064 18472 24070
rect 18420 24006 18472 24012
rect 18328 23112 18380 23118
rect 18328 23054 18380 23060
rect 18236 22976 18288 22982
rect 18236 22918 18288 22924
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 18340 22778 18368 23054
rect 18328 22772 18380 22778
rect 18328 22714 18380 22720
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 17960 19916 18012 19922
rect 17880 19876 17960 19904
rect 17776 19858 17828 19864
rect 17960 19858 18012 19864
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 17776 18828 17828 18834
rect 17776 18770 17828 18776
rect 17684 18692 17736 18698
rect 17684 18634 17736 18640
rect 17592 18624 17644 18630
rect 17644 18572 17724 18578
rect 17592 18566 17724 18572
rect 17604 18550 17724 18566
rect 17592 18080 17644 18086
rect 17592 18022 17644 18028
rect 17408 17740 17460 17746
rect 17408 17682 17460 17688
rect 17500 17740 17552 17746
rect 17500 17682 17552 17688
rect 17316 17672 17368 17678
rect 17316 17614 17368 17620
rect 17224 17536 17276 17542
rect 17420 17490 17448 17682
rect 17224 17478 17276 17484
rect 17132 17060 17184 17066
rect 17132 17002 17184 17008
rect 17144 16697 17172 17002
rect 17130 16688 17186 16697
rect 17130 16623 17186 16632
rect 17040 14952 17092 14958
rect 17040 14894 17092 14900
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16868 12434 16896 13806
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 16868 12406 16988 12434
rect 16960 12170 16988 12406
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 16672 11688 16724 11694
rect 16672 11630 16724 11636
rect 16488 11620 16540 11626
rect 16488 11562 16540 11568
rect 16684 11286 16712 11630
rect 16764 11620 16816 11626
rect 16764 11562 16816 11568
rect 16776 11286 16804 11562
rect 16672 11280 16724 11286
rect 16672 11222 16724 11228
rect 16764 11280 16816 11286
rect 16764 11222 16816 11228
rect 16488 10600 16540 10606
rect 16488 10542 16540 10548
rect 16500 9042 16528 10542
rect 16488 9036 16540 9042
rect 16488 8978 16540 8984
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16500 7750 16528 8026
rect 16488 7744 16540 7750
rect 16488 7686 16540 7692
rect 16396 7404 16448 7410
rect 16396 7346 16448 7352
rect 16684 7342 16712 11222
rect 16960 11218 16988 12106
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 16856 10464 16908 10470
rect 16856 10406 16908 10412
rect 16868 10266 16896 10406
rect 16856 10260 16908 10266
rect 16856 10202 16908 10208
rect 16960 10062 16988 11154
rect 17040 10464 17092 10470
rect 17040 10406 17092 10412
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16396 6792 16448 6798
rect 16224 6718 16344 6746
rect 16396 6734 16448 6740
rect 16120 6248 16172 6254
rect 16120 6190 16172 6196
rect 16028 4072 16080 4078
rect 16028 4014 16080 4020
rect 15936 3732 15988 3738
rect 15936 3674 15988 3680
rect 16040 3670 16068 4014
rect 16028 3664 16080 3670
rect 16028 3606 16080 3612
rect 15856 3454 16068 3482
rect 15844 2984 15896 2990
rect 15844 2926 15896 2932
rect 15660 2304 15712 2310
rect 15660 2246 15712 2252
rect 15568 1964 15620 1970
rect 15568 1906 15620 1912
rect 15856 800 15884 2926
rect 16040 2446 16068 3454
rect 16132 2582 16160 6190
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16120 2576 16172 2582
rect 16120 2518 16172 2524
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 16224 800 16252 4014
rect 16316 2922 16344 6718
rect 16408 6118 16436 6734
rect 16580 6724 16632 6730
rect 16580 6666 16632 6672
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16592 4706 16620 6666
rect 16592 4678 16712 4706
rect 16580 3120 16632 3126
rect 16580 3062 16632 3068
rect 16304 2916 16356 2922
rect 16304 2858 16356 2864
rect 16302 2408 16358 2417
rect 16302 2343 16304 2352
rect 16356 2343 16358 2352
rect 16304 2314 16356 2320
rect 16592 800 16620 3062
rect 16684 2378 16712 4678
rect 16776 2446 16804 9862
rect 16960 9518 16988 9998
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16854 8936 16910 8945
rect 16854 8871 16910 8880
rect 16868 8838 16896 8871
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 16868 8537 16896 8570
rect 16854 8528 16910 8537
rect 16854 8463 16910 8472
rect 16856 7744 16908 7750
rect 16856 7686 16908 7692
rect 16868 7002 16896 7686
rect 16856 6996 16908 7002
rect 16856 6938 16908 6944
rect 16960 6798 16988 9454
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16868 5574 16896 6190
rect 16960 5778 16988 6734
rect 16948 5772 17000 5778
rect 16948 5714 17000 5720
rect 16856 5568 16908 5574
rect 16856 5510 16908 5516
rect 17052 3534 17080 10406
rect 17144 7750 17172 13670
rect 17236 12986 17264 17478
rect 17328 17462 17448 17490
rect 17328 15994 17356 17462
rect 17406 17368 17462 17377
rect 17406 17303 17408 17312
rect 17460 17303 17462 17312
rect 17408 17274 17460 17280
rect 17328 15966 17448 15994
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17328 15337 17356 15846
rect 17314 15328 17370 15337
rect 17314 15263 17370 15272
rect 17420 13682 17448 15966
rect 17512 13734 17540 17682
rect 17328 13654 17448 13682
rect 17500 13728 17552 13734
rect 17500 13670 17552 13676
rect 17328 13530 17356 13654
rect 17406 13560 17462 13569
rect 17316 13524 17368 13530
rect 17604 13546 17632 18022
rect 17696 15978 17724 18550
rect 17788 15994 17816 18770
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 18328 18080 18380 18086
rect 18328 18022 18380 18028
rect 18340 17746 18368 18022
rect 18328 17740 18380 17746
rect 18328 17682 18380 17688
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17868 17128 17920 17134
rect 17868 17070 17920 17076
rect 17880 16658 17908 17070
rect 17868 16652 17920 16658
rect 17868 16594 17920 16600
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17684 15972 17736 15978
rect 17788 15966 17908 15994
rect 17684 15914 17736 15920
rect 17776 15904 17828 15910
rect 17776 15846 17828 15852
rect 17684 15700 17736 15706
rect 17684 15642 17736 15648
rect 17406 13495 17408 13504
rect 17316 13466 17368 13472
rect 17460 13495 17462 13504
rect 17512 13518 17632 13546
rect 17408 13466 17460 13472
rect 17328 13394 17356 13466
rect 17316 13388 17368 13394
rect 17316 13330 17368 13336
rect 17420 13258 17448 13466
rect 17408 13252 17460 13258
rect 17408 13194 17460 13200
rect 17224 12980 17276 12986
rect 17224 12922 17276 12928
rect 17224 12844 17276 12850
rect 17224 12786 17276 12792
rect 17236 8294 17264 12786
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17328 12238 17356 12378
rect 17316 12232 17368 12238
rect 17316 12174 17368 12180
rect 17316 11212 17368 11218
rect 17316 11154 17368 11160
rect 17224 8288 17276 8294
rect 17224 8230 17276 8236
rect 17132 7744 17184 7750
rect 17132 7686 17184 7692
rect 17224 7200 17276 7206
rect 17224 7142 17276 7148
rect 17132 6996 17184 7002
rect 17132 6938 17184 6944
rect 17144 4214 17172 6938
rect 17236 6662 17264 7142
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17236 6202 17264 6598
rect 17328 6322 17356 11154
rect 17420 9382 17448 12582
rect 17512 11830 17540 13518
rect 17592 12368 17644 12374
rect 17592 12310 17644 12316
rect 17500 11824 17552 11830
rect 17500 11766 17552 11772
rect 17512 11218 17540 11766
rect 17500 11212 17552 11218
rect 17500 11154 17552 11160
rect 17604 10742 17632 12310
rect 17696 11558 17724 15642
rect 17684 11552 17736 11558
rect 17684 11494 17736 11500
rect 17684 11076 17736 11082
rect 17684 11018 17736 11024
rect 17592 10736 17644 10742
rect 17592 10678 17644 10684
rect 17696 10588 17724 11018
rect 17604 10560 17724 10588
rect 17788 10577 17816 15846
rect 17880 15706 17908 15966
rect 18236 15972 18288 15978
rect 18236 15914 18288 15920
rect 17868 15700 17920 15706
rect 17868 15642 17920 15648
rect 18248 15450 18276 15914
rect 18340 15570 18368 17682
rect 18432 16114 18460 24006
rect 18616 23186 18644 24822
rect 18696 24812 18748 24818
rect 18696 24754 18748 24760
rect 18708 23866 18736 24754
rect 18696 23860 18748 23866
rect 18696 23802 18748 23808
rect 18800 23338 18828 27950
rect 18984 26790 19012 28562
rect 18972 26784 19024 26790
rect 18972 26726 19024 26732
rect 18984 24274 19012 26726
rect 18972 24268 19024 24274
rect 18972 24210 19024 24216
rect 18880 24132 18932 24138
rect 18880 24074 18932 24080
rect 18892 23866 18920 24074
rect 18880 23860 18932 23866
rect 18880 23802 18932 23808
rect 18892 23497 18920 23802
rect 18878 23488 18934 23497
rect 18878 23423 18934 23432
rect 18800 23310 18920 23338
rect 18696 23248 18748 23254
rect 18696 23190 18748 23196
rect 18512 23180 18564 23186
rect 18512 23122 18564 23128
rect 18604 23180 18656 23186
rect 18604 23122 18656 23128
rect 18524 20398 18552 23122
rect 18604 22976 18656 22982
rect 18604 22918 18656 22924
rect 18616 22710 18644 22918
rect 18604 22704 18656 22710
rect 18604 22646 18656 22652
rect 18604 22568 18656 22574
rect 18604 22510 18656 22516
rect 18616 20942 18644 22510
rect 18604 20936 18656 20942
rect 18604 20878 18656 20884
rect 18512 20392 18564 20398
rect 18512 20334 18564 20340
rect 18512 19712 18564 19718
rect 18512 19654 18564 19660
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 18524 15994 18552 19654
rect 18708 17610 18736 23190
rect 18788 23180 18840 23186
rect 18788 23122 18840 23128
rect 18800 22098 18828 23122
rect 18788 22092 18840 22098
rect 18788 22034 18840 22040
rect 18788 20800 18840 20806
rect 18788 20742 18840 20748
rect 18800 20534 18828 20742
rect 18788 20528 18840 20534
rect 18788 20470 18840 20476
rect 18696 17604 18748 17610
rect 18696 17546 18748 17552
rect 18604 17264 18656 17270
rect 18892 17218 18920 23310
rect 18972 22772 19024 22778
rect 18972 22714 19024 22720
rect 18984 20806 19012 22714
rect 19076 21486 19104 28970
rect 19352 28558 19380 29650
rect 19444 29306 19472 29838
rect 19432 29300 19484 29306
rect 19432 29242 19484 29248
rect 19340 28552 19392 28558
rect 19340 28494 19392 28500
rect 19352 27146 19380 28494
rect 19524 28416 19576 28422
rect 19524 28358 19576 28364
rect 19708 28416 19760 28422
rect 19708 28358 19760 28364
rect 19260 27130 19472 27146
rect 19248 27124 19472 27130
rect 19300 27118 19472 27124
rect 19248 27066 19300 27072
rect 19444 26450 19472 27118
rect 19432 26444 19484 26450
rect 19432 26386 19484 26392
rect 19156 26036 19208 26042
rect 19156 25978 19208 25984
rect 19168 25702 19196 25978
rect 19156 25696 19208 25702
rect 19156 25638 19208 25644
rect 19156 25220 19208 25226
rect 19156 25162 19208 25168
rect 19168 23866 19196 25162
rect 19444 24818 19472 26386
rect 19432 24812 19484 24818
rect 19432 24754 19484 24760
rect 19444 24274 19472 24754
rect 19432 24268 19484 24274
rect 19432 24210 19484 24216
rect 19156 23860 19208 23866
rect 19156 23802 19208 23808
rect 19340 23656 19392 23662
rect 19340 23598 19392 23604
rect 19352 23526 19380 23598
rect 19156 23520 19208 23526
rect 19156 23462 19208 23468
rect 19248 23520 19300 23526
rect 19248 23462 19300 23468
rect 19340 23520 19392 23526
rect 19340 23462 19392 23468
rect 19168 22574 19196 23462
rect 19260 23118 19288 23462
rect 19248 23112 19300 23118
rect 19248 23054 19300 23060
rect 19248 22976 19300 22982
rect 19248 22918 19300 22924
rect 19156 22568 19208 22574
rect 19156 22510 19208 22516
rect 19154 22400 19210 22409
rect 19154 22335 19210 22344
rect 19168 21486 19196 22335
rect 19064 21480 19116 21486
rect 19064 21422 19116 21428
rect 19156 21480 19208 21486
rect 19156 21422 19208 21428
rect 19168 21350 19196 21422
rect 19156 21344 19208 21350
rect 19156 21286 19208 21292
rect 18972 20800 19024 20806
rect 18972 20742 19024 20748
rect 19260 20448 19288 22918
rect 19444 20602 19472 24210
rect 19536 22658 19564 28358
rect 19720 28218 19748 28358
rect 19708 28212 19760 28218
rect 19708 28154 19760 28160
rect 19708 24132 19760 24138
rect 19708 24074 19760 24080
rect 19720 23798 19748 24074
rect 19708 23792 19760 23798
rect 19708 23734 19760 23740
rect 19616 23724 19668 23730
rect 19616 23666 19668 23672
rect 19628 22778 19656 23666
rect 19708 23656 19760 23662
rect 19708 23598 19760 23604
rect 19720 23254 19748 23598
rect 19708 23248 19760 23254
rect 19708 23190 19760 23196
rect 19616 22772 19668 22778
rect 19616 22714 19668 22720
rect 19536 22630 19656 22658
rect 19524 22568 19576 22574
rect 19524 22510 19576 22516
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19536 20466 19564 22510
rect 18984 20420 19288 20448
rect 19524 20460 19576 20466
rect 18984 17338 19012 20420
rect 19524 20402 19576 20408
rect 19156 20324 19208 20330
rect 19156 20266 19208 20272
rect 19064 20256 19116 20262
rect 19064 20198 19116 20204
rect 18972 17332 19024 17338
rect 18972 17274 19024 17280
rect 18604 17206 18656 17212
rect 18432 15966 18552 15994
rect 18328 15564 18380 15570
rect 18328 15506 18380 15512
rect 18248 15422 18368 15450
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 18340 13530 18368 15422
rect 18328 13524 18380 13530
rect 18328 13466 18380 13472
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 17880 11200 17908 13330
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 18052 12912 18104 12918
rect 18052 12854 18104 12860
rect 18064 12646 18092 12854
rect 18052 12640 18104 12646
rect 18052 12582 18104 12588
rect 18432 12306 18460 15966
rect 18512 15904 18564 15910
rect 18512 15846 18564 15852
rect 18420 12300 18472 12306
rect 18420 12242 18472 12248
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 18432 11898 18460 12038
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 18236 11688 18288 11694
rect 18236 11630 18288 11636
rect 17960 11212 18012 11218
rect 17880 11172 17960 11200
rect 17960 11154 18012 11160
rect 18248 11014 18276 11630
rect 18524 11200 18552 15846
rect 18616 14074 18644 17206
rect 18708 17190 18920 17218
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18604 13388 18656 13394
rect 18604 13330 18656 13336
rect 18340 11172 18552 11200
rect 18236 11008 18288 11014
rect 18236 10950 18288 10956
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 18340 10724 18368 11172
rect 18512 11076 18564 11082
rect 18512 11018 18564 11024
rect 18248 10696 18368 10724
rect 17774 10568 17830 10577
rect 17604 9738 17632 10560
rect 17774 10503 17830 10512
rect 17788 10130 17816 10503
rect 17684 10124 17736 10130
rect 17684 10066 17736 10072
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 17696 9926 17724 10066
rect 18248 10010 18276 10696
rect 18420 10668 18472 10674
rect 18420 10610 18472 10616
rect 18328 10192 18380 10198
rect 18328 10134 18380 10140
rect 17880 9982 18276 10010
rect 17684 9920 17736 9926
rect 17684 9862 17736 9868
rect 17604 9710 17724 9738
rect 17592 9512 17644 9518
rect 17592 9454 17644 9460
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17408 9036 17460 9042
rect 17408 8978 17460 8984
rect 17420 8514 17448 8978
rect 17500 8832 17552 8838
rect 17500 8774 17552 8780
rect 17512 8634 17540 8774
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17420 8486 17540 8514
rect 17408 8424 17460 8430
rect 17408 8366 17460 8372
rect 17420 6730 17448 8366
rect 17512 7954 17540 8486
rect 17500 7948 17552 7954
rect 17500 7890 17552 7896
rect 17604 7342 17632 9454
rect 17696 8838 17724 9710
rect 17880 9654 17908 9982
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17868 9648 17920 9654
rect 17774 9616 17830 9625
rect 17920 9596 18000 9602
rect 17868 9590 18000 9596
rect 17880 9574 18000 9590
rect 17774 9551 17830 9560
rect 17684 8832 17736 8838
rect 17684 8774 17736 8780
rect 17696 8430 17724 8774
rect 17788 8537 17816 9551
rect 17972 9518 18000 9574
rect 17960 9512 18012 9518
rect 17960 9454 18012 9460
rect 17868 9104 17920 9110
rect 17868 9046 17920 9052
rect 17774 8528 17830 8537
rect 17774 8463 17776 8472
rect 17828 8463 17830 8472
rect 17776 8434 17828 8440
rect 17684 8424 17736 8430
rect 17684 8366 17736 8372
rect 17776 7812 17828 7818
rect 17776 7754 17828 7760
rect 17788 7546 17816 7754
rect 17880 7750 17908 9046
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 17960 8288 18012 8294
rect 17960 8230 18012 8236
rect 17972 7886 18000 8230
rect 17960 7880 18012 7886
rect 18248 7857 18276 8434
rect 17960 7822 18012 7828
rect 18234 7848 18290 7857
rect 18340 7818 18368 10134
rect 18432 8022 18460 10610
rect 18524 9178 18552 11018
rect 18512 9172 18564 9178
rect 18512 9114 18564 9120
rect 18512 9036 18564 9042
rect 18512 8978 18564 8984
rect 18420 8016 18472 8022
rect 18420 7958 18472 7964
rect 18234 7783 18290 7792
rect 18328 7812 18380 7818
rect 18328 7754 18380 7760
rect 17868 7744 17920 7750
rect 17868 7686 17920 7692
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 18524 7410 18552 8978
rect 17684 7404 17736 7410
rect 17684 7346 17736 7352
rect 18512 7404 18564 7410
rect 18512 7346 18564 7352
rect 17592 7336 17644 7342
rect 17592 7278 17644 7284
rect 17604 7177 17632 7278
rect 17590 7168 17646 7177
rect 17590 7103 17646 7112
rect 17696 7041 17724 7346
rect 18328 7268 18380 7274
rect 18328 7210 18380 7216
rect 17776 7200 17828 7206
rect 17776 7142 17828 7148
rect 17682 7032 17738 7041
rect 17682 6967 17738 6976
rect 17408 6724 17460 6730
rect 17408 6666 17460 6672
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17236 6174 17356 6202
rect 17224 5772 17276 5778
rect 17224 5714 17276 5720
rect 17236 4826 17264 5714
rect 17328 5710 17356 6174
rect 17420 5914 17448 6666
rect 17592 6112 17644 6118
rect 17592 6054 17644 6060
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17604 5710 17632 6054
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 17316 4752 17368 4758
rect 17316 4694 17368 4700
rect 17132 4208 17184 4214
rect 17132 4150 17184 4156
rect 17328 4049 17356 4694
rect 17408 4684 17460 4690
rect 17408 4626 17460 4632
rect 17500 4684 17552 4690
rect 17500 4626 17552 4632
rect 17420 4214 17448 4626
rect 17408 4208 17460 4214
rect 17408 4150 17460 4156
rect 17314 4040 17370 4049
rect 17314 3975 17370 3984
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 16948 2916 17000 2922
rect 16948 2858 17000 2864
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 16672 2372 16724 2378
rect 16672 2314 16724 2320
rect 16960 800 16988 2858
rect 17316 2848 17368 2854
rect 17316 2790 17368 2796
rect 17328 2514 17356 2790
rect 17316 2508 17368 2514
rect 17316 2450 17368 2456
rect 17512 2258 17540 4626
rect 17684 3596 17736 3602
rect 17684 3538 17736 3544
rect 17328 2230 17540 2258
rect 17328 800 17356 2230
rect 17696 800 17724 3538
rect 17788 2310 17816 7142
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 18340 6322 18368 7210
rect 18328 6316 18380 6322
rect 18328 6258 18380 6264
rect 18328 5568 18380 5574
rect 18328 5510 18380 5516
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 18144 5160 18196 5166
rect 18144 5102 18196 5108
rect 17960 5092 18012 5098
rect 17960 5034 18012 5040
rect 17972 4468 18000 5034
rect 18156 4486 18184 5102
rect 17880 4440 18000 4468
rect 18144 4480 18196 4486
rect 17880 4162 17908 4440
rect 18144 4422 18196 4428
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 18340 4282 18368 5510
rect 18524 5234 18552 7346
rect 18512 5228 18564 5234
rect 18512 5170 18564 5176
rect 18524 4690 18552 5170
rect 18512 4684 18564 4690
rect 18512 4626 18564 4632
rect 18328 4276 18380 4282
rect 18328 4218 18380 4224
rect 17880 4134 18000 4162
rect 17972 3738 18000 4134
rect 18328 4072 18380 4078
rect 18328 4014 18380 4020
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 17776 2304 17828 2310
rect 17776 2246 17828 2252
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18064 870 18184 898
rect 18064 800 18092 870
rect 7852 734 8064 762
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18156 762 18184 870
rect 18340 762 18368 4014
rect 18616 3058 18644 13330
rect 18708 9926 18736 17190
rect 18972 17128 19024 17134
rect 18972 17070 19024 17076
rect 18984 16794 19012 17070
rect 18972 16788 19024 16794
rect 18972 16730 19024 16736
rect 18880 14884 18932 14890
rect 18880 14826 18932 14832
rect 18788 14068 18840 14074
rect 18788 14010 18840 14016
rect 18800 12782 18828 14010
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 18892 12442 18920 14826
rect 18984 14074 19012 16730
rect 18972 14068 19024 14074
rect 18972 14010 19024 14016
rect 18972 13252 19024 13258
rect 18972 13194 19024 13200
rect 18880 12436 18932 12442
rect 18880 12378 18932 12384
rect 18984 12186 19012 13194
rect 18800 12158 19012 12186
rect 18696 9920 18748 9926
rect 18696 9862 18748 9868
rect 18708 9625 18736 9862
rect 18694 9616 18750 9625
rect 18694 9551 18750 9560
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18708 8906 18736 9114
rect 18696 8900 18748 8906
rect 18696 8842 18748 8848
rect 18800 7562 18828 12158
rect 18972 12096 19024 12102
rect 18972 12038 19024 12044
rect 18880 10464 18932 10470
rect 18880 10406 18932 10412
rect 18892 10305 18920 10406
rect 18878 10296 18934 10305
rect 18878 10231 18934 10240
rect 18880 10124 18932 10130
rect 18880 10066 18932 10072
rect 18708 7534 18828 7562
rect 18708 4146 18736 7534
rect 18788 7472 18840 7478
rect 18788 7414 18840 7420
rect 18800 4146 18828 7414
rect 18892 7342 18920 10066
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 18892 5370 18920 7278
rect 18880 5364 18932 5370
rect 18880 5306 18932 5312
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 18788 4140 18840 4146
rect 18788 4082 18840 4088
rect 18880 3460 18932 3466
rect 18880 3402 18932 3408
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18420 2848 18472 2854
rect 18420 2790 18472 2796
rect 18432 800 18460 2790
rect 18892 1714 18920 3402
rect 18984 3058 19012 12038
rect 19076 9994 19104 20198
rect 19168 19378 19196 20266
rect 19524 20256 19576 20262
rect 19524 20198 19576 20204
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 19156 19372 19208 19378
rect 19156 19314 19208 19320
rect 19156 18080 19208 18086
rect 19156 18022 19208 18028
rect 19168 15706 19196 18022
rect 19156 15700 19208 15706
rect 19156 15642 19208 15648
rect 19168 14226 19196 15642
rect 19260 15094 19288 19450
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19352 17678 19380 19246
rect 19340 17672 19392 17678
rect 19340 17614 19392 17620
rect 19340 16652 19392 16658
rect 19340 16594 19392 16600
rect 19352 16114 19380 16594
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 19248 15088 19300 15094
rect 19248 15030 19300 15036
rect 19168 14198 19288 14226
rect 19156 14068 19208 14074
rect 19156 14010 19208 14016
rect 19168 13190 19196 14010
rect 19260 14006 19288 14198
rect 19248 14000 19300 14006
rect 19248 13942 19300 13948
rect 19352 13326 19380 16050
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19340 13320 19392 13326
rect 19340 13262 19392 13268
rect 19156 13184 19208 13190
rect 19156 13126 19208 13132
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 19168 12306 19196 12786
rect 19248 12436 19300 12442
rect 19248 12378 19300 12384
rect 19156 12300 19208 12306
rect 19156 12242 19208 12248
rect 19260 10849 19288 12378
rect 19444 11830 19472 14962
rect 19536 12374 19564 20198
rect 19628 19854 19656 22630
rect 19720 22409 19748 23190
rect 19812 22574 19840 29990
rect 19996 29510 20024 30262
rect 20548 30190 20576 33390
rect 20640 31414 20668 34954
rect 20720 34740 20772 34746
rect 20720 34682 20772 34688
rect 20628 31408 20680 31414
rect 20628 31350 20680 31356
rect 20628 31272 20680 31278
rect 20628 31214 20680 31220
rect 20640 31142 20668 31214
rect 20628 31136 20680 31142
rect 20628 31078 20680 31084
rect 20260 30184 20312 30190
rect 20260 30126 20312 30132
rect 20536 30184 20588 30190
rect 20536 30126 20588 30132
rect 20272 29782 20300 30126
rect 20260 29776 20312 29782
rect 20260 29718 20312 29724
rect 20732 29578 20760 34682
rect 21100 34406 21128 43658
rect 22100 43648 22152 43654
rect 22100 43590 22152 43596
rect 21916 39296 21968 39302
rect 21916 39238 21968 39244
rect 21824 35692 21876 35698
rect 21824 35634 21876 35640
rect 21272 35624 21324 35630
rect 21272 35566 21324 35572
rect 21088 34400 21140 34406
rect 21088 34342 21140 34348
rect 21284 33946 21312 35566
rect 21836 34950 21864 35634
rect 21824 34944 21876 34950
rect 21744 34904 21824 34932
rect 21364 34400 21416 34406
rect 21364 34342 21416 34348
rect 21376 34202 21404 34342
rect 21364 34196 21416 34202
rect 21364 34138 21416 34144
rect 21192 33918 21312 33946
rect 21192 33862 21220 33918
rect 21180 33856 21232 33862
rect 21180 33798 21232 33804
rect 21272 33856 21324 33862
rect 21376 33810 21404 34138
rect 21324 33804 21404 33810
rect 21272 33798 21404 33804
rect 21192 32366 21220 33798
rect 21284 33782 21404 33798
rect 21284 33590 21312 33782
rect 21272 33584 21324 33590
rect 21272 33526 21324 33532
rect 21284 33318 21312 33526
rect 21272 33312 21324 33318
rect 21272 33254 21324 33260
rect 21284 32570 21312 33254
rect 21272 32564 21324 32570
rect 21272 32506 21324 32512
rect 21180 32360 21232 32366
rect 21180 32302 21232 32308
rect 20904 32224 20956 32230
rect 20904 32166 20956 32172
rect 20720 29572 20772 29578
rect 20720 29514 20772 29520
rect 19984 29504 20036 29510
rect 19984 29446 20036 29452
rect 19996 29306 20024 29446
rect 19984 29300 20036 29306
rect 19984 29242 20036 29248
rect 20168 29300 20220 29306
rect 20168 29242 20220 29248
rect 20076 27056 20128 27062
rect 20076 26998 20128 27004
rect 20088 26790 20116 26998
rect 20076 26784 20128 26790
rect 20076 26726 20128 26732
rect 19984 25764 20036 25770
rect 19984 25706 20036 25712
rect 19892 25152 19944 25158
rect 19892 25094 19944 25100
rect 19904 24993 19932 25094
rect 19890 24984 19946 24993
rect 19890 24919 19946 24928
rect 19996 23186 20024 25706
rect 20076 25492 20128 25498
rect 20076 25434 20128 25440
rect 19984 23180 20036 23186
rect 19984 23122 20036 23128
rect 19800 22568 19852 22574
rect 19800 22510 19852 22516
rect 19706 22400 19762 22409
rect 19706 22335 19762 22344
rect 20088 21894 20116 25434
rect 20180 23730 20208 29242
rect 20916 29102 20944 32166
rect 20996 31680 21048 31686
rect 20996 31622 21048 31628
rect 21008 30666 21036 31622
rect 21284 31482 21312 32506
rect 21744 31686 21772 34904
rect 21824 34886 21876 34892
rect 21824 32768 21876 32774
rect 21824 32710 21876 32716
rect 21836 32434 21864 32710
rect 21824 32428 21876 32434
rect 21824 32370 21876 32376
rect 21836 32230 21864 32370
rect 21824 32224 21876 32230
rect 21824 32166 21876 32172
rect 21640 31680 21692 31686
rect 21640 31622 21692 31628
rect 21732 31680 21784 31686
rect 21732 31622 21784 31628
rect 21272 31476 21324 31482
rect 21272 31418 21324 31424
rect 21284 30666 21312 31418
rect 21364 31408 21416 31414
rect 21364 31350 21416 31356
rect 20996 30660 21048 30666
rect 20996 30602 21048 30608
rect 21272 30660 21324 30666
rect 21272 30602 21324 30608
rect 20904 29096 20956 29102
rect 20904 29038 20956 29044
rect 20628 28552 20680 28558
rect 20628 28494 20680 28500
rect 20640 28150 20668 28494
rect 20916 28490 20944 29038
rect 21008 28626 21036 30602
rect 21088 28756 21140 28762
rect 21088 28698 21140 28704
rect 20996 28620 21048 28626
rect 20996 28562 21048 28568
rect 20904 28484 20956 28490
rect 20904 28426 20956 28432
rect 20628 28144 20680 28150
rect 20628 28086 20680 28092
rect 20720 27872 20772 27878
rect 20720 27814 20772 27820
rect 20444 24744 20496 24750
rect 20444 24686 20496 24692
rect 20456 24410 20484 24686
rect 20444 24404 20496 24410
rect 20444 24346 20496 24352
rect 20168 23724 20220 23730
rect 20168 23666 20220 23672
rect 20260 23520 20312 23526
rect 20260 23462 20312 23468
rect 20168 22568 20220 22574
rect 20168 22510 20220 22516
rect 19892 21888 19944 21894
rect 19892 21830 19944 21836
rect 20076 21888 20128 21894
rect 20076 21830 20128 21836
rect 19708 21004 19760 21010
rect 19708 20946 19760 20952
rect 19616 19848 19668 19854
rect 19616 19790 19668 19796
rect 19616 16448 19668 16454
rect 19616 16390 19668 16396
rect 19524 12368 19576 12374
rect 19524 12310 19576 12316
rect 19432 11824 19484 11830
rect 19338 11792 19394 11801
rect 19432 11766 19484 11772
rect 19338 11727 19340 11736
rect 19392 11727 19394 11736
rect 19340 11698 19392 11704
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19246 10840 19302 10849
rect 19246 10775 19302 10784
rect 19248 10668 19300 10674
rect 19248 10610 19300 10616
rect 19064 9988 19116 9994
rect 19064 9930 19116 9936
rect 19064 9512 19116 9518
rect 19064 9454 19116 9460
rect 19076 4826 19104 9454
rect 19156 9376 19208 9382
rect 19156 9318 19208 9324
rect 19168 9110 19196 9318
rect 19156 9104 19208 9110
rect 19156 9046 19208 9052
rect 19260 8945 19288 10610
rect 19444 10606 19472 11290
rect 19628 11200 19656 16390
rect 19720 15434 19748 20946
rect 19800 19780 19852 19786
rect 19800 19722 19852 19728
rect 19812 17746 19840 19722
rect 19800 17740 19852 17746
rect 19800 17682 19852 17688
rect 19800 16584 19852 16590
rect 19800 16526 19852 16532
rect 19812 15978 19840 16526
rect 19904 16046 19932 21830
rect 20088 21690 20116 21830
rect 20076 21684 20128 21690
rect 20076 21626 20128 21632
rect 20180 21486 20208 22510
rect 20168 21480 20220 21486
rect 20168 21422 20220 21428
rect 20076 21072 20128 21078
rect 20076 21014 20128 21020
rect 19892 16040 19944 16046
rect 19892 15982 19944 15988
rect 19800 15972 19852 15978
rect 19800 15914 19852 15920
rect 19708 15428 19760 15434
rect 19708 15370 19760 15376
rect 19720 12374 19748 15370
rect 20088 15162 20116 21014
rect 20180 19786 20208 21422
rect 20272 20874 20300 23462
rect 20456 23186 20484 24346
rect 20732 24070 20760 27814
rect 21100 26568 21128 28698
rect 21376 27282 21404 31350
rect 21456 28620 21508 28626
rect 21456 28562 21508 28568
rect 21468 28490 21496 28562
rect 21456 28484 21508 28490
rect 21456 28426 21508 28432
rect 21468 27402 21496 28426
rect 21652 28422 21680 31622
rect 21836 29034 21864 32166
rect 21928 31890 21956 39238
rect 22008 35488 22060 35494
rect 22008 35430 22060 35436
rect 21916 31884 21968 31890
rect 21916 31826 21968 31832
rect 22020 31754 22048 35430
rect 22112 32978 22140 43590
rect 22100 32972 22152 32978
rect 22100 32914 22152 32920
rect 22100 32224 22152 32230
rect 22100 32166 22152 32172
rect 22112 32026 22140 32166
rect 22100 32020 22152 32026
rect 22100 31962 22152 31968
rect 21928 31726 22048 31754
rect 21928 30326 21956 31726
rect 22008 31680 22060 31686
rect 22008 31622 22060 31628
rect 22020 31278 22048 31622
rect 22008 31272 22060 31278
rect 22008 31214 22060 31220
rect 22100 31272 22152 31278
rect 22100 31214 22152 31220
rect 21916 30320 21968 30326
rect 21916 30262 21968 30268
rect 21916 30048 21968 30054
rect 21916 29990 21968 29996
rect 21824 29028 21876 29034
rect 21824 28970 21876 28976
rect 21640 28416 21692 28422
rect 21640 28358 21692 28364
rect 21836 28082 21864 28970
rect 21824 28076 21876 28082
rect 21824 28018 21876 28024
rect 21456 27396 21508 27402
rect 21456 27338 21508 27344
rect 21824 27396 21876 27402
rect 21824 27338 21876 27344
rect 21640 27328 21692 27334
rect 21376 27254 21496 27282
rect 21640 27270 21692 27276
rect 20916 26540 21128 26568
rect 20720 24064 20772 24070
rect 20720 24006 20772 24012
rect 20812 23724 20864 23730
rect 20812 23666 20864 23672
rect 20628 23520 20680 23526
rect 20628 23462 20680 23468
rect 20444 23180 20496 23186
rect 20444 23122 20496 23128
rect 20444 22636 20496 22642
rect 20444 22578 20496 22584
rect 20456 22438 20484 22578
rect 20444 22432 20496 22438
rect 20442 22400 20444 22409
rect 20496 22400 20498 22409
rect 20442 22335 20498 22344
rect 20352 22092 20404 22098
rect 20352 22034 20404 22040
rect 20260 20868 20312 20874
rect 20260 20810 20312 20816
rect 20260 19916 20312 19922
rect 20260 19858 20312 19864
rect 20168 19780 20220 19786
rect 20168 19722 20220 19728
rect 20180 17338 20208 19722
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 20272 16658 20300 19858
rect 20260 16652 20312 16658
rect 20260 16594 20312 16600
rect 20272 16250 20300 16594
rect 20260 16244 20312 16250
rect 20260 16186 20312 16192
rect 20272 15570 20300 16186
rect 20364 16182 20392 22034
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20456 19514 20484 21286
rect 20640 19904 20668 23462
rect 20824 23186 20852 23666
rect 20916 23662 20944 26540
rect 20996 26444 21048 26450
rect 20996 26386 21048 26392
rect 21008 23662 21036 26386
rect 21088 26308 21140 26314
rect 21088 26250 21140 26256
rect 21100 24818 21128 26250
rect 21468 25906 21496 27254
rect 21652 26450 21680 27270
rect 21836 26790 21864 27338
rect 21824 26784 21876 26790
rect 21824 26726 21876 26732
rect 21640 26444 21692 26450
rect 21640 26386 21692 26392
rect 21836 26314 21864 26726
rect 21824 26308 21876 26314
rect 21824 26250 21876 26256
rect 21456 25900 21508 25906
rect 21456 25842 21508 25848
rect 21468 25702 21496 25842
rect 21456 25696 21508 25702
rect 21456 25638 21508 25644
rect 21088 24812 21140 24818
rect 21088 24754 21140 24760
rect 21100 24138 21128 24754
rect 21088 24132 21140 24138
rect 21088 24074 21140 24080
rect 20904 23656 20956 23662
rect 20904 23598 20956 23604
rect 20996 23656 21048 23662
rect 20996 23598 21048 23604
rect 20812 23180 20864 23186
rect 20812 23122 20864 23128
rect 20904 22704 20956 22710
rect 20904 22646 20956 22652
rect 20720 22432 20772 22438
rect 20720 22374 20772 22380
rect 20548 19876 20668 19904
rect 20444 19508 20496 19514
rect 20444 19450 20496 19456
rect 20548 19394 20576 19876
rect 20732 19514 20760 22374
rect 20916 21146 20944 22646
rect 21468 22642 21496 25638
rect 21548 24064 21600 24070
rect 21548 24006 21600 24012
rect 21560 23526 21588 24006
rect 21548 23520 21600 23526
rect 21548 23462 21600 23468
rect 21456 22636 21508 22642
rect 21456 22578 21508 22584
rect 21364 22024 21416 22030
rect 21364 21966 21416 21972
rect 21376 21690 21404 21966
rect 21560 21962 21588 23462
rect 21928 22094 21956 29990
rect 22112 28966 22140 31214
rect 22100 28960 22152 28966
rect 22100 28902 22152 28908
rect 22204 27554 22232 53926
rect 22468 35624 22520 35630
rect 22468 35566 22520 35572
rect 22376 35556 22428 35562
rect 22376 35498 22428 35504
rect 22284 34060 22336 34066
rect 22284 34002 22336 34008
rect 22296 33590 22324 34002
rect 22284 33584 22336 33590
rect 22284 33526 22336 33532
rect 22388 33538 22416 35498
rect 22480 33658 22508 35566
rect 22560 34944 22612 34950
rect 22560 34886 22612 34892
rect 22468 33652 22520 33658
rect 22468 33594 22520 33600
rect 22296 32978 22324 33526
rect 22388 33510 22508 33538
rect 22376 33448 22428 33454
rect 22376 33390 22428 33396
rect 22388 33114 22416 33390
rect 22376 33108 22428 33114
rect 22376 33050 22428 33056
rect 22284 32972 22336 32978
rect 22284 32914 22336 32920
rect 22296 32502 22324 32914
rect 22376 32768 22428 32774
rect 22376 32710 22428 32716
rect 22284 32496 22336 32502
rect 22284 32438 22336 32444
rect 22296 31346 22324 32438
rect 22284 31340 22336 31346
rect 22284 31282 22336 31288
rect 22388 30274 22416 32710
rect 22480 32026 22508 33510
rect 22468 32020 22520 32026
rect 22468 31962 22520 31968
rect 22468 31680 22520 31686
rect 22468 31622 22520 31628
rect 22296 30246 22416 30274
rect 22296 30190 22324 30246
rect 22284 30184 22336 30190
rect 22284 30126 22336 30132
rect 22480 30122 22508 31622
rect 22572 30326 22600 34886
rect 22664 31686 22692 53926
rect 22950 53884 23258 53893
rect 22950 53882 22956 53884
rect 23012 53882 23036 53884
rect 23092 53882 23116 53884
rect 23172 53882 23196 53884
rect 23252 53882 23258 53884
rect 23012 53830 23014 53882
rect 23194 53830 23196 53882
rect 22950 53828 22956 53830
rect 23012 53828 23036 53830
rect 23092 53828 23116 53830
rect 23172 53828 23196 53830
rect 23252 53828 23258 53830
rect 22950 53819 23258 53828
rect 23400 53582 23428 56063
rect 24504 54194 24532 56200
rect 24766 55448 24822 55457
rect 24766 55383 24822 55392
rect 24582 54632 24638 54641
rect 24582 54567 24638 54576
rect 24492 54188 24544 54194
rect 24492 54130 24544 54136
rect 24596 53786 24624 54567
rect 24676 53984 24728 53990
rect 24676 53926 24728 53932
rect 24584 53780 24636 53786
rect 24584 53722 24636 53728
rect 23388 53576 23440 53582
rect 23388 53518 23440 53524
rect 22836 53440 22888 53446
rect 22836 53382 22888 53388
rect 22744 33448 22796 33454
rect 22744 33390 22796 33396
rect 22756 32586 22784 33390
rect 22848 32774 22876 53382
rect 23400 53242 23428 53518
rect 23940 53440 23992 53446
rect 23940 53382 23992 53388
rect 23388 53236 23440 53242
rect 23388 53178 23440 53184
rect 22950 52796 23258 52805
rect 22950 52794 22956 52796
rect 23012 52794 23036 52796
rect 23092 52794 23116 52796
rect 23172 52794 23196 52796
rect 23252 52794 23258 52796
rect 23012 52742 23014 52794
rect 23194 52742 23196 52794
rect 22950 52740 22956 52742
rect 23012 52740 23036 52742
rect 23092 52740 23116 52742
rect 23172 52740 23196 52742
rect 23252 52740 23258 52742
rect 22950 52731 23258 52740
rect 22950 51708 23258 51717
rect 22950 51706 22956 51708
rect 23012 51706 23036 51708
rect 23092 51706 23116 51708
rect 23172 51706 23196 51708
rect 23252 51706 23258 51708
rect 23012 51654 23014 51706
rect 23194 51654 23196 51706
rect 22950 51652 22956 51654
rect 23012 51652 23036 51654
rect 23092 51652 23116 51654
rect 23172 51652 23196 51654
rect 23252 51652 23258 51654
rect 22950 51643 23258 51652
rect 22950 50620 23258 50629
rect 22950 50618 22956 50620
rect 23012 50618 23036 50620
rect 23092 50618 23116 50620
rect 23172 50618 23196 50620
rect 23252 50618 23258 50620
rect 23012 50566 23014 50618
rect 23194 50566 23196 50618
rect 22950 50564 22956 50566
rect 23012 50564 23036 50566
rect 23092 50564 23116 50566
rect 23172 50564 23196 50566
rect 23252 50564 23258 50566
rect 22950 50555 23258 50564
rect 23664 49768 23716 49774
rect 23664 49710 23716 49716
rect 22950 49532 23258 49541
rect 22950 49530 22956 49532
rect 23012 49530 23036 49532
rect 23092 49530 23116 49532
rect 23172 49530 23196 49532
rect 23252 49530 23258 49532
rect 23012 49478 23014 49530
rect 23194 49478 23196 49530
rect 22950 49476 22956 49478
rect 23012 49476 23036 49478
rect 23092 49476 23116 49478
rect 23172 49476 23196 49478
rect 23252 49476 23258 49478
rect 22950 49467 23258 49476
rect 22950 48444 23258 48453
rect 22950 48442 22956 48444
rect 23012 48442 23036 48444
rect 23092 48442 23116 48444
rect 23172 48442 23196 48444
rect 23252 48442 23258 48444
rect 23012 48390 23014 48442
rect 23194 48390 23196 48442
rect 22950 48388 22956 48390
rect 23012 48388 23036 48390
rect 23092 48388 23116 48390
rect 23172 48388 23196 48390
rect 23252 48388 23258 48390
rect 22950 48379 23258 48388
rect 22950 47356 23258 47365
rect 22950 47354 22956 47356
rect 23012 47354 23036 47356
rect 23092 47354 23116 47356
rect 23172 47354 23196 47356
rect 23252 47354 23258 47356
rect 23012 47302 23014 47354
rect 23194 47302 23196 47354
rect 22950 47300 22956 47302
rect 23012 47300 23036 47302
rect 23092 47300 23116 47302
rect 23172 47300 23196 47302
rect 23252 47300 23258 47302
rect 22950 47291 23258 47300
rect 22950 46268 23258 46277
rect 22950 46266 22956 46268
rect 23012 46266 23036 46268
rect 23092 46266 23116 46268
rect 23172 46266 23196 46268
rect 23252 46266 23258 46268
rect 23012 46214 23014 46266
rect 23194 46214 23196 46266
rect 22950 46212 22956 46214
rect 23012 46212 23036 46214
rect 23092 46212 23116 46214
rect 23172 46212 23196 46214
rect 23252 46212 23258 46214
rect 22950 46203 23258 46212
rect 22950 45180 23258 45189
rect 22950 45178 22956 45180
rect 23012 45178 23036 45180
rect 23092 45178 23116 45180
rect 23172 45178 23196 45180
rect 23252 45178 23258 45180
rect 23012 45126 23014 45178
rect 23194 45126 23196 45178
rect 22950 45124 22956 45126
rect 23012 45124 23036 45126
rect 23092 45124 23116 45126
rect 23172 45124 23196 45126
rect 23252 45124 23258 45126
rect 22950 45115 23258 45124
rect 22950 44092 23258 44101
rect 22950 44090 22956 44092
rect 23012 44090 23036 44092
rect 23092 44090 23116 44092
rect 23172 44090 23196 44092
rect 23252 44090 23258 44092
rect 23012 44038 23014 44090
rect 23194 44038 23196 44090
rect 22950 44036 22956 44038
rect 23012 44036 23036 44038
rect 23092 44036 23116 44038
rect 23172 44036 23196 44038
rect 23252 44036 23258 44038
rect 22950 44027 23258 44036
rect 22950 43004 23258 43013
rect 22950 43002 22956 43004
rect 23012 43002 23036 43004
rect 23092 43002 23116 43004
rect 23172 43002 23196 43004
rect 23252 43002 23258 43004
rect 23012 42950 23014 43002
rect 23194 42950 23196 43002
rect 22950 42948 22956 42950
rect 23012 42948 23036 42950
rect 23092 42948 23116 42950
rect 23172 42948 23196 42950
rect 23252 42948 23258 42950
rect 22950 42939 23258 42948
rect 22950 41916 23258 41925
rect 22950 41914 22956 41916
rect 23012 41914 23036 41916
rect 23092 41914 23116 41916
rect 23172 41914 23196 41916
rect 23252 41914 23258 41916
rect 23012 41862 23014 41914
rect 23194 41862 23196 41914
rect 22950 41860 22956 41862
rect 23012 41860 23036 41862
rect 23092 41860 23116 41862
rect 23172 41860 23196 41862
rect 23252 41860 23258 41862
rect 22950 41851 23258 41860
rect 22950 40828 23258 40837
rect 22950 40826 22956 40828
rect 23012 40826 23036 40828
rect 23092 40826 23116 40828
rect 23172 40826 23196 40828
rect 23252 40826 23258 40828
rect 23012 40774 23014 40826
rect 23194 40774 23196 40826
rect 22950 40772 22956 40774
rect 23012 40772 23036 40774
rect 23092 40772 23116 40774
rect 23172 40772 23196 40774
rect 23252 40772 23258 40774
rect 22950 40763 23258 40772
rect 23388 40180 23440 40186
rect 23388 40122 23440 40128
rect 22950 39740 23258 39749
rect 22950 39738 22956 39740
rect 23012 39738 23036 39740
rect 23092 39738 23116 39740
rect 23172 39738 23196 39740
rect 23252 39738 23258 39740
rect 23012 39686 23014 39738
rect 23194 39686 23196 39738
rect 22950 39684 22956 39686
rect 23012 39684 23036 39686
rect 23092 39684 23116 39686
rect 23172 39684 23196 39686
rect 23252 39684 23258 39686
rect 22950 39675 23258 39684
rect 22950 38652 23258 38661
rect 22950 38650 22956 38652
rect 23012 38650 23036 38652
rect 23092 38650 23116 38652
rect 23172 38650 23196 38652
rect 23252 38650 23258 38652
rect 23012 38598 23014 38650
rect 23194 38598 23196 38650
rect 22950 38596 22956 38598
rect 23012 38596 23036 38598
rect 23092 38596 23116 38598
rect 23172 38596 23196 38598
rect 23252 38596 23258 38598
rect 22950 38587 23258 38596
rect 22950 37564 23258 37573
rect 22950 37562 22956 37564
rect 23012 37562 23036 37564
rect 23092 37562 23116 37564
rect 23172 37562 23196 37564
rect 23252 37562 23258 37564
rect 23012 37510 23014 37562
rect 23194 37510 23196 37562
rect 22950 37508 22956 37510
rect 23012 37508 23036 37510
rect 23092 37508 23116 37510
rect 23172 37508 23196 37510
rect 23252 37508 23258 37510
rect 22950 37499 23258 37508
rect 22950 36476 23258 36485
rect 22950 36474 22956 36476
rect 23012 36474 23036 36476
rect 23092 36474 23116 36476
rect 23172 36474 23196 36476
rect 23252 36474 23258 36476
rect 23012 36422 23014 36474
rect 23194 36422 23196 36474
rect 22950 36420 22956 36422
rect 23012 36420 23036 36422
rect 23092 36420 23116 36422
rect 23172 36420 23196 36422
rect 23252 36420 23258 36422
rect 22950 36411 23258 36420
rect 22950 35388 23258 35397
rect 22950 35386 22956 35388
rect 23012 35386 23036 35388
rect 23092 35386 23116 35388
rect 23172 35386 23196 35388
rect 23252 35386 23258 35388
rect 23012 35334 23014 35386
rect 23194 35334 23196 35386
rect 22950 35332 22956 35334
rect 23012 35332 23036 35334
rect 23092 35332 23116 35334
rect 23172 35332 23196 35334
rect 23252 35332 23258 35334
rect 22950 35323 23258 35332
rect 23296 35148 23348 35154
rect 23296 35090 23348 35096
rect 22950 34300 23258 34309
rect 22950 34298 22956 34300
rect 23012 34298 23036 34300
rect 23092 34298 23116 34300
rect 23172 34298 23196 34300
rect 23252 34298 23258 34300
rect 23012 34246 23014 34298
rect 23194 34246 23196 34298
rect 22950 34244 22956 34246
rect 23012 34244 23036 34246
rect 23092 34244 23116 34246
rect 23172 34244 23196 34246
rect 23252 34244 23258 34246
rect 22950 34235 23258 34244
rect 22928 33856 22980 33862
rect 22928 33798 22980 33804
rect 23204 33856 23256 33862
rect 23204 33798 23256 33804
rect 22940 33454 22968 33798
rect 23216 33658 23244 33798
rect 23204 33652 23256 33658
rect 23204 33594 23256 33600
rect 22928 33448 22980 33454
rect 22928 33390 22980 33396
rect 22950 33212 23258 33221
rect 22950 33210 22956 33212
rect 23012 33210 23036 33212
rect 23092 33210 23116 33212
rect 23172 33210 23196 33212
rect 23252 33210 23258 33212
rect 23012 33158 23014 33210
rect 23194 33158 23196 33210
rect 22950 33156 22956 33158
rect 23012 33156 23036 33158
rect 23092 33156 23116 33158
rect 23172 33156 23196 33158
rect 23252 33156 23258 33158
rect 22950 33147 23258 33156
rect 23308 33114 23336 35090
rect 23296 33108 23348 33114
rect 23296 33050 23348 33056
rect 22836 32768 22888 32774
rect 22836 32710 22888 32716
rect 22756 32558 22876 32586
rect 22744 31952 22796 31958
rect 22744 31894 22796 31900
rect 22652 31680 22704 31686
rect 22652 31622 22704 31628
rect 22652 31408 22704 31414
rect 22652 31350 22704 31356
rect 22664 30938 22692 31350
rect 22652 30932 22704 30938
rect 22652 30874 22704 30880
rect 22652 30388 22704 30394
rect 22652 30330 22704 30336
rect 22560 30320 22612 30326
rect 22560 30262 22612 30268
rect 22468 30116 22520 30122
rect 22468 30058 22520 30064
rect 22664 29594 22692 30330
rect 22572 29566 22692 29594
rect 22468 28960 22520 28966
rect 22468 28902 22520 28908
rect 22480 28422 22508 28902
rect 22572 28694 22600 29566
rect 22652 29504 22704 29510
rect 22652 29446 22704 29452
rect 22560 28688 22612 28694
rect 22560 28630 22612 28636
rect 22468 28416 22520 28422
rect 22468 28358 22520 28364
rect 22376 27872 22428 27878
rect 22376 27814 22428 27820
rect 22204 27526 22324 27554
rect 22100 26920 22152 26926
rect 22100 26862 22152 26868
rect 22112 26586 22140 26862
rect 22192 26784 22244 26790
rect 22192 26726 22244 26732
rect 22100 26580 22152 26586
rect 22100 26522 22152 26528
rect 22204 24834 22232 26726
rect 22296 26042 22324 27526
rect 22388 27402 22416 27814
rect 22376 27396 22428 27402
rect 22376 27338 22428 27344
rect 22388 26602 22416 27338
rect 22480 26858 22508 28358
rect 22572 28150 22600 28630
rect 22560 28144 22612 28150
rect 22560 28086 22612 28092
rect 22560 28008 22612 28014
rect 22560 27950 22612 27956
rect 22572 26926 22600 27950
rect 22560 26920 22612 26926
rect 22560 26862 22612 26868
rect 22468 26852 22520 26858
rect 22468 26794 22520 26800
rect 22388 26574 22600 26602
rect 22468 26512 22520 26518
rect 22468 26454 22520 26460
rect 22376 26444 22428 26450
rect 22376 26386 22428 26392
rect 22284 26036 22336 26042
rect 22284 25978 22336 25984
rect 22112 24806 22232 24834
rect 22112 23066 22140 24806
rect 22388 24750 22416 26386
rect 22376 24744 22428 24750
rect 22296 24692 22376 24698
rect 22296 24686 22428 24692
rect 22192 24676 22244 24682
rect 22192 24618 22244 24624
rect 22296 24670 22416 24686
rect 22204 24274 22232 24618
rect 22192 24268 22244 24274
rect 22192 24210 22244 24216
rect 22204 23662 22232 24210
rect 22296 24138 22324 24670
rect 22376 24608 22428 24614
rect 22376 24550 22428 24556
rect 22284 24132 22336 24138
rect 22284 24074 22336 24080
rect 22284 23724 22336 23730
rect 22284 23666 22336 23672
rect 22192 23656 22244 23662
rect 22192 23598 22244 23604
rect 22020 23038 22140 23066
rect 22020 22522 22048 23038
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 22112 22642 22140 22918
rect 22100 22636 22152 22642
rect 22100 22578 22152 22584
rect 22020 22494 22140 22522
rect 21836 22066 21956 22094
rect 21548 21956 21600 21962
rect 21548 21898 21600 21904
rect 21364 21684 21416 21690
rect 21364 21626 21416 21632
rect 21088 21412 21140 21418
rect 21088 21354 21140 21360
rect 20904 21140 20956 21146
rect 20904 21082 20956 21088
rect 20916 20602 20944 21082
rect 20904 20596 20956 20602
rect 20904 20538 20956 20544
rect 21100 20534 21128 21354
rect 21560 21350 21588 21898
rect 21548 21344 21600 21350
rect 21548 21286 21600 21292
rect 21732 21344 21784 21350
rect 21732 21286 21784 21292
rect 21088 20528 21140 20534
rect 21088 20470 21140 20476
rect 21272 20256 21324 20262
rect 21272 20198 21324 20204
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 20456 19366 20576 19394
rect 20352 16176 20404 16182
rect 20352 16118 20404 16124
rect 20456 16114 20484 19366
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 20904 17536 20956 17542
rect 20904 17478 20956 17484
rect 20536 16516 20588 16522
rect 20536 16458 20588 16464
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 20548 15366 20576 16458
rect 20628 16176 20680 16182
rect 20628 16118 20680 16124
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20076 15156 20128 15162
rect 20076 15098 20128 15104
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 20180 14414 20208 15098
rect 20548 14958 20576 15302
rect 20536 14952 20588 14958
rect 20536 14894 20588 14900
rect 20352 14544 20404 14550
rect 20352 14486 20404 14492
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 19892 13864 19944 13870
rect 19892 13806 19944 13812
rect 19800 13456 19852 13462
rect 19800 13398 19852 13404
rect 19812 12986 19840 13398
rect 19800 12980 19852 12986
rect 19800 12922 19852 12928
rect 19708 12368 19760 12374
rect 19708 12310 19760 12316
rect 19720 11694 19748 12310
rect 19708 11688 19760 11694
rect 19708 11630 19760 11636
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 19536 11172 19656 11200
rect 19536 10713 19564 11172
rect 19616 11076 19668 11082
rect 19616 11018 19668 11024
rect 19522 10704 19578 10713
rect 19522 10639 19578 10648
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 19536 10305 19564 10639
rect 19522 10296 19578 10305
rect 19522 10231 19578 10240
rect 19524 10124 19576 10130
rect 19524 10066 19576 10072
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19246 8936 19302 8945
rect 19246 8871 19302 8880
rect 19248 8356 19300 8362
rect 19248 8298 19300 8304
rect 19156 7540 19208 7546
rect 19156 7482 19208 7488
rect 19168 6730 19196 7482
rect 19260 7342 19288 8298
rect 19248 7336 19300 7342
rect 19248 7278 19300 7284
rect 19248 7200 19300 7206
rect 19246 7168 19248 7177
rect 19300 7168 19302 7177
rect 19246 7103 19302 7112
rect 19246 7032 19302 7041
rect 19246 6967 19248 6976
rect 19300 6967 19302 6976
rect 19248 6938 19300 6944
rect 19156 6724 19208 6730
rect 19156 6666 19208 6672
rect 19352 6474 19380 9522
rect 19444 9382 19472 9590
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19432 8900 19484 8906
rect 19432 8842 19484 8848
rect 19168 6446 19380 6474
rect 19168 5302 19196 6446
rect 19248 6384 19300 6390
rect 19248 6326 19300 6332
rect 19156 5296 19208 5302
rect 19156 5238 19208 5244
rect 19064 4820 19116 4826
rect 19064 4762 19116 4768
rect 19260 3534 19288 6326
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 19352 2774 19380 5714
rect 19444 3534 19472 8842
rect 19536 4554 19564 10066
rect 19628 5710 19656 11018
rect 19616 5704 19668 5710
rect 19616 5646 19668 5652
rect 19524 4548 19576 4554
rect 19524 4490 19576 4496
rect 19616 4208 19668 4214
rect 19616 4150 19668 4156
rect 19524 4140 19576 4146
rect 19524 4082 19576 4088
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 18800 1686 18920 1714
rect 19168 2746 19380 2774
rect 18800 800 18828 1686
rect 19168 800 19196 2746
rect 19536 800 19564 4082
rect 19628 2650 19656 4150
rect 19616 2644 19668 2650
rect 19616 2586 19668 2592
rect 19720 2446 19748 11494
rect 19800 10192 19852 10198
rect 19800 10134 19852 10140
rect 19812 7886 19840 10134
rect 19904 7886 19932 13806
rect 20180 13274 20208 14350
rect 20260 14272 20312 14278
rect 20260 14214 20312 14220
rect 20088 13246 20208 13274
rect 20088 12442 20116 13246
rect 20168 13184 20220 13190
rect 20168 13126 20220 13132
rect 20180 12850 20208 13126
rect 20168 12844 20220 12850
rect 20168 12786 20220 12792
rect 20076 12436 20128 12442
rect 20076 12378 20128 12384
rect 19982 12336 20038 12345
rect 19982 12271 20038 12280
rect 19996 11830 20024 12271
rect 20088 12238 20116 12378
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 19984 11824 20036 11830
rect 19984 11766 20036 11772
rect 19984 11688 20036 11694
rect 19984 11630 20036 11636
rect 19996 11150 20024 11630
rect 19984 11144 20036 11150
rect 19984 11086 20036 11092
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 20168 10600 20220 10606
rect 20168 10542 20220 10548
rect 19996 10198 20024 10542
rect 19984 10192 20036 10198
rect 19984 10134 20036 10140
rect 20180 10033 20208 10542
rect 20166 10024 20222 10033
rect 20166 9959 20222 9968
rect 19984 8900 20036 8906
rect 19984 8842 20036 8848
rect 19800 7880 19852 7886
rect 19800 7822 19852 7828
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 19996 7290 20024 8842
rect 20272 8634 20300 14214
rect 20364 13938 20392 14486
rect 20352 13932 20404 13938
rect 20352 13874 20404 13880
rect 20444 13252 20496 13258
rect 20444 13194 20496 13200
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20364 10538 20392 12786
rect 20456 12306 20484 13194
rect 20640 12782 20668 16118
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 20628 12776 20680 12782
rect 20628 12718 20680 12724
rect 20732 12628 20760 14758
rect 20824 12714 20852 16050
rect 20916 14346 20944 17478
rect 21008 17270 21036 19110
rect 20996 17264 21048 17270
rect 20996 17206 21048 17212
rect 21008 16794 21036 17206
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 21008 16522 21036 16730
rect 20996 16516 21048 16522
rect 20996 16458 21048 16464
rect 21088 15428 21140 15434
rect 21088 15370 21140 15376
rect 21100 15094 21128 15370
rect 21088 15088 21140 15094
rect 21088 15030 21140 15036
rect 21284 14482 21312 20198
rect 21560 19854 21588 21286
rect 21548 19848 21600 19854
rect 21548 19790 21600 19796
rect 21640 19712 21692 19718
rect 21640 19654 21692 19660
rect 21548 19440 21600 19446
rect 21548 19382 21600 19388
rect 21560 18766 21588 19382
rect 21652 19310 21680 19654
rect 21640 19304 21692 19310
rect 21640 19246 21692 19252
rect 21548 18760 21600 18766
rect 21548 18702 21600 18708
rect 21364 18624 21416 18630
rect 21364 18566 21416 18572
rect 21272 14476 21324 14482
rect 21272 14418 21324 14424
rect 20904 14340 20956 14346
rect 20904 14282 20956 14288
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 20904 13456 20956 13462
rect 20904 13398 20956 13404
rect 20812 12708 20864 12714
rect 20812 12650 20864 12656
rect 20640 12600 20760 12628
rect 20444 12300 20496 12306
rect 20444 12242 20496 12248
rect 20352 10532 20404 10538
rect 20352 10474 20404 10480
rect 20456 9450 20484 12242
rect 20640 10810 20668 12600
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20628 10804 20680 10810
rect 20628 10746 20680 10752
rect 20640 10713 20668 10746
rect 20626 10704 20682 10713
rect 20626 10639 20682 10648
rect 20626 9480 20682 9489
rect 20444 9444 20496 9450
rect 20626 9415 20682 9424
rect 20444 9386 20496 9392
rect 20352 9376 20404 9382
rect 20352 9318 20404 9324
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 20076 8492 20128 8498
rect 20076 8434 20128 8440
rect 19904 7274 20024 7290
rect 19892 7268 20024 7274
rect 19944 7262 20024 7268
rect 19892 7210 19944 7216
rect 19904 6866 19932 7210
rect 19892 6860 19944 6866
rect 19892 6802 19944 6808
rect 19984 6860 20036 6866
rect 19984 6802 20036 6808
rect 19892 6656 19944 6662
rect 19892 6598 19944 6604
rect 19904 6322 19932 6598
rect 19892 6316 19944 6322
rect 19892 6258 19944 6264
rect 19996 4808 20024 6802
rect 19812 4780 20024 4808
rect 19812 4690 19840 4780
rect 19800 4684 19852 4690
rect 19800 4626 19852 4632
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 19904 2774 19932 4626
rect 20088 2990 20116 8434
rect 20364 8022 20392 9318
rect 20456 9042 20484 9386
rect 20444 9036 20496 9042
rect 20444 8978 20496 8984
rect 20640 8838 20668 9415
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20536 8424 20588 8430
rect 20536 8366 20588 8372
rect 20352 8016 20404 8022
rect 20352 7958 20404 7964
rect 20260 7948 20312 7954
rect 20260 7890 20312 7896
rect 20168 7880 20220 7886
rect 20168 7822 20220 7828
rect 20180 3942 20208 7822
rect 20272 7546 20300 7890
rect 20260 7540 20312 7546
rect 20260 7482 20312 7488
rect 20364 7478 20392 7958
rect 20352 7472 20404 7478
rect 20352 7414 20404 7420
rect 20364 6798 20392 7414
rect 20352 6792 20404 6798
rect 20352 6734 20404 6740
rect 20260 6316 20312 6322
rect 20260 6258 20312 6264
rect 20272 5914 20300 6258
rect 20260 5908 20312 5914
rect 20260 5850 20312 5856
rect 20272 5358 20484 5386
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 20076 2984 20128 2990
rect 20076 2926 20128 2932
rect 19812 2746 19932 2774
rect 19708 2440 19760 2446
rect 19708 2382 19760 2388
rect 19812 1442 19840 2746
rect 19812 1414 19932 1442
rect 19904 800 19932 1414
rect 20272 800 20300 5358
rect 20456 5302 20484 5358
rect 20352 5296 20404 5302
rect 20352 5238 20404 5244
rect 20444 5296 20496 5302
rect 20444 5238 20496 5244
rect 20364 4554 20392 5238
rect 20444 5024 20496 5030
rect 20444 4966 20496 4972
rect 20352 4548 20404 4554
rect 20352 4490 20404 4496
rect 20364 4282 20392 4490
rect 20352 4276 20404 4282
rect 20352 4218 20404 4224
rect 20456 3194 20484 4966
rect 20548 4078 20576 8366
rect 20628 6180 20680 6186
rect 20628 6122 20680 6128
rect 20640 5846 20668 6122
rect 20732 5930 20760 11494
rect 20812 11144 20864 11150
rect 20812 11086 20864 11092
rect 20824 10130 20852 11086
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 20824 8838 20852 10066
rect 20812 8832 20864 8838
rect 20812 8774 20864 8780
rect 20812 7744 20864 7750
rect 20812 7686 20864 7692
rect 20824 6458 20852 7686
rect 20916 6798 20944 13398
rect 21100 13394 21128 14010
rect 21180 13524 21232 13530
rect 21180 13466 21232 13472
rect 20996 13388 21048 13394
rect 20996 13330 21048 13336
rect 21088 13388 21140 13394
rect 21088 13330 21140 13336
rect 21008 13274 21036 13330
rect 21008 13246 21128 13274
rect 20996 12096 21048 12102
rect 20996 12038 21048 12044
rect 21008 10266 21036 12038
rect 21100 11150 21128 13246
rect 21192 12986 21220 13466
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 21376 12434 21404 18566
rect 21548 18080 21600 18086
rect 21548 18022 21600 18028
rect 21456 15904 21508 15910
rect 21456 15846 21508 15852
rect 21468 15706 21496 15846
rect 21456 15700 21508 15706
rect 21456 15642 21508 15648
rect 21192 12406 21404 12434
rect 21088 11144 21140 11150
rect 21088 11086 21140 11092
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 20996 10260 21048 10266
rect 20996 10202 21048 10208
rect 21100 9722 21128 10610
rect 21192 9926 21220 12406
rect 21272 12300 21324 12306
rect 21272 12242 21324 12248
rect 21284 10606 21312 12242
rect 21364 11280 21416 11286
rect 21364 11222 21416 11228
rect 21376 10742 21404 11222
rect 21364 10736 21416 10742
rect 21364 10678 21416 10684
rect 21272 10600 21324 10606
rect 21272 10542 21324 10548
rect 21284 10441 21312 10542
rect 21364 10464 21416 10470
rect 21270 10432 21326 10441
rect 21364 10406 21416 10412
rect 21270 10367 21326 10376
rect 21180 9920 21232 9926
rect 21180 9862 21232 9868
rect 20996 9716 21048 9722
rect 20996 9658 21048 9664
rect 21088 9716 21140 9722
rect 21088 9658 21140 9664
rect 21008 7478 21036 9658
rect 21272 8628 21324 8634
rect 21272 8570 21324 8576
rect 21088 7812 21140 7818
rect 21088 7754 21140 7760
rect 20996 7472 21048 7478
rect 20996 7414 21048 7420
rect 20904 6792 20956 6798
rect 20904 6734 20956 6740
rect 20996 6724 21048 6730
rect 20996 6666 21048 6672
rect 20812 6452 20864 6458
rect 20812 6394 20864 6400
rect 20732 5902 20852 5930
rect 20628 5840 20680 5846
rect 20628 5782 20680 5788
rect 20720 5772 20772 5778
rect 20720 5714 20772 5720
rect 20536 4072 20588 4078
rect 20536 4014 20588 4020
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 20444 3188 20496 3194
rect 20444 3130 20496 3136
rect 20352 2916 20404 2922
rect 20352 2858 20404 2864
rect 20364 2446 20392 2858
rect 20548 2514 20576 3878
rect 20732 2774 20760 5714
rect 20824 3534 20852 5902
rect 21008 4146 21036 6666
rect 21100 5710 21128 7754
rect 21180 7472 21232 7478
rect 21180 7414 21232 7420
rect 21192 6934 21220 7414
rect 21180 6928 21232 6934
rect 21180 6870 21232 6876
rect 21180 6656 21232 6662
rect 21180 6598 21232 6604
rect 21088 5704 21140 5710
rect 21088 5646 21140 5652
rect 21192 5370 21220 6598
rect 21180 5364 21232 5370
rect 21180 5306 21232 5312
rect 21088 5228 21140 5234
rect 21088 5170 21140 5176
rect 21100 4826 21128 5170
rect 21180 5160 21232 5166
rect 21180 5102 21232 5108
rect 21192 4826 21220 5102
rect 21088 4820 21140 4826
rect 21088 4762 21140 4768
rect 21180 4820 21232 4826
rect 21180 4762 21232 4768
rect 20904 4140 20956 4146
rect 20904 4082 20956 4088
rect 20996 4140 21048 4146
rect 20996 4082 21048 4088
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 20812 3392 20864 3398
rect 20812 3334 20864 3340
rect 20824 3058 20852 3334
rect 20916 3194 20944 4082
rect 21192 4078 21220 4762
rect 21180 4072 21232 4078
rect 21180 4014 21232 4020
rect 20996 4004 21048 4010
rect 20996 3946 21048 3952
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 20812 3052 20864 3058
rect 20812 2994 20864 3000
rect 20640 2746 20760 2774
rect 20536 2508 20588 2514
rect 20536 2450 20588 2456
rect 20352 2440 20404 2446
rect 20352 2382 20404 2388
rect 20640 800 20668 2746
rect 21008 800 21036 3946
rect 21284 3398 21312 8570
rect 21376 6662 21404 10406
rect 21560 9178 21588 18022
rect 21744 14414 21772 21286
rect 21836 20466 21864 22066
rect 22008 21548 22060 21554
rect 22008 21490 22060 21496
rect 22020 21010 22048 21490
rect 22008 21004 22060 21010
rect 22008 20946 22060 20952
rect 21824 20460 21876 20466
rect 21824 20402 21876 20408
rect 22112 19938 22140 22494
rect 22204 22098 22232 23598
rect 22296 22506 22324 23666
rect 22284 22500 22336 22506
rect 22284 22442 22336 22448
rect 22192 22092 22244 22098
rect 22192 22034 22244 22040
rect 22204 21622 22232 22034
rect 22192 21616 22244 21622
rect 22192 21558 22244 21564
rect 22192 20460 22244 20466
rect 22192 20402 22244 20408
rect 22204 20058 22232 20402
rect 22192 20052 22244 20058
rect 22192 19994 22244 20000
rect 22112 19910 22232 19938
rect 21824 19848 21876 19854
rect 21824 19790 21876 19796
rect 21836 19718 21864 19790
rect 21824 19712 21876 19718
rect 21824 19654 21876 19660
rect 21836 19174 21864 19654
rect 21824 19168 21876 19174
rect 21824 19110 21876 19116
rect 22100 18624 22152 18630
rect 22100 18566 22152 18572
rect 22112 18290 22140 18566
rect 22204 18358 22232 19910
rect 22192 18352 22244 18358
rect 22192 18294 22244 18300
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 22388 18170 22416 24550
rect 22480 21690 22508 26454
rect 22572 25922 22600 26574
rect 22664 26042 22692 29446
rect 22756 27130 22784 31894
rect 22848 30190 22876 32558
rect 22950 32124 23258 32133
rect 22950 32122 22956 32124
rect 23012 32122 23036 32124
rect 23092 32122 23116 32124
rect 23172 32122 23196 32124
rect 23252 32122 23258 32124
rect 23012 32070 23014 32122
rect 23194 32070 23196 32122
rect 22950 32068 22956 32070
rect 23012 32068 23036 32070
rect 23092 32068 23116 32070
rect 23172 32068 23196 32070
rect 23252 32068 23258 32070
rect 22950 32059 23258 32068
rect 23204 32020 23256 32026
rect 23204 31962 23256 31968
rect 23020 31816 23072 31822
rect 23020 31758 23072 31764
rect 23032 31414 23060 31758
rect 23216 31754 23244 31962
rect 23400 31958 23428 40122
rect 23572 33992 23624 33998
rect 23572 33934 23624 33940
rect 23584 33590 23612 33934
rect 23572 33584 23624 33590
rect 23572 33526 23624 33532
rect 23584 32842 23612 33526
rect 23572 32836 23624 32842
rect 23572 32778 23624 32784
rect 23584 32570 23612 32778
rect 23572 32564 23624 32570
rect 23572 32506 23624 32512
rect 23388 31952 23440 31958
rect 23388 31894 23440 31900
rect 23204 31748 23256 31754
rect 23204 31690 23256 31696
rect 23020 31408 23072 31414
rect 23020 31350 23072 31356
rect 23216 31226 23244 31690
rect 23584 31482 23612 32506
rect 23676 31754 23704 49710
rect 23952 34474 23980 53382
rect 24492 52896 24544 52902
rect 24492 52838 24544 52844
rect 24504 52698 24532 52838
rect 24492 52692 24544 52698
rect 24492 52634 24544 52640
rect 24688 41414 24716 53926
rect 24780 53786 24808 55383
rect 25044 54052 25096 54058
rect 25044 53994 25096 54000
rect 25056 53825 25084 53994
rect 25136 53984 25188 53990
rect 25136 53926 25188 53932
rect 25042 53816 25098 53825
rect 24768 53780 24820 53786
rect 25042 53751 25098 53760
rect 24768 53722 24820 53728
rect 24780 53106 24808 53722
rect 25056 53582 25084 53751
rect 25044 53576 25096 53582
rect 25044 53518 25096 53524
rect 25148 53394 25176 53926
rect 25056 53366 25176 53394
rect 25056 53106 25084 53366
rect 24768 53100 24820 53106
rect 24768 53042 24820 53048
rect 25044 53100 25096 53106
rect 25044 53042 25096 53048
rect 25056 53009 25084 53042
rect 25042 53000 25098 53009
rect 25042 52935 25098 52944
rect 24952 52420 25004 52426
rect 24952 52362 25004 52368
rect 24964 52193 24992 52362
rect 24950 52184 25006 52193
rect 24950 52119 25006 52128
rect 25884 52018 25912 56200
rect 26516 53440 26568 53446
rect 26516 53382 26568 53388
rect 25872 52012 25924 52018
rect 25872 51954 25924 51960
rect 24860 51808 24912 51814
rect 24860 51750 24912 51756
rect 24872 45914 24900 51750
rect 24950 51368 25006 51377
rect 24950 51303 24952 51312
rect 25004 51303 25006 51312
rect 24952 51274 25004 51280
rect 24952 50924 25004 50930
rect 24952 50866 25004 50872
rect 24964 50561 24992 50866
rect 25044 50720 25096 50726
rect 25044 50662 25096 50668
rect 24950 50552 25006 50561
rect 25056 50522 25084 50662
rect 24950 50487 25006 50496
rect 25044 50516 25096 50522
rect 25044 50458 25096 50464
rect 25504 50176 25556 50182
rect 25504 50118 25556 50124
rect 25516 49842 25544 50118
rect 25504 49836 25556 49842
rect 25504 49778 25556 49784
rect 25516 49745 25544 49778
rect 25502 49736 25558 49745
rect 25502 49671 25558 49680
rect 25136 49156 25188 49162
rect 25136 49098 25188 49104
rect 25148 48929 25176 49098
rect 25228 49088 25280 49094
rect 25228 49030 25280 49036
rect 25134 48920 25190 48929
rect 25134 48855 25190 48864
rect 25136 48544 25188 48550
rect 25136 48486 25188 48492
rect 25148 48142 25176 48486
rect 25136 48136 25188 48142
rect 25134 48104 25136 48113
rect 25188 48104 25190 48113
rect 25134 48039 25190 48048
rect 24872 45886 24992 45914
rect 24860 45824 24912 45830
rect 24860 45766 24912 45772
rect 24768 44396 24820 44402
rect 24768 44338 24820 44344
rect 24780 44033 24808 44338
rect 24766 44024 24822 44033
rect 24766 43959 24822 43968
rect 24504 41386 24716 41414
rect 23940 34468 23992 34474
rect 23940 34410 23992 34416
rect 24504 32774 24532 41386
rect 24872 35834 24900 45766
rect 24964 43994 24992 45886
rect 25044 44736 25096 44742
rect 25044 44678 25096 44684
rect 24952 43988 25004 43994
rect 24952 43930 25004 43936
rect 25056 38298 25084 44678
rect 25136 42628 25188 42634
rect 25136 42570 25188 42576
rect 25148 42401 25176 42570
rect 25134 42392 25190 42401
rect 25134 42327 25190 42336
rect 25136 42016 25188 42022
rect 25136 41958 25188 41964
rect 25148 41614 25176 41958
rect 25136 41608 25188 41614
rect 25134 41576 25136 41585
rect 25188 41576 25190 41585
rect 25134 41511 25190 41520
rect 24964 38270 25084 38298
rect 24860 35828 24912 35834
rect 24860 35770 24912 35776
rect 24964 35086 24992 38270
rect 25044 38208 25096 38214
rect 25044 38150 25096 38156
rect 24952 35080 25004 35086
rect 24952 35022 25004 35028
rect 25056 34932 25084 38150
rect 25136 37868 25188 37874
rect 25136 37810 25188 37816
rect 25148 37505 25176 37810
rect 25134 37496 25190 37505
rect 25134 37431 25190 37440
rect 25056 34904 25176 34932
rect 24584 33312 24636 33318
rect 24584 33254 24636 33260
rect 24596 32910 24624 33254
rect 24952 33040 25004 33046
rect 24952 32982 25004 32988
rect 24584 32904 24636 32910
rect 24584 32846 24636 32852
rect 24768 32904 24820 32910
rect 24768 32846 24820 32852
rect 24492 32768 24544 32774
rect 24492 32710 24544 32716
rect 24584 32768 24636 32774
rect 24584 32710 24636 32716
rect 23676 31726 23888 31754
rect 23572 31476 23624 31482
rect 23572 31418 23624 31424
rect 23216 31198 23336 31226
rect 22950 31036 23258 31045
rect 22950 31034 22956 31036
rect 23012 31034 23036 31036
rect 23092 31034 23116 31036
rect 23172 31034 23196 31036
rect 23252 31034 23258 31036
rect 23012 30982 23014 31034
rect 23194 30982 23196 31034
rect 22950 30980 22956 30982
rect 23012 30980 23036 30982
rect 23092 30980 23116 30982
rect 23172 30980 23196 30982
rect 23252 30980 23258 30982
rect 22950 30971 23258 30980
rect 22928 30592 22980 30598
rect 22928 30534 22980 30540
rect 22836 30184 22888 30190
rect 22836 30126 22888 30132
rect 22940 30036 22968 30534
rect 23308 30394 23336 31198
rect 23756 31204 23808 31210
rect 23756 31146 23808 31152
rect 23768 31090 23796 31146
rect 23676 31062 23796 31090
rect 23296 30388 23348 30394
rect 23296 30330 23348 30336
rect 23676 30190 23704 31062
rect 23296 30184 23348 30190
rect 23296 30126 23348 30132
rect 23664 30184 23716 30190
rect 23664 30126 23716 30132
rect 22848 30008 22968 30036
rect 22848 27554 22876 30008
rect 22950 29948 23258 29957
rect 22950 29946 22956 29948
rect 23012 29946 23036 29948
rect 23092 29946 23116 29948
rect 23172 29946 23196 29948
rect 23252 29946 23258 29948
rect 23012 29894 23014 29946
rect 23194 29894 23196 29946
rect 22950 29892 22956 29894
rect 23012 29892 23036 29894
rect 23092 29892 23116 29894
rect 23172 29892 23196 29894
rect 23252 29892 23258 29894
rect 22950 29883 23258 29892
rect 23204 29776 23256 29782
rect 23204 29718 23256 29724
rect 23216 29016 23244 29718
rect 23308 29186 23336 30126
rect 23308 29158 23428 29186
rect 23400 29102 23428 29158
rect 23388 29096 23440 29102
rect 23388 29038 23440 29044
rect 23216 28988 23336 29016
rect 22950 28860 23258 28869
rect 22950 28858 22956 28860
rect 23012 28858 23036 28860
rect 23092 28858 23116 28860
rect 23172 28858 23196 28860
rect 23252 28858 23258 28860
rect 23012 28806 23014 28858
rect 23194 28806 23196 28858
rect 22950 28804 22956 28806
rect 23012 28804 23036 28806
rect 23092 28804 23116 28806
rect 23172 28804 23196 28806
rect 23252 28804 23258 28806
rect 22950 28795 23258 28804
rect 22950 27772 23258 27781
rect 22950 27770 22956 27772
rect 23012 27770 23036 27772
rect 23092 27770 23116 27772
rect 23172 27770 23196 27772
rect 23252 27770 23258 27772
rect 23012 27718 23014 27770
rect 23194 27718 23196 27770
rect 22950 27716 22956 27718
rect 23012 27716 23036 27718
rect 23092 27716 23116 27718
rect 23172 27716 23196 27718
rect 23252 27716 23258 27718
rect 22950 27707 23258 27716
rect 22848 27526 22968 27554
rect 22744 27124 22796 27130
rect 22744 27066 22796 27072
rect 22940 26994 22968 27526
rect 22928 26988 22980 26994
rect 22928 26930 22980 26936
rect 22836 26852 22888 26858
rect 22836 26794 22888 26800
rect 22848 26314 22876 26794
rect 22950 26684 23258 26693
rect 22950 26682 22956 26684
rect 23012 26682 23036 26684
rect 23092 26682 23116 26684
rect 23172 26682 23196 26684
rect 23252 26682 23258 26684
rect 23012 26630 23014 26682
rect 23194 26630 23196 26682
rect 22950 26628 22956 26630
rect 23012 26628 23036 26630
rect 23092 26628 23116 26630
rect 23172 26628 23196 26630
rect 23252 26628 23258 26630
rect 22950 26619 23258 26628
rect 23308 26382 23336 28988
rect 23400 28150 23428 29038
rect 23572 28620 23624 28626
rect 23572 28562 23624 28568
rect 23388 28144 23440 28150
rect 23388 28086 23440 28092
rect 23400 27538 23428 28086
rect 23480 28008 23532 28014
rect 23480 27950 23532 27956
rect 23492 27606 23520 27950
rect 23584 27674 23612 28562
rect 23572 27668 23624 27674
rect 23572 27610 23624 27616
rect 23480 27600 23532 27606
rect 23480 27542 23532 27548
rect 23388 27532 23440 27538
rect 23388 27474 23440 27480
rect 23400 26926 23428 27474
rect 23676 27130 23704 30126
rect 23664 27124 23716 27130
rect 23664 27066 23716 27072
rect 23388 26920 23440 26926
rect 23388 26862 23440 26868
rect 23296 26376 23348 26382
rect 23296 26318 23348 26324
rect 22836 26308 22888 26314
rect 22836 26250 22888 26256
rect 22652 26036 22704 26042
rect 22652 25978 22704 25984
rect 22572 25894 22692 25922
rect 22560 25832 22612 25838
rect 22560 25774 22612 25780
rect 22572 23798 22600 25774
rect 22664 24750 22692 25894
rect 22652 24744 22704 24750
rect 22652 24686 22704 24692
rect 22848 24290 22876 26250
rect 23296 25696 23348 25702
rect 23296 25638 23348 25644
rect 22950 25596 23258 25605
rect 22950 25594 22956 25596
rect 23012 25594 23036 25596
rect 23092 25594 23116 25596
rect 23172 25594 23196 25596
rect 23252 25594 23258 25596
rect 23012 25542 23014 25594
rect 23194 25542 23196 25594
rect 22950 25540 22956 25542
rect 23012 25540 23036 25542
rect 23092 25540 23116 25542
rect 23172 25540 23196 25542
rect 23252 25540 23258 25542
rect 22950 25531 23258 25540
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 22664 24262 22876 24290
rect 22560 23792 22612 23798
rect 22560 23734 22612 23740
rect 22560 22976 22612 22982
rect 22560 22918 22612 22924
rect 22468 21684 22520 21690
rect 22468 21626 22520 21632
rect 22572 19514 22600 22918
rect 22664 21690 22692 24262
rect 23308 23882 23336 25638
rect 23400 24682 23428 26862
rect 23480 26308 23532 26314
rect 23480 26250 23532 26256
rect 23492 24818 23520 26250
rect 23860 25378 23888 31726
rect 24492 29640 24544 29646
rect 24492 29582 24544 29588
rect 24504 29510 24532 29582
rect 24308 29504 24360 29510
rect 24308 29446 24360 29452
rect 24492 29504 24544 29510
rect 24492 29446 24544 29452
rect 24124 29300 24176 29306
rect 24124 29242 24176 29248
rect 23940 28552 23992 28558
rect 23940 28494 23992 28500
rect 23952 28150 23980 28494
rect 23940 28144 23992 28150
rect 23940 28086 23992 28092
rect 23952 28014 23980 28086
rect 23940 28008 23992 28014
rect 23940 27950 23992 27956
rect 23952 27470 23980 27950
rect 24030 27704 24086 27713
rect 24030 27639 24086 27648
rect 23940 27464 23992 27470
rect 23940 27406 23992 27412
rect 23952 27062 23980 27406
rect 23940 27056 23992 27062
rect 23940 26998 23992 27004
rect 24044 26382 24072 27639
rect 24136 27538 24164 29242
rect 24216 29096 24268 29102
rect 24216 29038 24268 29044
rect 24228 28490 24256 29038
rect 24216 28484 24268 28490
rect 24216 28426 24268 28432
rect 24124 27532 24176 27538
rect 24124 27474 24176 27480
rect 24032 26376 24084 26382
rect 24032 26318 24084 26324
rect 23940 25900 23992 25906
rect 23940 25842 23992 25848
rect 23952 25498 23980 25842
rect 23940 25492 23992 25498
rect 23940 25434 23992 25440
rect 24044 25430 24072 26318
rect 23768 25350 23888 25378
rect 24032 25424 24084 25430
rect 24032 25366 24084 25372
rect 23768 25158 23796 25350
rect 23848 25220 23900 25226
rect 23848 25162 23900 25168
rect 23756 25152 23808 25158
rect 23756 25094 23808 25100
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 23388 24676 23440 24682
rect 23388 24618 23440 24624
rect 23860 24449 23888 25162
rect 24124 24880 24176 24886
rect 24124 24822 24176 24828
rect 23846 24440 23902 24449
rect 23846 24375 23902 24384
rect 24136 24274 24164 24822
rect 24124 24268 24176 24274
rect 24124 24210 24176 24216
rect 23572 24064 23624 24070
rect 23572 24006 23624 24012
rect 22756 23854 23336 23882
rect 22652 21684 22704 21690
rect 22652 21626 22704 21632
rect 22756 21162 22784 23854
rect 23584 23662 23612 24006
rect 23572 23656 23624 23662
rect 23572 23598 23624 23604
rect 22836 23520 22888 23526
rect 22836 23462 22888 23468
rect 22848 22642 22876 23462
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 22836 22636 22888 22642
rect 22836 22578 22888 22584
rect 23388 22568 23440 22574
rect 23388 22510 23440 22516
rect 22836 22500 22888 22506
rect 22836 22442 22888 22448
rect 22848 22098 22876 22442
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23296 22228 23348 22234
rect 23296 22170 23348 22176
rect 22836 22092 22888 22098
rect 22836 22034 22888 22040
rect 23308 21690 23336 22170
rect 23400 22001 23428 22510
rect 23386 21992 23442 22001
rect 23386 21927 23442 21936
rect 22836 21684 22888 21690
rect 22836 21626 22888 21632
rect 23296 21684 23348 21690
rect 23296 21626 23348 21632
rect 22664 21134 22784 21162
rect 22468 19508 22520 19514
rect 22468 19450 22520 19456
rect 22560 19508 22612 19514
rect 22560 19450 22612 19456
rect 22112 18142 22416 18170
rect 21824 17876 21876 17882
rect 21824 17818 21876 17824
rect 21916 17876 21968 17882
rect 21916 17818 21968 17824
rect 21836 15502 21864 17818
rect 21928 17134 21956 17818
rect 21916 17128 21968 17134
rect 21916 17070 21968 17076
rect 21914 16552 21970 16561
rect 21914 16487 21970 16496
rect 21928 16454 21956 16487
rect 21916 16448 21968 16454
rect 21916 16390 21968 16396
rect 21928 16182 21956 16390
rect 21916 16176 21968 16182
rect 21916 16118 21968 16124
rect 22112 15994 22140 18142
rect 22192 17604 22244 17610
rect 22192 17546 22244 17552
rect 22020 15978 22140 15994
rect 22008 15972 22140 15978
rect 22060 15966 22140 15972
rect 22008 15914 22060 15920
rect 21824 15496 21876 15502
rect 21824 15438 21876 15444
rect 22100 15020 22152 15026
rect 22100 14962 22152 14968
rect 21732 14408 21784 14414
rect 21732 14350 21784 14356
rect 21824 14272 21876 14278
rect 22008 14272 22060 14278
rect 21824 14214 21876 14220
rect 21928 14232 22008 14260
rect 21836 12434 21864 14214
rect 21928 13938 21956 14232
rect 22008 14214 22060 14220
rect 21916 13932 21968 13938
rect 21916 13874 21968 13880
rect 21916 13796 21968 13802
rect 21916 13738 21968 13744
rect 21928 13274 21956 13738
rect 22112 13462 22140 14962
rect 22100 13456 22152 13462
rect 22100 13398 22152 13404
rect 21928 13246 22140 13274
rect 21916 12640 21968 12646
rect 21916 12582 21968 12588
rect 21652 12406 21864 12434
rect 21928 12434 21956 12582
rect 21928 12406 22048 12434
rect 21652 11354 21680 12406
rect 21824 12232 21876 12238
rect 21876 12192 21956 12220
rect 21824 12174 21876 12180
rect 21732 11620 21784 11626
rect 21732 11562 21784 11568
rect 21640 11348 21692 11354
rect 21640 11290 21692 11296
rect 21744 11150 21772 11562
rect 21732 11144 21784 11150
rect 21732 11086 21784 11092
rect 21928 10606 21956 12192
rect 21916 10600 21968 10606
rect 21916 10542 21968 10548
rect 21824 10464 21876 10470
rect 21824 10406 21876 10412
rect 21732 9444 21784 9450
rect 21732 9386 21784 9392
rect 21640 9376 21692 9382
rect 21640 9318 21692 9324
rect 21652 9178 21680 9318
rect 21548 9172 21600 9178
rect 21548 9114 21600 9120
rect 21640 9172 21692 9178
rect 21640 9114 21692 9120
rect 21652 8974 21680 9114
rect 21640 8968 21692 8974
rect 21640 8910 21692 8916
rect 21640 8424 21692 8430
rect 21640 8366 21692 8372
rect 21456 7812 21508 7818
rect 21456 7754 21508 7760
rect 21364 6656 21416 6662
rect 21364 6598 21416 6604
rect 21364 5160 21416 5166
rect 21364 5102 21416 5108
rect 21272 3392 21324 3398
rect 21272 3334 21324 3340
rect 21376 800 21404 5102
rect 21468 3398 21496 7754
rect 21548 4140 21600 4146
rect 21548 4082 21600 4088
rect 21560 3942 21588 4082
rect 21548 3936 21600 3942
rect 21548 3878 21600 3884
rect 21456 3392 21508 3398
rect 21456 3334 21508 3340
rect 21652 1290 21680 8366
rect 21744 7886 21772 9386
rect 21836 8090 21864 10406
rect 21928 10062 21956 10542
rect 22020 10130 22048 12406
rect 22008 10124 22060 10130
rect 22008 10066 22060 10072
rect 21916 10056 21968 10062
rect 21916 9998 21968 10004
rect 22008 9512 22060 9518
rect 22112 9489 22140 13246
rect 22008 9454 22060 9460
rect 22098 9480 22154 9489
rect 22020 8974 22048 9454
rect 22098 9415 22154 9424
rect 22008 8968 22060 8974
rect 22008 8910 22060 8916
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 21732 7880 21784 7886
rect 21732 7822 21784 7828
rect 21744 6916 21772 7822
rect 21836 7018 21864 8026
rect 21836 6990 22048 7018
rect 21744 6888 21864 6916
rect 21836 6322 21864 6888
rect 22020 6338 22048 6990
rect 22204 6458 22232 17546
rect 22284 16788 22336 16794
rect 22284 16730 22336 16736
rect 22296 16454 22324 16730
rect 22376 16584 22428 16590
rect 22376 16526 22428 16532
rect 22284 16448 22336 16454
rect 22284 16390 22336 16396
rect 22284 16244 22336 16250
rect 22284 16186 22336 16192
rect 22296 15570 22324 16186
rect 22284 15564 22336 15570
rect 22284 15506 22336 15512
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 22296 12918 22324 13874
rect 22388 13870 22416 16526
rect 22480 14278 22508 19450
rect 22560 16992 22612 16998
rect 22560 16934 22612 16940
rect 22468 14272 22520 14278
rect 22468 14214 22520 14220
rect 22376 13864 22428 13870
rect 22376 13806 22428 13812
rect 22468 13728 22520 13734
rect 22468 13670 22520 13676
rect 22284 12912 22336 12918
rect 22284 12854 22336 12860
rect 22376 12912 22428 12918
rect 22376 12854 22428 12860
rect 22388 12238 22416 12854
rect 22376 12232 22428 12238
rect 22376 12174 22428 12180
rect 22480 11218 22508 13670
rect 22572 13190 22600 16934
rect 22664 14006 22692 21134
rect 22744 20256 22796 20262
rect 22744 20198 22796 20204
rect 22756 18766 22784 20198
rect 22848 19922 22876 21626
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 22836 19916 22888 19922
rect 22836 19858 22888 19864
rect 23112 19916 23164 19922
rect 23112 19858 23164 19864
rect 23124 19825 23152 19858
rect 23110 19816 23166 19825
rect 23110 19751 23166 19760
rect 23308 19310 23336 21626
rect 23584 21350 23612 23598
rect 23940 23520 23992 23526
rect 23940 23462 23992 23468
rect 23756 23112 23808 23118
rect 23756 23054 23808 23060
rect 23768 22234 23796 23054
rect 23756 22228 23808 22234
rect 23756 22170 23808 22176
rect 23952 22030 23980 23462
rect 23940 22024 23992 22030
rect 23940 21966 23992 21972
rect 24032 21888 24084 21894
rect 24032 21830 24084 21836
rect 23572 21344 23624 21350
rect 23572 21286 23624 21292
rect 23940 20936 23992 20942
rect 23940 20878 23992 20884
rect 23388 20392 23440 20398
rect 23388 20334 23440 20340
rect 23572 20392 23624 20398
rect 23572 20334 23624 20340
rect 23296 19304 23348 19310
rect 23296 19246 23348 19252
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 22744 18760 22796 18766
rect 22744 18702 22796 18708
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 22836 17128 22888 17134
rect 22836 17070 22888 17076
rect 22848 16574 22876 17070
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 23400 16574 23428 20334
rect 23584 19446 23612 20334
rect 23664 20256 23716 20262
rect 23664 20198 23716 20204
rect 23572 19440 23624 19446
rect 23492 19400 23572 19428
rect 23492 17202 23520 19400
rect 23572 19382 23624 19388
rect 23676 18290 23704 20198
rect 23952 20058 23980 20878
rect 23940 20052 23992 20058
rect 23940 19994 23992 20000
rect 23846 19544 23902 19553
rect 23846 19479 23902 19488
rect 23860 18834 23888 19479
rect 23952 19446 23980 19994
rect 23940 19440 23992 19446
rect 23940 19382 23992 19388
rect 23848 18828 23900 18834
rect 23848 18770 23900 18776
rect 23664 18284 23716 18290
rect 23664 18226 23716 18232
rect 23572 17536 23624 17542
rect 23572 17478 23624 17484
rect 23480 17196 23532 17202
rect 23480 17138 23532 17144
rect 22742 16552 22798 16561
rect 22848 16546 23152 16574
rect 22742 16487 22798 16496
rect 22756 16046 22784 16487
rect 22744 16040 22796 16046
rect 22744 15982 22796 15988
rect 22836 16040 22888 16046
rect 22836 15982 22888 15988
rect 23124 15994 23152 16546
rect 23216 16546 23428 16574
rect 23216 16130 23244 16546
rect 23492 16402 23520 17138
rect 23308 16374 23520 16402
rect 23308 16250 23336 16374
rect 23296 16244 23348 16250
rect 23296 16186 23348 16192
rect 23216 16114 23336 16130
rect 23216 16108 23348 16114
rect 23216 16102 23296 16108
rect 23296 16050 23348 16056
rect 22744 15700 22796 15706
rect 22744 15642 22796 15648
rect 22848 15688 22876 15982
rect 23124 15966 23428 15994
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 22928 15700 22980 15706
rect 22848 15660 22928 15688
rect 22652 14000 22704 14006
rect 22652 13942 22704 13948
rect 22652 13864 22704 13870
rect 22652 13806 22704 13812
rect 22560 13184 22612 13190
rect 22560 13126 22612 13132
rect 22664 12782 22692 13806
rect 22652 12776 22704 12782
rect 22652 12718 22704 12724
rect 22468 11212 22520 11218
rect 22468 11154 22520 11160
rect 22664 10674 22692 12718
rect 22652 10668 22704 10674
rect 22652 10610 22704 10616
rect 22282 10432 22338 10441
rect 22282 10367 22338 10376
rect 22296 10198 22324 10367
rect 22558 10296 22614 10305
rect 22558 10231 22614 10240
rect 22284 10192 22336 10198
rect 22284 10134 22336 10140
rect 22374 10024 22430 10033
rect 22374 9959 22430 9968
rect 22388 9722 22416 9959
rect 22376 9716 22428 9722
rect 22376 9658 22428 9664
rect 22284 8492 22336 8498
rect 22284 8434 22336 8440
rect 22192 6452 22244 6458
rect 22192 6394 22244 6400
rect 21824 6316 21876 6322
rect 22020 6310 22232 6338
rect 21824 6258 21876 6264
rect 21732 6248 21784 6254
rect 21732 6190 21784 6196
rect 21640 1284 21692 1290
rect 21640 1226 21692 1232
rect 21744 800 21772 6190
rect 22008 6180 22060 6186
rect 22008 6122 22060 6128
rect 22020 5137 22048 6122
rect 22100 6112 22152 6118
rect 22100 6054 22152 6060
rect 22112 5234 22140 6054
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 22006 5128 22062 5137
rect 22006 5063 22062 5072
rect 21824 4276 21876 4282
rect 21824 4218 21876 4224
rect 21836 3466 21864 4218
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 22112 3738 22140 4082
rect 22100 3732 22152 3738
rect 22100 3674 22152 3680
rect 21824 3460 21876 3466
rect 21824 3402 21876 3408
rect 22204 3126 22232 6310
rect 22296 4570 22324 8434
rect 22388 7954 22416 9658
rect 22468 9580 22520 9586
rect 22468 9522 22520 9528
rect 22480 8634 22508 9522
rect 22468 8628 22520 8634
rect 22468 8570 22520 8576
rect 22468 8424 22520 8430
rect 22468 8366 22520 8372
rect 22376 7948 22428 7954
rect 22376 7890 22428 7896
rect 22376 6452 22428 6458
rect 22376 6394 22428 6400
rect 22388 4690 22416 6394
rect 22376 4684 22428 4690
rect 22376 4626 22428 4632
rect 22296 4542 22416 4570
rect 22284 4480 22336 4486
rect 22284 4422 22336 4428
rect 22192 3120 22244 3126
rect 22192 3062 22244 3068
rect 22100 2916 22152 2922
rect 22100 2858 22152 2864
rect 22112 2774 22140 2858
rect 22296 2774 22324 4422
rect 22388 4146 22416 4542
rect 22376 4140 22428 4146
rect 22376 4082 22428 4088
rect 22376 3936 22428 3942
rect 22376 3878 22428 3884
rect 22388 3233 22416 3878
rect 22374 3224 22430 3233
rect 22374 3159 22430 3168
rect 22112 2746 22232 2774
rect 22296 2746 22416 2774
rect 22204 2514 22232 2746
rect 22284 2576 22336 2582
rect 22284 2518 22336 2524
rect 22192 2508 22244 2514
rect 22192 2450 22244 2456
rect 22098 2408 22154 2417
rect 22098 2343 22154 2352
rect 22112 1834 22140 2343
rect 22100 1828 22152 1834
rect 22100 1770 22152 1776
rect 22296 1601 22324 2518
rect 22282 1592 22338 1601
rect 22282 1527 22338 1536
rect 22112 870 22232 898
rect 22112 800 22140 870
rect 18156 734 18368 762
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 21730 0 21786 800
rect 22098 0 22154 800
rect 22204 762 22232 870
rect 22388 762 22416 2746
rect 22480 800 22508 8366
rect 22572 8242 22600 10231
rect 22664 9518 22692 10610
rect 22652 9512 22704 9518
rect 22652 9454 22704 9460
rect 22756 9382 22784 15642
rect 22848 13734 22876 15660
rect 22928 15642 22980 15648
rect 23294 15464 23350 15473
rect 23294 15399 23350 15408
rect 23308 15094 23336 15399
rect 23296 15088 23348 15094
rect 23296 15030 23348 15036
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 23400 14634 23428 15966
rect 23308 14606 23428 14634
rect 23204 14476 23256 14482
rect 23204 14418 23256 14424
rect 23216 13870 23244 14418
rect 23204 13864 23256 13870
rect 23204 13806 23256 13812
rect 22836 13728 22888 13734
rect 22836 13670 22888 13676
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 22836 13456 22888 13462
rect 22836 13398 22888 13404
rect 22848 12646 22876 13398
rect 22836 12640 22888 12646
rect 22836 12582 22888 12588
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22836 12232 22888 12238
rect 22836 12174 22888 12180
rect 22848 11354 22876 12174
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 22836 11348 22888 11354
rect 22836 11290 22888 11296
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 23308 10146 23336 14606
rect 23388 14476 23440 14482
rect 23388 14418 23440 14424
rect 23400 12918 23428 14418
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 23492 13326 23520 14010
rect 23480 13320 23532 13326
rect 23480 13262 23532 13268
rect 23388 12912 23440 12918
rect 23388 12854 23440 12860
rect 23388 12640 23440 12646
rect 23388 12582 23440 12588
rect 23400 10742 23428 12582
rect 23480 11144 23532 11150
rect 23480 11086 23532 11092
rect 23388 10736 23440 10742
rect 23388 10678 23440 10684
rect 23388 10464 23440 10470
rect 23388 10406 23440 10412
rect 22848 10118 23336 10146
rect 23400 10130 23428 10406
rect 23388 10124 23440 10130
rect 22744 9376 22796 9382
rect 22744 9318 22796 9324
rect 22744 9172 22796 9178
rect 22744 9114 22796 9120
rect 22652 8968 22704 8974
rect 22652 8910 22704 8916
rect 22664 8401 22692 8910
rect 22756 8838 22784 9114
rect 22744 8832 22796 8838
rect 22744 8774 22796 8780
rect 22650 8392 22706 8401
rect 22650 8327 22706 8336
rect 22848 8294 22876 10118
rect 23388 10066 23440 10072
rect 23296 9988 23348 9994
rect 23296 9930 23348 9936
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22836 8288 22888 8294
rect 22572 8214 22784 8242
rect 22836 8230 22888 8236
rect 22560 7200 22612 7206
rect 22560 7142 22612 7148
rect 22572 3534 22600 7142
rect 22652 6792 22704 6798
rect 22652 6734 22704 6740
rect 22560 3528 22612 3534
rect 22560 3470 22612 3476
rect 22664 2582 22692 6734
rect 22756 5710 22784 8214
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22836 6724 22888 6730
rect 22836 6666 22888 6672
rect 22744 5704 22796 5710
rect 22848 5681 22876 6666
rect 23308 6168 23336 9930
rect 23400 9518 23428 10066
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 23492 8090 23520 11086
rect 23584 10810 23612 17478
rect 23846 17096 23902 17105
rect 23846 17031 23902 17040
rect 23860 16590 23888 17031
rect 23848 16584 23900 16590
rect 23848 16526 23900 16532
rect 23664 16448 23716 16454
rect 23664 16390 23716 16396
rect 23676 16182 23704 16390
rect 23664 16176 23716 16182
rect 23664 16118 23716 16124
rect 23676 15502 23704 16118
rect 23848 16108 23900 16114
rect 23848 16050 23900 16056
rect 23756 15904 23808 15910
rect 23756 15846 23808 15852
rect 23768 15570 23796 15846
rect 23756 15564 23808 15570
rect 23756 15506 23808 15512
rect 23664 15496 23716 15502
rect 23664 15438 23716 15444
rect 23676 14006 23704 15438
rect 23664 14000 23716 14006
rect 23860 13954 23888 16050
rect 24044 14958 24072 21830
rect 24124 21616 24176 21622
rect 24124 21558 24176 21564
rect 24136 21350 24164 21558
rect 24124 21344 24176 21350
rect 24124 21286 24176 21292
rect 24136 20534 24164 21286
rect 24124 20528 24176 20534
rect 24124 20470 24176 20476
rect 24136 19718 24164 20470
rect 24124 19712 24176 19718
rect 24124 19654 24176 19660
rect 24136 19446 24164 19654
rect 24124 19440 24176 19446
rect 24124 19382 24176 19388
rect 24228 17134 24256 28426
rect 24320 23186 24348 29446
rect 24400 29028 24452 29034
rect 24400 28970 24452 28976
rect 24308 23180 24360 23186
rect 24308 23122 24360 23128
rect 24308 17808 24360 17814
rect 24308 17750 24360 17756
rect 24216 17128 24268 17134
rect 24216 17070 24268 17076
rect 24124 15020 24176 15026
rect 24124 14962 24176 14968
rect 24032 14952 24084 14958
rect 24032 14894 24084 14900
rect 24032 14816 24084 14822
rect 24032 14758 24084 14764
rect 23664 13942 23716 13948
rect 23676 13462 23704 13942
rect 23768 13926 23888 13954
rect 23664 13456 23716 13462
rect 23664 13398 23716 13404
rect 23676 12986 23704 13398
rect 23664 12980 23716 12986
rect 23664 12922 23716 12928
rect 23768 11558 23796 13926
rect 23846 13832 23902 13841
rect 23846 13767 23902 13776
rect 23860 13394 23888 13767
rect 23848 13388 23900 13394
rect 23848 13330 23900 13336
rect 23940 11756 23992 11762
rect 23940 11698 23992 11704
rect 23756 11552 23808 11558
rect 23756 11494 23808 11500
rect 23756 11280 23808 11286
rect 23756 11222 23808 11228
rect 23572 10804 23624 10810
rect 23572 10746 23624 10752
rect 23662 10704 23718 10713
rect 23662 10639 23718 10648
rect 23572 8900 23624 8906
rect 23572 8842 23624 8848
rect 23480 8084 23532 8090
rect 23480 8026 23532 8032
rect 23308 6140 23428 6168
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22744 5646 22796 5652
rect 22834 5672 22890 5681
rect 22834 5607 22890 5616
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 22742 4040 22798 4049
rect 22742 3975 22798 3984
rect 22756 3738 22784 3975
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 22744 3732 22796 3738
rect 22744 3674 22796 3680
rect 22836 3392 22888 3398
rect 22836 3334 22888 3340
rect 22652 2576 22704 2582
rect 22652 2518 22704 2524
rect 22848 800 22876 3334
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 23400 2446 23428 6140
rect 23584 5778 23612 8842
rect 23572 5772 23624 5778
rect 23572 5714 23624 5720
rect 23676 5710 23704 10639
rect 23768 8974 23796 11222
rect 23848 11076 23900 11082
rect 23848 11018 23900 11024
rect 23860 10577 23888 11018
rect 23846 10568 23902 10577
rect 23846 10503 23902 10512
rect 23952 9178 23980 11698
rect 24044 10062 24072 14758
rect 24136 12442 24164 14962
rect 24320 14550 24348 17750
rect 24412 17338 24440 28970
rect 24504 28529 24532 29446
rect 24596 28558 24624 32710
rect 24676 31680 24728 31686
rect 24676 31622 24728 31628
rect 24688 31414 24716 31622
rect 24676 31408 24728 31414
rect 24676 31350 24728 31356
rect 24688 31142 24716 31350
rect 24676 31136 24728 31142
rect 24676 31078 24728 31084
rect 24688 30258 24716 31078
rect 24676 30252 24728 30258
rect 24676 30194 24728 30200
rect 24780 29306 24808 32846
rect 24964 32366 24992 32982
rect 25044 32768 25096 32774
rect 25044 32710 25096 32716
rect 25056 32570 25084 32710
rect 25044 32564 25096 32570
rect 25044 32506 25096 32512
rect 24952 32360 25004 32366
rect 24952 32302 25004 32308
rect 24860 32292 24912 32298
rect 24860 32234 24912 32240
rect 24768 29300 24820 29306
rect 24768 29242 24820 29248
rect 24872 28626 24900 32234
rect 24964 30190 24992 32302
rect 25056 32298 25084 32506
rect 25044 32292 25096 32298
rect 25044 32234 25096 32240
rect 25044 31952 25096 31958
rect 25044 31894 25096 31900
rect 24952 30184 25004 30190
rect 24952 30126 25004 30132
rect 24952 29572 25004 29578
rect 24952 29514 25004 29520
rect 24964 29345 24992 29514
rect 24950 29336 25006 29345
rect 24950 29271 25006 29280
rect 24952 29096 25004 29102
rect 24952 29038 25004 29044
rect 24860 28620 24912 28626
rect 24860 28562 24912 28568
rect 24964 28558 24992 29038
rect 24584 28552 24636 28558
rect 24490 28520 24546 28529
rect 24584 28494 24636 28500
rect 24952 28552 25004 28558
rect 24952 28494 25004 28500
rect 24490 28455 24546 28464
rect 24492 28416 24544 28422
rect 24492 28358 24544 28364
rect 24504 18902 24532 28358
rect 24768 27600 24820 27606
rect 24768 27542 24820 27548
rect 24584 27328 24636 27334
rect 24584 27270 24636 27276
rect 24596 26314 24624 27270
rect 24780 27130 24808 27542
rect 25056 27538 25084 31894
rect 25148 31278 25176 34904
rect 25136 31272 25188 31278
rect 25136 31214 25188 31220
rect 25136 31136 25188 31142
rect 25136 31078 25188 31084
rect 25044 27532 25096 27538
rect 25044 27474 25096 27480
rect 24860 27328 24912 27334
rect 24860 27270 24912 27276
rect 24768 27124 24820 27130
rect 24768 27066 24820 27072
rect 24584 26308 24636 26314
rect 24584 26250 24636 26256
rect 24872 26194 24900 27270
rect 24952 26580 25004 26586
rect 24952 26522 25004 26528
rect 24780 26166 24900 26194
rect 24780 25770 24808 26166
rect 24858 26072 24914 26081
rect 24858 26007 24914 26016
rect 24872 25974 24900 26007
rect 24860 25968 24912 25974
rect 24860 25910 24912 25916
rect 24768 25764 24820 25770
rect 24768 25706 24820 25712
rect 24872 25498 24900 25910
rect 24860 25492 24912 25498
rect 24860 25434 24912 25440
rect 24964 24970 24992 26522
rect 25044 26512 25096 26518
rect 25044 26454 25096 26460
rect 24872 24942 24992 24970
rect 24872 24154 24900 24942
rect 24872 24126 24992 24154
rect 24766 23624 24822 23633
rect 24766 23559 24822 23568
rect 24780 22574 24808 23559
rect 24860 23044 24912 23050
rect 24860 22986 24912 22992
rect 24872 22817 24900 22986
rect 24858 22808 24914 22817
rect 24858 22743 24914 22752
rect 24768 22568 24820 22574
rect 24768 22510 24820 22516
rect 24858 21176 24914 21185
rect 24858 21111 24914 21120
rect 24872 21010 24900 21111
rect 24964 21010 24992 24126
rect 25056 22098 25084 26454
rect 25148 26314 25176 31078
rect 25240 29050 25268 49030
rect 26332 48068 26384 48074
rect 26332 48010 26384 48016
rect 25320 47660 25372 47666
rect 25320 47602 25372 47608
rect 25332 47297 25360 47602
rect 25318 47288 25374 47297
rect 25318 47223 25374 47232
rect 25320 46912 25372 46918
rect 25320 46854 25372 46860
rect 25332 46578 25360 46854
rect 25320 46572 25372 46578
rect 25320 46514 25372 46520
rect 25332 46481 25360 46514
rect 25318 46472 25374 46481
rect 25318 46407 25374 46416
rect 25412 46368 25464 46374
rect 25412 46310 25464 46316
rect 25320 45960 25372 45966
rect 25320 45902 25372 45908
rect 25332 45665 25360 45902
rect 25318 45656 25374 45665
rect 25318 45591 25374 45600
rect 25320 45280 25372 45286
rect 25320 45222 25372 45228
rect 25332 44878 25360 45222
rect 25320 44872 25372 44878
rect 25318 44840 25320 44849
rect 25372 44840 25374 44849
rect 25318 44775 25374 44784
rect 25320 41132 25372 41138
rect 25320 41074 25372 41080
rect 25332 40769 25360 41074
rect 25318 40760 25374 40769
rect 25318 40695 25374 40704
rect 25320 39432 25372 39438
rect 25320 39374 25372 39380
rect 25332 39137 25360 39374
rect 25318 39128 25374 39137
rect 25318 39063 25374 39072
rect 25320 38752 25372 38758
rect 25320 38694 25372 38700
rect 25332 38350 25360 38694
rect 25320 38344 25372 38350
rect 25318 38312 25320 38321
rect 25372 38312 25374 38321
rect 25318 38247 25374 38256
rect 25320 36168 25372 36174
rect 25320 36110 25372 36116
rect 25332 35873 25360 36110
rect 25318 35864 25374 35873
rect 25318 35799 25374 35808
rect 25424 35766 25452 46310
rect 25872 44260 25924 44266
rect 25872 44202 25924 44208
rect 25504 43648 25556 43654
rect 25504 43590 25556 43596
rect 25516 43382 25544 43590
rect 25504 43376 25556 43382
rect 25504 43318 25556 43324
rect 25516 43217 25544 43318
rect 25502 43208 25558 43217
rect 25502 43143 25558 43152
rect 25688 42628 25740 42634
rect 25688 42570 25740 42576
rect 25596 40928 25648 40934
rect 25596 40870 25648 40876
rect 25504 40384 25556 40390
rect 25504 40326 25556 40332
rect 25516 40118 25544 40326
rect 25504 40112 25556 40118
rect 25504 40054 25556 40060
rect 25516 39953 25544 40054
rect 25502 39944 25558 39953
rect 25502 39879 25558 39888
rect 25504 37120 25556 37126
rect 25504 37062 25556 37068
rect 25516 36854 25544 37062
rect 25504 36848 25556 36854
rect 25504 36790 25556 36796
rect 25516 36689 25544 36790
rect 25502 36680 25558 36689
rect 25502 36615 25558 36624
rect 25412 35760 25464 35766
rect 25412 35702 25464 35708
rect 25320 35488 25372 35494
rect 25320 35430 25372 35436
rect 25332 35086 25360 35430
rect 25320 35080 25372 35086
rect 25318 35048 25320 35057
rect 25372 35048 25374 35057
rect 25318 34983 25374 34992
rect 25320 34604 25372 34610
rect 25320 34546 25372 34552
rect 25332 34241 25360 34546
rect 25318 34232 25374 34241
rect 25318 34167 25374 34176
rect 25320 33992 25372 33998
rect 25320 33934 25372 33940
rect 25332 33425 25360 33934
rect 25504 33516 25556 33522
rect 25504 33458 25556 33464
rect 25318 33416 25374 33425
rect 25318 33351 25374 33360
rect 25412 33312 25464 33318
rect 25412 33254 25464 33260
rect 25320 31816 25372 31822
rect 25318 31784 25320 31793
rect 25372 31784 25374 31793
rect 25318 31719 25374 31728
rect 25318 30152 25374 30161
rect 25318 30087 25374 30096
rect 25332 29646 25360 30087
rect 25320 29640 25372 29646
rect 25320 29582 25372 29588
rect 25332 29306 25360 29582
rect 25320 29300 25372 29306
rect 25320 29242 25372 29248
rect 25240 29022 25360 29050
rect 25228 28960 25280 28966
rect 25228 28902 25280 28908
rect 25240 28014 25268 28902
rect 25228 28008 25280 28014
rect 25228 27950 25280 27956
rect 25332 27334 25360 29022
rect 25424 28694 25452 33254
rect 25516 32609 25544 33458
rect 25608 32910 25636 40870
rect 25596 32904 25648 32910
rect 25596 32846 25648 32852
rect 25502 32600 25558 32609
rect 25502 32535 25558 32544
rect 25504 32496 25556 32502
rect 25504 32438 25556 32444
rect 25516 31754 25544 32438
rect 25516 31726 25636 31754
rect 25504 31340 25556 31346
rect 25504 31282 25556 31288
rect 25516 30977 25544 31282
rect 25502 30968 25558 30977
rect 25502 30903 25504 30912
rect 25556 30903 25558 30912
rect 25504 30874 25556 30880
rect 25504 28756 25556 28762
rect 25504 28698 25556 28704
rect 25412 28688 25464 28694
rect 25412 28630 25464 28636
rect 25412 27872 25464 27878
rect 25412 27814 25464 27820
rect 25424 27470 25452 27814
rect 25412 27464 25464 27470
rect 25412 27406 25464 27412
rect 25320 27328 25372 27334
rect 25320 27270 25372 27276
rect 25228 27056 25280 27062
rect 25228 26998 25280 27004
rect 25240 26586 25268 26998
rect 25318 26888 25374 26897
rect 25318 26823 25374 26832
rect 25228 26580 25280 26586
rect 25228 26522 25280 26528
rect 25228 26444 25280 26450
rect 25228 26386 25280 26392
rect 25136 26308 25188 26314
rect 25136 26250 25188 26256
rect 25136 25832 25188 25838
rect 25136 25774 25188 25780
rect 25148 25265 25176 25774
rect 25134 25256 25190 25265
rect 25134 25191 25190 25200
rect 25136 25152 25188 25158
rect 25136 25094 25188 25100
rect 25148 22778 25176 25094
rect 25240 24750 25268 26386
rect 25332 25294 25360 26823
rect 25424 26042 25452 27406
rect 25516 27062 25544 28698
rect 25504 27056 25556 27062
rect 25504 26998 25556 27004
rect 25504 26920 25556 26926
rect 25504 26862 25556 26868
rect 25412 26036 25464 26042
rect 25412 25978 25464 25984
rect 25320 25288 25372 25294
rect 25320 25230 25372 25236
rect 25228 24744 25280 24750
rect 25228 24686 25280 24692
rect 25240 23866 25268 24686
rect 25332 24410 25360 25230
rect 25412 25220 25464 25226
rect 25412 25162 25464 25168
rect 25424 24886 25452 25162
rect 25412 24880 25464 24886
rect 25412 24822 25464 24828
rect 25320 24404 25372 24410
rect 25320 24346 25372 24352
rect 25424 24290 25452 24822
rect 25516 24750 25544 26862
rect 25608 26586 25636 31726
rect 25596 26580 25648 26586
rect 25596 26522 25648 26528
rect 25596 26376 25648 26382
rect 25596 26318 25648 26324
rect 25504 24744 25556 24750
rect 25504 24686 25556 24692
rect 25332 24262 25452 24290
rect 25332 24070 25360 24262
rect 25320 24064 25372 24070
rect 25320 24006 25372 24012
rect 25228 23860 25280 23866
rect 25228 23802 25280 23808
rect 25332 23746 25360 24006
rect 25240 23730 25360 23746
rect 25228 23724 25360 23730
rect 25280 23718 25360 23724
rect 25228 23666 25280 23672
rect 25240 23526 25268 23666
rect 25228 23520 25280 23526
rect 25228 23462 25280 23468
rect 25136 22772 25188 22778
rect 25136 22714 25188 22720
rect 25044 22092 25096 22098
rect 25240 22094 25268 23462
rect 25320 23180 25372 23186
rect 25320 23122 25372 23128
rect 25044 22034 25096 22040
rect 25148 22066 25268 22094
rect 25148 21350 25176 22066
rect 25332 21486 25360 23122
rect 25516 22166 25544 24686
rect 25608 24342 25636 26318
rect 25596 24336 25648 24342
rect 25596 24278 25648 24284
rect 25608 23866 25636 24278
rect 25596 23860 25648 23866
rect 25596 23802 25648 23808
rect 25608 23118 25636 23802
rect 25596 23112 25648 23118
rect 25596 23054 25648 23060
rect 25504 22160 25556 22166
rect 25504 22102 25556 22108
rect 25320 21480 25372 21486
rect 25320 21422 25372 21428
rect 25136 21344 25188 21350
rect 25136 21286 25188 21292
rect 24860 21004 24912 21010
rect 24860 20946 24912 20952
rect 24952 21004 25004 21010
rect 24952 20946 25004 20952
rect 24584 20800 24636 20806
rect 24584 20742 24636 20748
rect 24860 20800 24912 20806
rect 24860 20742 24912 20748
rect 24492 18896 24544 18902
rect 24492 18838 24544 18844
rect 24596 17814 24624 20742
rect 24674 20360 24730 20369
rect 24674 20295 24730 20304
rect 24688 18222 24716 20295
rect 24872 19922 24900 20742
rect 25332 20602 25360 21422
rect 25320 20596 25372 20602
rect 25320 20538 25372 20544
rect 25136 20392 25188 20398
rect 25136 20334 25188 20340
rect 24860 19916 24912 19922
rect 24860 19858 24912 19864
rect 25148 19514 25176 20334
rect 25412 19712 25464 19718
rect 25412 19654 25464 19660
rect 25424 19514 25452 19654
rect 25136 19508 25188 19514
rect 25136 19450 25188 19456
rect 25412 19508 25464 19514
rect 25412 19450 25464 19456
rect 24858 18728 24914 18737
rect 24858 18663 24914 18672
rect 24872 18358 24900 18663
rect 24860 18352 24912 18358
rect 24860 18294 24912 18300
rect 24676 18216 24728 18222
rect 24676 18158 24728 18164
rect 24950 17912 25006 17921
rect 24950 17847 25006 17856
rect 24584 17808 24636 17814
rect 24584 17750 24636 17756
rect 24964 17746 24992 17847
rect 25148 17746 25176 19450
rect 25412 18692 25464 18698
rect 25412 18634 25464 18640
rect 24952 17740 25004 17746
rect 24952 17682 25004 17688
rect 25136 17740 25188 17746
rect 25136 17682 25188 17688
rect 24584 17672 24636 17678
rect 24584 17614 24636 17620
rect 24400 17332 24452 17338
rect 24400 17274 24452 17280
rect 24596 16794 24624 17614
rect 24676 17536 24728 17542
rect 24676 17478 24728 17484
rect 24584 16788 24636 16794
rect 24584 16730 24636 16736
rect 24584 16040 24636 16046
rect 24584 15982 24636 15988
rect 24308 14544 24360 14550
rect 24308 14486 24360 14492
rect 24492 14408 24544 14414
rect 24492 14350 24544 14356
rect 24400 14340 24452 14346
rect 24400 14282 24452 14288
rect 24412 13938 24440 14282
rect 24400 13932 24452 13938
rect 24400 13874 24452 13880
rect 24504 13530 24532 14350
rect 24492 13524 24544 13530
rect 24492 13466 24544 13472
rect 24124 12436 24176 12442
rect 24124 12378 24176 12384
rect 24124 11552 24176 11558
rect 24124 11494 24176 11500
rect 24032 10056 24084 10062
rect 24032 9998 24084 10004
rect 24032 9580 24084 9586
rect 24032 9522 24084 9528
rect 24044 9450 24072 9522
rect 24032 9444 24084 9450
rect 24032 9386 24084 9392
rect 23940 9172 23992 9178
rect 23940 9114 23992 9120
rect 24044 9058 24072 9386
rect 23952 9030 24072 9058
rect 23756 8968 23808 8974
rect 23756 8910 23808 8916
rect 23952 8838 23980 9030
rect 23940 8832 23992 8838
rect 23940 8774 23992 8780
rect 23952 7886 23980 8774
rect 24032 8016 24084 8022
rect 24032 7958 24084 7964
rect 23940 7880 23992 7886
rect 23940 7822 23992 7828
rect 23952 7750 23980 7822
rect 23848 7744 23900 7750
rect 23848 7686 23900 7692
rect 23940 7744 23992 7750
rect 23940 7686 23992 7692
rect 23860 6934 23888 7686
rect 23940 6996 23992 7002
rect 23940 6938 23992 6944
rect 23848 6928 23900 6934
rect 23848 6870 23900 6876
rect 23756 6860 23808 6866
rect 23756 6802 23808 6808
rect 23768 6254 23796 6802
rect 23860 6322 23888 6870
rect 23848 6316 23900 6322
rect 23848 6258 23900 6264
rect 23756 6248 23808 6254
rect 23756 6190 23808 6196
rect 23664 5704 23716 5710
rect 23664 5646 23716 5652
rect 23756 5636 23808 5642
rect 23756 5578 23808 5584
rect 23768 5234 23796 5578
rect 23756 5228 23808 5234
rect 23756 5170 23808 5176
rect 23848 5024 23900 5030
rect 23848 4966 23900 4972
rect 23754 4584 23810 4593
rect 23754 4519 23810 4528
rect 23768 4486 23796 4519
rect 23756 4480 23808 4486
rect 23756 4422 23808 4428
rect 23860 4146 23888 4966
rect 23848 4140 23900 4146
rect 23848 4082 23900 4088
rect 23480 3664 23532 3670
rect 23480 3606 23532 3612
rect 23388 2440 23440 2446
rect 23388 2382 23440 2388
rect 23492 1850 23520 3606
rect 23952 3602 23980 6938
rect 24044 4826 24072 7958
rect 24136 7274 24164 11494
rect 24306 10840 24362 10849
rect 24306 10775 24362 10784
rect 24216 9920 24268 9926
rect 24216 9862 24268 9868
rect 24124 7268 24176 7274
rect 24124 7210 24176 7216
rect 24228 6390 24256 9862
rect 24216 6384 24268 6390
rect 24216 6326 24268 6332
rect 24032 4820 24084 4826
rect 24032 4762 24084 4768
rect 24320 4622 24348 10775
rect 24400 10600 24452 10606
rect 24400 10542 24452 10548
rect 24412 9450 24440 10542
rect 24596 10266 24624 15982
rect 24688 15570 24716 17478
rect 24860 17196 24912 17202
rect 24860 17138 24912 17144
rect 24872 16454 24900 17138
rect 24860 16448 24912 16454
rect 24860 16390 24912 16396
rect 25136 16448 25188 16454
rect 25136 16390 25188 16396
rect 24766 16280 24822 16289
rect 24872 16250 24900 16390
rect 24766 16215 24822 16224
rect 24860 16244 24912 16250
rect 24676 15564 24728 15570
rect 24676 15506 24728 15512
rect 24780 14958 24808 16215
rect 24860 16186 24912 16192
rect 25148 15706 25176 16390
rect 25136 15700 25188 15706
rect 25136 15642 25188 15648
rect 25228 15428 25280 15434
rect 25228 15370 25280 15376
rect 24768 14952 24820 14958
rect 24768 14894 24820 14900
rect 24858 14648 24914 14657
rect 24858 14583 24914 14592
rect 25044 14612 25096 14618
rect 24872 14482 24900 14583
rect 25044 14554 25096 14560
rect 24860 14476 24912 14482
rect 24860 14418 24912 14424
rect 24860 14272 24912 14278
rect 24860 14214 24912 14220
rect 24766 13016 24822 13025
rect 24766 12951 24822 12960
rect 24780 11694 24808 12951
rect 24872 11914 24900 14214
rect 24950 12200 25006 12209
rect 24950 12135 24952 12144
rect 25004 12135 25006 12144
rect 24952 12106 25004 12112
rect 24872 11886 24992 11914
rect 24860 11824 24912 11830
rect 24860 11766 24912 11772
rect 24768 11688 24820 11694
rect 24768 11630 24820 11636
rect 24872 11393 24900 11766
rect 24964 11762 24992 11886
rect 24952 11756 25004 11762
rect 24952 11698 25004 11704
rect 24858 11384 24914 11393
rect 24858 11319 24914 11328
rect 24584 10260 24636 10266
rect 24584 10202 24636 10208
rect 24766 9752 24822 9761
rect 24766 9687 24822 9696
rect 24490 9480 24546 9489
rect 24400 9444 24452 9450
rect 24490 9415 24546 9424
rect 24400 9386 24452 9392
rect 24400 8628 24452 8634
rect 24400 8570 24452 8576
rect 24308 4616 24360 4622
rect 24308 4558 24360 4564
rect 24412 4049 24440 8570
rect 24504 4622 24532 9415
rect 24780 8430 24808 9687
rect 24860 9376 24912 9382
rect 24860 9318 24912 9324
rect 24768 8424 24820 8430
rect 24768 8366 24820 8372
rect 24768 7744 24820 7750
rect 24768 7686 24820 7692
rect 24584 6656 24636 6662
rect 24584 6598 24636 6604
rect 24676 6656 24728 6662
rect 24676 6598 24728 6604
rect 24596 6458 24624 6598
rect 24584 6452 24636 6458
rect 24584 6394 24636 6400
rect 24492 4616 24544 4622
rect 24492 4558 24544 4564
rect 24398 4040 24454 4049
rect 24398 3975 24454 3984
rect 23940 3596 23992 3602
rect 23940 3538 23992 3544
rect 23938 3496 23994 3505
rect 23938 3431 23994 3440
rect 23572 3052 23624 3058
rect 23572 2994 23624 3000
rect 23584 2650 23612 2994
rect 23572 2644 23624 2650
rect 23572 2586 23624 2592
rect 23848 2304 23900 2310
rect 23848 2246 23900 2252
rect 23860 2038 23888 2246
rect 23848 2032 23900 2038
rect 23848 1974 23900 1980
rect 23492 1822 23612 1850
rect 23204 1284 23256 1290
rect 23204 1226 23256 1232
rect 23216 800 23244 1226
rect 23584 800 23612 1822
rect 23952 800 23980 3431
rect 24688 3194 24716 6598
rect 24780 6322 24808 7686
rect 24872 7426 24900 9318
rect 24950 8936 25006 8945
rect 24950 8871 24952 8880
rect 25004 8871 25006 8880
rect 24952 8842 25004 8848
rect 24872 7398 24992 7426
rect 24860 7336 24912 7342
rect 24858 7304 24860 7313
rect 24912 7304 24914 7313
rect 24858 7239 24914 7248
rect 24964 6882 24992 7398
rect 24872 6854 24992 6882
rect 24768 6316 24820 6322
rect 24768 6258 24820 6264
rect 24780 6118 24808 6258
rect 24768 6112 24820 6118
rect 24768 6054 24820 6060
rect 24780 4486 24808 6054
rect 24768 4480 24820 4486
rect 24768 4422 24820 4428
rect 24780 3466 24808 4422
rect 24768 3460 24820 3466
rect 24768 3402 24820 3408
rect 24780 3194 24808 3402
rect 24676 3188 24728 3194
rect 24676 3130 24728 3136
rect 24768 3188 24820 3194
rect 24768 3130 24820 3136
rect 24872 2774 24900 6854
rect 24952 6792 25004 6798
rect 24952 6734 25004 6740
rect 24964 6497 24992 6734
rect 24950 6488 25006 6497
rect 24950 6423 25006 6432
rect 25056 6322 25084 14554
rect 25136 13252 25188 13258
rect 25136 13194 25188 13200
rect 25148 8242 25176 13194
rect 25240 11150 25268 15370
rect 25228 11144 25280 11150
rect 25228 11086 25280 11092
rect 25148 8214 25268 8242
rect 25134 8120 25190 8129
rect 25134 8055 25190 8064
rect 25148 7478 25176 8055
rect 25136 7472 25188 7478
rect 25136 7414 25188 7420
rect 25240 6458 25268 8214
rect 25320 7540 25372 7546
rect 25320 7482 25372 7488
rect 25228 6452 25280 6458
rect 25228 6394 25280 6400
rect 25044 6316 25096 6322
rect 25044 6258 25096 6264
rect 25136 5568 25188 5574
rect 25136 5510 25188 5516
rect 24952 3664 25004 3670
rect 24950 3632 24952 3641
rect 25004 3632 25006 3641
rect 24950 3567 25006 3576
rect 25148 3534 25176 5510
rect 25136 3528 25188 3534
rect 25136 3470 25188 3476
rect 24872 2746 24992 2774
rect 24308 2644 24360 2650
rect 24308 2586 24360 2592
rect 24320 800 24348 2586
rect 24964 2446 24992 2746
rect 24952 2440 25004 2446
rect 24952 2382 25004 2388
rect 22204 734 22416 762
rect 22466 0 22522 800
rect 22834 0 22890 800
rect 23202 0 23258 800
rect 23570 0 23626 800
rect 23938 0 23994 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 25042 0 25098 800
rect 25332 785 25360 7482
rect 25424 4146 25452 18634
rect 25700 15162 25728 42570
rect 25780 34944 25832 34950
rect 25780 34886 25832 34892
rect 25792 32502 25820 34886
rect 25780 32496 25832 32502
rect 25780 32438 25832 32444
rect 25780 26988 25832 26994
rect 25780 26930 25832 26936
rect 25688 15156 25740 15162
rect 25688 15098 25740 15104
rect 25792 11898 25820 26930
rect 25884 26772 25912 44202
rect 25964 43172 26016 43178
rect 25964 43114 26016 43120
rect 25976 26874 26004 43114
rect 26148 41540 26200 41546
rect 26148 41482 26200 41488
rect 26056 37732 26108 37738
rect 26056 37674 26108 37680
rect 26068 26994 26096 37674
rect 26056 26988 26108 26994
rect 26056 26930 26108 26936
rect 25976 26846 26096 26874
rect 25884 26744 26004 26772
rect 25872 26580 25924 26586
rect 25872 26522 25924 26528
rect 25884 17610 25912 26522
rect 25976 18970 26004 26744
rect 25964 18964 26016 18970
rect 25964 18906 26016 18912
rect 26068 17882 26096 26846
rect 26056 17876 26108 17882
rect 26056 17818 26108 17824
rect 25872 17604 25924 17610
rect 25872 17546 25924 17552
rect 25780 11892 25832 11898
rect 25780 11834 25832 11840
rect 26160 11626 26188 41482
rect 26240 33856 26292 33862
rect 26240 33798 26292 33804
rect 26252 28218 26280 33798
rect 26240 28212 26292 28218
rect 26240 28154 26292 28160
rect 26344 23322 26372 48010
rect 26424 47456 26476 47462
rect 26424 47398 26476 47404
rect 26436 29238 26464 47398
rect 26528 29850 26556 53382
rect 26792 52488 26844 52494
rect 26792 52430 26844 52436
rect 26700 36644 26752 36650
rect 26700 36586 26752 36592
rect 26608 36032 26660 36038
rect 26608 35974 26660 35980
rect 26516 29844 26568 29850
rect 26516 29786 26568 29792
rect 26424 29232 26476 29238
rect 26424 29174 26476 29180
rect 26332 23316 26384 23322
rect 26332 23258 26384 23264
rect 26620 18766 26648 35974
rect 26608 18760 26660 18766
rect 26608 18702 26660 18708
rect 26148 11620 26200 11626
rect 26148 11562 26200 11568
rect 26712 11218 26740 36586
rect 26804 32230 26832 52430
rect 26884 51332 26936 51338
rect 26884 51274 26936 51280
rect 26792 32224 26844 32230
rect 26792 32166 26844 32172
rect 26896 29170 26924 51274
rect 26884 29164 26936 29170
rect 26884 29106 26936 29112
rect 26700 11212 26752 11218
rect 26700 11154 26752 11160
rect 25412 4140 25464 4146
rect 25412 4082 25464 4088
rect 25318 776 25374 785
rect 25318 711 25374 720
<< via2 >>
rect 2956 53882 3012 53884
rect 3036 53882 3092 53884
rect 3116 53882 3172 53884
rect 3196 53882 3252 53884
rect 2956 53830 3002 53882
rect 3002 53830 3012 53882
rect 3036 53830 3066 53882
rect 3066 53830 3078 53882
rect 3078 53830 3092 53882
rect 3116 53830 3130 53882
rect 3130 53830 3142 53882
rect 3142 53830 3172 53882
rect 3196 53830 3206 53882
rect 3206 53830 3252 53882
rect 2956 53828 3012 53830
rect 3036 53828 3092 53830
rect 3116 53828 3172 53830
rect 3196 53828 3252 53830
rect 2956 52794 3012 52796
rect 3036 52794 3092 52796
rect 3116 52794 3172 52796
rect 3196 52794 3252 52796
rect 2956 52742 3002 52794
rect 3002 52742 3012 52794
rect 3036 52742 3066 52794
rect 3066 52742 3078 52794
rect 3078 52742 3092 52794
rect 3116 52742 3130 52794
rect 3130 52742 3142 52794
rect 3142 52742 3172 52794
rect 3196 52742 3206 52794
rect 3206 52742 3252 52794
rect 2956 52740 3012 52742
rect 3036 52740 3092 52742
rect 3116 52740 3172 52742
rect 3196 52740 3252 52742
rect 2956 51706 3012 51708
rect 3036 51706 3092 51708
rect 3116 51706 3172 51708
rect 3196 51706 3252 51708
rect 2956 51654 3002 51706
rect 3002 51654 3012 51706
rect 3036 51654 3066 51706
rect 3066 51654 3078 51706
rect 3078 51654 3092 51706
rect 3116 51654 3130 51706
rect 3130 51654 3142 51706
rect 3142 51654 3172 51706
rect 3196 51654 3206 51706
rect 3206 51654 3252 51706
rect 2956 51652 3012 51654
rect 3036 51652 3092 51654
rect 3116 51652 3172 51654
rect 3196 51652 3252 51654
rect 2956 50618 3012 50620
rect 3036 50618 3092 50620
rect 3116 50618 3172 50620
rect 3196 50618 3252 50620
rect 2956 50566 3002 50618
rect 3002 50566 3012 50618
rect 3036 50566 3066 50618
rect 3066 50566 3078 50618
rect 3078 50566 3092 50618
rect 3116 50566 3130 50618
rect 3130 50566 3142 50618
rect 3142 50566 3172 50618
rect 3196 50566 3206 50618
rect 3206 50566 3252 50618
rect 2956 50564 3012 50566
rect 3036 50564 3092 50566
rect 3116 50564 3172 50566
rect 3196 50564 3252 50566
rect 7956 54426 8012 54428
rect 8036 54426 8092 54428
rect 8116 54426 8172 54428
rect 8196 54426 8252 54428
rect 7956 54374 8002 54426
rect 8002 54374 8012 54426
rect 8036 54374 8066 54426
rect 8066 54374 8078 54426
rect 8078 54374 8092 54426
rect 8116 54374 8130 54426
rect 8130 54374 8142 54426
rect 8142 54374 8172 54426
rect 8196 54374 8206 54426
rect 8206 54374 8252 54426
rect 7956 54372 8012 54374
rect 8036 54372 8092 54374
rect 8116 54372 8172 54374
rect 8196 54372 8252 54374
rect 7956 53338 8012 53340
rect 8036 53338 8092 53340
rect 8116 53338 8172 53340
rect 8196 53338 8252 53340
rect 7956 53286 8002 53338
rect 8002 53286 8012 53338
rect 8036 53286 8066 53338
rect 8066 53286 8078 53338
rect 8078 53286 8092 53338
rect 8116 53286 8130 53338
rect 8130 53286 8142 53338
rect 8142 53286 8172 53338
rect 8196 53286 8206 53338
rect 8206 53286 8252 53338
rect 7956 53284 8012 53286
rect 8036 53284 8092 53286
rect 8116 53284 8172 53286
rect 8196 53284 8252 53286
rect 7956 52250 8012 52252
rect 8036 52250 8092 52252
rect 8116 52250 8172 52252
rect 8196 52250 8252 52252
rect 7956 52198 8002 52250
rect 8002 52198 8012 52250
rect 8036 52198 8066 52250
rect 8066 52198 8078 52250
rect 8078 52198 8092 52250
rect 8116 52198 8130 52250
rect 8130 52198 8142 52250
rect 8142 52198 8172 52250
rect 8196 52198 8206 52250
rect 8206 52198 8252 52250
rect 7956 52196 8012 52198
rect 8036 52196 8092 52198
rect 8116 52196 8172 52198
rect 8196 52196 8252 52198
rect 7956 51162 8012 51164
rect 8036 51162 8092 51164
rect 8116 51162 8172 51164
rect 8196 51162 8252 51164
rect 7956 51110 8002 51162
rect 8002 51110 8012 51162
rect 8036 51110 8066 51162
rect 8066 51110 8078 51162
rect 8078 51110 8092 51162
rect 8116 51110 8130 51162
rect 8130 51110 8142 51162
rect 8142 51110 8172 51162
rect 8196 51110 8206 51162
rect 8206 51110 8252 51162
rect 7956 51108 8012 51110
rect 8036 51108 8092 51110
rect 8116 51108 8172 51110
rect 8196 51108 8252 51110
rect 2956 49530 3012 49532
rect 3036 49530 3092 49532
rect 3116 49530 3172 49532
rect 3196 49530 3252 49532
rect 2956 49478 3002 49530
rect 3002 49478 3012 49530
rect 3036 49478 3066 49530
rect 3066 49478 3078 49530
rect 3078 49478 3092 49530
rect 3116 49478 3130 49530
rect 3130 49478 3142 49530
rect 3142 49478 3172 49530
rect 3196 49478 3206 49530
rect 3206 49478 3252 49530
rect 2956 49476 3012 49478
rect 3036 49476 3092 49478
rect 3116 49476 3172 49478
rect 3196 49476 3252 49478
rect 2956 48442 3012 48444
rect 3036 48442 3092 48444
rect 3116 48442 3172 48444
rect 3196 48442 3252 48444
rect 2956 48390 3002 48442
rect 3002 48390 3012 48442
rect 3036 48390 3066 48442
rect 3066 48390 3078 48442
rect 3078 48390 3092 48442
rect 3116 48390 3130 48442
rect 3130 48390 3142 48442
rect 3142 48390 3172 48442
rect 3196 48390 3206 48442
rect 3206 48390 3252 48442
rect 2956 48388 3012 48390
rect 3036 48388 3092 48390
rect 3116 48388 3172 48390
rect 3196 48388 3252 48390
rect 7956 50074 8012 50076
rect 8036 50074 8092 50076
rect 8116 50074 8172 50076
rect 8196 50074 8252 50076
rect 7956 50022 8002 50074
rect 8002 50022 8012 50074
rect 8036 50022 8066 50074
rect 8066 50022 8078 50074
rect 8078 50022 8092 50074
rect 8116 50022 8130 50074
rect 8130 50022 8142 50074
rect 8142 50022 8172 50074
rect 8196 50022 8206 50074
rect 8206 50022 8252 50074
rect 7956 50020 8012 50022
rect 8036 50020 8092 50022
rect 8116 50020 8172 50022
rect 8196 50020 8252 50022
rect 7956 48986 8012 48988
rect 8036 48986 8092 48988
rect 8116 48986 8172 48988
rect 8196 48986 8252 48988
rect 7956 48934 8002 48986
rect 8002 48934 8012 48986
rect 8036 48934 8066 48986
rect 8066 48934 8078 48986
rect 8078 48934 8092 48986
rect 8116 48934 8130 48986
rect 8130 48934 8142 48986
rect 8142 48934 8172 48986
rect 8196 48934 8206 48986
rect 8206 48934 8252 48986
rect 7956 48932 8012 48934
rect 8036 48932 8092 48934
rect 8116 48932 8172 48934
rect 8196 48932 8252 48934
rect 2956 47354 3012 47356
rect 3036 47354 3092 47356
rect 3116 47354 3172 47356
rect 3196 47354 3252 47356
rect 2956 47302 3002 47354
rect 3002 47302 3012 47354
rect 3036 47302 3066 47354
rect 3066 47302 3078 47354
rect 3078 47302 3092 47354
rect 3116 47302 3130 47354
rect 3130 47302 3142 47354
rect 3142 47302 3172 47354
rect 3196 47302 3206 47354
rect 3206 47302 3252 47354
rect 2956 47300 3012 47302
rect 3036 47300 3092 47302
rect 3116 47300 3172 47302
rect 3196 47300 3252 47302
rect 2956 46266 3012 46268
rect 3036 46266 3092 46268
rect 3116 46266 3172 46268
rect 3196 46266 3252 46268
rect 2956 46214 3002 46266
rect 3002 46214 3012 46266
rect 3036 46214 3066 46266
rect 3066 46214 3078 46266
rect 3078 46214 3092 46266
rect 3116 46214 3130 46266
rect 3130 46214 3142 46266
rect 3142 46214 3172 46266
rect 3196 46214 3206 46266
rect 3206 46214 3252 46266
rect 2956 46212 3012 46214
rect 3036 46212 3092 46214
rect 3116 46212 3172 46214
rect 3196 46212 3252 46214
rect 7956 47898 8012 47900
rect 8036 47898 8092 47900
rect 8116 47898 8172 47900
rect 8196 47898 8252 47900
rect 7956 47846 8002 47898
rect 8002 47846 8012 47898
rect 8036 47846 8066 47898
rect 8066 47846 8078 47898
rect 8078 47846 8092 47898
rect 8116 47846 8130 47898
rect 8130 47846 8142 47898
rect 8142 47846 8172 47898
rect 8196 47846 8206 47898
rect 8206 47846 8252 47898
rect 7956 47844 8012 47846
rect 8036 47844 8092 47846
rect 8116 47844 8172 47846
rect 8196 47844 8252 47846
rect 7956 46810 8012 46812
rect 8036 46810 8092 46812
rect 8116 46810 8172 46812
rect 8196 46810 8252 46812
rect 7956 46758 8002 46810
rect 8002 46758 8012 46810
rect 8036 46758 8066 46810
rect 8066 46758 8078 46810
rect 8078 46758 8092 46810
rect 8116 46758 8130 46810
rect 8130 46758 8142 46810
rect 8142 46758 8172 46810
rect 8196 46758 8206 46810
rect 8206 46758 8252 46810
rect 7956 46756 8012 46758
rect 8036 46756 8092 46758
rect 8116 46756 8172 46758
rect 8196 46756 8252 46758
rect 2956 45178 3012 45180
rect 3036 45178 3092 45180
rect 3116 45178 3172 45180
rect 3196 45178 3252 45180
rect 2956 45126 3002 45178
rect 3002 45126 3012 45178
rect 3036 45126 3066 45178
rect 3066 45126 3078 45178
rect 3078 45126 3092 45178
rect 3116 45126 3130 45178
rect 3130 45126 3142 45178
rect 3142 45126 3172 45178
rect 3196 45126 3206 45178
rect 3206 45126 3252 45178
rect 2956 45124 3012 45126
rect 3036 45124 3092 45126
rect 3116 45124 3172 45126
rect 3196 45124 3252 45126
rect 2956 44090 3012 44092
rect 3036 44090 3092 44092
rect 3116 44090 3172 44092
rect 3196 44090 3252 44092
rect 2956 44038 3002 44090
rect 3002 44038 3012 44090
rect 3036 44038 3066 44090
rect 3066 44038 3078 44090
rect 3078 44038 3092 44090
rect 3116 44038 3130 44090
rect 3130 44038 3142 44090
rect 3142 44038 3172 44090
rect 3196 44038 3206 44090
rect 3206 44038 3252 44090
rect 2956 44036 3012 44038
rect 3036 44036 3092 44038
rect 3116 44036 3172 44038
rect 3196 44036 3252 44038
rect 2956 43002 3012 43004
rect 3036 43002 3092 43004
rect 3116 43002 3172 43004
rect 3196 43002 3252 43004
rect 2956 42950 3002 43002
rect 3002 42950 3012 43002
rect 3036 42950 3066 43002
rect 3066 42950 3078 43002
rect 3078 42950 3092 43002
rect 3116 42950 3130 43002
rect 3130 42950 3142 43002
rect 3142 42950 3172 43002
rect 3196 42950 3206 43002
rect 3206 42950 3252 43002
rect 2956 42948 3012 42950
rect 3036 42948 3092 42950
rect 3116 42948 3172 42950
rect 3196 42948 3252 42950
rect 2956 41914 3012 41916
rect 3036 41914 3092 41916
rect 3116 41914 3172 41916
rect 3196 41914 3252 41916
rect 2956 41862 3002 41914
rect 3002 41862 3012 41914
rect 3036 41862 3066 41914
rect 3066 41862 3078 41914
rect 3078 41862 3092 41914
rect 3116 41862 3130 41914
rect 3130 41862 3142 41914
rect 3142 41862 3172 41914
rect 3196 41862 3206 41914
rect 3206 41862 3252 41914
rect 2956 41860 3012 41862
rect 3036 41860 3092 41862
rect 3116 41860 3172 41862
rect 3196 41860 3252 41862
rect 2956 40826 3012 40828
rect 3036 40826 3092 40828
rect 3116 40826 3172 40828
rect 3196 40826 3252 40828
rect 2956 40774 3002 40826
rect 3002 40774 3012 40826
rect 3036 40774 3066 40826
rect 3066 40774 3078 40826
rect 3078 40774 3092 40826
rect 3116 40774 3130 40826
rect 3130 40774 3142 40826
rect 3142 40774 3172 40826
rect 3196 40774 3206 40826
rect 3206 40774 3252 40826
rect 2956 40772 3012 40774
rect 3036 40772 3092 40774
rect 3116 40772 3172 40774
rect 3196 40772 3252 40774
rect 2956 39738 3012 39740
rect 3036 39738 3092 39740
rect 3116 39738 3172 39740
rect 3196 39738 3252 39740
rect 2956 39686 3002 39738
rect 3002 39686 3012 39738
rect 3036 39686 3066 39738
rect 3066 39686 3078 39738
rect 3078 39686 3092 39738
rect 3116 39686 3130 39738
rect 3130 39686 3142 39738
rect 3142 39686 3172 39738
rect 3196 39686 3206 39738
rect 3206 39686 3252 39738
rect 2956 39684 3012 39686
rect 3036 39684 3092 39686
rect 3116 39684 3172 39686
rect 3196 39684 3252 39686
rect 2956 38650 3012 38652
rect 3036 38650 3092 38652
rect 3116 38650 3172 38652
rect 3196 38650 3252 38652
rect 2956 38598 3002 38650
rect 3002 38598 3012 38650
rect 3036 38598 3066 38650
rect 3066 38598 3078 38650
rect 3078 38598 3092 38650
rect 3116 38598 3130 38650
rect 3130 38598 3142 38650
rect 3142 38598 3172 38650
rect 3196 38598 3206 38650
rect 3206 38598 3252 38650
rect 2956 38596 3012 38598
rect 3036 38596 3092 38598
rect 3116 38596 3172 38598
rect 3196 38596 3252 38598
rect 7956 45722 8012 45724
rect 8036 45722 8092 45724
rect 8116 45722 8172 45724
rect 8196 45722 8252 45724
rect 7956 45670 8002 45722
rect 8002 45670 8012 45722
rect 8036 45670 8066 45722
rect 8066 45670 8078 45722
rect 8078 45670 8092 45722
rect 8116 45670 8130 45722
rect 8130 45670 8142 45722
rect 8142 45670 8172 45722
rect 8196 45670 8206 45722
rect 8206 45670 8252 45722
rect 7956 45668 8012 45670
rect 8036 45668 8092 45670
rect 8116 45668 8172 45670
rect 8196 45668 8252 45670
rect 7956 44634 8012 44636
rect 8036 44634 8092 44636
rect 8116 44634 8172 44636
rect 8196 44634 8252 44636
rect 7956 44582 8002 44634
rect 8002 44582 8012 44634
rect 8036 44582 8066 44634
rect 8066 44582 8078 44634
rect 8078 44582 8092 44634
rect 8116 44582 8130 44634
rect 8130 44582 8142 44634
rect 8142 44582 8172 44634
rect 8196 44582 8206 44634
rect 8206 44582 8252 44634
rect 7956 44580 8012 44582
rect 8036 44580 8092 44582
rect 8116 44580 8172 44582
rect 8196 44580 8252 44582
rect 7956 43546 8012 43548
rect 8036 43546 8092 43548
rect 8116 43546 8172 43548
rect 8196 43546 8252 43548
rect 7956 43494 8002 43546
rect 8002 43494 8012 43546
rect 8036 43494 8066 43546
rect 8066 43494 8078 43546
rect 8078 43494 8092 43546
rect 8116 43494 8130 43546
rect 8130 43494 8142 43546
rect 8142 43494 8172 43546
rect 8196 43494 8206 43546
rect 8206 43494 8252 43546
rect 7956 43492 8012 43494
rect 8036 43492 8092 43494
rect 8116 43492 8172 43494
rect 8196 43492 8252 43494
rect 7956 42458 8012 42460
rect 8036 42458 8092 42460
rect 8116 42458 8172 42460
rect 8196 42458 8252 42460
rect 7956 42406 8002 42458
rect 8002 42406 8012 42458
rect 8036 42406 8066 42458
rect 8066 42406 8078 42458
rect 8078 42406 8092 42458
rect 8116 42406 8130 42458
rect 8130 42406 8142 42458
rect 8142 42406 8172 42458
rect 8196 42406 8206 42458
rect 8206 42406 8252 42458
rect 7956 42404 8012 42406
rect 8036 42404 8092 42406
rect 8116 42404 8172 42406
rect 8196 42404 8252 42406
rect 7956 41370 8012 41372
rect 8036 41370 8092 41372
rect 8116 41370 8172 41372
rect 8196 41370 8252 41372
rect 7956 41318 8002 41370
rect 8002 41318 8012 41370
rect 8036 41318 8066 41370
rect 8066 41318 8078 41370
rect 8078 41318 8092 41370
rect 8116 41318 8130 41370
rect 8130 41318 8142 41370
rect 8142 41318 8172 41370
rect 8196 41318 8206 41370
rect 8206 41318 8252 41370
rect 7956 41316 8012 41318
rect 8036 41316 8092 41318
rect 8116 41316 8172 41318
rect 8196 41316 8252 41318
rect 7956 40282 8012 40284
rect 8036 40282 8092 40284
rect 8116 40282 8172 40284
rect 8196 40282 8252 40284
rect 7956 40230 8002 40282
rect 8002 40230 8012 40282
rect 8036 40230 8066 40282
rect 8066 40230 8078 40282
rect 8078 40230 8092 40282
rect 8116 40230 8130 40282
rect 8130 40230 8142 40282
rect 8142 40230 8172 40282
rect 8196 40230 8206 40282
rect 8206 40230 8252 40282
rect 7956 40228 8012 40230
rect 8036 40228 8092 40230
rect 8116 40228 8172 40230
rect 8196 40228 8252 40230
rect 7956 39194 8012 39196
rect 8036 39194 8092 39196
rect 8116 39194 8172 39196
rect 8196 39194 8252 39196
rect 7956 39142 8002 39194
rect 8002 39142 8012 39194
rect 8036 39142 8066 39194
rect 8066 39142 8078 39194
rect 8078 39142 8092 39194
rect 8116 39142 8130 39194
rect 8130 39142 8142 39194
rect 8142 39142 8172 39194
rect 8196 39142 8206 39194
rect 8206 39142 8252 39194
rect 7956 39140 8012 39142
rect 8036 39140 8092 39142
rect 8116 39140 8172 39142
rect 8196 39140 8252 39142
rect 7956 38106 8012 38108
rect 8036 38106 8092 38108
rect 8116 38106 8172 38108
rect 8196 38106 8252 38108
rect 7956 38054 8002 38106
rect 8002 38054 8012 38106
rect 8036 38054 8066 38106
rect 8066 38054 8078 38106
rect 8078 38054 8092 38106
rect 8116 38054 8130 38106
rect 8130 38054 8142 38106
rect 8142 38054 8172 38106
rect 8196 38054 8206 38106
rect 8206 38054 8252 38106
rect 7956 38052 8012 38054
rect 8036 38052 8092 38054
rect 8116 38052 8172 38054
rect 8196 38052 8252 38054
rect 2956 37562 3012 37564
rect 3036 37562 3092 37564
rect 3116 37562 3172 37564
rect 3196 37562 3252 37564
rect 2956 37510 3002 37562
rect 3002 37510 3012 37562
rect 3036 37510 3066 37562
rect 3066 37510 3078 37562
rect 3078 37510 3092 37562
rect 3116 37510 3130 37562
rect 3130 37510 3142 37562
rect 3142 37510 3172 37562
rect 3196 37510 3206 37562
rect 3206 37510 3252 37562
rect 2956 37508 3012 37510
rect 3036 37508 3092 37510
rect 3116 37508 3172 37510
rect 3196 37508 3252 37510
rect 7956 37018 8012 37020
rect 8036 37018 8092 37020
rect 8116 37018 8172 37020
rect 8196 37018 8252 37020
rect 7956 36966 8002 37018
rect 8002 36966 8012 37018
rect 8036 36966 8066 37018
rect 8066 36966 8078 37018
rect 8078 36966 8092 37018
rect 8116 36966 8130 37018
rect 8130 36966 8142 37018
rect 8142 36966 8172 37018
rect 8196 36966 8206 37018
rect 8206 36966 8252 37018
rect 7956 36964 8012 36966
rect 8036 36964 8092 36966
rect 8116 36964 8172 36966
rect 8196 36964 8252 36966
rect 2956 36474 3012 36476
rect 3036 36474 3092 36476
rect 3116 36474 3172 36476
rect 3196 36474 3252 36476
rect 2956 36422 3002 36474
rect 3002 36422 3012 36474
rect 3036 36422 3066 36474
rect 3066 36422 3078 36474
rect 3078 36422 3092 36474
rect 3116 36422 3130 36474
rect 3130 36422 3142 36474
rect 3142 36422 3172 36474
rect 3196 36422 3206 36474
rect 3206 36422 3252 36474
rect 2956 36420 3012 36422
rect 3036 36420 3092 36422
rect 3116 36420 3172 36422
rect 3196 36420 3252 36422
rect 7956 35930 8012 35932
rect 8036 35930 8092 35932
rect 8116 35930 8172 35932
rect 8196 35930 8252 35932
rect 7956 35878 8002 35930
rect 8002 35878 8012 35930
rect 8036 35878 8066 35930
rect 8066 35878 8078 35930
rect 8078 35878 8092 35930
rect 8116 35878 8130 35930
rect 8130 35878 8142 35930
rect 8142 35878 8172 35930
rect 8196 35878 8206 35930
rect 8206 35878 8252 35930
rect 7956 35876 8012 35878
rect 8036 35876 8092 35878
rect 8116 35876 8172 35878
rect 8196 35876 8252 35878
rect 2956 35386 3012 35388
rect 3036 35386 3092 35388
rect 3116 35386 3172 35388
rect 3196 35386 3252 35388
rect 2956 35334 3002 35386
rect 3002 35334 3012 35386
rect 3036 35334 3066 35386
rect 3066 35334 3078 35386
rect 3078 35334 3092 35386
rect 3116 35334 3130 35386
rect 3130 35334 3142 35386
rect 3142 35334 3172 35386
rect 3196 35334 3206 35386
rect 3206 35334 3252 35386
rect 2956 35332 3012 35334
rect 3036 35332 3092 35334
rect 3116 35332 3172 35334
rect 3196 35332 3252 35334
rect 7956 34842 8012 34844
rect 8036 34842 8092 34844
rect 8116 34842 8172 34844
rect 8196 34842 8252 34844
rect 7956 34790 8002 34842
rect 8002 34790 8012 34842
rect 8036 34790 8066 34842
rect 8066 34790 8078 34842
rect 8078 34790 8092 34842
rect 8116 34790 8130 34842
rect 8130 34790 8142 34842
rect 8142 34790 8172 34842
rect 8196 34790 8206 34842
rect 8206 34790 8252 34842
rect 7956 34788 8012 34790
rect 8036 34788 8092 34790
rect 8116 34788 8172 34790
rect 8196 34788 8252 34790
rect 2956 34298 3012 34300
rect 3036 34298 3092 34300
rect 3116 34298 3172 34300
rect 3196 34298 3252 34300
rect 2956 34246 3002 34298
rect 3002 34246 3012 34298
rect 3036 34246 3066 34298
rect 3066 34246 3078 34298
rect 3078 34246 3092 34298
rect 3116 34246 3130 34298
rect 3130 34246 3142 34298
rect 3142 34246 3172 34298
rect 3196 34246 3206 34298
rect 3206 34246 3252 34298
rect 2956 34244 3012 34246
rect 3036 34244 3092 34246
rect 3116 34244 3172 34246
rect 3196 34244 3252 34246
rect 7956 33754 8012 33756
rect 8036 33754 8092 33756
rect 8116 33754 8172 33756
rect 8196 33754 8252 33756
rect 7956 33702 8002 33754
rect 8002 33702 8012 33754
rect 8036 33702 8066 33754
rect 8066 33702 8078 33754
rect 8078 33702 8092 33754
rect 8116 33702 8130 33754
rect 8130 33702 8142 33754
rect 8142 33702 8172 33754
rect 8196 33702 8206 33754
rect 8206 33702 8252 33754
rect 7956 33700 8012 33702
rect 8036 33700 8092 33702
rect 8116 33700 8172 33702
rect 8196 33700 8252 33702
rect 2956 33210 3012 33212
rect 3036 33210 3092 33212
rect 3116 33210 3172 33212
rect 3196 33210 3252 33212
rect 2956 33158 3002 33210
rect 3002 33158 3012 33210
rect 3036 33158 3066 33210
rect 3066 33158 3078 33210
rect 3078 33158 3092 33210
rect 3116 33158 3130 33210
rect 3130 33158 3142 33210
rect 3142 33158 3172 33210
rect 3196 33158 3206 33210
rect 3206 33158 3252 33210
rect 2956 33156 3012 33158
rect 3036 33156 3092 33158
rect 3116 33156 3172 33158
rect 3196 33156 3252 33158
rect 7956 32666 8012 32668
rect 8036 32666 8092 32668
rect 8116 32666 8172 32668
rect 8196 32666 8252 32668
rect 7956 32614 8002 32666
rect 8002 32614 8012 32666
rect 8036 32614 8066 32666
rect 8066 32614 8078 32666
rect 8078 32614 8092 32666
rect 8116 32614 8130 32666
rect 8130 32614 8142 32666
rect 8142 32614 8172 32666
rect 8196 32614 8206 32666
rect 8206 32614 8252 32666
rect 7956 32612 8012 32614
rect 8036 32612 8092 32614
rect 8116 32612 8172 32614
rect 8196 32612 8252 32614
rect 2956 32122 3012 32124
rect 3036 32122 3092 32124
rect 3116 32122 3172 32124
rect 3196 32122 3252 32124
rect 2956 32070 3002 32122
rect 3002 32070 3012 32122
rect 3036 32070 3066 32122
rect 3066 32070 3078 32122
rect 3078 32070 3092 32122
rect 3116 32070 3130 32122
rect 3130 32070 3142 32122
rect 3142 32070 3172 32122
rect 3196 32070 3206 32122
rect 3206 32070 3252 32122
rect 2956 32068 3012 32070
rect 3036 32068 3092 32070
rect 3116 32068 3172 32070
rect 3196 32068 3252 32070
rect 7956 31578 8012 31580
rect 8036 31578 8092 31580
rect 8116 31578 8172 31580
rect 8196 31578 8252 31580
rect 7956 31526 8002 31578
rect 8002 31526 8012 31578
rect 8036 31526 8066 31578
rect 8066 31526 8078 31578
rect 8078 31526 8092 31578
rect 8116 31526 8130 31578
rect 8130 31526 8142 31578
rect 8142 31526 8172 31578
rect 8196 31526 8206 31578
rect 8206 31526 8252 31578
rect 7956 31524 8012 31526
rect 8036 31524 8092 31526
rect 8116 31524 8172 31526
rect 8196 31524 8252 31526
rect 2956 31034 3012 31036
rect 3036 31034 3092 31036
rect 3116 31034 3172 31036
rect 3196 31034 3252 31036
rect 2956 30982 3002 31034
rect 3002 30982 3012 31034
rect 3036 30982 3066 31034
rect 3066 30982 3078 31034
rect 3078 30982 3092 31034
rect 3116 30982 3130 31034
rect 3130 30982 3142 31034
rect 3142 30982 3172 31034
rect 3196 30982 3206 31034
rect 3206 30982 3252 31034
rect 2956 30980 3012 30982
rect 3036 30980 3092 30982
rect 3116 30980 3172 30982
rect 3196 30980 3252 30982
rect 7956 30490 8012 30492
rect 8036 30490 8092 30492
rect 8116 30490 8172 30492
rect 8196 30490 8252 30492
rect 7956 30438 8002 30490
rect 8002 30438 8012 30490
rect 8036 30438 8066 30490
rect 8066 30438 8078 30490
rect 8078 30438 8092 30490
rect 8116 30438 8130 30490
rect 8130 30438 8142 30490
rect 8142 30438 8172 30490
rect 8196 30438 8206 30490
rect 8206 30438 8252 30490
rect 7956 30436 8012 30438
rect 8036 30436 8092 30438
rect 8116 30436 8172 30438
rect 8196 30436 8252 30438
rect 2956 29946 3012 29948
rect 3036 29946 3092 29948
rect 3116 29946 3172 29948
rect 3196 29946 3252 29948
rect 2956 29894 3002 29946
rect 3002 29894 3012 29946
rect 3036 29894 3066 29946
rect 3066 29894 3078 29946
rect 3078 29894 3092 29946
rect 3116 29894 3130 29946
rect 3130 29894 3142 29946
rect 3142 29894 3172 29946
rect 3196 29894 3206 29946
rect 3206 29894 3252 29946
rect 2956 29892 3012 29894
rect 3036 29892 3092 29894
rect 3116 29892 3172 29894
rect 3196 29892 3252 29894
rect 7956 29402 8012 29404
rect 8036 29402 8092 29404
rect 8116 29402 8172 29404
rect 8196 29402 8252 29404
rect 7956 29350 8002 29402
rect 8002 29350 8012 29402
rect 8036 29350 8066 29402
rect 8066 29350 8078 29402
rect 8078 29350 8092 29402
rect 8116 29350 8130 29402
rect 8130 29350 8142 29402
rect 8142 29350 8172 29402
rect 8196 29350 8206 29402
rect 8206 29350 8252 29402
rect 7956 29348 8012 29350
rect 8036 29348 8092 29350
rect 8116 29348 8172 29350
rect 8196 29348 8252 29350
rect 2956 28858 3012 28860
rect 3036 28858 3092 28860
rect 3116 28858 3172 28860
rect 3196 28858 3252 28860
rect 2956 28806 3002 28858
rect 3002 28806 3012 28858
rect 3036 28806 3066 28858
rect 3066 28806 3078 28858
rect 3078 28806 3092 28858
rect 3116 28806 3130 28858
rect 3130 28806 3142 28858
rect 3142 28806 3172 28858
rect 3196 28806 3206 28858
rect 3206 28806 3252 28858
rect 2956 28804 3012 28806
rect 3036 28804 3092 28806
rect 3116 28804 3172 28806
rect 3196 28804 3252 28806
rect 7956 28314 8012 28316
rect 8036 28314 8092 28316
rect 8116 28314 8172 28316
rect 8196 28314 8252 28316
rect 7956 28262 8002 28314
rect 8002 28262 8012 28314
rect 8036 28262 8066 28314
rect 8066 28262 8078 28314
rect 8078 28262 8092 28314
rect 8116 28262 8130 28314
rect 8130 28262 8142 28314
rect 8142 28262 8172 28314
rect 8196 28262 8206 28314
rect 8206 28262 8252 28314
rect 7956 28260 8012 28262
rect 8036 28260 8092 28262
rect 8116 28260 8172 28262
rect 8196 28260 8252 28262
rect 2956 27770 3012 27772
rect 3036 27770 3092 27772
rect 3116 27770 3172 27772
rect 3196 27770 3252 27772
rect 2956 27718 3002 27770
rect 3002 27718 3012 27770
rect 3036 27718 3066 27770
rect 3066 27718 3078 27770
rect 3078 27718 3092 27770
rect 3116 27718 3130 27770
rect 3130 27718 3142 27770
rect 3142 27718 3172 27770
rect 3196 27718 3206 27770
rect 3206 27718 3252 27770
rect 2956 27716 3012 27718
rect 3036 27716 3092 27718
rect 3116 27716 3172 27718
rect 3196 27716 3252 27718
rect 2956 26682 3012 26684
rect 3036 26682 3092 26684
rect 3116 26682 3172 26684
rect 3196 26682 3252 26684
rect 2956 26630 3002 26682
rect 3002 26630 3012 26682
rect 3036 26630 3066 26682
rect 3066 26630 3078 26682
rect 3078 26630 3092 26682
rect 3116 26630 3130 26682
rect 3130 26630 3142 26682
rect 3142 26630 3172 26682
rect 3196 26630 3206 26682
rect 3206 26630 3252 26682
rect 2956 26628 3012 26630
rect 3036 26628 3092 26630
rect 3116 26628 3172 26630
rect 3196 26628 3252 26630
rect 2956 25594 3012 25596
rect 3036 25594 3092 25596
rect 3116 25594 3172 25596
rect 3196 25594 3252 25596
rect 2956 25542 3002 25594
rect 3002 25542 3012 25594
rect 3036 25542 3066 25594
rect 3066 25542 3078 25594
rect 3078 25542 3092 25594
rect 3116 25542 3130 25594
rect 3130 25542 3142 25594
rect 3142 25542 3172 25594
rect 3196 25542 3206 25594
rect 3206 25542 3252 25594
rect 2956 25540 3012 25542
rect 3036 25540 3092 25542
rect 3116 25540 3172 25542
rect 3196 25540 3252 25542
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 7956 27226 8012 27228
rect 8036 27226 8092 27228
rect 8116 27226 8172 27228
rect 8196 27226 8252 27228
rect 7956 27174 8002 27226
rect 8002 27174 8012 27226
rect 8036 27174 8066 27226
rect 8066 27174 8078 27226
rect 8078 27174 8092 27226
rect 8116 27174 8130 27226
rect 8130 27174 8142 27226
rect 8142 27174 8172 27226
rect 8196 27174 8206 27226
rect 8206 27174 8252 27226
rect 7956 27172 8012 27174
rect 8036 27172 8092 27174
rect 8116 27172 8172 27174
rect 8196 27172 8252 27174
rect 7956 26138 8012 26140
rect 8036 26138 8092 26140
rect 8116 26138 8172 26140
rect 8196 26138 8252 26140
rect 7956 26086 8002 26138
rect 8002 26086 8012 26138
rect 8036 26086 8066 26138
rect 8066 26086 8078 26138
rect 8078 26086 8092 26138
rect 8116 26086 8130 26138
rect 8130 26086 8142 26138
rect 8142 26086 8172 26138
rect 8196 26086 8206 26138
rect 8206 26086 8252 26138
rect 7956 26084 8012 26086
rect 8036 26084 8092 26086
rect 8116 26084 8172 26086
rect 8196 26084 8252 26086
rect 7956 25050 8012 25052
rect 8036 25050 8092 25052
rect 8116 25050 8172 25052
rect 8196 25050 8252 25052
rect 7956 24998 8002 25050
rect 8002 24998 8012 25050
rect 8036 24998 8066 25050
rect 8066 24998 8078 25050
rect 8078 24998 8092 25050
rect 8116 24998 8130 25050
rect 8130 24998 8142 25050
rect 8142 24998 8172 25050
rect 8196 24998 8206 25050
rect 8206 24998 8252 25050
rect 7956 24996 8012 24998
rect 8036 24996 8092 24998
rect 8116 24996 8172 24998
rect 8196 24996 8252 24998
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 3514 8744 3570 8800
rect 3422 6432 3478 6488
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 5170 3596 5226 3632
rect 5170 3576 5172 3596
rect 5172 3576 5224 3596
rect 5224 3576 5226 3596
rect 5446 2508 5502 2544
rect 5446 2488 5448 2508
rect 5448 2488 5500 2508
rect 5500 2488 5502 2508
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 17956 54426 18012 54428
rect 18036 54426 18092 54428
rect 18116 54426 18172 54428
rect 18196 54426 18252 54428
rect 17956 54374 18002 54426
rect 18002 54374 18012 54426
rect 18036 54374 18066 54426
rect 18066 54374 18078 54426
rect 18078 54374 18092 54426
rect 18116 54374 18130 54426
rect 18130 54374 18142 54426
rect 18142 54374 18172 54426
rect 18196 54374 18206 54426
rect 18206 54374 18252 54426
rect 17956 54372 18012 54374
rect 18036 54372 18092 54374
rect 18116 54372 18172 54374
rect 18196 54372 18252 54374
rect 23386 56072 23442 56128
rect 12956 53882 13012 53884
rect 13036 53882 13092 53884
rect 13116 53882 13172 53884
rect 13196 53882 13252 53884
rect 12956 53830 13002 53882
rect 13002 53830 13012 53882
rect 13036 53830 13066 53882
rect 13066 53830 13078 53882
rect 13078 53830 13092 53882
rect 13116 53830 13130 53882
rect 13130 53830 13142 53882
rect 13142 53830 13172 53882
rect 13196 53830 13206 53882
rect 13206 53830 13252 53882
rect 12956 53828 13012 53830
rect 13036 53828 13092 53830
rect 13116 53828 13172 53830
rect 13196 53828 13252 53830
rect 12956 52794 13012 52796
rect 13036 52794 13092 52796
rect 13116 52794 13172 52796
rect 13196 52794 13252 52796
rect 12956 52742 13002 52794
rect 13002 52742 13012 52794
rect 13036 52742 13066 52794
rect 13066 52742 13078 52794
rect 13078 52742 13092 52794
rect 13116 52742 13130 52794
rect 13130 52742 13142 52794
rect 13142 52742 13172 52794
rect 13196 52742 13206 52794
rect 13206 52742 13252 52794
rect 12956 52740 13012 52742
rect 13036 52740 13092 52742
rect 13116 52740 13172 52742
rect 13196 52740 13252 52742
rect 12956 51706 13012 51708
rect 13036 51706 13092 51708
rect 13116 51706 13172 51708
rect 13196 51706 13252 51708
rect 12956 51654 13002 51706
rect 13002 51654 13012 51706
rect 13036 51654 13066 51706
rect 13066 51654 13078 51706
rect 13078 51654 13092 51706
rect 13116 51654 13130 51706
rect 13130 51654 13142 51706
rect 13142 51654 13172 51706
rect 13196 51654 13206 51706
rect 13206 51654 13252 51706
rect 12956 51652 13012 51654
rect 13036 51652 13092 51654
rect 13116 51652 13172 51654
rect 13196 51652 13252 51654
rect 12956 50618 13012 50620
rect 13036 50618 13092 50620
rect 13116 50618 13172 50620
rect 13196 50618 13252 50620
rect 12956 50566 13002 50618
rect 13002 50566 13012 50618
rect 13036 50566 13066 50618
rect 13066 50566 13078 50618
rect 13078 50566 13092 50618
rect 13116 50566 13130 50618
rect 13130 50566 13142 50618
rect 13142 50566 13172 50618
rect 13196 50566 13206 50618
rect 13206 50566 13252 50618
rect 12956 50564 13012 50566
rect 13036 50564 13092 50566
rect 13116 50564 13172 50566
rect 13196 50564 13252 50566
rect 12956 49530 13012 49532
rect 13036 49530 13092 49532
rect 13116 49530 13172 49532
rect 13196 49530 13252 49532
rect 12956 49478 13002 49530
rect 13002 49478 13012 49530
rect 13036 49478 13066 49530
rect 13066 49478 13078 49530
rect 13078 49478 13092 49530
rect 13116 49478 13130 49530
rect 13130 49478 13142 49530
rect 13142 49478 13172 49530
rect 13196 49478 13206 49530
rect 13206 49478 13252 49530
rect 12956 49476 13012 49478
rect 13036 49476 13092 49478
rect 13116 49476 13172 49478
rect 13196 49476 13252 49478
rect 12956 48442 13012 48444
rect 13036 48442 13092 48444
rect 13116 48442 13172 48444
rect 13196 48442 13252 48444
rect 12956 48390 13002 48442
rect 13002 48390 13012 48442
rect 13036 48390 13066 48442
rect 13066 48390 13078 48442
rect 13078 48390 13092 48442
rect 13116 48390 13130 48442
rect 13130 48390 13142 48442
rect 13142 48390 13172 48442
rect 13196 48390 13206 48442
rect 13206 48390 13252 48442
rect 12956 48388 13012 48390
rect 13036 48388 13092 48390
rect 13116 48388 13172 48390
rect 13196 48388 13252 48390
rect 12956 47354 13012 47356
rect 13036 47354 13092 47356
rect 13116 47354 13172 47356
rect 13196 47354 13252 47356
rect 12956 47302 13002 47354
rect 13002 47302 13012 47354
rect 13036 47302 13066 47354
rect 13066 47302 13078 47354
rect 13078 47302 13092 47354
rect 13116 47302 13130 47354
rect 13130 47302 13142 47354
rect 13142 47302 13172 47354
rect 13196 47302 13206 47354
rect 13206 47302 13252 47354
rect 12956 47300 13012 47302
rect 13036 47300 13092 47302
rect 13116 47300 13172 47302
rect 13196 47300 13252 47302
rect 12956 46266 13012 46268
rect 13036 46266 13092 46268
rect 13116 46266 13172 46268
rect 13196 46266 13252 46268
rect 12956 46214 13002 46266
rect 13002 46214 13012 46266
rect 13036 46214 13066 46266
rect 13066 46214 13078 46266
rect 13078 46214 13092 46266
rect 13116 46214 13130 46266
rect 13130 46214 13142 46266
rect 13142 46214 13172 46266
rect 13196 46214 13206 46266
rect 13206 46214 13252 46266
rect 12956 46212 13012 46214
rect 13036 46212 13092 46214
rect 13116 46212 13172 46214
rect 13196 46212 13252 46214
rect 12956 45178 13012 45180
rect 13036 45178 13092 45180
rect 13116 45178 13172 45180
rect 13196 45178 13252 45180
rect 12956 45126 13002 45178
rect 13002 45126 13012 45178
rect 13036 45126 13066 45178
rect 13066 45126 13078 45178
rect 13078 45126 13092 45178
rect 13116 45126 13130 45178
rect 13130 45126 13142 45178
rect 13142 45126 13172 45178
rect 13196 45126 13206 45178
rect 13206 45126 13252 45178
rect 12956 45124 13012 45126
rect 13036 45124 13092 45126
rect 13116 45124 13172 45126
rect 13196 45124 13252 45126
rect 12956 44090 13012 44092
rect 13036 44090 13092 44092
rect 13116 44090 13172 44092
rect 13196 44090 13252 44092
rect 12956 44038 13002 44090
rect 13002 44038 13012 44090
rect 13036 44038 13066 44090
rect 13066 44038 13078 44090
rect 13078 44038 13092 44090
rect 13116 44038 13130 44090
rect 13130 44038 13142 44090
rect 13142 44038 13172 44090
rect 13196 44038 13206 44090
rect 13206 44038 13252 44090
rect 12956 44036 13012 44038
rect 13036 44036 13092 44038
rect 13116 44036 13172 44038
rect 13196 44036 13252 44038
rect 12956 43002 13012 43004
rect 13036 43002 13092 43004
rect 13116 43002 13172 43004
rect 13196 43002 13252 43004
rect 12956 42950 13002 43002
rect 13002 42950 13012 43002
rect 13036 42950 13066 43002
rect 13066 42950 13078 43002
rect 13078 42950 13092 43002
rect 13116 42950 13130 43002
rect 13130 42950 13142 43002
rect 13142 42950 13172 43002
rect 13196 42950 13206 43002
rect 13206 42950 13252 43002
rect 12956 42948 13012 42950
rect 13036 42948 13092 42950
rect 13116 42948 13172 42950
rect 13196 42948 13252 42950
rect 12956 41914 13012 41916
rect 13036 41914 13092 41916
rect 13116 41914 13172 41916
rect 13196 41914 13252 41916
rect 12956 41862 13002 41914
rect 13002 41862 13012 41914
rect 13036 41862 13066 41914
rect 13066 41862 13078 41914
rect 13078 41862 13092 41914
rect 13116 41862 13130 41914
rect 13130 41862 13142 41914
rect 13142 41862 13172 41914
rect 13196 41862 13206 41914
rect 13206 41862 13252 41914
rect 12956 41860 13012 41862
rect 13036 41860 13092 41862
rect 13116 41860 13172 41862
rect 13196 41860 13252 41862
rect 12956 40826 13012 40828
rect 13036 40826 13092 40828
rect 13116 40826 13172 40828
rect 13196 40826 13252 40828
rect 12956 40774 13002 40826
rect 13002 40774 13012 40826
rect 13036 40774 13066 40826
rect 13066 40774 13078 40826
rect 13078 40774 13092 40826
rect 13116 40774 13130 40826
rect 13130 40774 13142 40826
rect 13142 40774 13172 40826
rect 13196 40774 13206 40826
rect 13206 40774 13252 40826
rect 12956 40772 13012 40774
rect 13036 40772 13092 40774
rect 13116 40772 13172 40774
rect 13196 40772 13252 40774
rect 12956 39738 13012 39740
rect 13036 39738 13092 39740
rect 13116 39738 13172 39740
rect 13196 39738 13252 39740
rect 12956 39686 13002 39738
rect 13002 39686 13012 39738
rect 13036 39686 13066 39738
rect 13066 39686 13078 39738
rect 13078 39686 13092 39738
rect 13116 39686 13130 39738
rect 13130 39686 13142 39738
rect 13142 39686 13172 39738
rect 13196 39686 13206 39738
rect 13206 39686 13252 39738
rect 12956 39684 13012 39686
rect 13036 39684 13092 39686
rect 13116 39684 13172 39686
rect 13196 39684 13252 39686
rect 12956 38650 13012 38652
rect 13036 38650 13092 38652
rect 13116 38650 13172 38652
rect 13196 38650 13252 38652
rect 12956 38598 13002 38650
rect 13002 38598 13012 38650
rect 13036 38598 13066 38650
rect 13066 38598 13078 38650
rect 13078 38598 13092 38650
rect 13116 38598 13130 38650
rect 13130 38598 13142 38650
rect 13142 38598 13172 38650
rect 13196 38598 13206 38650
rect 13206 38598 13252 38650
rect 12956 38596 13012 38598
rect 13036 38596 13092 38598
rect 13116 38596 13172 38598
rect 13196 38596 13252 38598
rect 12956 37562 13012 37564
rect 13036 37562 13092 37564
rect 13116 37562 13172 37564
rect 13196 37562 13252 37564
rect 12956 37510 13002 37562
rect 13002 37510 13012 37562
rect 13036 37510 13066 37562
rect 13066 37510 13078 37562
rect 13078 37510 13092 37562
rect 13116 37510 13130 37562
rect 13130 37510 13142 37562
rect 13142 37510 13172 37562
rect 13196 37510 13206 37562
rect 13206 37510 13252 37562
rect 12956 37508 13012 37510
rect 13036 37508 13092 37510
rect 13116 37508 13172 37510
rect 13196 37508 13252 37510
rect 12956 36474 13012 36476
rect 13036 36474 13092 36476
rect 13116 36474 13172 36476
rect 13196 36474 13252 36476
rect 12956 36422 13002 36474
rect 13002 36422 13012 36474
rect 13036 36422 13066 36474
rect 13066 36422 13078 36474
rect 13078 36422 13092 36474
rect 13116 36422 13130 36474
rect 13130 36422 13142 36474
rect 13142 36422 13172 36474
rect 13196 36422 13206 36474
rect 13206 36422 13252 36474
rect 12956 36420 13012 36422
rect 13036 36420 13092 36422
rect 13116 36420 13172 36422
rect 13196 36420 13252 36422
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 12956 35386 13012 35388
rect 13036 35386 13092 35388
rect 13116 35386 13172 35388
rect 13196 35386 13252 35388
rect 12956 35334 13002 35386
rect 13002 35334 13012 35386
rect 13036 35334 13066 35386
rect 13066 35334 13078 35386
rect 13078 35334 13092 35386
rect 13116 35334 13130 35386
rect 13130 35334 13142 35386
rect 13142 35334 13172 35386
rect 13196 35334 13206 35386
rect 13206 35334 13252 35386
rect 12956 35332 13012 35334
rect 13036 35332 13092 35334
rect 13116 35332 13172 35334
rect 13196 35332 13252 35334
rect 12956 34298 13012 34300
rect 13036 34298 13092 34300
rect 13116 34298 13172 34300
rect 13196 34298 13252 34300
rect 12956 34246 13002 34298
rect 13002 34246 13012 34298
rect 13036 34246 13066 34298
rect 13066 34246 13078 34298
rect 13078 34246 13092 34298
rect 13116 34246 13130 34298
rect 13130 34246 13142 34298
rect 13142 34246 13172 34298
rect 13196 34246 13206 34298
rect 13206 34246 13252 34298
rect 12956 34244 13012 34246
rect 13036 34244 13092 34246
rect 13116 34244 13172 34246
rect 13196 34244 13252 34246
rect 12956 33210 13012 33212
rect 13036 33210 13092 33212
rect 13116 33210 13172 33212
rect 13196 33210 13252 33212
rect 12956 33158 13002 33210
rect 13002 33158 13012 33210
rect 13036 33158 13066 33210
rect 13066 33158 13078 33210
rect 13078 33158 13092 33210
rect 13116 33158 13130 33210
rect 13130 33158 13142 33210
rect 13142 33158 13172 33210
rect 13196 33158 13206 33210
rect 13206 33158 13252 33210
rect 12956 33156 13012 33158
rect 13036 33156 13092 33158
rect 13116 33156 13172 33158
rect 13196 33156 13252 33158
rect 12956 32122 13012 32124
rect 13036 32122 13092 32124
rect 13116 32122 13172 32124
rect 13196 32122 13252 32124
rect 12956 32070 13002 32122
rect 13002 32070 13012 32122
rect 13036 32070 13066 32122
rect 13066 32070 13078 32122
rect 13078 32070 13092 32122
rect 13116 32070 13130 32122
rect 13130 32070 13142 32122
rect 13142 32070 13172 32122
rect 13196 32070 13206 32122
rect 13206 32070 13252 32122
rect 12956 32068 13012 32070
rect 13036 32068 13092 32070
rect 13116 32068 13172 32070
rect 13196 32068 13252 32070
rect 12956 31034 13012 31036
rect 13036 31034 13092 31036
rect 13116 31034 13172 31036
rect 13196 31034 13252 31036
rect 12956 30982 13002 31034
rect 13002 30982 13012 31034
rect 13036 30982 13066 31034
rect 13066 30982 13078 31034
rect 13078 30982 13092 31034
rect 13116 30982 13130 31034
rect 13130 30982 13142 31034
rect 13142 30982 13172 31034
rect 13196 30982 13206 31034
rect 13206 30982 13252 31034
rect 12956 30980 13012 30982
rect 13036 30980 13092 30982
rect 13116 30980 13172 30982
rect 13196 30980 13252 30982
rect 12956 29946 13012 29948
rect 13036 29946 13092 29948
rect 13116 29946 13172 29948
rect 13196 29946 13252 29948
rect 12956 29894 13002 29946
rect 13002 29894 13012 29946
rect 13036 29894 13066 29946
rect 13066 29894 13078 29946
rect 13078 29894 13092 29946
rect 13116 29894 13130 29946
rect 13130 29894 13142 29946
rect 13142 29894 13172 29946
rect 13196 29894 13206 29946
rect 13206 29894 13252 29946
rect 12956 29892 13012 29894
rect 13036 29892 13092 29894
rect 13116 29892 13172 29894
rect 13196 29892 13252 29894
rect 12956 28858 13012 28860
rect 13036 28858 13092 28860
rect 13116 28858 13172 28860
rect 13196 28858 13252 28860
rect 12956 28806 13002 28858
rect 13002 28806 13012 28858
rect 13036 28806 13066 28858
rect 13066 28806 13078 28858
rect 13078 28806 13092 28858
rect 13116 28806 13130 28858
rect 13130 28806 13142 28858
rect 13142 28806 13172 28858
rect 13196 28806 13206 28858
rect 13206 28806 13252 28858
rect 12956 28804 13012 28806
rect 13036 28804 13092 28806
rect 13116 28804 13172 28806
rect 13196 28804 13252 28806
rect 12956 27770 13012 27772
rect 13036 27770 13092 27772
rect 13116 27770 13172 27772
rect 13196 27770 13252 27772
rect 12956 27718 13002 27770
rect 13002 27718 13012 27770
rect 13036 27718 13066 27770
rect 13066 27718 13078 27770
rect 13078 27718 13092 27770
rect 13116 27718 13130 27770
rect 13130 27718 13142 27770
rect 13142 27718 13172 27770
rect 13196 27718 13206 27770
rect 13206 27718 13252 27770
rect 12956 27716 13012 27718
rect 13036 27716 13092 27718
rect 13116 27716 13172 27718
rect 13196 27716 13252 27718
rect 12956 26682 13012 26684
rect 13036 26682 13092 26684
rect 13116 26682 13172 26684
rect 13196 26682 13252 26684
rect 12956 26630 13002 26682
rect 13002 26630 13012 26682
rect 13036 26630 13066 26682
rect 13066 26630 13078 26682
rect 13078 26630 13092 26682
rect 13116 26630 13130 26682
rect 13130 26630 13142 26682
rect 13142 26630 13172 26682
rect 13196 26630 13206 26682
rect 13206 26630 13252 26682
rect 12956 26628 13012 26630
rect 13036 26628 13092 26630
rect 13116 26628 13172 26630
rect 13196 26628 13252 26630
rect 12956 25594 13012 25596
rect 13036 25594 13092 25596
rect 13116 25594 13172 25596
rect 13196 25594 13252 25596
rect 12956 25542 13002 25594
rect 13002 25542 13012 25594
rect 13036 25542 13066 25594
rect 13066 25542 13078 25594
rect 13078 25542 13092 25594
rect 13116 25542 13130 25594
rect 13130 25542 13142 25594
rect 13142 25542 13172 25594
rect 13196 25542 13206 25594
rect 13206 25542 13252 25594
rect 12956 25540 13012 25542
rect 13036 25540 13092 25542
rect 13116 25540 13172 25542
rect 13196 25540 13252 25542
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 10874 6196 10876 6216
rect 10876 6196 10928 6216
rect 10928 6196 10930 6216
rect 10874 6160 10930 6196
rect 11794 11872 11850 11928
rect 11886 11212 11942 11248
rect 11886 11192 11888 11212
rect 11888 11192 11940 11212
rect 11940 11192 11942 11212
rect 10966 3984 11022 4040
rect 12070 11756 12126 11792
rect 12070 11736 12072 11756
rect 12072 11736 12124 11756
rect 12124 11736 12126 11756
rect 12438 12416 12494 12472
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12714 17484 12716 17504
rect 12716 17484 12768 17504
rect 12768 17484 12770 17504
rect 12714 17448 12770 17484
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 17956 53338 18012 53340
rect 18036 53338 18092 53340
rect 18116 53338 18172 53340
rect 18196 53338 18252 53340
rect 17956 53286 18002 53338
rect 18002 53286 18012 53338
rect 18036 53286 18066 53338
rect 18066 53286 18078 53338
rect 18078 53286 18092 53338
rect 18116 53286 18130 53338
rect 18130 53286 18142 53338
rect 18142 53286 18172 53338
rect 18196 53286 18206 53338
rect 18206 53286 18252 53338
rect 17956 53284 18012 53286
rect 18036 53284 18092 53286
rect 18116 53284 18172 53286
rect 18196 53284 18252 53286
rect 17956 52250 18012 52252
rect 18036 52250 18092 52252
rect 18116 52250 18172 52252
rect 18196 52250 18252 52252
rect 17956 52198 18002 52250
rect 18002 52198 18012 52250
rect 18036 52198 18066 52250
rect 18066 52198 18078 52250
rect 18078 52198 18092 52250
rect 18116 52198 18130 52250
rect 18130 52198 18142 52250
rect 18142 52198 18172 52250
rect 18196 52198 18206 52250
rect 18206 52198 18252 52250
rect 17956 52196 18012 52198
rect 18036 52196 18092 52198
rect 18116 52196 18172 52198
rect 18196 52196 18252 52198
rect 17956 51162 18012 51164
rect 18036 51162 18092 51164
rect 18116 51162 18172 51164
rect 18196 51162 18252 51164
rect 17956 51110 18002 51162
rect 18002 51110 18012 51162
rect 18036 51110 18066 51162
rect 18066 51110 18078 51162
rect 18078 51110 18092 51162
rect 18116 51110 18130 51162
rect 18130 51110 18142 51162
rect 18142 51110 18172 51162
rect 18196 51110 18206 51162
rect 18206 51110 18252 51162
rect 17956 51108 18012 51110
rect 18036 51108 18092 51110
rect 18116 51108 18172 51110
rect 18196 51108 18252 51110
rect 17956 50074 18012 50076
rect 18036 50074 18092 50076
rect 18116 50074 18172 50076
rect 18196 50074 18252 50076
rect 17956 50022 18002 50074
rect 18002 50022 18012 50074
rect 18036 50022 18066 50074
rect 18066 50022 18078 50074
rect 18078 50022 18092 50074
rect 18116 50022 18130 50074
rect 18130 50022 18142 50074
rect 18142 50022 18172 50074
rect 18196 50022 18206 50074
rect 18206 50022 18252 50074
rect 17956 50020 18012 50022
rect 18036 50020 18092 50022
rect 18116 50020 18172 50022
rect 18196 50020 18252 50022
rect 17956 48986 18012 48988
rect 18036 48986 18092 48988
rect 18116 48986 18172 48988
rect 18196 48986 18252 48988
rect 17956 48934 18002 48986
rect 18002 48934 18012 48986
rect 18036 48934 18066 48986
rect 18066 48934 18078 48986
rect 18078 48934 18092 48986
rect 18116 48934 18130 48986
rect 18130 48934 18142 48986
rect 18142 48934 18172 48986
rect 18196 48934 18206 48986
rect 18206 48934 18252 48986
rect 17956 48932 18012 48934
rect 18036 48932 18092 48934
rect 18116 48932 18172 48934
rect 18196 48932 18252 48934
rect 17956 47898 18012 47900
rect 18036 47898 18092 47900
rect 18116 47898 18172 47900
rect 18196 47898 18252 47900
rect 17956 47846 18002 47898
rect 18002 47846 18012 47898
rect 18036 47846 18066 47898
rect 18066 47846 18078 47898
rect 18078 47846 18092 47898
rect 18116 47846 18130 47898
rect 18130 47846 18142 47898
rect 18142 47846 18172 47898
rect 18196 47846 18206 47898
rect 18206 47846 18252 47898
rect 17956 47844 18012 47846
rect 18036 47844 18092 47846
rect 18116 47844 18172 47846
rect 18196 47844 18252 47846
rect 17956 46810 18012 46812
rect 18036 46810 18092 46812
rect 18116 46810 18172 46812
rect 18196 46810 18252 46812
rect 17956 46758 18002 46810
rect 18002 46758 18012 46810
rect 18036 46758 18066 46810
rect 18066 46758 18078 46810
rect 18078 46758 18092 46810
rect 18116 46758 18130 46810
rect 18130 46758 18142 46810
rect 18142 46758 18172 46810
rect 18196 46758 18206 46810
rect 18206 46758 18252 46810
rect 17956 46756 18012 46758
rect 18036 46756 18092 46758
rect 18116 46756 18172 46758
rect 18196 46756 18252 46758
rect 17956 45722 18012 45724
rect 18036 45722 18092 45724
rect 18116 45722 18172 45724
rect 18196 45722 18252 45724
rect 17956 45670 18002 45722
rect 18002 45670 18012 45722
rect 18036 45670 18066 45722
rect 18066 45670 18078 45722
rect 18078 45670 18092 45722
rect 18116 45670 18130 45722
rect 18130 45670 18142 45722
rect 18142 45670 18172 45722
rect 18196 45670 18206 45722
rect 18206 45670 18252 45722
rect 17956 45668 18012 45670
rect 18036 45668 18092 45670
rect 18116 45668 18172 45670
rect 18196 45668 18252 45670
rect 17956 44634 18012 44636
rect 18036 44634 18092 44636
rect 18116 44634 18172 44636
rect 18196 44634 18252 44636
rect 17956 44582 18002 44634
rect 18002 44582 18012 44634
rect 18036 44582 18066 44634
rect 18066 44582 18078 44634
rect 18078 44582 18092 44634
rect 18116 44582 18130 44634
rect 18130 44582 18142 44634
rect 18142 44582 18172 44634
rect 18196 44582 18206 44634
rect 18206 44582 18252 44634
rect 17956 44580 18012 44582
rect 18036 44580 18092 44582
rect 18116 44580 18172 44582
rect 18196 44580 18252 44582
rect 17956 43546 18012 43548
rect 18036 43546 18092 43548
rect 18116 43546 18172 43548
rect 18196 43546 18252 43548
rect 17956 43494 18002 43546
rect 18002 43494 18012 43546
rect 18036 43494 18066 43546
rect 18066 43494 18078 43546
rect 18078 43494 18092 43546
rect 18116 43494 18130 43546
rect 18130 43494 18142 43546
rect 18142 43494 18172 43546
rect 18196 43494 18206 43546
rect 18206 43494 18252 43546
rect 17956 43492 18012 43494
rect 18036 43492 18092 43494
rect 18116 43492 18172 43494
rect 18196 43492 18252 43494
rect 17956 42458 18012 42460
rect 18036 42458 18092 42460
rect 18116 42458 18172 42460
rect 18196 42458 18252 42460
rect 17956 42406 18002 42458
rect 18002 42406 18012 42458
rect 18036 42406 18066 42458
rect 18066 42406 18078 42458
rect 18078 42406 18092 42458
rect 18116 42406 18130 42458
rect 18130 42406 18142 42458
rect 18142 42406 18172 42458
rect 18196 42406 18206 42458
rect 18206 42406 18252 42458
rect 17956 42404 18012 42406
rect 18036 42404 18092 42406
rect 18116 42404 18172 42406
rect 18196 42404 18252 42406
rect 17956 41370 18012 41372
rect 18036 41370 18092 41372
rect 18116 41370 18172 41372
rect 18196 41370 18252 41372
rect 17956 41318 18002 41370
rect 18002 41318 18012 41370
rect 18036 41318 18066 41370
rect 18066 41318 18078 41370
rect 18078 41318 18092 41370
rect 18116 41318 18130 41370
rect 18130 41318 18142 41370
rect 18142 41318 18172 41370
rect 18196 41318 18206 41370
rect 18206 41318 18252 41370
rect 17956 41316 18012 41318
rect 18036 41316 18092 41318
rect 18116 41316 18172 41318
rect 18196 41316 18252 41318
rect 17956 40282 18012 40284
rect 18036 40282 18092 40284
rect 18116 40282 18172 40284
rect 18196 40282 18252 40284
rect 17956 40230 18002 40282
rect 18002 40230 18012 40282
rect 18036 40230 18066 40282
rect 18066 40230 18078 40282
rect 18078 40230 18092 40282
rect 18116 40230 18130 40282
rect 18130 40230 18142 40282
rect 18142 40230 18172 40282
rect 18196 40230 18206 40282
rect 18206 40230 18252 40282
rect 17956 40228 18012 40230
rect 18036 40228 18092 40230
rect 18116 40228 18172 40230
rect 18196 40228 18252 40230
rect 17956 39194 18012 39196
rect 18036 39194 18092 39196
rect 18116 39194 18172 39196
rect 18196 39194 18252 39196
rect 17956 39142 18002 39194
rect 18002 39142 18012 39194
rect 18036 39142 18066 39194
rect 18066 39142 18078 39194
rect 18078 39142 18092 39194
rect 18116 39142 18130 39194
rect 18130 39142 18142 39194
rect 18142 39142 18172 39194
rect 18196 39142 18206 39194
rect 18206 39142 18252 39194
rect 17956 39140 18012 39142
rect 18036 39140 18092 39142
rect 18116 39140 18172 39142
rect 18196 39140 18252 39142
rect 17956 38106 18012 38108
rect 18036 38106 18092 38108
rect 18116 38106 18172 38108
rect 18196 38106 18252 38108
rect 17956 38054 18002 38106
rect 18002 38054 18012 38106
rect 18036 38054 18066 38106
rect 18066 38054 18078 38106
rect 18078 38054 18092 38106
rect 18116 38054 18130 38106
rect 18130 38054 18142 38106
rect 18142 38054 18172 38106
rect 18196 38054 18206 38106
rect 18206 38054 18252 38106
rect 17956 38052 18012 38054
rect 18036 38052 18092 38054
rect 18116 38052 18172 38054
rect 18196 38052 18252 38054
rect 17956 37018 18012 37020
rect 18036 37018 18092 37020
rect 18116 37018 18172 37020
rect 18196 37018 18252 37020
rect 17956 36966 18002 37018
rect 18002 36966 18012 37018
rect 18036 36966 18066 37018
rect 18066 36966 18078 37018
rect 18078 36966 18092 37018
rect 18116 36966 18130 37018
rect 18130 36966 18142 37018
rect 18142 36966 18172 37018
rect 18196 36966 18206 37018
rect 18206 36966 18252 37018
rect 17956 36964 18012 36966
rect 18036 36964 18092 36966
rect 18116 36964 18172 36966
rect 18196 36964 18252 36966
rect 17956 35930 18012 35932
rect 18036 35930 18092 35932
rect 18116 35930 18172 35932
rect 18196 35930 18252 35932
rect 17956 35878 18002 35930
rect 18002 35878 18012 35930
rect 18036 35878 18066 35930
rect 18066 35878 18078 35930
rect 18078 35878 18092 35930
rect 18116 35878 18130 35930
rect 18130 35878 18142 35930
rect 18142 35878 18172 35930
rect 18196 35878 18206 35930
rect 18206 35878 18252 35930
rect 17956 35876 18012 35878
rect 18036 35876 18092 35878
rect 18116 35876 18172 35878
rect 18196 35876 18252 35878
rect 17956 34842 18012 34844
rect 18036 34842 18092 34844
rect 18116 34842 18172 34844
rect 18196 34842 18252 34844
rect 17956 34790 18002 34842
rect 18002 34790 18012 34842
rect 18036 34790 18066 34842
rect 18066 34790 18078 34842
rect 18078 34790 18092 34842
rect 18116 34790 18130 34842
rect 18130 34790 18142 34842
rect 18142 34790 18172 34842
rect 18196 34790 18206 34842
rect 18206 34790 18252 34842
rect 17956 34788 18012 34790
rect 18036 34788 18092 34790
rect 18116 34788 18172 34790
rect 18196 34788 18252 34790
rect 17956 33754 18012 33756
rect 18036 33754 18092 33756
rect 18116 33754 18172 33756
rect 18196 33754 18252 33756
rect 17956 33702 18002 33754
rect 18002 33702 18012 33754
rect 18036 33702 18066 33754
rect 18066 33702 18078 33754
rect 18078 33702 18092 33754
rect 18116 33702 18130 33754
rect 18130 33702 18142 33754
rect 18142 33702 18172 33754
rect 18196 33702 18206 33754
rect 18206 33702 18252 33754
rect 17956 33700 18012 33702
rect 18036 33700 18092 33702
rect 18116 33700 18172 33702
rect 18196 33700 18252 33702
rect 15842 29008 15898 29064
rect 15566 25064 15622 25120
rect 12346 11772 12348 11792
rect 12348 11772 12400 11792
rect 12400 11772 12402 11792
rect 12346 11736 12402 11772
rect 12254 4700 12256 4720
rect 12256 4700 12308 4720
rect 12308 4700 12310 4720
rect 12254 4664 12310 4700
rect 12254 4528 12310 4584
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 13082 12688 13138 12744
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 13174 11228 13176 11248
rect 13176 11228 13228 11248
rect 13228 11228 13230 11248
rect 13174 11192 13230 11228
rect 13542 14220 13544 14240
rect 13544 14220 13596 14240
rect 13596 14220 13598 14240
rect 13542 14184 13598 14220
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 13266 6840 13322 6896
rect 12898 6196 12900 6216
rect 12900 6196 12952 6216
rect 12952 6196 12954 6216
rect 12898 6160 12954 6196
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 13542 8880 13598 8936
rect 13910 7792 13966 7848
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 13174 3052 13230 3088
rect 13174 3032 13176 3052
rect 13176 3032 13228 3052
rect 13228 3032 13230 3052
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 14738 14220 14740 14240
rect 14740 14220 14792 14240
rect 14792 14220 14794 14240
rect 14738 14184 14794 14220
rect 14554 12416 14610 12472
rect 14922 12416 14978 12472
rect 14186 10512 14242 10568
rect 15290 11872 15346 11928
rect 15014 10648 15070 10704
rect 14554 7948 14610 7984
rect 14554 7928 14556 7948
rect 14556 7928 14608 7948
rect 14608 7928 14610 7948
rect 14462 3576 14518 3632
rect 15198 7928 15254 7984
rect 14830 3712 14886 3768
rect 15474 7248 15530 7304
rect 15474 6160 15530 6216
rect 17956 32666 18012 32668
rect 18036 32666 18092 32668
rect 18116 32666 18172 32668
rect 18196 32666 18252 32668
rect 17956 32614 18002 32666
rect 18002 32614 18012 32666
rect 18036 32614 18066 32666
rect 18066 32614 18078 32666
rect 18078 32614 18092 32666
rect 18116 32614 18130 32666
rect 18130 32614 18142 32666
rect 18142 32614 18172 32666
rect 18196 32614 18206 32666
rect 18206 32614 18252 32666
rect 17956 32612 18012 32614
rect 18036 32612 18092 32614
rect 18116 32612 18172 32614
rect 18196 32612 18252 32614
rect 17956 31578 18012 31580
rect 18036 31578 18092 31580
rect 18116 31578 18172 31580
rect 18196 31578 18252 31580
rect 17956 31526 18002 31578
rect 18002 31526 18012 31578
rect 18036 31526 18066 31578
rect 18066 31526 18078 31578
rect 18078 31526 18092 31578
rect 18116 31526 18130 31578
rect 18130 31526 18142 31578
rect 18142 31526 18172 31578
rect 18196 31526 18206 31578
rect 18206 31526 18252 31578
rect 17956 31524 18012 31526
rect 18036 31524 18092 31526
rect 18116 31524 18172 31526
rect 18196 31524 18252 31526
rect 17406 29044 17408 29064
rect 17408 29044 17460 29064
rect 17460 29044 17462 29064
rect 16762 22752 16818 22808
rect 16026 11192 16082 11248
rect 16302 12416 16358 12472
rect 16302 11192 16358 11248
rect 15934 8880 15990 8936
rect 17406 29008 17462 29044
rect 16854 17992 16910 18048
rect 16854 16244 16910 16280
rect 16854 16224 16856 16244
rect 16856 16224 16908 16244
rect 16908 16224 16910 16244
rect 17590 25900 17646 25936
rect 17590 25880 17592 25900
rect 17592 25880 17644 25900
rect 17644 25880 17646 25900
rect 17956 30490 18012 30492
rect 18036 30490 18092 30492
rect 18116 30490 18172 30492
rect 18196 30490 18252 30492
rect 17956 30438 18002 30490
rect 18002 30438 18012 30490
rect 18036 30438 18066 30490
rect 18066 30438 18078 30490
rect 18078 30438 18092 30490
rect 18116 30438 18130 30490
rect 18130 30438 18142 30490
rect 18142 30438 18172 30490
rect 18196 30438 18206 30490
rect 18206 30438 18252 30490
rect 17956 30436 18012 30438
rect 18036 30436 18092 30438
rect 18116 30436 18172 30438
rect 18196 30436 18252 30438
rect 17956 29402 18012 29404
rect 18036 29402 18092 29404
rect 18116 29402 18172 29404
rect 18196 29402 18252 29404
rect 17956 29350 18002 29402
rect 18002 29350 18012 29402
rect 18036 29350 18066 29402
rect 18066 29350 18078 29402
rect 18078 29350 18092 29402
rect 18116 29350 18130 29402
rect 18130 29350 18142 29402
rect 18142 29350 18172 29402
rect 18196 29350 18206 29402
rect 18206 29350 18252 29402
rect 17956 29348 18012 29350
rect 18036 29348 18092 29350
rect 18116 29348 18172 29350
rect 18196 29348 18252 29350
rect 17956 28314 18012 28316
rect 18036 28314 18092 28316
rect 18116 28314 18172 28316
rect 18196 28314 18252 28316
rect 17956 28262 18002 28314
rect 18002 28262 18012 28314
rect 18036 28262 18066 28314
rect 18066 28262 18078 28314
rect 18078 28262 18092 28314
rect 18116 28262 18130 28314
rect 18130 28262 18142 28314
rect 18142 28262 18172 28314
rect 18196 28262 18206 28314
rect 18206 28262 18252 28314
rect 17956 28260 18012 28262
rect 18036 28260 18092 28262
rect 18116 28260 18172 28262
rect 18196 28260 18252 28262
rect 17956 27226 18012 27228
rect 18036 27226 18092 27228
rect 18116 27226 18172 27228
rect 18196 27226 18252 27228
rect 17956 27174 18002 27226
rect 18002 27174 18012 27226
rect 18036 27174 18066 27226
rect 18066 27174 18078 27226
rect 18078 27174 18092 27226
rect 18116 27174 18130 27226
rect 18130 27174 18142 27226
rect 18142 27174 18172 27226
rect 18196 27174 18206 27226
rect 18206 27174 18252 27226
rect 17956 27172 18012 27174
rect 18036 27172 18092 27174
rect 18116 27172 18172 27174
rect 18196 27172 18252 27174
rect 17956 26138 18012 26140
rect 18036 26138 18092 26140
rect 18116 26138 18172 26140
rect 18196 26138 18252 26140
rect 17956 26086 18002 26138
rect 18002 26086 18012 26138
rect 18036 26086 18066 26138
rect 18066 26086 18078 26138
rect 18078 26086 18092 26138
rect 18116 26086 18130 26138
rect 18130 26086 18142 26138
rect 18142 26086 18172 26138
rect 18196 26086 18206 26138
rect 18206 26086 18252 26138
rect 17956 26084 18012 26086
rect 18036 26084 18092 26086
rect 18116 26084 18172 26086
rect 18196 26084 18252 26086
rect 17956 25050 18012 25052
rect 18036 25050 18092 25052
rect 18116 25050 18172 25052
rect 18196 25050 18252 25052
rect 17956 24998 18002 25050
rect 18002 24998 18012 25050
rect 18036 24998 18066 25050
rect 18066 24998 18078 25050
rect 18078 24998 18092 25050
rect 18116 24998 18130 25050
rect 18130 24998 18142 25050
rect 18142 24998 18172 25050
rect 18196 24998 18206 25050
rect 18206 24998 18252 25050
rect 17956 24996 18012 24998
rect 18036 24996 18092 24998
rect 18116 24996 18172 24998
rect 18196 24996 18252 24998
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17130 16632 17186 16688
rect 16302 2372 16358 2408
rect 16302 2352 16304 2372
rect 16304 2352 16356 2372
rect 16356 2352 16358 2372
rect 16854 8880 16910 8936
rect 16854 8472 16910 8528
rect 17406 17332 17462 17368
rect 17406 17312 17408 17332
rect 17408 17312 17460 17332
rect 17460 17312 17462 17332
rect 17314 15272 17370 15328
rect 17406 13524 17462 13560
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17406 13504 17408 13524
rect 17408 13504 17460 13524
rect 17460 13504 17462 13524
rect 18878 23432 18934 23488
rect 19154 22344 19210 22400
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17774 10512 17830 10568
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17774 9560 17830 9616
rect 17774 8492 17830 8528
rect 17774 8472 17776 8492
rect 17776 8472 17828 8492
rect 17828 8472 17830 8492
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18234 7792 18290 7848
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17590 7112 17646 7168
rect 17682 6976 17738 7032
rect 17314 3984 17370 4040
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18694 9560 18750 9616
rect 18878 10240 18934 10296
rect 19890 24928 19946 24984
rect 19706 22344 19762 22400
rect 19338 11756 19394 11792
rect 19338 11736 19340 11756
rect 19340 11736 19392 11756
rect 19392 11736 19394 11756
rect 19246 10784 19302 10840
rect 20442 22380 20444 22400
rect 20444 22380 20496 22400
rect 20496 22380 20498 22400
rect 20442 22344 20498 22380
rect 22956 53882 23012 53884
rect 23036 53882 23092 53884
rect 23116 53882 23172 53884
rect 23196 53882 23252 53884
rect 22956 53830 23002 53882
rect 23002 53830 23012 53882
rect 23036 53830 23066 53882
rect 23066 53830 23078 53882
rect 23078 53830 23092 53882
rect 23116 53830 23130 53882
rect 23130 53830 23142 53882
rect 23142 53830 23172 53882
rect 23196 53830 23206 53882
rect 23206 53830 23252 53882
rect 22956 53828 23012 53830
rect 23036 53828 23092 53830
rect 23116 53828 23172 53830
rect 23196 53828 23252 53830
rect 24766 55392 24822 55448
rect 24582 54576 24638 54632
rect 22956 52794 23012 52796
rect 23036 52794 23092 52796
rect 23116 52794 23172 52796
rect 23196 52794 23252 52796
rect 22956 52742 23002 52794
rect 23002 52742 23012 52794
rect 23036 52742 23066 52794
rect 23066 52742 23078 52794
rect 23078 52742 23092 52794
rect 23116 52742 23130 52794
rect 23130 52742 23142 52794
rect 23142 52742 23172 52794
rect 23196 52742 23206 52794
rect 23206 52742 23252 52794
rect 22956 52740 23012 52742
rect 23036 52740 23092 52742
rect 23116 52740 23172 52742
rect 23196 52740 23252 52742
rect 22956 51706 23012 51708
rect 23036 51706 23092 51708
rect 23116 51706 23172 51708
rect 23196 51706 23252 51708
rect 22956 51654 23002 51706
rect 23002 51654 23012 51706
rect 23036 51654 23066 51706
rect 23066 51654 23078 51706
rect 23078 51654 23092 51706
rect 23116 51654 23130 51706
rect 23130 51654 23142 51706
rect 23142 51654 23172 51706
rect 23196 51654 23206 51706
rect 23206 51654 23252 51706
rect 22956 51652 23012 51654
rect 23036 51652 23092 51654
rect 23116 51652 23172 51654
rect 23196 51652 23252 51654
rect 22956 50618 23012 50620
rect 23036 50618 23092 50620
rect 23116 50618 23172 50620
rect 23196 50618 23252 50620
rect 22956 50566 23002 50618
rect 23002 50566 23012 50618
rect 23036 50566 23066 50618
rect 23066 50566 23078 50618
rect 23078 50566 23092 50618
rect 23116 50566 23130 50618
rect 23130 50566 23142 50618
rect 23142 50566 23172 50618
rect 23196 50566 23206 50618
rect 23206 50566 23252 50618
rect 22956 50564 23012 50566
rect 23036 50564 23092 50566
rect 23116 50564 23172 50566
rect 23196 50564 23252 50566
rect 22956 49530 23012 49532
rect 23036 49530 23092 49532
rect 23116 49530 23172 49532
rect 23196 49530 23252 49532
rect 22956 49478 23002 49530
rect 23002 49478 23012 49530
rect 23036 49478 23066 49530
rect 23066 49478 23078 49530
rect 23078 49478 23092 49530
rect 23116 49478 23130 49530
rect 23130 49478 23142 49530
rect 23142 49478 23172 49530
rect 23196 49478 23206 49530
rect 23206 49478 23252 49530
rect 22956 49476 23012 49478
rect 23036 49476 23092 49478
rect 23116 49476 23172 49478
rect 23196 49476 23252 49478
rect 22956 48442 23012 48444
rect 23036 48442 23092 48444
rect 23116 48442 23172 48444
rect 23196 48442 23252 48444
rect 22956 48390 23002 48442
rect 23002 48390 23012 48442
rect 23036 48390 23066 48442
rect 23066 48390 23078 48442
rect 23078 48390 23092 48442
rect 23116 48390 23130 48442
rect 23130 48390 23142 48442
rect 23142 48390 23172 48442
rect 23196 48390 23206 48442
rect 23206 48390 23252 48442
rect 22956 48388 23012 48390
rect 23036 48388 23092 48390
rect 23116 48388 23172 48390
rect 23196 48388 23252 48390
rect 22956 47354 23012 47356
rect 23036 47354 23092 47356
rect 23116 47354 23172 47356
rect 23196 47354 23252 47356
rect 22956 47302 23002 47354
rect 23002 47302 23012 47354
rect 23036 47302 23066 47354
rect 23066 47302 23078 47354
rect 23078 47302 23092 47354
rect 23116 47302 23130 47354
rect 23130 47302 23142 47354
rect 23142 47302 23172 47354
rect 23196 47302 23206 47354
rect 23206 47302 23252 47354
rect 22956 47300 23012 47302
rect 23036 47300 23092 47302
rect 23116 47300 23172 47302
rect 23196 47300 23252 47302
rect 22956 46266 23012 46268
rect 23036 46266 23092 46268
rect 23116 46266 23172 46268
rect 23196 46266 23252 46268
rect 22956 46214 23002 46266
rect 23002 46214 23012 46266
rect 23036 46214 23066 46266
rect 23066 46214 23078 46266
rect 23078 46214 23092 46266
rect 23116 46214 23130 46266
rect 23130 46214 23142 46266
rect 23142 46214 23172 46266
rect 23196 46214 23206 46266
rect 23206 46214 23252 46266
rect 22956 46212 23012 46214
rect 23036 46212 23092 46214
rect 23116 46212 23172 46214
rect 23196 46212 23252 46214
rect 22956 45178 23012 45180
rect 23036 45178 23092 45180
rect 23116 45178 23172 45180
rect 23196 45178 23252 45180
rect 22956 45126 23002 45178
rect 23002 45126 23012 45178
rect 23036 45126 23066 45178
rect 23066 45126 23078 45178
rect 23078 45126 23092 45178
rect 23116 45126 23130 45178
rect 23130 45126 23142 45178
rect 23142 45126 23172 45178
rect 23196 45126 23206 45178
rect 23206 45126 23252 45178
rect 22956 45124 23012 45126
rect 23036 45124 23092 45126
rect 23116 45124 23172 45126
rect 23196 45124 23252 45126
rect 22956 44090 23012 44092
rect 23036 44090 23092 44092
rect 23116 44090 23172 44092
rect 23196 44090 23252 44092
rect 22956 44038 23002 44090
rect 23002 44038 23012 44090
rect 23036 44038 23066 44090
rect 23066 44038 23078 44090
rect 23078 44038 23092 44090
rect 23116 44038 23130 44090
rect 23130 44038 23142 44090
rect 23142 44038 23172 44090
rect 23196 44038 23206 44090
rect 23206 44038 23252 44090
rect 22956 44036 23012 44038
rect 23036 44036 23092 44038
rect 23116 44036 23172 44038
rect 23196 44036 23252 44038
rect 22956 43002 23012 43004
rect 23036 43002 23092 43004
rect 23116 43002 23172 43004
rect 23196 43002 23252 43004
rect 22956 42950 23002 43002
rect 23002 42950 23012 43002
rect 23036 42950 23066 43002
rect 23066 42950 23078 43002
rect 23078 42950 23092 43002
rect 23116 42950 23130 43002
rect 23130 42950 23142 43002
rect 23142 42950 23172 43002
rect 23196 42950 23206 43002
rect 23206 42950 23252 43002
rect 22956 42948 23012 42950
rect 23036 42948 23092 42950
rect 23116 42948 23172 42950
rect 23196 42948 23252 42950
rect 22956 41914 23012 41916
rect 23036 41914 23092 41916
rect 23116 41914 23172 41916
rect 23196 41914 23252 41916
rect 22956 41862 23002 41914
rect 23002 41862 23012 41914
rect 23036 41862 23066 41914
rect 23066 41862 23078 41914
rect 23078 41862 23092 41914
rect 23116 41862 23130 41914
rect 23130 41862 23142 41914
rect 23142 41862 23172 41914
rect 23196 41862 23206 41914
rect 23206 41862 23252 41914
rect 22956 41860 23012 41862
rect 23036 41860 23092 41862
rect 23116 41860 23172 41862
rect 23196 41860 23252 41862
rect 22956 40826 23012 40828
rect 23036 40826 23092 40828
rect 23116 40826 23172 40828
rect 23196 40826 23252 40828
rect 22956 40774 23002 40826
rect 23002 40774 23012 40826
rect 23036 40774 23066 40826
rect 23066 40774 23078 40826
rect 23078 40774 23092 40826
rect 23116 40774 23130 40826
rect 23130 40774 23142 40826
rect 23142 40774 23172 40826
rect 23196 40774 23206 40826
rect 23206 40774 23252 40826
rect 22956 40772 23012 40774
rect 23036 40772 23092 40774
rect 23116 40772 23172 40774
rect 23196 40772 23252 40774
rect 22956 39738 23012 39740
rect 23036 39738 23092 39740
rect 23116 39738 23172 39740
rect 23196 39738 23252 39740
rect 22956 39686 23002 39738
rect 23002 39686 23012 39738
rect 23036 39686 23066 39738
rect 23066 39686 23078 39738
rect 23078 39686 23092 39738
rect 23116 39686 23130 39738
rect 23130 39686 23142 39738
rect 23142 39686 23172 39738
rect 23196 39686 23206 39738
rect 23206 39686 23252 39738
rect 22956 39684 23012 39686
rect 23036 39684 23092 39686
rect 23116 39684 23172 39686
rect 23196 39684 23252 39686
rect 22956 38650 23012 38652
rect 23036 38650 23092 38652
rect 23116 38650 23172 38652
rect 23196 38650 23252 38652
rect 22956 38598 23002 38650
rect 23002 38598 23012 38650
rect 23036 38598 23066 38650
rect 23066 38598 23078 38650
rect 23078 38598 23092 38650
rect 23116 38598 23130 38650
rect 23130 38598 23142 38650
rect 23142 38598 23172 38650
rect 23196 38598 23206 38650
rect 23206 38598 23252 38650
rect 22956 38596 23012 38598
rect 23036 38596 23092 38598
rect 23116 38596 23172 38598
rect 23196 38596 23252 38598
rect 22956 37562 23012 37564
rect 23036 37562 23092 37564
rect 23116 37562 23172 37564
rect 23196 37562 23252 37564
rect 22956 37510 23002 37562
rect 23002 37510 23012 37562
rect 23036 37510 23066 37562
rect 23066 37510 23078 37562
rect 23078 37510 23092 37562
rect 23116 37510 23130 37562
rect 23130 37510 23142 37562
rect 23142 37510 23172 37562
rect 23196 37510 23206 37562
rect 23206 37510 23252 37562
rect 22956 37508 23012 37510
rect 23036 37508 23092 37510
rect 23116 37508 23172 37510
rect 23196 37508 23252 37510
rect 22956 36474 23012 36476
rect 23036 36474 23092 36476
rect 23116 36474 23172 36476
rect 23196 36474 23252 36476
rect 22956 36422 23002 36474
rect 23002 36422 23012 36474
rect 23036 36422 23066 36474
rect 23066 36422 23078 36474
rect 23078 36422 23092 36474
rect 23116 36422 23130 36474
rect 23130 36422 23142 36474
rect 23142 36422 23172 36474
rect 23196 36422 23206 36474
rect 23206 36422 23252 36474
rect 22956 36420 23012 36422
rect 23036 36420 23092 36422
rect 23116 36420 23172 36422
rect 23196 36420 23252 36422
rect 22956 35386 23012 35388
rect 23036 35386 23092 35388
rect 23116 35386 23172 35388
rect 23196 35386 23252 35388
rect 22956 35334 23002 35386
rect 23002 35334 23012 35386
rect 23036 35334 23066 35386
rect 23066 35334 23078 35386
rect 23078 35334 23092 35386
rect 23116 35334 23130 35386
rect 23130 35334 23142 35386
rect 23142 35334 23172 35386
rect 23196 35334 23206 35386
rect 23206 35334 23252 35386
rect 22956 35332 23012 35334
rect 23036 35332 23092 35334
rect 23116 35332 23172 35334
rect 23196 35332 23252 35334
rect 22956 34298 23012 34300
rect 23036 34298 23092 34300
rect 23116 34298 23172 34300
rect 23196 34298 23252 34300
rect 22956 34246 23002 34298
rect 23002 34246 23012 34298
rect 23036 34246 23066 34298
rect 23066 34246 23078 34298
rect 23078 34246 23092 34298
rect 23116 34246 23130 34298
rect 23130 34246 23142 34298
rect 23142 34246 23172 34298
rect 23196 34246 23206 34298
rect 23206 34246 23252 34298
rect 22956 34244 23012 34246
rect 23036 34244 23092 34246
rect 23116 34244 23172 34246
rect 23196 34244 23252 34246
rect 22956 33210 23012 33212
rect 23036 33210 23092 33212
rect 23116 33210 23172 33212
rect 23196 33210 23252 33212
rect 22956 33158 23002 33210
rect 23002 33158 23012 33210
rect 23036 33158 23066 33210
rect 23066 33158 23078 33210
rect 23078 33158 23092 33210
rect 23116 33158 23130 33210
rect 23130 33158 23142 33210
rect 23142 33158 23172 33210
rect 23196 33158 23206 33210
rect 23206 33158 23252 33210
rect 22956 33156 23012 33158
rect 23036 33156 23092 33158
rect 23116 33156 23172 33158
rect 23196 33156 23252 33158
rect 19522 10648 19578 10704
rect 19522 10240 19578 10296
rect 19246 8880 19302 8936
rect 19246 7148 19248 7168
rect 19248 7148 19300 7168
rect 19300 7148 19302 7168
rect 19246 7112 19302 7148
rect 19246 6996 19302 7032
rect 19246 6976 19248 6996
rect 19248 6976 19300 6996
rect 19300 6976 19302 6996
rect 19982 12280 20038 12336
rect 20166 9968 20222 10024
rect 20626 10648 20682 10704
rect 20626 9424 20682 9480
rect 21270 10376 21326 10432
rect 22956 32122 23012 32124
rect 23036 32122 23092 32124
rect 23116 32122 23172 32124
rect 23196 32122 23252 32124
rect 22956 32070 23002 32122
rect 23002 32070 23012 32122
rect 23036 32070 23066 32122
rect 23066 32070 23078 32122
rect 23078 32070 23092 32122
rect 23116 32070 23130 32122
rect 23130 32070 23142 32122
rect 23142 32070 23172 32122
rect 23196 32070 23206 32122
rect 23206 32070 23252 32122
rect 22956 32068 23012 32070
rect 23036 32068 23092 32070
rect 23116 32068 23172 32070
rect 23196 32068 23252 32070
rect 25042 53760 25098 53816
rect 25042 52944 25098 53000
rect 24950 52128 25006 52184
rect 24950 51332 25006 51368
rect 24950 51312 24952 51332
rect 24952 51312 25004 51332
rect 25004 51312 25006 51332
rect 24950 50496 25006 50552
rect 25502 49680 25558 49736
rect 25134 48864 25190 48920
rect 25134 48084 25136 48104
rect 25136 48084 25188 48104
rect 25188 48084 25190 48104
rect 25134 48048 25190 48084
rect 24766 43968 24822 44024
rect 25134 42336 25190 42392
rect 25134 41556 25136 41576
rect 25136 41556 25188 41576
rect 25188 41556 25190 41576
rect 25134 41520 25190 41556
rect 25134 37440 25190 37496
rect 22956 31034 23012 31036
rect 23036 31034 23092 31036
rect 23116 31034 23172 31036
rect 23196 31034 23252 31036
rect 22956 30982 23002 31034
rect 23002 30982 23012 31034
rect 23036 30982 23066 31034
rect 23066 30982 23078 31034
rect 23078 30982 23092 31034
rect 23116 30982 23130 31034
rect 23130 30982 23142 31034
rect 23142 30982 23172 31034
rect 23196 30982 23206 31034
rect 23206 30982 23252 31034
rect 22956 30980 23012 30982
rect 23036 30980 23092 30982
rect 23116 30980 23172 30982
rect 23196 30980 23252 30982
rect 22956 29946 23012 29948
rect 23036 29946 23092 29948
rect 23116 29946 23172 29948
rect 23196 29946 23252 29948
rect 22956 29894 23002 29946
rect 23002 29894 23012 29946
rect 23036 29894 23066 29946
rect 23066 29894 23078 29946
rect 23078 29894 23092 29946
rect 23116 29894 23130 29946
rect 23130 29894 23142 29946
rect 23142 29894 23172 29946
rect 23196 29894 23206 29946
rect 23206 29894 23252 29946
rect 22956 29892 23012 29894
rect 23036 29892 23092 29894
rect 23116 29892 23172 29894
rect 23196 29892 23252 29894
rect 22956 28858 23012 28860
rect 23036 28858 23092 28860
rect 23116 28858 23172 28860
rect 23196 28858 23252 28860
rect 22956 28806 23002 28858
rect 23002 28806 23012 28858
rect 23036 28806 23066 28858
rect 23066 28806 23078 28858
rect 23078 28806 23092 28858
rect 23116 28806 23130 28858
rect 23130 28806 23142 28858
rect 23142 28806 23172 28858
rect 23196 28806 23206 28858
rect 23206 28806 23252 28858
rect 22956 28804 23012 28806
rect 23036 28804 23092 28806
rect 23116 28804 23172 28806
rect 23196 28804 23252 28806
rect 22956 27770 23012 27772
rect 23036 27770 23092 27772
rect 23116 27770 23172 27772
rect 23196 27770 23252 27772
rect 22956 27718 23002 27770
rect 23002 27718 23012 27770
rect 23036 27718 23066 27770
rect 23066 27718 23078 27770
rect 23078 27718 23092 27770
rect 23116 27718 23130 27770
rect 23130 27718 23142 27770
rect 23142 27718 23172 27770
rect 23196 27718 23206 27770
rect 23206 27718 23252 27770
rect 22956 27716 23012 27718
rect 23036 27716 23092 27718
rect 23116 27716 23172 27718
rect 23196 27716 23252 27718
rect 22956 26682 23012 26684
rect 23036 26682 23092 26684
rect 23116 26682 23172 26684
rect 23196 26682 23252 26684
rect 22956 26630 23002 26682
rect 23002 26630 23012 26682
rect 23036 26630 23066 26682
rect 23066 26630 23078 26682
rect 23078 26630 23092 26682
rect 23116 26630 23130 26682
rect 23130 26630 23142 26682
rect 23142 26630 23172 26682
rect 23196 26630 23206 26682
rect 23206 26630 23252 26682
rect 22956 26628 23012 26630
rect 23036 26628 23092 26630
rect 23116 26628 23172 26630
rect 23196 26628 23252 26630
rect 22956 25594 23012 25596
rect 23036 25594 23092 25596
rect 23116 25594 23172 25596
rect 23196 25594 23252 25596
rect 22956 25542 23002 25594
rect 23002 25542 23012 25594
rect 23036 25542 23066 25594
rect 23066 25542 23078 25594
rect 23078 25542 23092 25594
rect 23116 25542 23130 25594
rect 23130 25542 23142 25594
rect 23142 25542 23172 25594
rect 23196 25542 23206 25594
rect 23206 25542 23252 25594
rect 22956 25540 23012 25542
rect 23036 25540 23092 25542
rect 23116 25540 23172 25542
rect 23196 25540 23252 25542
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 24030 27648 24086 27704
rect 23846 24384 23902 24440
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 23386 21936 23442 21992
rect 21914 16496 21970 16552
rect 22098 9424 22154 9480
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 23110 19760 23166 19816
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 23846 19488 23902 19544
rect 22742 16496 22798 16552
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22282 10376 22338 10432
rect 22558 10240 22614 10296
rect 22374 9968 22430 10024
rect 22006 5072 22062 5128
rect 22374 3168 22430 3224
rect 22098 2352 22154 2408
rect 22282 1536 22338 1592
rect 23294 15408 23350 15464
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22650 8336 22706 8392
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 23846 17040 23902 17096
rect 23846 13776 23902 13832
rect 23662 10648 23718 10704
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22834 5616 22890 5672
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22742 3984 22798 4040
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 23846 10512 23902 10568
rect 24950 29280 25006 29336
rect 24490 28464 24546 28520
rect 24858 26016 24914 26072
rect 24766 23568 24822 23624
rect 24858 22752 24914 22808
rect 24858 21120 24914 21176
rect 25318 47232 25374 47288
rect 25318 46416 25374 46472
rect 25318 45600 25374 45656
rect 25318 44820 25320 44840
rect 25320 44820 25372 44840
rect 25372 44820 25374 44840
rect 25318 44784 25374 44820
rect 25318 40704 25374 40760
rect 25318 39072 25374 39128
rect 25318 38292 25320 38312
rect 25320 38292 25372 38312
rect 25372 38292 25374 38312
rect 25318 38256 25374 38292
rect 25318 35808 25374 35864
rect 25502 43152 25558 43208
rect 25502 39888 25558 39944
rect 25502 36624 25558 36680
rect 25318 35028 25320 35048
rect 25320 35028 25372 35048
rect 25372 35028 25374 35048
rect 25318 34992 25374 35028
rect 25318 34176 25374 34232
rect 25318 33360 25374 33416
rect 25318 31764 25320 31784
rect 25320 31764 25372 31784
rect 25372 31764 25374 31784
rect 25318 31728 25374 31764
rect 25318 30096 25374 30152
rect 25502 32544 25558 32600
rect 25502 30932 25558 30968
rect 25502 30912 25504 30932
rect 25504 30912 25556 30932
rect 25556 30912 25558 30932
rect 25318 26832 25374 26888
rect 25134 25200 25190 25256
rect 24674 20304 24730 20360
rect 24858 18672 24914 18728
rect 24950 17856 25006 17912
rect 23754 4528 23810 4584
rect 24306 10784 24362 10840
rect 24766 16224 24822 16280
rect 24858 14592 24914 14648
rect 24766 12960 24822 13016
rect 24950 12164 25006 12200
rect 24950 12144 24952 12164
rect 24952 12144 25004 12164
rect 25004 12144 25006 12164
rect 24858 11328 24914 11384
rect 24766 9696 24822 9752
rect 24490 9424 24546 9480
rect 24398 3984 24454 4040
rect 23938 3440 23994 3496
rect 24950 8900 25006 8936
rect 24950 8880 24952 8900
rect 24952 8880 25004 8900
rect 25004 8880 25006 8900
rect 24858 7284 24860 7304
rect 24860 7284 24912 7304
rect 24912 7284 24914 7304
rect 24858 7248 24914 7284
rect 24950 6432 25006 6488
rect 25134 8064 25190 8120
rect 24950 3612 24952 3632
rect 24952 3612 25004 3632
rect 25004 3612 25006 3632
rect 24950 3576 25006 3612
rect 25318 720 25374 776
<< metal3 >>
rect 26200 56266 27000 56296
rect 23430 56206 27000 56266
rect 23430 56133 23490 56206
rect 26200 56176 27000 56206
rect 23381 56128 23490 56133
rect 23381 56072 23386 56128
rect 23442 56072 23490 56128
rect 23381 56070 23490 56072
rect 23381 56067 23447 56070
rect 24761 55450 24827 55453
rect 26200 55450 27000 55480
rect 24761 55448 27000 55450
rect 24761 55392 24766 55448
rect 24822 55392 27000 55448
rect 24761 55390 27000 55392
rect 24761 55387 24827 55390
rect 26200 55360 27000 55390
rect 24577 54634 24643 54637
rect 26200 54634 27000 54664
rect 24577 54632 27000 54634
rect 24577 54576 24582 54632
rect 24638 54576 27000 54632
rect 24577 54574 27000 54576
rect 24577 54571 24643 54574
rect 26200 54544 27000 54574
rect 7946 54432 8262 54433
rect 7946 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8262 54432
rect 7946 54367 8262 54368
rect 17946 54432 18262 54433
rect 17946 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18262 54432
rect 17946 54367 18262 54368
rect 2946 53888 3262 53889
rect 2946 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3262 53888
rect 2946 53823 3262 53824
rect 12946 53888 13262 53889
rect 12946 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13262 53888
rect 12946 53823 13262 53824
rect 22946 53888 23262 53889
rect 22946 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23262 53888
rect 22946 53823 23262 53824
rect 25037 53818 25103 53821
rect 26200 53818 27000 53848
rect 25037 53816 27000 53818
rect 25037 53760 25042 53816
rect 25098 53760 27000 53816
rect 25037 53758 27000 53760
rect 25037 53755 25103 53758
rect 26200 53728 27000 53758
rect 7946 53344 8262 53345
rect 7946 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8262 53344
rect 7946 53279 8262 53280
rect 17946 53344 18262 53345
rect 17946 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18262 53344
rect 17946 53279 18262 53280
rect 25037 53002 25103 53005
rect 26200 53002 27000 53032
rect 25037 53000 27000 53002
rect 25037 52944 25042 53000
rect 25098 52944 27000 53000
rect 25037 52942 27000 52944
rect 25037 52939 25103 52942
rect 26200 52912 27000 52942
rect 2946 52800 3262 52801
rect 2946 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3262 52800
rect 2946 52735 3262 52736
rect 12946 52800 13262 52801
rect 12946 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13262 52800
rect 12946 52735 13262 52736
rect 22946 52800 23262 52801
rect 22946 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23262 52800
rect 22946 52735 23262 52736
rect 7946 52256 8262 52257
rect 7946 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8262 52256
rect 7946 52191 8262 52192
rect 17946 52256 18262 52257
rect 17946 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18262 52256
rect 17946 52191 18262 52192
rect 24945 52186 25011 52189
rect 26200 52186 27000 52216
rect 24945 52184 27000 52186
rect 24945 52128 24950 52184
rect 25006 52128 27000 52184
rect 24945 52126 27000 52128
rect 24945 52123 25011 52126
rect 26200 52096 27000 52126
rect 2946 51712 3262 51713
rect 2946 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3262 51712
rect 2946 51647 3262 51648
rect 12946 51712 13262 51713
rect 12946 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13262 51712
rect 12946 51647 13262 51648
rect 22946 51712 23262 51713
rect 22946 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23262 51712
rect 22946 51647 23262 51648
rect 24945 51370 25011 51373
rect 26200 51370 27000 51400
rect 24945 51368 27000 51370
rect 24945 51312 24950 51368
rect 25006 51312 27000 51368
rect 24945 51310 27000 51312
rect 24945 51307 25011 51310
rect 26200 51280 27000 51310
rect 7946 51168 8262 51169
rect 7946 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8262 51168
rect 7946 51103 8262 51104
rect 17946 51168 18262 51169
rect 17946 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18262 51168
rect 17946 51103 18262 51104
rect 2946 50624 3262 50625
rect 2946 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3262 50624
rect 2946 50559 3262 50560
rect 12946 50624 13262 50625
rect 12946 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13262 50624
rect 12946 50559 13262 50560
rect 22946 50624 23262 50625
rect 22946 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23262 50624
rect 22946 50559 23262 50560
rect 24945 50554 25011 50557
rect 26200 50554 27000 50584
rect 24945 50552 27000 50554
rect 24945 50496 24950 50552
rect 25006 50496 27000 50552
rect 24945 50494 27000 50496
rect 24945 50491 25011 50494
rect 26200 50464 27000 50494
rect 7946 50080 8262 50081
rect 7946 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8262 50080
rect 7946 50015 8262 50016
rect 17946 50080 18262 50081
rect 17946 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18262 50080
rect 17946 50015 18262 50016
rect 25497 49738 25563 49741
rect 26200 49738 27000 49768
rect 25497 49736 27000 49738
rect 25497 49680 25502 49736
rect 25558 49680 27000 49736
rect 25497 49678 27000 49680
rect 25497 49675 25563 49678
rect 26200 49648 27000 49678
rect 2946 49536 3262 49537
rect 2946 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3262 49536
rect 2946 49471 3262 49472
rect 12946 49536 13262 49537
rect 12946 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13262 49536
rect 12946 49471 13262 49472
rect 22946 49536 23262 49537
rect 22946 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23262 49536
rect 22946 49471 23262 49472
rect 7946 48992 8262 48993
rect 7946 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8262 48992
rect 7946 48927 8262 48928
rect 17946 48992 18262 48993
rect 17946 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18262 48992
rect 17946 48927 18262 48928
rect 25129 48922 25195 48925
rect 26200 48922 27000 48952
rect 25129 48920 27000 48922
rect 25129 48864 25134 48920
rect 25190 48864 27000 48920
rect 25129 48862 27000 48864
rect 25129 48859 25195 48862
rect 26200 48832 27000 48862
rect 2946 48448 3262 48449
rect 2946 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3262 48448
rect 2946 48383 3262 48384
rect 12946 48448 13262 48449
rect 12946 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13262 48448
rect 12946 48383 13262 48384
rect 22946 48448 23262 48449
rect 22946 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23262 48448
rect 22946 48383 23262 48384
rect 25129 48106 25195 48109
rect 26200 48106 27000 48136
rect 25129 48104 27000 48106
rect 25129 48048 25134 48104
rect 25190 48048 27000 48104
rect 25129 48046 27000 48048
rect 25129 48043 25195 48046
rect 26200 48016 27000 48046
rect 7946 47904 8262 47905
rect 7946 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8262 47904
rect 7946 47839 8262 47840
rect 17946 47904 18262 47905
rect 17946 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18262 47904
rect 17946 47839 18262 47840
rect 2946 47360 3262 47361
rect 2946 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3262 47360
rect 2946 47295 3262 47296
rect 12946 47360 13262 47361
rect 12946 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13262 47360
rect 12946 47295 13262 47296
rect 22946 47360 23262 47361
rect 22946 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23262 47360
rect 22946 47295 23262 47296
rect 25313 47290 25379 47293
rect 26200 47290 27000 47320
rect 25313 47288 27000 47290
rect 25313 47232 25318 47288
rect 25374 47232 27000 47288
rect 25313 47230 27000 47232
rect 25313 47227 25379 47230
rect 26200 47200 27000 47230
rect 7946 46816 8262 46817
rect 7946 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8262 46816
rect 7946 46751 8262 46752
rect 17946 46816 18262 46817
rect 17946 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18262 46816
rect 17946 46751 18262 46752
rect 25313 46474 25379 46477
rect 26200 46474 27000 46504
rect 25313 46472 27000 46474
rect 25313 46416 25318 46472
rect 25374 46416 27000 46472
rect 25313 46414 27000 46416
rect 25313 46411 25379 46414
rect 26200 46384 27000 46414
rect 2946 46272 3262 46273
rect 2946 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3262 46272
rect 2946 46207 3262 46208
rect 12946 46272 13262 46273
rect 12946 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13262 46272
rect 12946 46207 13262 46208
rect 22946 46272 23262 46273
rect 22946 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23262 46272
rect 22946 46207 23262 46208
rect 7946 45728 8262 45729
rect 7946 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8262 45728
rect 7946 45663 8262 45664
rect 17946 45728 18262 45729
rect 17946 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18262 45728
rect 17946 45663 18262 45664
rect 25313 45658 25379 45661
rect 26200 45658 27000 45688
rect 25313 45656 27000 45658
rect 25313 45600 25318 45656
rect 25374 45600 27000 45656
rect 25313 45598 27000 45600
rect 25313 45595 25379 45598
rect 26200 45568 27000 45598
rect 2946 45184 3262 45185
rect 2946 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3262 45184
rect 2946 45119 3262 45120
rect 12946 45184 13262 45185
rect 12946 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13262 45184
rect 12946 45119 13262 45120
rect 22946 45184 23262 45185
rect 22946 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23262 45184
rect 22946 45119 23262 45120
rect 25313 44842 25379 44845
rect 26200 44842 27000 44872
rect 25313 44840 27000 44842
rect 25313 44784 25318 44840
rect 25374 44784 27000 44840
rect 25313 44782 27000 44784
rect 25313 44779 25379 44782
rect 26200 44752 27000 44782
rect 7946 44640 8262 44641
rect 7946 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8262 44640
rect 7946 44575 8262 44576
rect 17946 44640 18262 44641
rect 17946 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18262 44640
rect 17946 44575 18262 44576
rect 2946 44096 3262 44097
rect 2946 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3262 44096
rect 2946 44031 3262 44032
rect 12946 44096 13262 44097
rect 12946 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13262 44096
rect 12946 44031 13262 44032
rect 22946 44096 23262 44097
rect 22946 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23262 44096
rect 22946 44031 23262 44032
rect 24761 44026 24827 44029
rect 26200 44026 27000 44056
rect 24761 44024 27000 44026
rect 24761 43968 24766 44024
rect 24822 43968 27000 44024
rect 24761 43966 27000 43968
rect 24761 43963 24827 43966
rect 26200 43936 27000 43966
rect 7946 43552 8262 43553
rect 7946 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8262 43552
rect 7946 43487 8262 43488
rect 17946 43552 18262 43553
rect 17946 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18262 43552
rect 17946 43487 18262 43488
rect 25497 43210 25563 43213
rect 26200 43210 27000 43240
rect 25497 43208 27000 43210
rect 25497 43152 25502 43208
rect 25558 43152 27000 43208
rect 25497 43150 27000 43152
rect 25497 43147 25563 43150
rect 26200 43120 27000 43150
rect 2946 43008 3262 43009
rect 2946 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3262 43008
rect 2946 42943 3262 42944
rect 12946 43008 13262 43009
rect 12946 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13262 43008
rect 12946 42943 13262 42944
rect 22946 43008 23262 43009
rect 22946 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23262 43008
rect 22946 42943 23262 42944
rect 7946 42464 8262 42465
rect 7946 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8262 42464
rect 7946 42399 8262 42400
rect 17946 42464 18262 42465
rect 17946 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18262 42464
rect 17946 42399 18262 42400
rect 25129 42394 25195 42397
rect 26200 42394 27000 42424
rect 25129 42392 27000 42394
rect 25129 42336 25134 42392
rect 25190 42336 27000 42392
rect 25129 42334 27000 42336
rect 25129 42331 25195 42334
rect 26200 42304 27000 42334
rect 2946 41920 3262 41921
rect 2946 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3262 41920
rect 2946 41855 3262 41856
rect 12946 41920 13262 41921
rect 12946 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13262 41920
rect 12946 41855 13262 41856
rect 22946 41920 23262 41921
rect 22946 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23262 41920
rect 22946 41855 23262 41856
rect 25129 41578 25195 41581
rect 26200 41578 27000 41608
rect 25129 41576 27000 41578
rect 25129 41520 25134 41576
rect 25190 41520 27000 41576
rect 25129 41518 27000 41520
rect 25129 41515 25195 41518
rect 26200 41488 27000 41518
rect 7946 41376 8262 41377
rect 7946 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8262 41376
rect 7946 41311 8262 41312
rect 17946 41376 18262 41377
rect 17946 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18262 41376
rect 17946 41311 18262 41312
rect 2946 40832 3262 40833
rect 2946 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3262 40832
rect 2946 40767 3262 40768
rect 12946 40832 13262 40833
rect 12946 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13262 40832
rect 12946 40767 13262 40768
rect 22946 40832 23262 40833
rect 22946 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23262 40832
rect 22946 40767 23262 40768
rect 25313 40762 25379 40765
rect 26200 40762 27000 40792
rect 25313 40760 27000 40762
rect 25313 40704 25318 40760
rect 25374 40704 27000 40760
rect 25313 40702 27000 40704
rect 25313 40699 25379 40702
rect 26200 40672 27000 40702
rect 7946 40288 8262 40289
rect 7946 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8262 40288
rect 7946 40223 8262 40224
rect 17946 40288 18262 40289
rect 17946 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18262 40288
rect 17946 40223 18262 40224
rect 25497 39946 25563 39949
rect 26200 39946 27000 39976
rect 25497 39944 27000 39946
rect 25497 39888 25502 39944
rect 25558 39888 27000 39944
rect 25497 39886 27000 39888
rect 25497 39883 25563 39886
rect 26200 39856 27000 39886
rect 2946 39744 3262 39745
rect 2946 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3262 39744
rect 2946 39679 3262 39680
rect 12946 39744 13262 39745
rect 12946 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13262 39744
rect 12946 39679 13262 39680
rect 22946 39744 23262 39745
rect 22946 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23262 39744
rect 22946 39679 23262 39680
rect 7946 39200 8262 39201
rect 7946 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8262 39200
rect 7946 39135 8262 39136
rect 17946 39200 18262 39201
rect 17946 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18262 39200
rect 17946 39135 18262 39136
rect 25313 39130 25379 39133
rect 26200 39130 27000 39160
rect 25313 39128 27000 39130
rect 25313 39072 25318 39128
rect 25374 39072 27000 39128
rect 25313 39070 27000 39072
rect 25313 39067 25379 39070
rect 26200 39040 27000 39070
rect 2946 38656 3262 38657
rect 2946 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3262 38656
rect 2946 38591 3262 38592
rect 12946 38656 13262 38657
rect 12946 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13262 38656
rect 12946 38591 13262 38592
rect 22946 38656 23262 38657
rect 22946 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23262 38656
rect 22946 38591 23262 38592
rect 25313 38314 25379 38317
rect 26200 38314 27000 38344
rect 25313 38312 27000 38314
rect 25313 38256 25318 38312
rect 25374 38256 27000 38312
rect 25313 38254 27000 38256
rect 25313 38251 25379 38254
rect 26200 38224 27000 38254
rect 7946 38112 8262 38113
rect 7946 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8262 38112
rect 7946 38047 8262 38048
rect 17946 38112 18262 38113
rect 17946 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18262 38112
rect 17946 38047 18262 38048
rect 2946 37568 3262 37569
rect 2946 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3262 37568
rect 2946 37503 3262 37504
rect 12946 37568 13262 37569
rect 12946 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13262 37568
rect 12946 37503 13262 37504
rect 22946 37568 23262 37569
rect 22946 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23262 37568
rect 22946 37503 23262 37504
rect 25129 37498 25195 37501
rect 26200 37498 27000 37528
rect 25129 37496 27000 37498
rect 25129 37440 25134 37496
rect 25190 37440 27000 37496
rect 25129 37438 27000 37440
rect 25129 37435 25195 37438
rect 26200 37408 27000 37438
rect 7946 37024 8262 37025
rect 7946 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8262 37024
rect 7946 36959 8262 36960
rect 17946 37024 18262 37025
rect 17946 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18262 37024
rect 17946 36959 18262 36960
rect 25497 36682 25563 36685
rect 26200 36682 27000 36712
rect 25497 36680 27000 36682
rect 25497 36624 25502 36680
rect 25558 36624 27000 36680
rect 25497 36622 27000 36624
rect 25497 36619 25563 36622
rect 26200 36592 27000 36622
rect 2946 36480 3262 36481
rect 2946 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3262 36480
rect 2946 36415 3262 36416
rect 12946 36480 13262 36481
rect 12946 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13262 36480
rect 12946 36415 13262 36416
rect 22946 36480 23262 36481
rect 22946 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23262 36480
rect 22946 36415 23262 36416
rect 7946 35936 8262 35937
rect 7946 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8262 35936
rect 7946 35871 8262 35872
rect 17946 35936 18262 35937
rect 17946 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18262 35936
rect 17946 35871 18262 35872
rect 25313 35866 25379 35869
rect 26200 35866 27000 35896
rect 25313 35864 27000 35866
rect 25313 35808 25318 35864
rect 25374 35808 27000 35864
rect 25313 35806 27000 35808
rect 25313 35803 25379 35806
rect 26200 35776 27000 35806
rect 2946 35392 3262 35393
rect 2946 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3262 35392
rect 2946 35327 3262 35328
rect 12946 35392 13262 35393
rect 12946 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13262 35392
rect 12946 35327 13262 35328
rect 22946 35392 23262 35393
rect 22946 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23262 35392
rect 22946 35327 23262 35328
rect 25313 35050 25379 35053
rect 26200 35050 27000 35080
rect 25313 35048 27000 35050
rect 25313 34992 25318 35048
rect 25374 34992 27000 35048
rect 25313 34990 27000 34992
rect 25313 34987 25379 34990
rect 26200 34960 27000 34990
rect 7946 34848 8262 34849
rect 7946 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8262 34848
rect 7946 34783 8262 34784
rect 17946 34848 18262 34849
rect 17946 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18262 34848
rect 17946 34783 18262 34784
rect 2946 34304 3262 34305
rect 2946 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3262 34304
rect 2946 34239 3262 34240
rect 12946 34304 13262 34305
rect 12946 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13262 34304
rect 12946 34239 13262 34240
rect 22946 34304 23262 34305
rect 22946 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23262 34304
rect 22946 34239 23262 34240
rect 25313 34234 25379 34237
rect 26200 34234 27000 34264
rect 25313 34232 27000 34234
rect 25313 34176 25318 34232
rect 25374 34176 27000 34232
rect 25313 34174 27000 34176
rect 25313 34171 25379 34174
rect 26200 34144 27000 34174
rect 7946 33760 8262 33761
rect 7946 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8262 33760
rect 7946 33695 8262 33696
rect 17946 33760 18262 33761
rect 17946 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18262 33760
rect 17946 33695 18262 33696
rect 25313 33418 25379 33421
rect 26200 33418 27000 33448
rect 25313 33416 27000 33418
rect 25313 33360 25318 33416
rect 25374 33360 27000 33416
rect 25313 33358 27000 33360
rect 25313 33355 25379 33358
rect 26200 33328 27000 33358
rect 2946 33216 3262 33217
rect 2946 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3262 33216
rect 2946 33151 3262 33152
rect 12946 33216 13262 33217
rect 12946 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13262 33216
rect 12946 33151 13262 33152
rect 22946 33216 23262 33217
rect 22946 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23262 33216
rect 22946 33151 23262 33152
rect 7946 32672 8262 32673
rect 7946 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8262 32672
rect 7946 32607 8262 32608
rect 17946 32672 18262 32673
rect 17946 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18262 32672
rect 17946 32607 18262 32608
rect 25497 32602 25563 32605
rect 26200 32602 27000 32632
rect 25497 32600 27000 32602
rect 25497 32544 25502 32600
rect 25558 32544 27000 32600
rect 25497 32542 27000 32544
rect 25497 32539 25563 32542
rect 26200 32512 27000 32542
rect 2946 32128 3262 32129
rect 2946 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3262 32128
rect 2946 32063 3262 32064
rect 12946 32128 13262 32129
rect 12946 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13262 32128
rect 12946 32063 13262 32064
rect 22946 32128 23262 32129
rect 22946 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23262 32128
rect 22946 32063 23262 32064
rect 25313 31786 25379 31789
rect 26200 31786 27000 31816
rect 25313 31784 27000 31786
rect 25313 31728 25318 31784
rect 25374 31728 27000 31784
rect 25313 31726 27000 31728
rect 25313 31723 25379 31726
rect 26200 31696 27000 31726
rect 7946 31584 8262 31585
rect 7946 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8262 31584
rect 7946 31519 8262 31520
rect 17946 31584 18262 31585
rect 17946 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18262 31584
rect 17946 31519 18262 31520
rect 2946 31040 3262 31041
rect 2946 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3262 31040
rect 2946 30975 3262 30976
rect 12946 31040 13262 31041
rect 12946 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13262 31040
rect 12946 30975 13262 30976
rect 22946 31040 23262 31041
rect 22946 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23262 31040
rect 22946 30975 23262 30976
rect 25497 30970 25563 30973
rect 26200 30970 27000 31000
rect 25497 30968 27000 30970
rect 25497 30912 25502 30968
rect 25558 30912 27000 30968
rect 25497 30910 27000 30912
rect 25497 30907 25563 30910
rect 26200 30880 27000 30910
rect 7946 30496 8262 30497
rect 7946 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8262 30496
rect 7946 30431 8262 30432
rect 17946 30496 18262 30497
rect 17946 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18262 30496
rect 17946 30431 18262 30432
rect 25313 30154 25379 30157
rect 26200 30154 27000 30184
rect 25313 30152 27000 30154
rect 25313 30096 25318 30152
rect 25374 30096 27000 30152
rect 25313 30094 27000 30096
rect 25313 30091 25379 30094
rect 26200 30064 27000 30094
rect 2946 29952 3262 29953
rect 2946 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3262 29952
rect 2946 29887 3262 29888
rect 12946 29952 13262 29953
rect 12946 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13262 29952
rect 12946 29887 13262 29888
rect 22946 29952 23262 29953
rect 22946 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23262 29952
rect 22946 29887 23262 29888
rect 7946 29408 8262 29409
rect 7946 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8262 29408
rect 7946 29343 8262 29344
rect 17946 29408 18262 29409
rect 17946 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18262 29408
rect 17946 29343 18262 29344
rect 24945 29338 25011 29341
rect 26200 29338 27000 29368
rect 24945 29336 27000 29338
rect 24945 29280 24950 29336
rect 25006 29280 27000 29336
rect 24945 29278 27000 29280
rect 24945 29275 25011 29278
rect 26200 29248 27000 29278
rect 15837 29066 15903 29069
rect 17401 29066 17467 29069
rect 15837 29064 17467 29066
rect 15837 29008 15842 29064
rect 15898 29008 17406 29064
rect 17462 29008 17467 29064
rect 15837 29006 17467 29008
rect 15837 29003 15903 29006
rect 17401 29003 17467 29006
rect 2946 28864 3262 28865
rect 2946 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3262 28864
rect 2946 28799 3262 28800
rect 12946 28864 13262 28865
rect 12946 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13262 28864
rect 12946 28799 13262 28800
rect 22946 28864 23262 28865
rect 22946 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23262 28864
rect 22946 28799 23262 28800
rect 24485 28522 24551 28525
rect 26200 28522 27000 28552
rect 24485 28520 27000 28522
rect 24485 28464 24490 28520
rect 24546 28464 27000 28520
rect 24485 28462 27000 28464
rect 24485 28459 24551 28462
rect 26200 28432 27000 28462
rect 7946 28320 8262 28321
rect 7946 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8262 28320
rect 7946 28255 8262 28256
rect 17946 28320 18262 28321
rect 17946 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18262 28320
rect 17946 28255 18262 28256
rect 2946 27776 3262 27777
rect 2946 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3262 27776
rect 2946 27711 3262 27712
rect 12946 27776 13262 27777
rect 12946 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13262 27776
rect 12946 27711 13262 27712
rect 22946 27776 23262 27777
rect 22946 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23262 27776
rect 22946 27711 23262 27712
rect 24025 27706 24091 27709
rect 26200 27706 27000 27736
rect 24025 27704 27000 27706
rect 24025 27648 24030 27704
rect 24086 27648 27000 27704
rect 24025 27646 27000 27648
rect 24025 27643 24091 27646
rect 26200 27616 27000 27646
rect 7946 27232 8262 27233
rect 7946 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8262 27232
rect 7946 27167 8262 27168
rect 17946 27232 18262 27233
rect 17946 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18262 27232
rect 17946 27167 18262 27168
rect 25313 26890 25379 26893
rect 26200 26890 27000 26920
rect 25313 26888 27000 26890
rect 25313 26832 25318 26888
rect 25374 26832 27000 26888
rect 25313 26830 27000 26832
rect 25313 26827 25379 26830
rect 26200 26800 27000 26830
rect 2946 26688 3262 26689
rect 2946 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3262 26688
rect 2946 26623 3262 26624
rect 12946 26688 13262 26689
rect 12946 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13262 26688
rect 12946 26623 13262 26624
rect 22946 26688 23262 26689
rect 22946 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23262 26688
rect 22946 26623 23262 26624
rect 7946 26144 8262 26145
rect 7946 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8262 26144
rect 7946 26079 8262 26080
rect 17946 26144 18262 26145
rect 17946 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18262 26144
rect 17946 26079 18262 26080
rect 24853 26074 24919 26077
rect 26200 26074 27000 26104
rect 24853 26072 27000 26074
rect 24853 26016 24858 26072
rect 24914 26016 27000 26072
rect 24853 26014 27000 26016
rect 24853 26011 24919 26014
rect 26200 25984 27000 26014
rect 17585 25940 17651 25941
rect 17534 25938 17540 25940
rect 17494 25878 17540 25938
rect 17604 25936 17651 25940
rect 17646 25880 17651 25936
rect 17534 25876 17540 25878
rect 17604 25876 17651 25880
rect 17585 25875 17651 25876
rect 2946 25600 3262 25601
rect 2946 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3262 25600
rect 2946 25535 3262 25536
rect 12946 25600 13262 25601
rect 12946 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13262 25600
rect 12946 25535 13262 25536
rect 22946 25600 23262 25601
rect 22946 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23262 25600
rect 22946 25535 23262 25536
rect 25129 25258 25195 25261
rect 26200 25258 27000 25288
rect 25129 25256 27000 25258
rect 25129 25200 25134 25256
rect 25190 25200 27000 25256
rect 25129 25198 27000 25200
rect 25129 25195 25195 25198
rect 26200 25168 27000 25198
rect 15326 25060 15332 25124
rect 15396 25122 15402 25124
rect 15561 25122 15627 25125
rect 15396 25120 15627 25122
rect 15396 25064 15566 25120
rect 15622 25064 15627 25120
rect 15396 25062 15627 25064
rect 15396 25060 15402 25062
rect 15561 25059 15627 25062
rect 7946 25056 8262 25057
rect 7946 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8262 25056
rect 7946 24991 8262 24992
rect 17946 25056 18262 25057
rect 17946 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18262 25056
rect 17946 24991 18262 24992
rect 19885 24988 19951 24989
rect 19885 24984 19932 24988
rect 19996 24986 20002 24988
rect 19885 24928 19890 24984
rect 19885 24924 19932 24928
rect 19996 24926 20042 24986
rect 19996 24924 20002 24926
rect 19885 24923 19951 24924
rect 2946 24512 3262 24513
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 23841 24442 23907 24445
rect 26200 24442 27000 24472
rect 23841 24440 27000 24442
rect 23841 24384 23846 24440
rect 23902 24384 27000 24440
rect 23841 24382 27000 24384
rect 23841 24379 23907 24382
rect 26200 24352 27000 24382
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 24761 23626 24827 23629
rect 26200 23626 27000 23656
rect 24761 23624 27000 23626
rect 24761 23568 24766 23624
rect 24822 23568 27000 23624
rect 24761 23566 27000 23568
rect 24761 23563 24827 23566
rect 26200 23536 27000 23566
rect 18873 23490 18939 23493
rect 19006 23490 19012 23492
rect 18873 23488 19012 23490
rect 18873 23432 18878 23488
rect 18934 23432 19012 23488
rect 18873 23430 19012 23432
rect 18873 23427 18939 23430
rect 19006 23428 19012 23430
rect 19076 23428 19082 23492
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 7946 22880 8262 22881
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 16757 22812 16823 22813
rect 16757 22808 16804 22812
rect 16868 22810 16874 22812
rect 24853 22810 24919 22813
rect 26200 22810 27000 22840
rect 16757 22752 16762 22808
rect 16757 22748 16804 22752
rect 16868 22750 16914 22810
rect 24853 22808 27000 22810
rect 24853 22752 24858 22808
rect 24914 22752 27000 22808
rect 24853 22750 27000 22752
rect 16868 22748 16874 22750
rect 16757 22747 16823 22748
rect 24853 22747 24919 22750
rect 26200 22720 27000 22750
rect 19149 22402 19215 22405
rect 19701 22402 19767 22405
rect 20437 22404 20503 22405
rect 20437 22402 20484 22404
rect 19149 22400 19767 22402
rect 19149 22344 19154 22400
rect 19210 22344 19706 22400
rect 19762 22344 19767 22400
rect 19149 22342 19767 22344
rect 20392 22400 20484 22402
rect 20392 22344 20442 22400
rect 20392 22342 20484 22344
rect 19149 22339 19215 22342
rect 19701 22339 19767 22342
rect 20437 22340 20484 22342
rect 20548 22340 20554 22404
rect 20437 22339 20503 22340
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 23381 21994 23447 21997
rect 26200 21994 27000 22024
rect 23381 21992 27000 21994
rect 23381 21936 23386 21992
rect 23442 21936 27000 21992
rect 23381 21934 27000 21936
rect 23381 21931 23447 21934
rect 26200 21904 27000 21934
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 2946 21248 3262 21249
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 24853 21178 24919 21181
rect 26200 21178 27000 21208
rect 24853 21176 27000 21178
rect 24853 21120 24858 21176
rect 24914 21120 27000 21176
rect 24853 21118 27000 21120
rect 24853 21115 24919 21118
rect 26200 21088 27000 21118
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 24669 20362 24735 20365
rect 26200 20362 27000 20392
rect 24669 20360 27000 20362
rect 24669 20304 24674 20360
rect 24730 20304 27000 20360
rect 24669 20302 27000 20304
rect 24669 20299 24735 20302
rect 26200 20272 27000 20302
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 22134 19756 22140 19820
rect 22204 19818 22210 19820
rect 23105 19818 23171 19821
rect 22204 19816 23171 19818
rect 22204 19760 23110 19816
rect 23166 19760 23171 19816
rect 22204 19758 23171 19760
rect 22204 19756 22210 19758
rect 23105 19755 23171 19758
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 23841 19546 23907 19549
rect 26200 19546 27000 19576
rect 23841 19544 27000 19546
rect 23841 19488 23846 19544
rect 23902 19488 27000 19544
rect 23841 19486 27000 19488
rect 23841 19483 23907 19486
rect 26200 19456 27000 19486
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 24853 18730 24919 18733
rect 26200 18730 27000 18760
rect 24853 18728 27000 18730
rect 24853 18672 24858 18728
rect 24914 18672 27000 18728
rect 24853 18670 27000 18672
rect 24853 18667 24919 18670
rect 26200 18640 27000 18670
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 16849 18050 16915 18053
rect 17350 18050 17356 18052
rect 16849 18048 17356 18050
rect 16849 17992 16854 18048
rect 16910 17992 17356 18048
rect 16849 17990 17356 17992
rect 16849 17987 16915 17990
rect 17350 17988 17356 17990
rect 17420 17988 17426 18052
rect 2946 17984 3262 17985
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 24945 17914 25011 17917
rect 26200 17914 27000 17944
rect 24945 17912 27000 17914
rect 24945 17856 24950 17912
rect 25006 17856 27000 17912
rect 24945 17854 27000 17856
rect 24945 17851 25011 17854
rect 26200 17824 27000 17854
rect 12566 17444 12572 17508
rect 12636 17506 12642 17508
rect 12709 17506 12775 17509
rect 12636 17504 12775 17506
rect 12636 17448 12714 17504
rect 12770 17448 12775 17504
rect 12636 17446 12775 17448
rect 12636 17444 12642 17446
rect 12709 17443 12775 17446
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 17401 17370 17467 17373
rect 17534 17370 17540 17372
rect 17401 17368 17540 17370
rect 17401 17312 17406 17368
rect 17462 17312 17540 17368
rect 17401 17310 17540 17312
rect 17401 17307 17467 17310
rect 17534 17308 17540 17310
rect 17604 17308 17610 17372
rect 23841 17098 23907 17101
rect 26200 17098 27000 17128
rect 23841 17096 27000 17098
rect 23841 17040 23846 17096
rect 23902 17040 27000 17096
rect 23841 17038 27000 17040
rect 23841 17035 23907 17038
rect 26200 17008 27000 17038
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 17125 16692 17191 16693
rect 17125 16688 17172 16692
rect 17236 16690 17242 16692
rect 17125 16632 17130 16688
rect 17125 16628 17172 16632
rect 17236 16630 17282 16690
rect 17236 16628 17242 16630
rect 17125 16627 17191 16628
rect 21909 16554 21975 16557
rect 22737 16554 22803 16557
rect 21909 16552 22803 16554
rect 21909 16496 21914 16552
rect 21970 16496 22742 16552
rect 22798 16496 22803 16552
rect 21909 16494 22803 16496
rect 21909 16491 21975 16494
rect 22737 16491 22803 16494
rect 7946 16352 8262 16353
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 16849 16284 16915 16285
rect 16798 16220 16804 16284
rect 16868 16282 16915 16284
rect 24761 16282 24827 16285
rect 26200 16282 27000 16312
rect 16868 16280 16960 16282
rect 16910 16224 16960 16280
rect 16868 16222 16960 16224
rect 24761 16280 27000 16282
rect 24761 16224 24766 16280
rect 24822 16224 27000 16280
rect 24761 16222 27000 16224
rect 16868 16220 16915 16222
rect 16849 16219 16915 16220
rect 24761 16219 24827 16222
rect 26200 16192 27000 16222
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 23289 15466 23355 15469
rect 26200 15466 27000 15496
rect 23289 15464 27000 15466
rect 23289 15408 23294 15464
rect 23350 15408 27000 15464
rect 23289 15406 27000 15408
rect 23289 15403 23355 15406
rect 26200 15376 27000 15406
rect 16982 15268 16988 15332
rect 17052 15330 17058 15332
rect 17309 15330 17375 15333
rect 17052 15328 17375 15330
rect 17052 15272 17314 15328
rect 17370 15272 17375 15328
rect 17052 15270 17375 15272
rect 17052 15268 17058 15270
rect 17309 15267 17375 15270
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 24853 14650 24919 14653
rect 26200 14650 27000 14680
rect 24853 14648 27000 14650
rect 24853 14592 24858 14648
rect 24914 14592 27000 14648
rect 24853 14590 27000 14592
rect 24853 14587 24919 14590
rect 26200 14560 27000 14590
rect 13537 14242 13603 14245
rect 14733 14244 14799 14245
rect 13670 14242 13676 14244
rect 13537 14240 13676 14242
rect 13537 14184 13542 14240
rect 13598 14184 13676 14240
rect 13537 14182 13676 14184
rect 13537 14179 13603 14182
rect 13670 14180 13676 14182
rect 13740 14180 13746 14244
rect 14733 14242 14780 14244
rect 14688 14240 14780 14242
rect 14688 14184 14738 14240
rect 14688 14182 14780 14184
rect 14733 14180 14780 14182
rect 14844 14180 14850 14244
rect 14733 14179 14799 14180
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 23841 13834 23907 13837
rect 26200 13834 27000 13864
rect 23841 13832 27000 13834
rect 23841 13776 23846 13832
rect 23902 13776 27000 13832
rect 23841 13774 27000 13776
rect 23841 13771 23907 13774
rect 26200 13744 27000 13774
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 17401 13564 17467 13565
rect 17350 13500 17356 13564
rect 17420 13562 17467 13564
rect 17420 13560 17512 13562
rect 17462 13504 17512 13560
rect 17420 13502 17512 13504
rect 17420 13500 17467 13502
rect 17401 13499 17467 13500
rect 7946 13088 8262 13089
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 24761 13018 24827 13021
rect 26200 13018 27000 13048
rect 24761 13016 27000 13018
rect 24761 12960 24766 13016
rect 24822 12960 27000 13016
rect 24761 12958 27000 12960
rect 24761 12955 24827 12958
rect 26200 12928 27000 12958
rect 13077 12746 13143 12749
rect 12758 12744 13143 12746
rect 12758 12688 13082 12744
rect 13138 12688 13143 12744
rect 12758 12686 13143 12688
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12433 12474 12499 12477
rect 12758 12474 12818 12686
rect 13077 12683 13143 12686
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 12433 12472 12818 12474
rect 12433 12416 12438 12472
rect 12494 12416 12818 12472
rect 12433 12414 12818 12416
rect 14549 12474 14615 12477
rect 14917 12474 14983 12477
rect 14549 12472 14983 12474
rect 14549 12416 14554 12472
rect 14610 12416 14922 12472
rect 14978 12416 14983 12472
rect 14549 12414 14983 12416
rect 12433 12411 12499 12414
rect 14549 12411 14615 12414
rect 14917 12411 14983 12414
rect 16297 12474 16363 12477
rect 16297 12472 16590 12474
rect 16297 12416 16302 12472
rect 16358 12416 16590 12472
rect 16297 12414 16590 12416
rect 16297 12411 16363 12414
rect 16530 12338 16590 12414
rect 19977 12338 20043 12341
rect 16530 12336 20043 12338
rect 16530 12280 19982 12336
rect 20038 12280 20043 12336
rect 16530 12278 20043 12280
rect 19977 12275 20043 12278
rect 24945 12202 25011 12205
rect 26200 12202 27000 12232
rect 24945 12200 27000 12202
rect 24945 12144 24950 12200
rect 25006 12144 27000 12200
rect 24945 12142 27000 12144
rect 24945 12139 25011 12142
rect 26200 12112 27000 12142
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 11789 11930 11855 11933
rect 15285 11930 15351 11933
rect 11789 11928 15351 11930
rect 11789 11872 11794 11928
rect 11850 11872 15290 11928
rect 15346 11872 15351 11928
rect 11789 11870 15351 11872
rect 11789 11867 11855 11870
rect 15285 11867 15351 11870
rect 12065 11794 12131 11797
rect 12341 11794 12407 11797
rect 12065 11792 12407 11794
rect 12065 11736 12070 11792
rect 12126 11736 12346 11792
rect 12402 11736 12407 11792
rect 12065 11734 12407 11736
rect 12065 11731 12131 11734
rect 12341 11731 12407 11734
rect 13670 11732 13676 11796
rect 13740 11794 13746 11796
rect 19333 11794 19399 11797
rect 13740 11792 19399 11794
rect 13740 11736 19338 11792
rect 19394 11736 19399 11792
rect 13740 11734 19399 11736
rect 13740 11732 13746 11734
rect 19333 11731 19399 11734
rect 2946 11456 3262 11457
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 24853 11386 24919 11389
rect 26200 11386 27000 11416
rect 24853 11384 27000 11386
rect 24853 11328 24858 11384
rect 24914 11328 27000 11384
rect 24853 11326 27000 11328
rect 24853 11323 24919 11326
rect 26200 11296 27000 11326
rect 11881 11250 11947 11253
rect 13169 11250 13235 11253
rect 16021 11250 16087 11253
rect 16297 11250 16363 11253
rect 11881 11248 16363 11250
rect 11881 11192 11886 11248
rect 11942 11192 13174 11248
rect 13230 11192 16026 11248
rect 16082 11192 16302 11248
rect 16358 11192 16363 11248
rect 11881 11190 16363 11192
rect 11881 11187 11947 11190
rect 13169 11187 13235 11190
rect 16021 11187 16087 11190
rect 16297 11187 16363 11190
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 19241 10842 19307 10845
rect 24301 10842 24367 10845
rect 19241 10840 24367 10842
rect 19241 10784 19246 10840
rect 19302 10784 24306 10840
rect 24362 10784 24367 10840
rect 19241 10782 24367 10784
rect 19241 10779 19307 10782
rect 24301 10779 24367 10782
rect 15009 10706 15075 10709
rect 19517 10706 19583 10709
rect 15009 10704 19583 10706
rect 15009 10648 15014 10704
rect 15070 10648 19522 10704
rect 19578 10648 19583 10704
rect 15009 10646 19583 10648
rect 15009 10643 15075 10646
rect 19517 10643 19583 10646
rect 20621 10706 20687 10709
rect 23657 10706 23723 10709
rect 20621 10704 23723 10706
rect 20621 10648 20626 10704
rect 20682 10648 23662 10704
rect 23718 10648 23723 10704
rect 20621 10646 23723 10648
rect 20621 10643 20687 10646
rect 23657 10643 23723 10646
rect 14181 10570 14247 10573
rect 17769 10570 17835 10573
rect 14181 10568 17835 10570
rect 14181 10512 14186 10568
rect 14242 10512 17774 10568
rect 17830 10512 17835 10568
rect 14181 10510 17835 10512
rect 14181 10507 14247 10510
rect 17769 10507 17835 10510
rect 23841 10570 23907 10573
rect 26200 10570 27000 10600
rect 23841 10568 27000 10570
rect 23841 10512 23846 10568
rect 23902 10512 27000 10568
rect 23841 10510 27000 10512
rect 23841 10507 23907 10510
rect 26200 10480 27000 10510
rect 21265 10434 21331 10437
rect 22277 10434 22343 10437
rect 21265 10432 22343 10434
rect 21265 10376 21270 10432
rect 21326 10376 22282 10432
rect 22338 10376 22343 10432
rect 21265 10374 22343 10376
rect 21265 10371 21331 10374
rect 22277 10371 22343 10374
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 18454 10236 18460 10300
rect 18524 10298 18530 10300
rect 18873 10298 18939 10301
rect 18524 10296 18939 10298
rect 18524 10240 18878 10296
rect 18934 10240 18939 10296
rect 18524 10238 18939 10240
rect 18524 10236 18530 10238
rect 18873 10235 18939 10238
rect 19517 10298 19583 10301
rect 22553 10298 22619 10301
rect 19517 10296 22619 10298
rect 19517 10240 19522 10296
rect 19578 10240 22558 10296
rect 22614 10240 22619 10296
rect 19517 10238 22619 10240
rect 19517 10235 19583 10238
rect 22553 10235 22619 10238
rect 20161 10026 20227 10029
rect 22369 10026 22435 10029
rect 20161 10024 22435 10026
rect 20161 9968 20166 10024
rect 20222 9968 22374 10024
rect 22430 9968 22435 10024
rect 20161 9966 22435 9968
rect 20161 9963 20227 9966
rect 22369 9963 22435 9966
rect 7946 9824 8262 9825
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 24761 9754 24827 9757
rect 26200 9754 27000 9784
rect 24761 9752 27000 9754
rect 24761 9696 24766 9752
rect 24822 9696 27000 9752
rect 24761 9694 27000 9696
rect 24761 9691 24827 9694
rect 26200 9664 27000 9694
rect 17769 9618 17835 9621
rect 18689 9618 18755 9621
rect 17769 9616 18755 9618
rect 17769 9560 17774 9616
rect 17830 9560 18694 9616
rect 18750 9560 18755 9616
rect 17769 9558 18755 9560
rect 17769 9555 17835 9558
rect 18689 9555 18755 9558
rect 20621 9482 20687 9485
rect 22093 9482 22159 9485
rect 24485 9482 24551 9485
rect 20621 9480 24551 9482
rect 20621 9424 20626 9480
rect 20682 9424 22098 9480
rect 22154 9424 24490 9480
rect 24546 9424 24551 9480
rect 20621 9422 24551 9424
rect 20621 9419 20687 9422
rect 22093 9419 22159 9422
rect 24485 9419 24551 9422
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 13537 8938 13603 8941
rect 15929 8938 15995 8941
rect 13537 8936 15995 8938
rect 13537 8880 13542 8936
rect 13598 8880 15934 8936
rect 15990 8880 15995 8936
rect 13537 8878 15995 8880
rect 13537 8875 13603 8878
rect 15929 8875 15995 8878
rect 16849 8938 16915 8941
rect 19241 8938 19307 8941
rect 16849 8936 19307 8938
rect 16849 8880 16854 8936
rect 16910 8880 19246 8936
rect 19302 8880 19307 8936
rect 16849 8878 19307 8880
rect 16849 8875 16915 8878
rect 19241 8875 19307 8878
rect 24945 8938 25011 8941
rect 26200 8938 27000 8968
rect 24945 8936 27000 8938
rect 24945 8880 24950 8936
rect 25006 8880 27000 8936
rect 24945 8878 27000 8880
rect 24945 8875 25011 8878
rect 26200 8848 27000 8878
rect 0 8802 800 8832
rect 3509 8802 3575 8805
rect 0 8800 3575 8802
rect 0 8744 3514 8800
rect 3570 8744 3575 8800
rect 0 8742 3575 8744
rect 0 8712 800 8742
rect 3509 8739 3575 8742
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 16849 8532 16915 8533
rect 16798 8468 16804 8532
rect 16868 8530 16915 8532
rect 17769 8530 17835 8533
rect 16868 8528 17835 8530
rect 16910 8472 17774 8528
rect 17830 8472 17835 8528
rect 16868 8470 17835 8472
rect 16868 8468 16915 8470
rect 16849 8467 16915 8468
rect 17769 8467 17835 8470
rect 22318 8332 22324 8396
rect 22388 8394 22394 8396
rect 22645 8394 22711 8397
rect 22388 8392 22711 8394
rect 22388 8336 22650 8392
rect 22706 8336 22711 8392
rect 22388 8334 22711 8336
rect 22388 8332 22394 8334
rect 22645 8331 22711 8334
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 25129 8122 25195 8125
rect 26200 8122 27000 8152
rect 25129 8120 27000 8122
rect 25129 8064 25134 8120
rect 25190 8064 27000 8120
rect 25129 8062 27000 8064
rect 25129 8059 25195 8062
rect 26200 8032 27000 8062
rect 14549 7986 14615 7989
rect 15193 7986 15259 7989
rect 14549 7984 15259 7986
rect 14549 7928 14554 7984
rect 14610 7928 15198 7984
rect 15254 7928 15259 7984
rect 14549 7926 15259 7928
rect 14549 7923 14615 7926
rect 15193 7923 15259 7926
rect 13905 7850 13971 7853
rect 18229 7850 18295 7853
rect 13905 7848 18295 7850
rect 13905 7792 13910 7848
rect 13966 7792 18234 7848
rect 18290 7792 18295 7848
rect 13905 7790 18295 7792
rect 13905 7787 13971 7790
rect 18229 7787 18295 7790
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 15326 7244 15332 7308
rect 15396 7306 15402 7308
rect 15469 7306 15535 7309
rect 15396 7304 15535 7306
rect 15396 7248 15474 7304
rect 15530 7248 15535 7304
rect 15396 7246 15535 7248
rect 15396 7244 15402 7246
rect 15469 7243 15535 7246
rect 24853 7306 24919 7309
rect 26200 7306 27000 7336
rect 24853 7304 27000 7306
rect 24853 7248 24858 7304
rect 24914 7248 27000 7304
rect 24853 7246 27000 7248
rect 24853 7243 24919 7246
rect 26200 7216 27000 7246
rect 17585 7170 17651 7173
rect 19241 7170 19307 7173
rect 17585 7168 19307 7170
rect 17585 7112 17590 7168
rect 17646 7112 19246 7168
rect 19302 7112 19307 7168
rect 17585 7110 19307 7112
rect 17585 7107 17651 7110
rect 19241 7107 19307 7110
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 17677 7034 17743 7037
rect 19241 7034 19307 7037
rect 17677 7032 19307 7034
rect 17677 6976 17682 7032
rect 17738 6976 19246 7032
rect 19302 6976 19307 7032
rect 17677 6974 19307 6976
rect 17677 6971 17743 6974
rect 19241 6971 19307 6974
rect 13261 6898 13327 6901
rect 16798 6898 16804 6900
rect 13261 6896 16804 6898
rect 13261 6840 13266 6896
rect 13322 6840 16804 6896
rect 13261 6838 16804 6840
rect 13261 6835 13327 6838
rect 16798 6836 16804 6838
rect 16868 6836 16874 6900
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 3417 6490 3483 6493
rect 0 6488 3483 6490
rect 0 6432 3422 6488
rect 3478 6432 3483 6488
rect 0 6430 3483 6432
rect 0 6400 800 6430
rect 3417 6427 3483 6430
rect 24945 6490 25011 6493
rect 26200 6490 27000 6520
rect 24945 6488 27000 6490
rect 24945 6432 24950 6488
rect 25006 6432 27000 6488
rect 24945 6430 27000 6432
rect 24945 6427 25011 6430
rect 26200 6400 27000 6430
rect 10869 6218 10935 6221
rect 12893 6218 12959 6221
rect 15469 6218 15535 6221
rect 10869 6216 15535 6218
rect 10869 6160 10874 6216
rect 10930 6160 12898 6216
rect 12954 6160 15474 6216
rect 15530 6160 15535 6216
rect 10869 6158 15535 6160
rect 10869 6155 10935 6158
rect 12893 6155 12959 6158
rect 15469 6155 15535 6158
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 22829 5674 22895 5677
rect 26200 5674 27000 5704
rect 22829 5672 27000 5674
rect 22829 5616 22834 5672
rect 22890 5616 27000 5672
rect 22829 5614 27000 5616
rect 22829 5611 22895 5614
rect 26200 5584 27000 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 22001 5130 22067 5133
rect 22001 5128 23858 5130
rect 22001 5072 22006 5128
rect 22062 5072 23858 5128
rect 22001 5070 23858 5072
rect 22001 5067 22067 5070
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 23798 4858 23858 5070
rect 26200 4858 27000 4888
rect 23798 4798 27000 4858
rect 26200 4768 27000 4798
rect 12249 4722 12315 4725
rect 22318 4722 22324 4724
rect 12249 4720 22324 4722
rect 12249 4664 12254 4720
rect 12310 4664 22324 4720
rect 12249 4662 22324 4664
rect 12249 4659 12315 4662
rect 22318 4660 22324 4662
rect 22388 4660 22394 4724
rect 12249 4586 12315 4589
rect 23749 4586 23815 4589
rect 12249 4584 23815 4586
rect 12249 4528 12254 4584
rect 12310 4528 23754 4584
rect 23810 4528 23815 4584
rect 12249 4526 23815 4528
rect 12249 4523 12315 4526
rect 23749 4523 23815 4526
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 0 4178 800 4208
rect 22134 4178 22140 4180
rect 0 4118 22140 4178
rect 0 4088 800 4118
rect 22134 4116 22140 4118
rect 22204 4116 22210 4180
rect 10961 4042 11027 4045
rect 17309 4042 17375 4045
rect 22737 4042 22803 4045
rect 10961 4040 15762 4042
rect 10961 3984 10966 4040
rect 11022 3984 15762 4040
rect 10961 3982 15762 3984
rect 10961 3979 11027 3982
rect 15702 3906 15762 3982
rect 17309 4040 22803 4042
rect 17309 3984 17314 4040
rect 17370 3984 22742 4040
rect 22798 3984 22803 4040
rect 17309 3982 22803 3984
rect 17309 3979 17375 3982
rect 22737 3979 22803 3982
rect 24393 4042 24459 4045
rect 26200 4042 27000 4072
rect 24393 4040 27000 4042
rect 24393 3984 24398 4040
rect 24454 3984 27000 4040
rect 24393 3982 27000 3984
rect 24393 3979 24459 3982
rect 26200 3952 27000 3982
rect 18454 3906 18460 3908
rect 15702 3846 18460 3906
rect 18454 3844 18460 3846
rect 18524 3844 18530 3908
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 14825 3770 14891 3773
rect 14825 3768 22110 3770
rect 14825 3712 14830 3768
rect 14886 3712 22110 3768
rect 14825 3710 22110 3712
rect 14825 3707 14891 3710
rect 5165 3634 5231 3637
rect 12566 3634 12572 3636
rect 5165 3632 12572 3634
rect 5165 3576 5170 3632
rect 5226 3576 12572 3632
rect 5165 3574 12572 3576
rect 5165 3571 5231 3574
rect 12566 3572 12572 3574
rect 12636 3572 12642 3636
rect 14457 3634 14523 3637
rect 16982 3634 16988 3636
rect 14457 3632 16988 3634
rect 14457 3576 14462 3632
rect 14518 3576 16988 3632
rect 14457 3574 16988 3576
rect 14457 3571 14523 3574
rect 16982 3572 16988 3574
rect 17052 3572 17058 3636
rect 22050 3634 22110 3710
rect 24945 3634 25011 3637
rect 22050 3632 25011 3634
rect 22050 3576 24950 3632
rect 25006 3576 25011 3632
rect 22050 3574 25011 3576
rect 24945 3571 25011 3574
rect 19006 3436 19012 3500
rect 19076 3498 19082 3500
rect 23933 3498 23999 3501
rect 19076 3496 23999 3498
rect 19076 3440 23938 3496
rect 23994 3440 23999 3496
rect 19076 3438 23999 3440
rect 19076 3436 19082 3438
rect 23933 3435 23999 3438
rect 7946 3296 8262 3297
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 22369 3226 22435 3229
rect 26200 3226 27000 3256
rect 22369 3224 27000 3226
rect 22369 3168 22374 3224
rect 22430 3168 27000 3224
rect 22369 3166 27000 3168
rect 22369 3163 22435 3166
rect 26200 3136 27000 3166
rect 13169 3090 13235 3093
rect 17166 3090 17172 3092
rect 13169 3088 17172 3090
rect 13169 3032 13174 3088
rect 13230 3032 17172 3088
rect 13169 3030 17172 3032
rect 13169 3027 13235 3030
rect 17166 3028 17172 3030
rect 17236 3028 17242 3092
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 5441 2546 5507 2549
rect 14774 2546 14780 2548
rect 5441 2544 14780 2546
rect 5441 2488 5446 2544
rect 5502 2488 14780 2544
rect 5441 2486 14780 2488
rect 5441 2483 5507 2486
rect 14774 2484 14780 2486
rect 14844 2484 14850 2548
rect 16297 2410 16363 2413
rect 19926 2410 19932 2412
rect 16297 2408 19932 2410
rect 16297 2352 16302 2408
rect 16358 2352 19932 2408
rect 16297 2350 19932 2352
rect 16297 2347 16363 2350
rect 19926 2348 19932 2350
rect 19996 2348 20002 2412
rect 22093 2410 22159 2413
rect 26200 2410 27000 2440
rect 22093 2408 27000 2410
rect 22093 2352 22098 2408
rect 22154 2352 27000 2408
rect 22093 2350 27000 2352
rect 22093 2347 22159 2350
rect 26200 2320 27000 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 0 1866 800 1896
rect 20478 1866 20484 1868
rect 0 1806 20484 1866
rect 0 1776 800 1806
rect 20478 1804 20484 1806
rect 20548 1804 20554 1868
rect 22277 1594 22343 1597
rect 26200 1594 27000 1624
rect 22277 1592 27000 1594
rect 22277 1536 22282 1592
rect 22338 1536 27000 1592
rect 22277 1534 27000 1536
rect 22277 1531 22343 1534
rect 26200 1504 27000 1534
rect 25313 778 25379 781
rect 26200 778 27000 808
rect 25313 776 27000 778
rect 25313 720 25318 776
rect 25374 720 27000 776
rect 25313 718 27000 720
rect 25313 715 25379 718
rect 26200 688 27000 718
<< via3 >>
rect 7952 54428 8016 54432
rect 7952 54372 7956 54428
rect 7956 54372 8012 54428
rect 8012 54372 8016 54428
rect 7952 54368 8016 54372
rect 8032 54428 8096 54432
rect 8032 54372 8036 54428
rect 8036 54372 8092 54428
rect 8092 54372 8096 54428
rect 8032 54368 8096 54372
rect 8112 54428 8176 54432
rect 8112 54372 8116 54428
rect 8116 54372 8172 54428
rect 8172 54372 8176 54428
rect 8112 54368 8176 54372
rect 8192 54428 8256 54432
rect 8192 54372 8196 54428
rect 8196 54372 8252 54428
rect 8252 54372 8256 54428
rect 8192 54368 8256 54372
rect 17952 54428 18016 54432
rect 17952 54372 17956 54428
rect 17956 54372 18012 54428
rect 18012 54372 18016 54428
rect 17952 54368 18016 54372
rect 18032 54428 18096 54432
rect 18032 54372 18036 54428
rect 18036 54372 18092 54428
rect 18092 54372 18096 54428
rect 18032 54368 18096 54372
rect 18112 54428 18176 54432
rect 18112 54372 18116 54428
rect 18116 54372 18172 54428
rect 18172 54372 18176 54428
rect 18112 54368 18176 54372
rect 18192 54428 18256 54432
rect 18192 54372 18196 54428
rect 18196 54372 18252 54428
rect 18252 54372 18256 54428
rect 18192 54368 18256 54372
rect 2952 53884 3016 53888
rect 2952 53828 2956 53884
rect 2956 53828 3012 53884
rect 3012 53828 3016 53884
rect 2952 53824 3016 53828
rect 3032 53884 3096 53888
rect 3032 53828 3036 53884
rect 3036 53828 3092 53884
rect 3092 53828 3096 53884
rect 3032 53824 3096 53828
rect 3112 53884 3176 53888
rect 3112 53828 3116 53884
rect 3116 53828 3172 53884
rect 3172 53828 3176 53884
rect 3112 53824 3176 53828
rect 3192 53884 3256 53888
rect 3192 53828 3196 53884
rect 3196 53828 3252 53884
rect 3252 53828 3256 53884
rect 3192 53824 3256 53828
rect 12952 53884 13016 53888
rect 12952 53828 12956 53884
rect 12956 53828 13012 53884
rect 13012 53828 13016 53884
rect 12952 53824 13016 53828
rect 13032 53884 13096 53888
rect 13032 53828 13036 53884
rect 13036 53828 13092 53884
rect 13092 53828 13096 53884
rect 13032 53824 13096 53828
rect 13112 53884 13176 53888
rect 13112 53828 13116 53884
rect 13116 53828 13172 53884
rect 13172 53828 13176 53884
rect 13112 53824 13176 53828
rect 13192 53884 13256 53888
rect 13192 53828 13196 53884
rect 13196 53828 13252 53884
rect 13252 53828 13256 53884
rect 13192 53824 13256 53828
rect 22952 53884 23016 53888
rect 22952 53828 22956 53884
rect 22956 53828 23012 53884
rect 23012 53828 23016 53884
rect 22952 53824 23016 53828
rect 23032 53884 23096 53888
rect 23032 53828 23036 53884
rect 23036 53828 23092 53884
rect 23092 53828 23096 53884
rect 23032 53824 23096 53828
rect 23112 53884 23176 53888
rect 23112 53828 23116 53884
rect 23116 53828 23172 53884
rect 23172 53828 23176 53884
rect 23112 53824 23176 53828
rect 23192 53884 23256 53888
rect 23192 53828 23196 53884
rect 23196 53828 23252 53884
rect 23252 53828 23256 53884
rect 23192 53824 23256 53828
rect 7952 53340 8016 53344
rect 7952 53284 7956 53340
rect 7956 53284 8012 53340
rect 8012 53284 8016 53340
rect 7952 53280 8016 53284
rect 8032 53340 8096 53344
rect 8032 53284 8036 53340
rect 8036 53284 8092 53340
rect 8092 53284 8096 53340
rect 8032 53280 8096 53284
rect 8112 53340 8176 53344
rect 8112 53284 8116 53340
rect 8116 53284 8172 53340
rect 8172 53284 8176 53340
rect 8112 53280 8176 53284
rect 8192 53340 8256 53344
rect 8192 53284 8196 53340
rect 8196 53284 8252 53340
rect 8252 53284 8256 53340
rect 8192 53280 8256 53284
rect 17952 53340 18016 53344
rect 17952 53284 17956 53340
rect 17956 53284 18012 53340
rect 18012 53284 18016 53340
rect 17952 53280 18016 53284
rect 18032 53340 18096 53344
rect 18032 53284 18036 53340
rect 18036 53284 18092 53340
rect 18092 53284 18096 53340
rect 18032 53280 18096 53284
rect 18112 53340 18176 53344
rect 18112 53284 18116 53340
rect 18116 53284 18172 53340
rect 18172 53284 18176 53340
rect 18112 53280 18176 53284
rect 18192 53340 18256 53344
rect 18192 53284 18196 53340
rect 18196 53284 18252 53340
rect 18252 53284 18256 53340
rect 18192 53280 18256 53284
rect 2952 52796 3016 52800
rect 2952 52740 2956 52796
rect 2956 52740 3012 52796
rect 3012 52740 3016 52796
rect 2952 52736 3016 52740
rect 3032 52796 3096 52800
rect 3032 52740 3036 52796
rect 3036 52740 3092 52796
rect 3092 52740 3096 52796
rect 3032 52736 3096 52740
rect 3112 52796 3176 52800
rect 3112 52740 3116 52796
rect 3116 52740 3172 52796
rect 3172 52740 3176 52796
rect 3112 52736 3176 52740
rect 3192 52796 3256 52800
rect 3192 52740 3196 52796
rect 3196 52740 3252 52796
rect 3252 52740 3256 52796
rect 3192 52736 3256 52740
rect 12952 52796 13016 52800
rect 12952 52740 12956 52796
rect 12956 52740 13012 52796
rect 13012 52740 13016 52796
rect 12952 52736 13016 52740
rect 13032 52796 13096 52800
rect 13032 52740 13036 52796
rect 13036 52740 13092 52796
rect 13092 52740 13096 52796
rect 13032 52736 13096 52740
rect 13112 52796 13176 52800
rect 13112 52740 13116 52796
rect 13116 52740 13172 52796
rect 13172 52740 13176 52796
rect 13112 52736 13176 52740
rect 13192 52796 13256 52800
rect 13192 52740 13196 52796
rect 13196 52740 13252 52796
rect 13252 52740 13256 52796
rect 13192 52736 13256 52740
rect 22952 52796 23016 52800
rect 22952 52740 22956 52796
rect 22956 52740 23012 52796
rect 23012 52740 23016 52796
rect 22952 52736 23016 52740
rect 23032 52796 23096 52800
rect 23032 52740 23036 52796
rect 23036 52740 23092 52796
rect 23092 52740 23096 52796
rect 23032 52736 23096 52740
rect 23112 52796 23176 52800
rect 23112 52740 23116 52796
rect 23116 52740 23172 52796
rect 23172 52740 23176 52796
rect 23112 52736 23176 52740
rect 23192 52796 23256 52800
rect 23192 52740 23196 52796
rect 23196 52740 23252 52796
rect 23252 52740 23256 52796
rect 23192 52736 23256 52740
rect 7952 52252 8016 52256
rect 7952 52196 7956 52252
rect 7956 52196 8012 52252
rect 8012 52196 8016 52252
rect 7952 52192 8016 52196
rect 8032 52252 8096 52256
rect 8032 52196 8036 52252
rect 8036 52196 8092 52252
rect 8092 52196 8096 52252
rect 8032 52192 8096 52196
rect 8112 52252 8176 52256
rect 8112 52196 8116 52252
rect 8116 52196 8172 52252
rect 8172 52196 8176 52252
rect 8112 52192 8176 52196
rect 8192 52252 8256 52256
rect 8192 52196 8196 52252
rect 8196 52196 8252 52252
rect 8252 52196 8256 52252
rect 8192 52192 8256 52196
rect 17952 52252 18016 52256
rect 17952 52196 17956 52252
rect 17956 52196 18012 52252
rect 18012 52196 18016 52252
rect 17952 52192 18016 52196
rect 18032 52252 18096 52256
rect 18032 52196 18036 52252
rect 18036 52196 18092 52252
rect 18092 52196 18096 52252
rect 18032 52192 18096 52196
rect 18112 52252 18176 52256
rect 18112 52196 18116 52252
rect 18116 52196 18172 52252
rect 18172 52196 18176 52252
rect 18112 52192 18176 52196
rect 18192 52252 18256 52256
rect 18192 52196 18196 52252
rect 18196 52196 18252 52252
rect 18252 52196 18256 52252
rect 18192 52192 18256 52196
rect 2952 51708 3016 51712
rect 2952 51652 2956 51708
rect 2956 51652 3012 51708
rect 3012 51652 3016 51708
rect 2952 51648 3016 51652
rect 3032 51708 3096 51712
rect 3032 51652 3036 51708
rect 3036 51652 3092 51708
rect 3092 51652 3096 51708
rect 3032 51648 3096 51652
rect 3112 51708 3176 51712
rect 3112 51652 3116 51708
rect 3116 51652 3172 51708
rect 3172 51652 3176 51708
rect 3112 51648 3176 51652
rect 3192 51708 3256 51712
rect 3192 51652 3196 51708
rect 3196 51652 3252 51708
rect 3252 51652 3256 51708
rect 3192 51648 3256 51652
rect 12952 51708 13016 51712
rect 12952 51652 12956 51708
rect 12956 51652 13012 51708
rect 13012 51652 13016 51708
rect 12952 51648 13016 51652
rect 13032 51708 13096 51712
rect 13032 51652 13036 51708
rect 13036 51652 13092 51708
rect 13092 51652 13096 51708
rect 13032 51648 13096 51652
rect 13112 51708 13176 51712
rect 13112 51652 13116 51708
rect 13116 51652 13172 51708
rect 13172 51652 13176 51708
rect 13112 51648 13176 51652
rect 13192 51708 13256 51712
rect 13192 51652 13196 51708
rect 13196 51652 13252 51708
rect 13252 51652 13256 51708
rect 13192 51648 13256 51652
rect 22952 51708 23016 51712
rect 22952 51652 22956 51708
rect 22956 51652 23012 51708
rect 23012 51652 23016 51708
rect 22952 51648 23016 51652
rect 23032 51708 23096 51712
rect 23032 51652 23036 51708
rect 23036 51652 23092 51708
rect 23092 51652 23096 51708
rect 23032 51648 23096 51652
rect 23112 51708 23176 51712
rect 23112 51652 23116 51708
rect 23116 51652 23172 51708
rect 23172 51652 23176 51708
rect 23112 51648 23176 51652
rect 23192 51708 23256 51712
rect 23192 51652 23196 51708
rect 23196 51652 23252 51708
rect 23252 51652 23256 51708
rect 23192 51648 23256 51652
rect 7952 51164 8016 51168
rect 7952 51108 7956 51164
rect 7956 51108 8012 51164
rect 8012 51108 8016 51164
rect 7952 51104 8016 51108
rect 8032 51164 8096 51168
rect 8032 51108 8036 51164
rect 8036 51108 8092 51164
rect 8092 51108 8096 51164
rect 8032 51104 8096 51108
rect 8112 51164 8176 51168
rect 8112 51108 8116 51164
rect 8116 51108 8172 51164
rect 8172 51108 8176 51164
rect 8112 51104 8176 51108
rect 8192 51164 8256 51168
rect 8192 51108 8196 51164
rect 8196 51108 8252 51164
rect 8252 51108 8256 51164
rect 8192 51104 8256 51108
rect 17952 51164 18016 51168
rect 17952 51108 17956 51164
rect 17956 51108 18012 51164
rect 18012 51108 18016 51164
rect 17952 51104 18016 51108
rect 18032 51164 18096 51168
rect 18032 51108 18036 51164
rect 18036 51108 18092 51164
rect 18092 51108 18096 51164
rect 18032 51104 18096 51108
rect 18112 51164 18176 51168
rect 18112 51108 18116 51164
rect 18116 51108 18172 51164
rect 18172 51108 18176 51164
rect 18112 51104 18176 51108
rect 18192 51164 18256 51168
rect 18192 51108 18196 51164
rect 18196 51108 18252 51164
rect 18252 51108 18256 51164
rect 18192 51104 18256 51108
rect 2952 50620 3016 50624
rect 2952 50564 2956 50620
rect 2956 50564 3012 50620
rect 3012 50564 3016 50620
rect 2952 50560 3016 50564
rect 3032 50620 3096 50624
rect 3032 50564 3036 50620
rect 3036 50564 3092 50620
rect 3092 50564 3096 50620
rect 3032 50560 3096 50564
rect 3112 50620 3176 50624
rect 3112 50564 3116 50620
rect 3116 50564 3172 50620
rect 3172 50564 3176 50620
rect 3112 50560 3176 50564
rect 3192 50620 3256 50624
rect 3192 50564 3196 50620
rect 3196 50564 3252 50620
rect 3252 50564 3256 50620
rect 3192 50560 3256 50564
rect 12952 50620 13016 50624
rect 12952 50564 12956 50620
rect 12956 50564 13012 50620
rect 13012 50564 13016 50620
rect 12952 50560 13016 50564
rect 13032 50620 13096 50624
rect 13032 50564 13036 50620
rect 13036 50564 13092 50620
rect 13092 50564 13096 50620
rect 13032 50560 13096 50564
rect 13112 50620 13176 50624
rect 13112 50564 13116 50620
rect 13116 50564 13172 50620
rect 13172 50564 13176 50620
rect 13112 50560 13176 50564
rect 13192 50620 13256 50624
rect 13192 50564 13196 50620
rect 13196 50564 13252 50620
rect 13252 50564 13256 50620
rect 13192 50560 13256 50564
rect 22952 50620 23016 50624
rect 22952 50564 22956 50620
rect 22956 50564 23012 50620
rect 23012 50564 23016 50620
rect 22952 50560 23016 50564
rect 23032 50620 23096 50624
rect 23032 50564 23036 50620
rect 23036 50564 23092 50620
rect 23092 50564 23096 50620
rect 23032 50560 23096 50564
rect 23112 50620 23176 50624
rect 23112 50564 23116 50620
rect 23116 50564 23172 50620
rect 23172 50564 23176 50620
rect 23112 50560 23176 50564
rect 23192 50620 23256 50624
rect 23192 50564 23196 50620
rect 23196 50564 23252 50620
rect 23252 50564 23256 50620
rect 23192 50560 23256 50564
rect 7952 50076 8016 50080
rect 7952 50020 7956 50076
rect 7956 50020 8012 50076
rect 8012 50020 8016 50076
rect 7952 50016 8016 50020
rect 8032 50076 8096 50080
rect 8032 50020 8036 50076
rect 8036 50020 8092 50076
rect 8092 50020 8096 50076
rect 8032 50016 8096 50020
rect 8112 50076 8176 50080
rect 8112 50020 8116 50076
rect 8116 50020 8172 50076
rect 8172 50020 8176 50076
rect 8112 50016 8176 50020
rect 8192 50076 8256 50080
rect 8192 50020 8196 50076
rect 8196 50020 8252 50076
rect 8252 50020 8256 50076
rect 8192 50016 8256 50020
rect 17952 50076 18016 50080
rect 17952 50020 17956 50076
rect 17956 50020 18012 50076
rect 18012 50020 18016 50076
rect 17952 50016 18016 50020
rect 18032 50076 18096 50080
rect 18032 50020 18036 50076
rect 18036 50020 18092 50076
rect 18092 50020 18096 50076
rect 18032 50016 18096 50020
rect 18112 50076 18176 50080
rect 18112 50020 18116 50076
rect 18116 50020 18172 50076
rect 18172 50020 18176 50076
rect 18112 50016 18176 50020
rect 18192 50076 18256 50080
rect 18192 50020 18196 50076
rect 18196 50020 18252 50076
rect 18252 50020 18256 50076
rect 18192 50016 18256 50020
rect 2952 49532 3016 49536
rect 2952 49476 2956 49532
rect 2956 49476 3012 49532
rect 3012 49476 3016 49532
rect 2952 49472 3016 49476
rect 3032 49532 3096 49536
rect 3032 49476 3036 49532
rect 3036 49476 3092 49532
rect 3092 49476 3096 49532
rect 3032 49472 3096 49476
rect 3112 49532 3176 49536
rect 3112 49476 3116 49532
rect 3116 49476 3172 49532
rect 3172 49476 3176 49532
rect 3112 49472 3176 49476
rect 3192 49532 3256 49536
rect 3192 49476 3196 49532
rect 3196 49476 3252 49532
rect 3252 49476 3256 49532
rect 3192 49472 3256 49476
rect 12952 49532 13016 49536
rect 12952 49476 12956 49532
rect 12956 49476 13012 49532
rect 13012 49476 13016 49532
rect 12952 49472 13016 49476
rect 13032 49532 13096 49536
rect 13032 49476 13036 49532
rect 13036 49476 13092 49532
rect 13092 49476 13096 49532
rect 13032 49472 13096 49476
rect 13112 49532 13176 49536
rect 13112 49476 13116 49532
rect 13116 49476 13172 49532
rect 13172 49476 13176 49532
rect 13112 49472 13176 49476
rect 13192 49532 13256 49536
rect 13192 49476 13196 49532
rect 13196 49476 13252 49532
rect 13252 49476 13256 49532
rect 13192 49472 13256 49476
rect 22952 49532 23016 49536
rect 22952 49476 22956 49532
rect 22956 49476 23012 49532
rect 23012 49476 23016 49532
rect 22952 49472 23016 49476
rect 23032 49532 23096 49536
rect 23032 49476 23036 49532
rect 23036 49476 23092 49532
rect 23092 49476 23096 49532
rect 23032 49472 23096 49476
rect 23112 49532 23176 49536
rect 23112 49476 23116 49532
rect 23116 49476 23172 49532
rect 23172 49476 23176 49532
rect 23112 49472 23176 49476
rect 23192 49532 23256 49536
rect 23192 49476 23196 49532
rect 23196 49476 23252 49532
rect 23252 49476 23256 49532
rect 23192 49472 23256 49476
rect 7952 48988 8016 48992
rect 7952 48932 7956 48988
rect 7956 48932 8012 48988
rect 8012 48932 8016 48988
rect 7952 48928 8016 48932
rect 8032 48988 8096 48992
rect 8032 48932 8036 48988
rect 8036 48932 8092 48988
rect 8092 48932 8096 48988
rect 8032 48928 8096 48932
rect 8112 48988 8176 48992
rect 8112 48932 8116 48988
rect 8116 48932 8172 48988
rect 8172 48932 8176 48988
rect 8112 48928 8176 48932
rect 8192 48988 8256 48992
rect 8192 48932 8196 48988
rect 8196 48932 8252 48988
rect 8252 48932 8256 48988
rect 8192 48928 8256 48932
rect 17952 48988 18016 48992
rect 17952 48932 17956 48988
rect 17956 48932 18012 48988
rect 18012 48932 18016 48988
rect 17952 48928 18016 48932
rect 18032 48988 18096 48992
rect 18032 48932 18036 48988
rect 18036 48932 18092 48988
rect 18092 48932 18096 48988
rect 18032 48928 18096 48932
rect 18112 48988 18176 48992
rect 18112 48932 18116 48988
rect 18116 48932 18172 48988
rect 18172 48932 18176 48988
rect 18112 48928 18176 48932
rect 18192 48988 18256 48992
rect 18192 48932 18196 48988
rect 18196 48932 18252 48988
rect 18252 48932 18256 48988
rect 18192 48928 18256 48932
rect 2952 48444 3016 48448
rect 2952 48388 2956 48444
rect 2956 48388 3012 48444
rect 3012 48388 3016 48444
rect 2952 48384 3016 48388
rect 3032 48444 3096 48448
rect 3032 48388 3036 48444
rect 3036 48388 3092 48444
rect 3092 48388 3096 48444
rect 3032 48384 3096 48388
rect 3112 48444 3176 48448
rect 3112 48388 3116 48444
rect 3116 48388 3172 48444
rect 3172 48388 3176 48444
rect 3112 48384 3176 48388
rect 3192 48444 3256 48448
rect 3192 48388 3196 48444
rect 3196 48388 3252 48444
rect 3252 48388 3256 48444
rect 3192 48384 3256 48388
rect 12952 48444 13016 48448
rect 12952 48388 12956 48444
rect 12956 48388 13012 48444
rect 13012 48388 13016 48444
rect 12952 48384 13016 48388
rect 13032 48444 13096 48448
rect 13032 48388 13036 48444
rect 13036 48388 13092 48444
rect 13092 48388 13096 48444
rect 13032 48384 13096 48388
rect 13112 48444 13176 48448
rect 13112 48388 13116 48444
rect 13116 48388 13172 48444
rect 13172 48388 13176 48444
rect 13112 48384 13176 48388
rect 13192 48444 13256 48448
rect 13192 48388 13196 48444
rect 13196 48388 13252 48444
rect 13252 48388 13256 48444
rect 13192 48384 13256 48388
rect 22952 48444 23016 48448
rect 22952 48388 22956 48444
rect 22956 48388 23012 48444
rect 23012 48388 23016 48444
rect 22952 48384 23016 48388
rect 23032 48444 23096 48448
rect 23032 48388 23036 48444
rect 23036 48388 23092 48444
rect 23092 48388 23096 48444
rect 23032 48384 23096 48388
rect 23112 48444 23176 48448
rect 23112 48388 23116 48444
rect 23116 48388 23172 48444
rect 23172 48388 23176 48444
rect 23112 48384 23176 48388
rect 23192 48444 23256 48448
rect 23192 48388 23196 48444
rect 23196 48388 23252 48444
rect 23252 48388 23256 48444
rect 23192 48384 23256 48388
rect 7952 47900 8016 47904
rect 7952 47844 7956 47900
rect 7956 47844 8012 47900
rect 8012 47844 8016 47900
rect 7952 47840 8016 47844
rect 8032 47900 8096 47904
rect 8032 47844 8036 47900
rect 8036 47844 8092 47900
rect 8092 47844 8096 47900
rect 8032 47840 8096 47844
rect 8112 47900 8176 47904
rect 8112 47844 8116 47900
rect 8116 47844 8172 47900
rect 8172 47844 8176 47900
rect 8112 47840 8176 47844
rect 8192 47900 8256 47904
rect 8192 47844 8196 47900
rect 8196 47844 8252 47900
rect 8252 47844 8256 47900
rect 8192 47840 8256 47844
rect 17952 47900 18016 47904
rect 17952 47844 17956 47900
rect 17956 47844 18012 47900
rect 18012 47844 18016 47900
rect 17952 47840 18016 47844
rect 18032 47900 18096 47904
rect 18032 47844 18036 47900
rect 18036 47844 18092 47900
rect 18092 47844 18096 47900
rect 18032 47840 18096 47844
rect 18112 47900 18176 47904
rect 18112 47844 18116 47900
rect 18116 47844 18172 47900
rect 18172 47844 18176 47900
rect 18112 47840 18176 47844
rect 18192 47900 18256 47904
rect 18192 47844 18196 47900
rect 18196 47844 18252 47900
rect 18252 47844 18256 47900
rect 18192 47840 18256 47844
rect 2952 47356 3016 47360
rect 2952 47300 2956 47356
rect 2956 47300 3012 47356
rect 3012 47300 3016 47356
rect 2952 47296 3016 47300
rect 3032 47356 3096 47360
rect 3032 47300 3036 47356
rect 3036 47300 3092 47356
rect 3092 47300 3096 47356
rect 3032 47296 3096 47300
rect 3112 47356 3176 47360
rect 3112 47300 3116 47356
rect 3116 47300 3172 47356
rect 3172 47300 3176 47356
rect 3112 47296 3176 47300
rect 3192 47356 3256 47360
rect 3192 47300 3196 47356
rect 3196 47300 3252 47356
rect 3252 47300 3256 47356
rect 3192 47296 3256 47300
rect 12952 47356 13016 47360
rect 12952 47300 12956 47356
rect 12956 47300 13012 47356
rect 13012 47300 13016 47356
rect 12952 47296 13016 47300
rect 13032 47356 13096 47360
rect 13032 47300 13036 47356
rect 13036 47300 13092 47356
rect 13092 47300 13096 47356
rect 13032 47296 13096 47300
rect 13112 47356 13176 47360
rect 13112 47300 13116 47356
rect 13116 47300 13172 47356
rect 13172 47300 13176 47356
rect 13112 47296 13176 47300
rect 13192 47356 13256 47360
rect 13192 47300 13196 47356
rect 13196 47300 13252 47356
rect 13252 47300 13256 47356
rect 13192 47296 13256 47300
rect 22952 47356 23016 47360
rect 22952 47300 22956 47356
rect 22956 47300 23012 47356
rect 23012 47300 23016 47356
rect 22952 47296 23016 47300
rect 23032 47356 23096 47360
rect 23032 47300 23036 47356
rect 23036 47300 23092 47356
rect 23092 47300 23096 47356
rect 23032 47296 23096 47300
rect 23112 47356 23176 47360
rect 23112 47300 23116 47356
rect 23116 47300 23172 47356
rect 23172 47300 23176 47356
rect 23112 47296 23176 47300
rect 23192 47356 23256 47360
rect 23192 47300 23196 47356
rect 23196 47300 23252 47356
rect 23252 47300 23256 47356
rect 23192 47296 23256 47300
rect 7952 46812 8016 46816
rect 7952 46756 7956 46812
rect 7956 46756 8012 46812
rect 8012 46756 8016 46812
rect 7952 46752 8016 46756
rect 8032 46812 8096 46816
rect 8032 46756 8036 46812
rect 8036 46756 8092 46812
rect 8092 46756 8096 46812
rect 8032 46752 8096 46756
rect 8112 46812 8176 46816
rect 8112 46756 8116 46812
rect 8116 46756 8172 46812
rect 8172 46756 8176 46812
rect 8112 46752 8176 46756
rect 8192 46812 8256 46816
rect 8192 46756 8196 46812
rect 8196 46756 8252 46812
rect 8252 46756 8256 46812
rect 8192 46752 8256 46756
rect 17952 46812 18016 46816
rect 17952 46756 17956 46812
rect 17956 46756 18012 46812
rect 18012 46756 18016 46812
rect 17952 46752 18016 46756
rect 18032 46812 18096 46816
rect 18032 46756 18036 46812
rect 18036 46756 18092 46812
rect 18092 46756 18096 46812
rect 18032 46752 18096 46756
rect 18112 46812 18176 46816
rect 18112 46756 18116 46812
rect 18116 46756 18172 46812
rect 18172 46756 18176 46812
rect 18112 46752 18176 46756
rect 18192 46812 18256 46816
rect 18192 46756 18196 46812
rect 18196 46756 18252 46812
rect 18252 46756 18256 46812
rect 18192 46752 18256 46756
rect 2952 46268 3016 46272
rect 2952 46212 2956 46268
rect 2956 46212 3012 46268
rect 3012 46212 3016 46268
rect 2952 46208 3016 46212
rect 3032 46268 3096 46272
rect 3032 46212 3036 46268
rect 3036 46212 3092 46268
rect 3092 46212 3096 46268
rect 3032 46208 3096 46212
rect 3112 46268 3176 46272
rect 3112 46212 3116 46268
rect 3116 46212 3172 46268
rect 3172 46212 3176 46268
rect 3112 46208 3176 46212
rect 3192 46268 3256 46272
rect 3192 46212 3196 46268
rect 3196 46212 3252 46268
rect 3252 46212 3256 46268
rect 3192 46208 3256 46212
rect 12952 46268 13016 46272
rect 12952 46212 12956 46268
rect 12956 46212 13012 46268
rect 13012 46212 13016 46268
rect 12952 46208 13016 46212
rect 13032 46268 13096 46272
rect 13032 46212 13036 46268
rect 13036 46212 13092 46268
rect 13092 46212 13096 46268
rect 13032 46208 13096 46212
rect 13112 46268 13176 46272
rect 13112 46212 13116 46268
rect 13116 46212 13172 46268
rect 13172 46212 13176 46268
rect 13112 46208 13176 46212
rect 13192 46268 13256 46272
rect 13192 46212 13196 46268
rect 13196 46212 13252 46268
rect 13252 46212 13256 46268
rect 13192 46208 13256 46212
rect 22952 46268 23016 46272
rect 22952 46212 22956 46268
rect 22956 46212 23012 46268
rect 23012 46212 23016 46268
rect 22952 46208 23016 46212
rect 23032 46268 23096 46272
rect 23032 46212 23036 46268
rect 23036 46212 23092 46268
rect 23092 46212 23096 46268
rect 23032 46208 23096 46212
rect 23112 46268 23176 46272
rect 23112 46212 23116 46268
rect 23116 46212 23172 46268
rect 23172 46212 23176 46268
rect 23112 46208 23176 46212
rect 23192 46268 23256 46272
rect 23192 46212 23196 46268
rect 23196 46212 23252 46268
rect 23252 46212 23256 46268
rect 23192 46208 23256 46212
rect 7952 45724 8016 45728
rect 7952 45668 7956 45724
rect 7956 45668 8012 45724
rect 8012 45668 8016 45724
rect 7952 45664 8016 45668
rect 8032 45724 8096 45728
rect 8032 45668 8036 45724
rect 8036 45668 8092 45724
rect 8092 45668 8096 45724
rect 8032 45664 8096 45668
rect 8112 45724 8176 45728
rect 8112 45668 8116 45724
rect 8116 45668 8172 45724
rect 8172 45668 8176 45724
rect 8112 45664 8176 45668
rect 8192 45724 8256 45728
rect 8192 45668 8196 45724
rect 8196 45668 8252 45724
rect 8252 45668 8256 45724
rect 8192 45664 8256 45668
rect 17952 45724 18016 45728
rect 17952 45668 17956 45724
rect 17956 45668 18012 45724
rect 18012 45668 18016 45724
rect 17952 45664 18016 45668
rect 18032 45724 18096 45728
rect 18032 45668 18036 45724
rect 18036 45668 18092 45724
rect 18092 45668 18096 45724
rect 18032 45664 18096 45668
rect 18112 45724 18176 45728
rect 18112 45668 18116 45724
rect 18116 45668 18172 45724
rect 18172 45668 18176 45724
rect 18112 45664 18176 45668
rect 18192 45724 18256 45728
rect 18192 45668 18196 45724
rect 18196 45668 18252 45724
rect 18252 45668 18256 45724
rect 18192 45664 18256 45668
rect 2952 45180 3016 45184
rect 2952 45124 2956 45180
rect 2956 45124 3012 45180
rect 3012 45124 3016 45180
rect 2952 45120 3016 45124
rect 3032 45180 3096 45184
rect 3032 45124 3036 45180
rect 3036 45124 3092 45180
rect 3092 45124 3096 45180
rect 3032 45120 3096 45124
rect 3112 45180 3176 45184
rect 3112 45124 3116 45180
rect 3116 45124 3172 45180
rect 3172 45124 3176 45180
rect 3112 45120 3176 45124
rect 3192 45180 3256 45184
rect 3192 45124 3196 45180
rect 3196 45124 3252 45180
rect 3252 45124 3256 45180
rect 3192 45120 3256 45124
rect 12952 45180 13016 45184
rect 12952 45124 12956 45180
rect 12956 45124 13012 45180
rect 13012 45124 13016 45180
rect 12952 45120 13016 45124
rect 13032 45180 13096 45184
rect 13032 45124 13036 45180
rect 13036 45124 13092 45180
rect 13092 45124 13096 45180
rect 13032 45120 13096 45124
rect 13112 45180 13176 45184
rect 13112 45124 13116 45180
rect 13116 45124 13172 45180
rect 13172 45124 13176 45180
rect 13112 45120 13176 45124
rect 13192 45180 13256 45184
rect 13192 45124 13196 45180
rect 13196 45124 13252 45180
rect 13252 45124 13256 45180
rect 13192 45120 13256 45124
rect 22952 45180 23016 45184
rect 22952 45124 22956 45180
rect 22956 45124 23012 45180
rect 23012 45124 23016 45180
rect 22952 45120 23016 45124
rect 23032 45180 23096 45184
rect 23032 45124 23036 45180
rect 23036 45124 23092 45180
rect 23092 45124 23096 45180
rect 23032 45120 23096 45124
rect 23112 45180 23176 45184
rect 23112 45124 23116 45180
rect 23116 45124 23172 45180
rect 23172 45124 23176 45180
rect 23112 45120 23176 45124
rect 23192 45180 23256 45184
rect 23192 45124 23196 45180
rect 23196 45124 23252 45180
rect 23252 45124 23256 45180
rect 23192 45120 23256 45124
rect 7952 44636 8016 44640
rect 7952 44580 7956 44636
rect 7956 44580 8012 44636
rect 8012 44580 8016 44636
rect 7952 44576 8016 44580
rect 8032 44636 8096 44640
rect 8032 44580 8036 44636
rect 8036 44580 8092 44636
rect 8092 44580 8096 44636
rect 8032 44576 8096 44580
rect 8112 44636 8176 44640
rect 8112 44580 8116 44636
rect 8116 44580 8172 44636
rect 8172 44580 8176 44636
rect 8112 44576 8176 44580
rect 8192 44636 8256 44640
rect 8192 44580 8196 44636
rect 8196 44580 8252 44636
rect 8252 44580 8256 44636
rect 8192 44576 8256 44580
rect 17952 44636 18016 44640
rect 17952 44580 17956 44636
rect 17956 44580 18012 44636
rect 18012 44580 18016 44636
rect 17952 44576 18016 44580
rect 18032 44636 18096 44640
rect 18032 44580 18036 44636
rect 18036 44580 18092 44636
rect 18092 44580 18096 44636
rect 18032 44576 18096 44580
rect 18112 44636 18176 44640
rect 18112 44580 18116 44636
rect 18116 44580 18172 44636
rect 18172 44580 18176 44636
rect 18112 44576 18176 44580
rect 18192 44636 18256 44640
rect 18192 44580 18196 44636
rect 18196 44580 18252 44636
rect 18252 44580 18256 44636
rect 18192 44576 18256 44580
rect 2952 44092 3016 44096
rect 2952 44036 2956 44092
rect 2956 44036 3012 44092
rect 3012 44036 3016 44092
rect 2952 44032 3016 44036
rect 3032 44092 3096 44096
rect 3032 44036 3036 44092
rect 3036 44036 3092 44092
rect 3092 44036 3096 44092
rect 3032 44032 3096 44036
rect 3112 44092 3176 44096
rect 3112 44036 3116 44092
rect 3116 44036 3172 44092
rect 3172 44036 3176 44092
rect 3112 44032 3176 44036
rect 3192 44092 3256 44096
rect 3192 44036 3196 44092
rect 3196 44036 3252 44092
rect 3252 44036 3256 44092
rect 3192 44032 3256 44036
rect 12952 44092 13016 44096
rect 12952 44036 12956 44092
rect 12956 44036 13012 44092
rect 13012 44036 13016 44092
rect 12952 44032 13016 44036
rect 13032 44092 13096 44096
rect 13032 44036 13036 44092
rect 13036 44036 13092 44092
rect 13092 44036 13096 44092
rect 13032 44032 13096 44036
rect 13112 44092 13176 44096
rect 13112 44036 13116 44092
rect 13116 44036 13172 44092
rect 13172 44036 13176 44092
rect 13112 44032 13176 44036
rect 13192 44092 13256 44096
rect 13192 44036 13196 44092
rect 13196 44036 13252 44092
rect 13252 44036 13256 44092
rect 13192 44032 13256 44036
rect 22952 44092 23016 44096
rect 22952 44036 22956 44092
rect 22956 44036 23012 44092
rect 23012 44036 23016 44092
rect 22952 44032 23016 44036
rect 23032 44092 23096 44096
rect 23032 44036 23036 44092
rect 23036 44036 23092 44092
rect 23092 44036 23096 44092
rect 23032 44032 23096 44036
rect 23112 44092 23176 44096
rect 23112 44036 23116 44092
rect 23116 44036 23172 44092
rect 23172 44036 23176 44092
rect 23112 44032 23176 44036
rect 23192 44092 23256 44096
rect 23192 44036 23196 44092
rect 23196 44036 23252 44092
rect 23252 44036 23256 44092
rect 23192 44032 23256 44036
rect 7952 43548 8016 43552
rect 7952 43492 7956 43548
rect 7956 43492 8012 43548
rect 8012 43492 8016 43548
rect 7952 43488 8016 43492
rect 8032 43548 8096 43552
rect 8032 43492 8036 43548
rect 8036 43492 8092 43548
rect 8092 43492 8096 43548
rect 8032 43488 8096 43492
rect 8112 43548 8176 43552
rect 8112 43492 8116 43548
rect 8116 43492 8172 43548
rect 8172 43492 8176 43548
rect 8112 43488 8176 43492
rect 8192 43548 8256 43552
rect 8192 43492 8196 43548
rect 8196 43492 8252 43548
rect 8252 43492 8256 43548
rect 8192 43488 8256 43492
rect 17952 43548 18016 43552
rect 17952 43492 17956 43548
rect 17956 43492 18012 43548
rect 18012 43492 18016 43548
rect 17952 43488 18016 43492
rect 18032 43548 18096 43552
rect 18032 43492 18036 43548
rect 18036 43492 18092 43548
rect 18092 43492 18096 43548
rect 18032 43488 18096 43492
rect 18112 43548 18176 43552
rect 18112 43492 18116 43548
rect 18116 43492 18172 43548
rect 18172 43492 18176 43548
rect 18112 43488 18176 43492
rect 18192 43548 18256 43552
rect 18192 43492 18196 43548
rect 18196 43492 18252 43548
rect 18252 43492 18256 43548
rect 18192 43488 18256 43492
rect 2952 43004 3016 43008
rect 2952 42948 2956 43004
rect 2956 42948 3012 43004
rect 3012 42948 3016 43004
rect 2952 42944 3016 42948
rect 3032 43004 3096 43008
rect 3032 42948 3036 43004
rect 3036 42948 3092 43004
rect 3092 42948 3096 43004
rect 3032 42944 3096 42948
rect 3112 43004 3176 43008
rect 3112 42948 3116 43004
rect 3116 42948 3172 43004
rect 3172 42948 3176 43004
rect 3112 42944 3176 42948
rect 3192 43004 3256 43008
rect 3192 42948 3196 43004
rect 3196 42948 3252 43004
rect 3252 42948 3256 43004
rect 3192 42944 3256 42948
rect 12952 43004 13016 43008
rect 12952 42948 12956 43004
rect 12956 42948 13012 43004
rect 13012 42948 13016 43004
rect 12952 42944 13016 42948
rect 13032 43004 13096 43008
rect 13032 42948 13036 43004
rect 13036 42948 13092 43004
rect 13092 42948 13096 43004
rect 13032 42944 13096 42948
rect 13112 43004 13176 43008
rect 13112 42948 13116 43004
rect 13116 42948 13172 43004
rect 13172 42948 13176 43004
rect 13112 42944 13176 42948
rect 13192 43004 13256 43008
rect 13192 42948 13196 43004
rect 13196 42948 13252 43004
rect 13252 42948 13256 43004
rect 13192 42944 13256 42948
rect 22952 43004 23016 43008
rect 22952 42948 22956 43004
rect 22956 42948 23012 43004
rect 23012 42948 23016 43004
rect 22952 42944 23016 42948
rect 23032 43004 23096 43008
rect 23032 42948 23036 43004
rect 23036 42948 23092 43004
rect 23092 42948 23096 43004
rect 23032 42944 23096 42948
rect 23112 43004 23176 43008
rect 23112 42948 23116 43004
rect 23116 42948 23172 43004
rect 23172 42948 23176 43004
rect 23112 42944 23176 42948
rect 23192 43004 23256 43008
rect 23192 42948 23196 43004
rect 23196 42948 23252 43004
rect 23252 42948 23256 43004
rect 23192 42944 23256 42948
rect 7952 42460 8016 42464
rect 7952 42404 7956 42460
rect 7956 42404 8012 42460
rect 8012 42404 8016 42460
rect 7952 42400 8016 42404
rect 8032 42460 8096 42464
rect 8032 42404 8036 42460
rect 8036 42404 8092 42460
rect 8092 42404 8096 42460
rect 8032 42400 8096 42404
rect 8112 42460 8176 42464
rect 8112 42404 8116 42460
rect 8116 42404 8172 42460
rect 8172 42404 8176 42460
rect 8112 42400 8176 42404
rect 8192 42460 8256 42464
rect 8192 42404 8196 42460
rect 8196 42404 8252 42460
rect 8252 42404 8256 42460
rect 8192 42400 8256 42404
rect 17952 42460 18016 42464
rect 17952 42404 17956 42460
rect 17956 42404 18012 42460
rect 18012 42404 18016 42460
rect 17952 42400 18016 42404
rect 18032 42460 18096 42464
rect 18032 42404 18036 42460
rect 18036 42404 18092 42460
rect 18092 42404 18096 42460
rect 18032 42400 18096 42404
rect 18112 42460 18176 42464
rect 18112 42404 18116 42460
rect 18116 42404 18172 42460
rect 18172 42404 18176 42460
rect 18112 42400 18176 42404
rect 18192 42460 18256 42464
rect 18192 42404 18196 42460
rect 18196 42404 18252 42460
rect 18252 42404 18256 42460
rect 18192 42400 18256 42404
rect 2952 41916 3016 41920
rect 2952 41860 2956 41916
rect 2956 41860 3012 41916
rect 3012 41860 3016 41916
rect 2952 41856 3016 41860
rect 3032 41916 3096 41920
rect 3032 41860 3036 41916
rect 3036 41860 3092 41916
rect 3092 41860 3096 41916
rect 3032 41856 3096 41860
rect 3112 41916 3176 41920
rect 3112 41860 3116 41916
rect 3116 41860 3172 41916
rect 3172 41860 3176 41916
rect 3112 41856 3176 41860
rect 3192 41916 3256 41920
rect 3192 41860 3196 41916
rect 3196 41860 3252 41916
rect 3252 41860 3256 41916
rect 3192 41856 3256 41860
rect 12952 41916 13016 41920
rect 12952 41860 12956 41916
rect 12956 41860 13012 41916
rect 13012 41860 13016 41916
rect 12952 41856 13016 41860
rect 13032 41916 13096 41920
rect 13032 41860 13036 41916
rect 13036 41860 13092 41916
rect 13092 41860 13096 41916
rect 13032 41856 13096 41860
rect 13112 41916 13176 41920
rect 13112 41860 13116 41916
rect 13116 41860 13172 41916
rect 13172 41860 13176 41916
rect 13112 41856 13176 41860
rect 13192 41916 13256 41920
rect 13192 41860 13196 41916
rect 13196 41860 13252 41916
rect 13252 41860 13256 41916
rect 13192 41856 13256 41860
rect 22952 41916 23016 41920
rect 22952 41860 22956 41916
rect 22956 41860 23012 41916
rect 23012 41860 23016 41916
rect 22952 41856 23016 41860
rect 23032 41916 23096 41920
rect 23032 41860 23036 41916
rect 23036 41860 23092 41916
rect 23092 41860 23096 41916
rect 23032 41856 23096 41860
rect 23112 41916 23176 41920
rect 23112 41860 23116 41916
rect 23116 41860 23172 41916
rect 23172 41860 23176 41916
rect 23112 41856 23176 41860
rect 23192 41916 23256 41920
rect 23192 41860 23196 41916
rect 23196 41860 23252 41916
rect 23252 41860 23256 41916
rect 23192 41856 23256 41860
rect 7952 41372 8016 41376
rect 7952 41316 7956 41372
rect 7956 41316 8012 41372
rect 8012 41316 8016 41372
rect 7952 41312 8016 41316
rect 8032 41372 8096 41376
rect 8032 41316 8036 41372
rect 8036 41316 8092 41372
rect 8092 41316 8096 41372
rect 8032 41312 8096 41316
rect 8112 41372 8176 41376
rect 8112 41316 8116 41372
rect 8116 41316 8172 41372
rect 8172 41316 8176 41372
rect 8112 41312 8176 41316
rect 8192 41372 8256 41376
rect 8192 41316 8196 41372
rect 8196 41316 8252 41372
rect 8252 41316 8256 41372
rect 8192 41312 8256 41316
rect 17952 41372 18016 41376
rect 17952 41316 17956 41372
rect 17956 41316 18012 41372
rect 18012 41316 18016 41372
rect 17952 41312 18016 41316
rect 18032 41372 18096 41376
rect 18032 41316 18036 41372
rect 18036 41316 18092 41372
rect 18092 41316 18096 41372
rect 18032 41312 18096 41316
rect 18112 41372 18176 41376
rect 18112 41316 18116 41372
rect 18116 41316 18172 41372
rect 18172 41316 18176 41372
rect 18112 41312 18176 41316
rect 18192 41372 18256 41376
rect 18192 41316 18196 41372
rect 18196 41316 18252 41372
rect 18252 41316 18256 41372
rect 18192 41312 18256 41316
rect 2952 40828 3016 40832
rect 2952 40772 2956 40828
rect 2956 40772 3012 40828
rect 3012 40772 3016 40828
rect 2952 40768 3016 40772
rect 3032 40828 3096 40832
rect 3032 40772 3036 40828
rect 3036 40772 3092 40828
rect 3092 40772 3096 40828
rect 3032 40768 3096 40772
rect 3112 40828 3176 40832
rect 3112 40772 3116 40828
rect 3116 40772 3172 40828
rect 3172 40772 3176 40828
rect 3112 40768 3176 40772
rect 3192 40828 3256 40832
rect 3192 40772 3196 40828
rect 3196 40772 3252 40828
rect 3252 40772 3256 40828
rect 3192 40768 3256 40772
rect 12952 40828 13016 40832
rect 12952 40772 12956 40828
rect 12956 40772 13012 40828
rect 13012 40772 13016 40828
rect 12952 40768 13016 40772
rect 13032 40828 13096 40832
rect 13032 40772 13036 40828
rect 13036 40772 13092 40828
rect 13092 40772 13096 40828
rect 13032 40768 13096 40772
rect 13112 40828 13176 40832
rect 13112 40772 13116 40828
rect 13116 40772 13172 40828
rect 13172 40772 13176 40828
rect 13112 40768 13176 40772
rect 13192 40828 13256 40832
rect 13192 40772 13196 40828
rect 13196 40772 13252 40828
rect 13252 40772 13256 40828
rect 13192 40768 13256 40772
rect 22952 40828 23016 40832
rect 22952 40772 22956 40828
rect 22956 40772 23012 40828
rect 23012 40772 23016 40828
rect 22952 40768 23016 40772
rect 23032 40828 23096 40832
rect 23032 40772 23036 40828
rect 23036 40772 23092 40828
rect 23092 40772 23096 40828
rect 23032 40768 23096 40772
rect 23112 40828 23176 40832
rect 23112 40772 23116 40828
rect 23116 40772 23172 40828
rect 23172 40772 23176 40828
rect 23112 40768 23176 40772
rect 23192 40828 23256 40832
rect 23192 40772 23196 40828
rect 23196 40772 23252 40828
rect 23252 40772 23256 40828
rect 23192 40768 23256 40772
rect 7952 40284 8016 40288
rect 7952 40228 7956 40284
rect 7956 40228 8012 40284
rect 8012 40228 8016 40284
rect 7952 40224 8016 40228
rect 8032 40284 8096 40288
rect 8032 40228 8036 40284
rect 8036 40228 8092 40284
rect 8092 40228 8096 40284
rect 8032 40224 8096 40228
rect 8112 40284 8176 40288
rect 8112 40228 8116 40284
rect 8116 40228 8172 40284
rect 8172 40228 8176 40284
rect 8112 40224 8176 40228
rect 8192 40284 8256 40288
rect 8192 40228 8196 40284
rect 8196 40228 8252 40284
rect 8252 40228 8256 40284
rect 8192 40224 8256 40228
rect 17952 40284 18016 40288
rect 17952 40228 17956 40284
rect 17956 40228 18012 40284
rect 18012 40228 18016 40284
rect 17952 40224 18016 40228
rect 18032 40284 18096 40288
rect 18032 40228 18036 40284
rect 18036 40228 18092 40284
rect 18092 40228 18096 40284
rect 18032 40224 18096 40228
rect 18112 40284 18176 40288
rect 18112 40228 18116 40284
rect 18116 40228 18172 40284
rect 18172 40228 18176 40284
rect 18112 40224 18176 40228
rect 18192 40284 18256 40288
rect 18192 40228 18196 40284
rect 18196 40228 18252 40284
rect 18252 40228 18256 40284
rect 18192 40224 18256 40228
rect 2952 39740 3016 39744
rect 2952 39684 2956 39740
rect 2956 39684 3012 39740
rect 3012 39684 3016 39740
rect 2952 39680 3016 39684
rect 3032 39740 3096 39744
rect 3032 39684 3036 39740
rect 3036 39684 3092 39740
rect 3092 39684 3096 39740
rect 3032 39680 3096 39684
rect 3112 39740 3176 39744
rect 3112 39684 3116 39740
rect 3116 39684 3172 39740
rect 3172 39684 3176 39740
rect 3112 39680 3176 39684
rect 3192 39740 3256 39744
rect 3192 39684 3196 39740
rect 3196 39684 3252 39740
rect 3252 39684 3256 39740
rect 3192 39680 3256 39684
rect 12952 39740 13016 39744
rect 12952 39684 12956 39740
rect 12956 39684 13012 39740
rect 13012 39684 13016 39740
rect 12952 39680 13016 39684
rect 13032 39740 13096 39744
rect 13032 39684 13036 39740
rect 13036 39684 13092 39740
rect 13092 39684 13096 39740
rect 13032 39680 13096 39684
rect 13112 39740 13176 39744
rect 13112 39684 13116 39740
rect 13116 39684 13172 39740
rect 13172 39684 13176 39740
rect 13112 39680 13176 39684
rect 13192 39740 13256 39744
rect 13192 39684 13196 39740
rect 13196 39684 13252 39740
rect 13252 39684 13256 39740
rect 13192 39680 13256 39684
rect 22952 39740 23016 39744
rect 22952 39684 22956 39740
rect 22956 39684 23012 39740
rect 23012 39684 23016 39740
rect 22952 39680 23016 39684
rect 23032 39740 23096 39744
rect 23032 39684 23036 39740
rect 23036 39684 23092 39740
rect 23092 39684 23096 39740
rect 23032 39680 23096 39684
rect 23112 39740 23176 39744
rect 23112 39684 23116 39740
rect 23116 39684 23172 39740
rect 23172 39684 23176 39740
rect 23112 39680 23176 39684
rect 23192 39740 23256 39744
rect 23192 39684 23196 39740
rect 23196 39684 23252 39740
rect 23252 39684 23256 39740
rect 23192 39680 23256 39684
rect 7952 39196 8016 39200
rect 7952 39140 7956 39196
rect 7956 39140 8012 39196
rect 8012 39140 8016 39196
rect 7952 39136 8016 39140
rect 8032 39196 8096 39200
rect 8032 39140 8036 39196
rect 8036 39140 8092 39196
rect 8092 39140 8096 39196
rect 8032 39136 8096 39140
rect 8112 39196 8176 39200
rect 8112 39140 8116 39196
rect 8116 39140 8172 39196
rect 8172 39140 8176 39196
rect 8112 39136 8176 39140
rect 8192 39196 8256 39200
rect 8192 39140 8196 39196
rect 8196 39140 8252 39196
rect 8252 39140 8256 39196
rect 8192 39136 8256 39140
rect 17952 39196 18016 39200
rect 17952 39140 17956 39196
rect 17956 39140 18012 39196
rect 18012 39140 18016 39196
rect 17952 39136 18016 39140
rect 18032 39196 18096 39200
rect 18032 39140 18036 39196
rect 18036 39140 18092 39196
rect 18092 39140 18096 39196
rect 18032 39136 18096 39140
rect 18112 39196 18176 39200
rect 18112 39140 18116 39196
rect 18116 39140 18172 39196
rect 18172 39140 18176 39196
rect 18112 39136 18176 39140
rect 18192 39196 18256 39200
rect 18192 39140 18196 39196
rect 18196 39140 18252 39196
rect 18252 39140 18256 39196
rect 18192 39136 18256 39140
rect 2952 38652 3016 38656
rect 2952 38596 2956 38652
rect 2956 38596 3012 38652
rect 3012 38596 3016 38652
rect 2952 38592 3016 38596
rect 3032 38652 3096 38656
rect 3032 38596 3036 38652
rect 3036 38596 3092 38652
rect 3092 38596 3096 38652
rect 3032 38592 3096 38596
rect 3112 38652 3176 38656
rect 3112 38596 3116 38652
rect 3116 38596 3172 38652
rect 3172 38596 3176 38652
rect 3112 38592 3176 38596
rect 3192 38652 3256 38656
rect 3192 38596 3196 38652
rect 3196 38596 3252 38652
rect 3252 38596 3256 38652
rect 3192 38592 3256 38596
rect 12952 38652 13016 38656
rect 12952 38596 12956 38652
rect 12956 38596 13012 38652
rect 13012 38596 13016 38652
rect 12952 38592 13016 38596
rect 13032 38652 13096 38656
rect 13032 38596 13036 38652
rect 13036 38596 13092 38652
rect 13092 38596 13096 38652
rect 13032 38592 13096 38596
rect 13112 38652 13176 38656
rect 13112 38596 13116 38652
rect 13116 38596 13172 38652
rect 13172 38596 13176 38652
rect 13112 38592 13176 38596
rect 13192 38652 13256 38656
rect 13192 38596 13196 38652
rect 13196 38596 13252 38652
rect 13252 38596 13256 38652
rect 13192 38592 13256 38596
rect 22952 38652 23016 38656
rect 22952 38596 22956 38652
rect 22956 38596 23012 38652
rect 23012 38596 23016 38652
rect 22952 38592 23016 38596
rect 23032 38652 23096 38656
rect 23032 38596 23036 38652
rect 23036 38596 23092 38652
rect 23092 38596 23096 38652
rect 23032 38592 23096 38596
rect 23112 38652 23176 38656
rect 23112 38596 23116 38652
rect 23116 38596 23172 38652
rect 23172 38596 23176 38652
rect 23112 38592 23176 38596
rect 23192 38652 23256 38656
rect 23192 38596 23196 38652
rect 23196 38596 23252 38652
rect 23252 38596 23256 38652
rect 23192 38592 23256 38596
rect 7952 38108 8016 38112
rect 7952 38052 7956 38108
rect 7956 38052 8012 38108
rect 8012 38052 8016 38108
rect 7952 38048 8016 38052
rect 8032 38108 8096 38112
rect 8032 38052 8036 38108
rect 8036 38052 8092 38108
rect 8092 38052 8096 38108
rect 8032 38048 8096 38052
rect 8112 38108 8176 38112
rect 8112 38052 8116 38108
rect 8116 38052 8172 38108
rect 8172 38052 8176 38108
rect 8112 38048 8176 38052
rect 8192 38108 8256 38112
rect 8192 38052 8196 38108
rect 8196 38052 8252 38108
rect 8252 38052 8256 38108
rect 8192 38048 8256 38052
rect 17952 38108 18016 38112
rect 17952 38052 17956 38108
rect 17956 38052 18012 38108
rect 18012 38052 18016 38108
rect 17952 38048 18016 38052
rect 18032 38108 18096 38112
rect 18032 38052 18036 38108
rect 18036 38052 18092 38108
rect 18092 38052 18096 38108
rect 18032 38048 18096 38052
rect 18112 38108 18176 38112
rect 18112 38052 18116 38108
rect 18116 38052 18172 38108
rect 18172 38052 18176 38108
rect 18112 38048 18176 38052
rect 18192 38108 18256 38112
rect 18192 38052 18196 38108
rect 18196 38052 18252 38108
rect 18252 38052 18256 38108
rect 18192 38048 18256 38052
rect 2952 37564 3016 37568
rect 2952 37508 2956 37564
rect 2956 37508 3012 37564
rect 3012 37508 3016 37564
rect 2952 37504 3016 37508
rect 3032 37564 3096 37568
rect 3032 37508 3036 37564
rect 3036 37508 3092 37564
rect 3092 37508 3096 37564
rect 3032 37504 3096 37508
rect 3112 37564 3176 37568
rect 3112 37508 3116 37564
rect 3116 37508 3172 37564
rect 3172 37508 3176 37564
rect 3112 37504 3176 37508
rect 3192 37564 3256 37568
rect 3192 37508 3196 37564
rect 3196 37508 3252 37564
rect 3252 37508 3256 37564
rect 3192 37504 3256 37508
rect 12952 37564 13016 37568
rect 12952 37508 12956 37564
rect 12956 37508 13012 37564
rect 13012 37508 13016 37564
rect 12952 37504 13016 37508
rect 13032 37564 13096 37568
rect 13032 37508 13036 37564
rect 13036 37508 13092 37564
rect 13092 37508 13096 37564
rect 13032 37504 13096 37508
rect 13112 37564 13176 37568
rect 13112 37508 13116 37564
rect 13116 37508 13172 37564
rect 13172 37508 13176 37564
rect 13112 37504 13176 37508
rect 13192 37564 13256 37568
rect 13192 37508 13196 37564
rect 13196 37508 13252 37564
rect 13252 37508 13256 37564
rect 13192 37504 13256 37508
rect 22952 37564 23016 37568
rect 22952 37508 22956 37564
rect 22956 37508 23012 37564
rect 23012 37508 23016 37564
rect 22952 37504 23016 37508
rect 23032 37564 23096 37568
rect 23032 37508 23036 37564
rect 23036 37508 23092 37564
rect 23092 37508 23096 37564
rect 23032 37504 23096 37508
rect 23112 37564 23176 37568
rect 23112 37508 23116 37564
rect 23116 37508 23172 37564
rect 23172 37508 23176 37564
rect 23112 37504 23176 37508
rect 23192 37564 23256 37568
rect 23192 37508 23196 37564
rect 23196 37508 23252 37564
rect 23252 37508 23256 37564
rect 23192 37504 23256 37508
rect 7952 37020 8016 37024
rect 7952 36964 7956 37020
rect 7956 36964 8012 37020
rect 8012 36964 8016 37020
rect 7952 36960 8016 36964
rect 8032 37020 8096 37024
rect 8032 36964 8036 37020
rect 8036 36964 8092 37020
rect 8092 36964 8096 37020
rect 8032 36960 8096 36964
rect 8112 37020 8176 37024
rect 8112 36964 8116 37020
rect 8116 36964 8172 37020
rect 8172 36964 8176 37020
rect 8112 36960 8176 36964
rect 8192 37020 8256 37024
rect 8192 36964 8196 37020
rect 8196 36964 8252 37020
rect 8252 36964 8256 37020
rect 8192 36960 8256 36964
rect 17952 37020 18016 37024
rect 17952 36964 17956 37020
rect 17956 36964 18012 37020
rect 18012 36964 18016 37020
rect 17952 36960 18016 36964
rect 18032 37020 18096 37024
rect 18032 36964 18036 37020
rect 18036 36964 18092 37020
rect 18092 36964 18096 37020
rect 18032 36960 18096 36964
rect 18112 37020 18176 37024
rect 18112 36964 18116 37020
rect 18116 36964 18172 37020
rect 18172 36964 18176 37020
rect 18112 36960 18176 36964
rect 18192 37020 18256 37024
rect 18192 36964 18196 37020
rect 18196 36964 18252 37020
rect 18252 36964 18256 37020
rect 18192 36960 18256 36964
rect 2952 36476 3016 36480
rect 2952 36420 2956 36476
rect 2956 36420 3012 36476
rect 3012 36420 3016 36476
rect 2952 36416 3016 36420
rect 3032 36476 3096 36480
rect 3032 36420 3036 36476
rect 3036 36420 3092 36476
rect 3092 36420 3096 36476
rect 3032 36416 3096 36420
rect 3112 36476 3176 36480
rect 3112 36420 3116 36476
rect 3116 36420 3172 36476
rect 3172 36420 3176 36476
rect 3112 36416 3176 36420
rect 3192 36476 3256 36480
rect 3192 36420 3196 36476
rect 3196 36420 3252 36476
rect 3252 36420 3256 36476
rect 3192 36416 3256 36420
rect 12952 36476 13016 36480
rect 12952 36420 12956 36476
rect 12956 36420 13012 36476
rect 13012 36420 13016 36476
rect 12952 36416 13016 36420
rect 13032 36476 13096 36480
rect 13032 36420 13036 36476
rect 13036 36420 13092 36476
rect 13092 36420 13096 36476
rect 13032 36416 13096 36420
rect 13112 36476 13176 36480
rect 13112 36420 13116 36476
rect 13116 36420 13172 36476
rect 13172 36420 13176 36476
rect 13112 36416 13176 36420
rect 13192 36476 13256 36480
rect 13192 36420 13196 36476
rect 13196 36420 13252 36476
rect 13252 36420 13256 36476
rect 13192 36416 13256 36420
rect 22952 36476 23016 36480
rect 22952 36420 22956 36476
rect 22956 36420 23012 36476
rect 23012 36420 23016 36476
rect 22952 36416 23016 36420
rect 23032 36476 23096 36480
rect 23032 36420 23036 36476
rect 23036 36420 23092 36476
rect 23092 36420 23096 36476
rect 23032 36416 23096 36420
rect 23112 36476 23176 36480
rect 23112 36420 23116 36476
rect 23116 36420 23172 36476
rect 23172 36420 23176 36476
rect 23112 36416 23176 36420
rect 23192 36476 23256 36480
rect 23192 36420 23196 36476
rect 23196 36420 23252 36476
rect 23252 36420 23256 36476
rect 23192 36416 23256 36420
rect 7952 35932 8016 35936
rect 7952 35876 7956 35932
rect 7956 35876 8012 35932
rect 8012 35876 8016 35932
rect 7952 35872 8016 35876
rect 8032 35932 8096 35936
rect 8032 35876 8036 35932
rect 8036 35876 8092 35932
rect 8092 35876 8096 35932
rect 8032 35872 8096 35876
rect 8112 35932 8176 35936
rect 8112 35876 8116 35932
rect 8116 35876 8172 35932
rect 8172 35876 8176 35932
rect 8112 35872 8176 35876
rect 8192 35932 8256 35936
rect 8192 35876 8196 35932
rect 8196 35876 8252 35932
rect 8252 35876 8256 35932
rect 8192 35872 8256 35876
rect 17952 35932 18016 35936
rect 17952 35876 17956 35932
rect 17956 35876 18012 35932
rect 18012 35876 18016 35932
rect 17952 35872 18016 35876
rect 18032 35932 18096 35936
rect 18032 35876 18036 35932
rect 18036 35876 18092 35932
rect 18092 35876 18096 35932
rect 18032 35872 18096 35876
rect 18112 35932 18176 35936
rect 18112 35876 18116 35932
rect 18116 35876 18172 35932
rect 18172 35876 18176 35932
rect 18112 35872 18176 35876
rect 18192 35932 18256 35936
rect 18192 35876 18196 35932
rect 18196 35876 18252 35932
rect 18252 35876 18256 35932
rect 18192 35872 18256 35876
rect 2952 35388 3016 35392
rect 2952 35332 2956 35388
rect 2956 35332 3012 35388
rect 3012 35332 3016 35388
rect 2952 35328 3016 35332
rect 3032 35388 3096 35392
rect 3032 35332 3036 35388
rect 3036 35332 3092 35388
rect 3092 35332 3096 35388
rect 3032 35328 3096 35332
rect 3112 35388 3176 35392
rect 3112 35332 3116 35388
rect 3116 35332 3172 35388
rect 3172 35332 3176 35388
rect 3112 35328 3176 35332
rect 3192 35388 3256 35392
rect 3192 35332 3196 35388
rect 3196 35332 3252 35388
rect 3252 35332 3256 35388
rect 3192 35328 3256 35332
rect 12952 35388 13016 35392
rect 12952 35332 12956 35388
rect 12956 35332 13012 35388
rect 13012 35332 13016 35388
rect 12952 35328 13016 35332
rect 13032 35388 13096 35392
rect 13032 35332 13036 35388
rect 13036 35332 13092 35388
rect 13092 35332 13096 35388
rect 13032 35328 13096 35332
rect 13112 35388 13176 35392
rect 13112 35332 13116 35388
rect 13116 35332 13172 35388
rect 13172 35332 13176 35388
rect 13112 35328 13176 35332
rect 13192 35388 13256 35392
rect 13192 35332 13196 35388
rect 13196 35332 13252 35388
rect 13252 35332 13256 35388
rect 13192 35328 13256 35332
rect 22952 35388 23016 35392
rect 22952 35332 22956 35388
rect 22956 35332 23012 35388
rect 23012 35332 23016 35388
rect 22952 35328 23016 35332
rect 23032 35388 23096 35392
rect 23032 35332 23036 35388
rect 23036 35332 23092 35388
rect 23092 35332 23096 35388
rect 23032 35328 23096 35332
rect 23112 35388 23176 35392
rect 23112 35332 23116 35388
rect 23116 35332 23172 35388
rect 23172 35332 23176 35388
rect 23112 35328 23176 35332
rect 23192 35388 23256 35392
rect 23192 35332 23196 35388
rect 23196 35332 23252 35388
rect 23252 35332 23256 35388
rect 23192 35328 23256 35332
rect 7952 34844 8016 34848
rect 7952 34788 7956 34844
rect 7956 34788 8012 34844
rect 8012 34788 8016 34844
rect 7952 34784 8016 34788
rect 8032 34844 8096 34848
rect 8032 34788 8036 34844
rect 8036 34788 8092 34844
rect 8092 34788 8096 34844
rect 8032 34784 8096 34788
rect 8112 34844 8176 34848
rect 8112 34788 8116 34844
rect 8116 34788 8172 34844
rect 8172 34788 8176 34844
rect 8112 34784 8176 34788
rect 8192 34844 8256 34848
rect 8192 34788 8196 34844
rect 8196 34788 8252 34844
rect 8252 34788 8256 34844
rect 8192 34784 8256 34788
rect 17952 34844 18016 34848
rect 17952 34788 17956 34844
rect 17956 34788 18012 34844
rect 18012 34788 18016 34844
rect 17952 34784 18016 34788
rect 18032 34844 18096 34848
rect 18032 34788 18036 34844
rect 18036 34788 18092 34844
rect 18092 34788 18096 34844
rect 18032 34784 18096 34788
rect 18112 34844 18176 34848
rect 18112 34788 18116 34844
rect 18116 34788 18172 34844
rect 18172 34788 18176 34844
rect 18112 34784 18176 34788
rect 18192 34844 18256 34848
rect 18192 34788 18196 34844
rect 18196 34788 18252 34844
rect 18252 34788 18256 34844
rect 18192 34784 18256 34788
rect 2952 34300 3016 34304
rect 2952 34244 2956 34300
rect 2956 34244 3012 34300
rect 3012 34244 3016 34300
rect 2952 34240 3016 34244
rect 3032 34300 3096 34304
rect 3032 34244 3036 34300
rect 3036 34244 3092 34300
rect 3092 34244 3096 34300
rect 3032 34240 3096 34244
rect 3112 34300 3176 34304
rect 3112 34244 3116 34300
rect 3116 34244 3172 34300
rect 3172 34244 3176 34300
rect 3112 34240 3176 34244
rect 3192 34300 3256 34304
rect 3192 34244 3196 34300
rect 3196 34244 3252 34300
rect 3252 34244 3256 34300
rect 3192 34240 3256 34244
rect 12952 34300 13016 34304
rect 12952 34244 12956 34300
rect 12956 34244 13012 34300
rect 13012 34244 13016 34300
rect 12952 34240 13016 34244
rect 13032 34300 13096 34304
rect 13032 34244 13036 34300
rect 13036 34244 13092 34300
rect 13092 34244 13096 34300
rect 13032 34240 13096 34244
rect 13112 34300 13176 34304
rect 13112 34244 13116 34300
rect 13116 34244 13172 34300
rect 13172 34244 13176 34300
rect 13112 34240 13176 34244
rect 13192 34300 13256 34304
rect 13192 34244 13196 34300
rect 13196 34244 13252 34300
rect 13252 34244 13256 34300
rect 13192 34240 13256 34244
rect 22952 34300 23016 34304
rect 22952 34244 22956 34300
rect 22956 34244 23012 34300
rect 23012 34244 23016 34300
rect 22952 34240 23016 34244
rect 23032 34300 23096 34304
rect 23032 34244 23036 34300
rect 23036 34244 23092 34300
rect 23092 34244 23096 34300
rect 23032 34240 23096 34244
rect 23112 34300 23176 34304
rect 23112 34244 23116 34300
rect 23116 34244 23172 34300
rect 23172 34244 23176 34300
rect 23112 34240 23176 34244
rect 23192 34300 23256 34304
rect 23192 34244 23196 34300
rect 23196 34244 23252 34300
rect 23252 34244 23256 34300
rect 23192 34240 23256 34244
rect 7952 33756 8016 33760
rect 7952 33700 7956 33756
rect 7956 33700 8012 33756
rect 8012 33700 8016 33756
rect 7952 33696 8016 33700
rect 8032 33756 8096 33760
rect 8032 33700 8036 33756
rect 8036 33700 8092 33756
rect 8092 33700 8096 33756
rect 8032 33696 8096 33700
rect 8112 33756 8176 33760
rect 8112 33700 8116 33756
rect 8116 33700 8172 33756
rect 8172 33700 8176 33756
rect 8112 33696 8176 33700
rect 8192 33756 8256 33760
rect 8192 33700 8196 33756
rect 8196 33700 8252 33756
rect 8252 33700 8256 33756
rect 8192 33696 8256 33700
rect 17952 33756 18016 33760
rect 17952 33700 17956 33756
rect 17956 33700 18012 33756
rect 18012 33700 18016 33756
rect 17952 33696 18016 33700
rect 18032 33756 18096 33760
rect 18032 33700 18036 33756
rect 18036 33700 18092 33756
rect 18092 33700 18096 33756
rect 18032 33696 18096 33700
rect 18112 33756 18176 33760
rect 18112 33700 18116 33756
rect 18116 33700 18172 33756
rect 18172 33700 18176 33756
rect 18112 33696 18176 33700
rect 18192 33756 18256 33760
rect 18192 33700 18196 33756
rect 18196 33700 18252 33756
rect 18252 33700 18256 33756
rect 18192 33696 18256 33700
rect 2952 33212 3016 33216
rect 2952 33156 2956 33212
rect 2956 33156 3012 33212
rect 3012 33156 3016 33212
rect 2952 33152 3016 33156
rect 3032 33212 3096 33216
rect 3032 33156 3036 33212
rect 3036 33156 3092 33212
rect 3092 33156 3096 33212
rect 3032 33152 3096 33156
rect 3112 33212 3176 33216
rect 3112 33156 3116 33212
rect 3116 33156 3172 33212
rect 3172 33156 3176 33212
rect 3112 33152 3176 33156
rect 3192 33212 3256 33216
rect 3192 33156 3196 33212
rect 3196 33156 3252 33212
rect 3252 33156 3256 33212
rect 3192 33152 3256 33156
rect 12952 33212 13016 33216
rect 12952 33156 12956 33212
rect 12956 33156 13012 33212
rect 13012 33156 13016 33212
rect 12952 33152 13016 33156
rect 13032 33212 13096 33216
rect 13032 33156 13036 33212
rect 13036 33156 13092 33212
rect 13092 33156 13096 33212
rect 13032 33152 13096 33156
rect 13112 33212 13176 33216
rect 13112 33156 13116 33212
rect 13116 33156 13172 33212
rect 13172 33156 13176 33212
rect 13112 33152 13176 33156
rect 13192 33212 13256 33216
rect 13192 33156 13196 33212
rect 13196 33156 13252 33212
rect 13252 33156 13256 33212
rect 13192 33152 13256 33156
rect 22952 33212 23016 33216
rect 22952 33156 22956 33212
rect 22956 33156 23012 33212
rect 23012 33156 23016 33212
rect 22952 33152 23016 33156
rect 23032 33212 23096 33216
rect 23032 33156 23036 33212
rect 23036 33156 23092 33212
rect 23092 33156 23096 33212
rect 23032 33152 23096 33156
rect 23112 33212 23176 33216
rect 23112 33156 23116 33212
rect 23116 33156 23172 33212
rect 23172 33156 23176 33212
rect 23112 33152 23176 33156
rect 23192 33212 23256 33216
rect 23192 33156 23196 33212
rect 23196 33156 23252 33212
rect 23252 33156 23256 33212
rect 23192 33152 23256 33156
rect 7952 32668 8016 32672
rect 7952 32612 7956 32668
rect 7956 32612 8012 32668
rect 8012 32612 8016 32668
rect 7952 32608 8016 32612
rect 8032 32668 8096 32672
rect 8032 32612 8036 32668
rect 8036 32612 8092 32668
rect 8092 32612 8096 32668
rect 8032 32608 8096 32612
rect 8112 32668 8176 32672
rect 8112 32612 8116 32668
rect 8116 32612 8172 32668
rect 8172 32612 8176 32668
rect 8112 32608 8176 32612
rect 8192 32668 8256 32672
rect 8192 32612 8196 32668
rect 8196 32612 8252 32668
rect 8252 32612 8256 32668
rect 8192 32608 8256 32612
rect 17952 32668 18016 32672
rect 17952 32612 17956 32668
rect 17956 32612 18012 32668
rect 18012 32612 18016 32668
rect 17952 32608 18016 32612
rect 18032 32668 18096 32672
rect 18032 32612 18036 32668
rect 18036 32612 18092 32668
rect 18092 32612 18096 32668
rect 18032 32608 18096 32612
rect 18112 32668 18176 32672
rect 18112 32612 18116 32668
rect 18116 32612 18172 32668
rect 18172 32612 18176 32668
rect 18112 32608 18176 32612
rect 18192 32668 18256 32672
rect 18192 32612 18196 32668
rect 18196 32612 18252 32668
rect 18252 32612 18256 32668
rect 18192 32608 18256 32612
rect 2952 32124 3016 32128
rect 2952 32068 2956 32124
rect 2956 32068 3012 32124
rect 3012 32068 3016 32124
rect 2952 32064 3016 32068
rect 3032 32124 3096 32128
rect 3032 32068 3036 32124
rect 3036 32068 3092 32124
rect 3092 32068 3096 32124
rect 3032 32064 3096 32068
rect 3112 32124 3176 32128
rect 3112 32068 3116 32124
rect 3116 32068 3172 32124
rect 3172 32068 3176 32124
rect 3112 32064 3176 32068
rect 3192 32124 3256 32128
rect 3192 32068 3196 32124
rect 3196 32068 3252 32124
rect 3252 32068 3256 32124
rect 3192 32064 3256 32068
rect 12952 32124 13016 32128
rect 12952 32068 12956 32124
rect 12956 32068 13012 32124
rect 13012 32068 13016 32124
rect 12952 32064 13016 32068
rect 13032 32124 13096 32128
rect 13032 32068 13036 32124
rect 13036 32068 13092 32124
rect 13092 32068 13096 32124
rect 13032 32064 13096 32068
rect 13112 32124 13176 32128
rect 13112 32068 13116 32124
rect 13116 32068 13172 32124
rect 13172 32068 13176 32124
rect 13112 32064 13176 32068
rect 13192 32124 13256 32128
rect 13192 32068 13196 32124
rect 13196 32068 13252 32124
rect 13252 32068 13256 32124
rect 13192 32064 13256 32068
rect 22952 32124 23016 32128
rect 22952 32068 22956 32124
rect 22956 32068 23012 32124
rect 23012 32068 23016 32124
rect 22952 32064 23016 32068
rect 23032 32124 23096 32128
rect 23032 32068 23036 32124
rect 23036 32068 23092 32124
rect 23092 32068 23096 32124
rect 23032 32064 23096 32068
rect 23112 32124 23176 32128
rect 23112 32068 23116 32124
rect 23116 32068 23172 32124
rect 23172 32068 23176 32124
rect 23112 32064 23176 32068
rect 23192 32124 23256 32128
rect 23192 32068 23196 32124
rect 23196 32068 23252 32124
rect 23252 32068 23256 32124
rect 23192 32064 23256 32068
rect 7952 31580 8016 31584
rect 7952 31524 7956 31580
rect 7956 31524 8012 31580
rect 8012 31524 8016 31580
rect 7952 31520 8016 31524
rect 8032 31580 8096 31584
rect 8032 31524 8036 31580
rect 8036 31524 8092 31580
rect 8092 31524 8096 31580
rect 8032 31520 8096 31524
rect 8112 31580 8176 31584
rect 8112 31524 8116 31580
rect 8116 31524 8172 31580
rect 8172 31524 8176 31580
rect 8112 31520 8176 31524
rect 8192 31580 8256 31584
rect 8192 31524 8196 31580
rect 8196 31524 8252 31580
rect 8252 31524 8256 31580
rect 8192 31520 8256 31524
rect 17952 31580 18016 31584
rect 17952 31524 17956 31580
rect 17956 31524 18012 31580
rect 18012 31524 18016 31580
rect 17952 31520 18016 31524
rect 18032 31580 18096 31584
rect 18032 31524 18036 31580
rect 18036 31524 18092 31580
rect 18092 31524 18096 31580
rect 18032 31520 18096 31524
rect 18112 31580 18176 31584
rect 18112 31524 18116 31580
rect 18116 31524 18172 31580
rect 18172 31524 18176 31580
rect 18112 31520 18176 31524
rect 18192 31580 18256 31584
rect 18192 31524 18196 31580
rect 18196 31524 18252 31580
rect 18252 31524 18256 31580
rect 18192 31520 18256 31524
rect 2952 31036 3016 31040
rect 2952 30980 2956 31036
rect 2956 30980 3012 31036
rect 3012 30980 3016 31036
rect 2952 30976 3016 30980
rect 3032 31036 3096 31040
rect 3032 30980 3036 31036
rect 3036 30980 3092 31036
rect 3092 30980 3096 31036
rect 3032 30976 3096 30980
rect 3112 31036 3176 31040
rect 3112 30980 3116 31036
rect 3116 30980 3172 31036
rect 3172 30980 3176 31036
rect 3112 30976 3176 30980
rect 3192 31036 3256 31040
rect 3192 30980 3196 31036
rect 3196 30980 3252 31036
rect 3252 30980 3256 31036
rect 3192 30976 3256 30980
rect 12952 31036 13016 31040
rect 12952 30980 12956 31036
rect 12956 30980 13012 31036
rect 13012 30980 13016 31036
rect 12952 30976 13016 30980
rect 13032 31036 13096 31040
rect 13032 30980 13036 31036
rect 13036 30980 13092 31036
rect 13092 30980 13096 31036
rect 13032 30976 13096 30980
rect 13112 31036 13176 31040
rect 13112 30980 13116 31036
rect 13116 30980 13172 31036
rect 13172 30980 13176 31036
rect 13112 30976 13176 30980
rect 13192 31036 13256 31040
rect 13192 30980 13196 31036
rect 13196 30980 13252 31036
rect 13252 30980 13256 31036
rect 13192 30976 13256 30980
rect 22952 31036 23016 31040
rect 22952 30980 22956 31036
rect 22956 30980 23012 31036
rect 23012 30980 23016 31036
rect 22952 30976 23016 30980
rect 23032 31036 23096 31040
rect 23032 30980 23036 31036
rect 23036 30980 23092 31036
rect 23092 30980 23096 31036
rect 23032 30976 23096 30980
rect 23112 31036 23176 31040
rect 23112 30980 23116 31036
rect 23116 30980 23172 31036
rect 23172 30980 23176 31036
rect 23112 30976 23176 30980
rect 23192 31036 23256 31040
rect 23192 30980 23196 31036
rect 23196 30980 23252 31036
rect 23252 30980 23256 31036
rect 23192 30976 23256 30980
rect 7952 30492 8016 30496
rect 7952 30436 7956 30492
rect 7956 30436 8012 30492
rect 8012 30436 8016 30492
rect 7952 30432 8016 30436
rect 8032 30492 8096 30496
rect 8032 30436 8036 30492
rect 8036 30436 8092 30492
rect 8092 30436 8096 30492
rect 8032 30432 8096 30436
rect 8112 30492 8176 30496
rect 8112 30436 8116 30492
rect 8116 30436 8172 30492
rect 8172 30436 8176 30492
rect 8112 30432 8176 30436
rect 8192 30492 8256 30496
rect 8192 30436 8196 30492
rect 8196 30436 8252 30492
rect 8252 30436 8256 30492
rect 8192 30432 8256 30436
rect 17952 30492 18016 30496
rect 17952 30436 17956 30492
rect 17956 30436 18012 30492
rect 18012 30436 18016 30492
rect 17952 30432 18016 30436
rect 18032 30492 18096 30496
rect 18032 30436 18036 30492
rect 18036 30436 18092 30492
rect 18092 30436 18096 30492
rect 18032 30432 18096 30436
rect 18112 30492 18176 30496
rect 18112 30436 18116 30492
rect 18116 30436 18172 30492
rect 18172 30436 18176 30492
rect 18112 30432 18176 30436
rect 18192 30492 18256 30496
rect 18192 30436 18196 30492
rect 18196 30436 18252 30492
rect 18252 30436 18256 30492
rect 18192 30432 18256 30436
rect 2952 29948 3016 29952
rect 2952 29892 2956 29948
rect 2956 29892 3012 29948
rect 3012 29892 3016 29948
rect 2952 29888 3016 29892
rect 3032 29948 3096 29952
rect 3032 29892 3036 29948
rect 3036 29892 3092 29948
rect 3092 29892 3096 29948
rect 3032 29888 3096 29892
rect 3112 29948 3176 29952
rect 3112 29892 3116 29948
rect 3116 29892 3172 29948
rect 3172 29892 3176 29948
rect 3112 29888 3176 29892
rect 3192 29948 3256 29952
rect 3192 29892 3196 29948
rect 3196 29892 3252 29948
rect 3252 29892 3256 29948
rect 3192 29888 3256 29892
rect 12952 29948 13016 29952
rect 12952 29892 12956 29948
rect 12956 29892 13012 29948
rect 13012 29892 13016 29948
rect 12952 29888 13016 29892
rect 13032 29948 13096 29952
rect 13032 29892 13036 29948
rect 13036 29892 13092 29948
rect 13092 29892 13096 29948
rect 13032 29888 13096 29892
rect 13112 29948 13176 29952
rect 13112 29892 13116 29948
rect 13116 29892 13172 29948
rect 13172 29892 13176 29948
rect 13112 29888 13176 29892
rect 13192 29948 13256 29952
rect 13192 29892 13196 29948
rect 13196 29892 13252 29948
rect 13252 29892 13256 29948
rect 13192 29888 13256 29892
rect 22952 29948 23016 29952
rect 22952 29892 22956 29948
rect 22956 29892 23012 29948
rect 23012 29892 23016 29948
rect 22952 29888 23016 29892
rect 23032 29948 23096 29952
rect 23032 29892 23036 29948
rect 23036 29892 23092 29948
rect 23092 29892 23096 29948
rect 23032 29888 23096 29892
rect 23112 29948 23176 29952
rect 23112 29892 23116 29948
rect 23116 29892 23172 29948
rect 23172 29892 23176 29948
rect 23112 29888 23176 29892
rect 23192 29948 23256 29952
rect 23192 29892 23196 29948
rect 23196 29892 23252 29948
rect 23252 29892 23256 29948
rect 23192 29888 23256 29892
rect 7952 29404 8016 29408
rect 7952 29348 7956 29404
rect 7956 29348 8012 29404
rect 8012 29348 8016 29404
rect 7952 29344 8016 29348
rect 8032 29404 8096 29408
rect 8032 29348 8036 29404
rect 8036 29348 8092 29404
rect 8092 29348 8096 29404
rect 8032 29344 8096 29348
rect 8112 29404 8176 29408
rect 8112 29348 8116 29404
rect 8116 29348 8172 29404
rect 8172 29348 8176 29404
rect 8112 29344 8176 29348
rect 8192 29404 8256 29408
rect 8192 29348 8196 29404
rect 8196 29348 8252 29404
rect 8252 29348 8256 29404
rect 8192 29344 8256 29348
rect 17952 29404 18016 29408
rect 17952 29348 17956 29404
rect 17956 29348 18012 29404
rect 18012 29348 18016 29404
rect 17952 29344 18016 29348
rect 18032 29404 18096 29408
rect 18032 29348 18036 29404
rect 18036 29348 18092 29404
rect 18092 29348 18096 29404
rect 18032 29344 18096 29348
rect 18112 29404 18176 29408
rect 18112 29348 18116 29404
rect 18116 29348 18172 29404
rect 18172 29348 18176 29404
rect 18112 29344 18176 29348
rect 18192 29404 18256 29408
rect 18192 29348 18196 29404
rect 18196 29348 18252 29404
rect 18252 29348 18256 29404
rect 18192 29344 18256 29348
rect 2952 28860 3016 28864
rect 2952 28804 2956 28860
rect 2956 28804 3012 28860
rect 3012 28804 3016 28860
rect 2952 28800 3016 28804
rect 3032 28860 3096 28864
rect 3032 28804 3036 28860
rect 3036 28804 3092 28860
rect 3092 28804 3096 28860
rect 3032 28800 3096 28804
rect 3112 28860 3176 28864
rect 3112 28804 3116 28860
rect 3116 28804 3172 28860
rect 3172 28804 3176 28860
rect 3112 28800 3176 28804
rect 3192 28860 3256 28864
rect 3192 28804 3196 28860
rect 3196 28804 3252 28860
rect 3252 28804 3256 28860
rect 3192 28800 3256 28804
rect 12952 28860 13016 28864
rect 12952 28804 12956 28860
rect 12956 28804 13012 28860
rect 13012 28804 13016 28860
rect 12952 28800 13016 28804
rect 13032 28860 13096 28864
rect 13032 28804 13036 28860
rect 13036 28804 13092 28860
rect 13092 28804 13096 28860
rect 13032 28800 13096 28804
rect 13112 28860 13176 28864
rect 13112 28804 13116 28860
rect 13116 28804 13172 28860
rect 13172 28804 13176 28860
rect 13112 28800 13176 28804
rect 13192 28860 13256 28864
rect 13192 28804 13196 28860
rect 13196 28804 13252 28860
rect 13252 28804 13256 28860
rect 13192 28800 13256 28804
rect 22952 28860 23016 28864
rect 22952 28804 22956 28860
rect 22956 28804 23012 28860
rect 23012 28804 23016 28860
rect 22952 28800 23016 28804
rect 23032 28860 23096 28864
rect 23032 28804 23036 28860
rect 23036 28804 23092 28860
rect 23092 28804 23096 28860
rect 23032 28800 23096 28804
rect 23112 28860 23176 28864
rect 23112 28804 23116 28860
rect 23116 28804 23172 28860
rect 23172 28804 23176 28860
rect 23112 28800 23176 28804
rect 23192 28860 23256 28864
rect 23192 28804 23196 28860
rect 23196 28804 23252 28860
rect 23252 28804 23256 28860
rect 23192 28800 23256 28804
rect 7952 28316 8016 28320
rect 7952 28260 7956 28316
rect 7956 28260 8012 28316
rect 8012 28260 8016 28316
rect 7952 28256 8016 28260
rect 8032 28316 8096 28320
rect 8032 28260 8036 28316
rect 8036 28260 8092 28316
rect 8092 28260 8096 28316
rect 8032 28256 8096 28260
rect 8112 28316 8176 28320
rect 8112 28260 8116 28316
rect 8116 28260 8172 28316
rect 8172 28260 8176 28316
rect 8112 28256 8176 28260
rect 8192 28316 8256 28320
rect 8192 28260 8196 28316
rect 8196 28260 8252 28316
rect 8252 28260 8256 28316
rect 8192 28256 8256 28260
rect 17952 28316 18016 28320
rect 17952 28260 17956 28316
rect 17956 28260 18012 28316
rect 18012 28260 18016 28316
rect 17952 28256 18016 28260
rect 18032 28316 18096 28320
rect 18032 28260 18036 28316
rect 18036 28260 18092 28316
rect 18092 28260 18096 28316
rect 18032 28256 18096 28260
rect 18112 28316 18176 28320
rect 18112 28260 18116 28316
rect 18116 28260 18172 28316
rect 18172 28260 18176 28316
rect 18112 28256 18176 28260
rect 18192 28316 18256 28320
rect 18192 28260 18196 28316
rect 18196 28260 18252 28316
rect 18252 28260 18256 28316
rect 18192 28256 18256 28260
rect 2952 27772 3016 27776
rect 2952 27716 2956 27772
rect 2956 27716 3012 27772
rect 3012 27716 3016 27772
rect 2952 27712 3016 27716
rect 3032 27772 3096 27776
rect 3032 27716 3036 27772
rect 3036 27716 3092 27772
rect 3092 27716 3096 27772
rect 3032 27712 3096 27716
rect 3112 27772 3176 27776
rect 3112 27716 3116 27772
rect 3116 27716 3172 27772
rect 3172 27716 3176 27772
rect 3112 27712 3176 27716
rect 3192 27772 3256 27776
rect 3192 27716 3196 27772
rect 3196 27716 3252 27772
rect 3252 27716 3256 27772
rect 3192 27712 3256 27716
rect 12952 27772 13016 27776
rect 12952 27716 12956 27772
rect 12956 27716 13012 27772
rect 13012 27716 13016 27772
rect 12952 27712 13016 27716
rect 13032 27772 13096 27776
rect 13032 27716 13036 27772
rect 13036 27716 13092 27772
rect 13092 27716 13096 27772
rect 13032 27712 13096 27716
rect 13112 27772 13176 27776
rect 13112 27716 13116 27772
rect 13116 27716 13172 27772
rect 13172 27716 13176 27772
rect 13112 27712 13176 27716
rect 13192 27772 13256 27776
rect 13192 27716 13196 27772
rect 13196 27716 13252 27772
rect 13252 27716 13256 27772
rect 13192 27712 13256 27716
rect 22952 27772 23016 27776
rect 22952 27716 22956 27772
rect 22956 27716 23012 27772
rect 23012 27716 23016 27772
rect 22952 27712 23016 27716
rect 23032 27772 23096 27776
rect 23032 27716 23036 27772
rect 23036 27716 23092 27772
rect 23092 27716 23096 27772
rect 23032 27712 23096 27716
rect 23112 27772 23176 27776
rect 23112 27716 23116 27772
rect 23116 27716 23172 27772
rect 23172 27716 23176 27772
rect 23112 27712 23176 27716
rect 23192 27772 23256 27776
rect 23192 27716 23196 27772
rect 23196 27716 23252 27772
rect 23252 27716 23256 27772
rect 23192 27712 23256 27716
rect 7952 27228 8016 27232
rect 7952 27172 7956 27228
rect 7956 27172 8012 27228
rect 8012 27172 8016 27228
rect 7952 27168 8016 27172
rect 8032 27228 8096 27232
rect 8032 27172 8036 27228
rect 8036 27172 8092 27228
rect 8092 27172 8096 27228
rect 8032 27168 8096 27172
rect 8112 27228 8176 27232
rect 8112 27172 8116 27228
rect 8116 27172 8172 27228
rect 8172 27172 8176 27228
rect 8112 27168 8176 27172
rect 8192 27228 8256 27232
rect 8192 27172 8196 27228
rect 8196 27172 8252 27228
rect 8252 27172 8256 27228
rect 8192 27168 8256 27172
rect 17952 27228 18016 27232
rect 17952 27172 17956 27228
rect 17956 27172 18012 27228
rect 18012 27172 18016 27228
rect 17952 27168 18016 27172
rect 18032 27228 18096 27232
rect 18032 27172 18036 27228
rect 18036 27172 18092 27228
rect 18092 27172 18096 27228
rect 18032 27168 18096 27172
rect 18112 27228 18176 27232
rect 18112 27172 18116 27228
rect 18116 27172 18172 27228
rect 18172 27172 18176 27228
rect 18112 27168 18176 27172
rect 18192 27228 18256 27232
rect 18192 27172 18196 27228
rect 18196 27172 18252 27228
rect 18252 27172 18256 27228
rect 18192 27168 18256 27172
rect 2952 26684 3016 26688
rect 2952 26628 2956 26684
rect 2956 26628 3012 26684
rect 3012 26628 3016 26684
rect 2952 26624 3016 26628
rect 3032 26684 3096 26688
rect 3032 26628 3036 26684
rect 3036 26628 3092 26684
rect 3092 26628 3096 26684
rect 3032 26624 3096 26628
rect 3112 26684 3176 26688
rect 3112 26628 3116 26684
rect 3116 26628 3172 26684
rect 3172 26628 3176 26684
rect 3112 26624 3176 26628
rect 3192 26684 3256 26688
rect 3192 26628 3196 26684
rect 3196 26628 3252 26684
rect 3252 26628 3256 26684
rect 3192 26624 3256 26628
rect 12952 26684 13016 26688
rect 12952 26628 12956 26684
rect 12956 26628 13012 26684
rect 13012 26628 13016 26684
rect 12952 26624 13016 26628
rect 13032 26684 13096 26688
rect 13032 26628 13036 26684
rect 13036 26628 13092 26684
rect 13092 26628 13096 26684
rect 13032 26624 13096 26628
rect 13112 26684 13176 26688
rect 13112 26628 13116 26684
rect 13116 26628 13172 26684
rect 13172 26628 13176 26684
rect 13112 26624 13176 26628
rect 13192 26684 13256 26688
rect 13192 26628 13196 26684
rect 13196 26628 13252 26684
rect 13252 26628 13256 26684
rect 13192 26624 13256 26628
rect 22952 26684 23016 26688
rect 22952 26628 22956 26684
rect 22956 26628 23012 26684
rect 23012 26628 23016 26684
rect 22952 26624 23016 26628
rect 23032 26684 23096 26688
rect 23032 26628 23036 26684
rect 23036 26628 23092 26684
rect 23092 26628 23096 26684
rect 23032 26624 23096 26628
rect 23112 26684 23176 26688
rect 23112 26628 23116 26684
rect 23116 26628 23172 26684
rect 23172 26628 23176 26684
rect 23112 26624 23176 26628
rect 23192 26684 23256 26688
rect 23192 26628 23196 26684
rect 23196 26628 23252 26684
rect 23252 26628 23256 26684
rect 23192 26624 23256 26628
rect 7952 26140 8016 26144
rect 7952 26084 7956 26140
rect 7956 26084 8012 26140
rect 8012 26084 8016 26140
rect 7952 26080 8016 26084
rect 8032 26140 8096 26144
rect 8032 26084 8036 26140
rect 8036 26084 8092 26140
rect 8092 26084 8096 26140
rect 8032 26080 8096 26084
rect 8112 26140 8176 26144
rect 8112 26084 8116 26140
rect 8116 26084 8172 26140
rect 8172 26084 8176 26140
rect 8112 26080 8176 26084
rect 8192 26140 8256 26144
rect 8192 26084 8196 26140
rect 8196 26084 8252 26140
rect 8252 26084 8256 26140
rect 8192 26080 8256 26084
rect 17952 26140 18016 26144
rect 17952 26084 17956 26140
rect 17956 26084 18012 26140
rect 18012 26084 18016 26140
rect 17952 26080 18016 26084
rect 18032 26140 18096 26144
rect 18032 26084 18036 26140
rect 18036 26084 18092 26140
rect 18092 26084 18096 26140
rect 18032 26080 18096 26084
rect 18112 26140 18176 26144
rect 18112 26084 18116 26140
rect 18116 26084 18172 26140
rect 18172 26084 18176 26140
rect 18112 26080 18176 26084
rect 18192 26140 18256 26144
rect 18192 26084 18196 26140
rect 18196 26084 18252 26140
rect 18252 26084 18256 26140
rect 18192 26080 18256 26084
rect 17540 25936 17604 25940
rect 17540 25880 17590 25936
rect 17590 25880 17604 25936
rect 17540 25876 17604 25880
rect 2952 25596 3016 25600
rect 2952 25540 2956 25596
rect 2956 25540 3012 25596
rect 3012 25540 3016 25596
rect 2952 25536 3016 25540
rect 3032 25596 3096 25600
rect 3032 25540 3036 25596
rect 3036 25540 3092 25596
rect 3092 25540 3096 25596
rect 3032 25536 3096 25540
rect 3112 25596 3176 25600
rect 3112 25540 3116 25596
rect 3116 25540 3172 25596
rect 3172 25540 3176 25596
rect 3112 25536 3176 25540
rect 3192 25596 3256 25600
rect 3192 25540 3196 25596
rect 3196 25540 3252 25596
rect 3252 25540 3256 25596
rect 3192 25536 3256 25540
rect 12952 25596 13016 25600
rect 12952 25540 12956 25596
rect 12956 25540 13012 25596
rect 13012 25540 13016 25596
rect 12952 25536 13016 25540
rect 13032 25596 13096 25600
rect 13032 25540 13036 25596
rect 13036 25540 13092 25596
rect 13092 25540 13096 25596
rect 13032 25536 13096 25540
rect 13112 25596 13176 25600
rect 13112 25540 13116 25596
rect 13116 25540 13172 25596
rect 13172 25540 13176 25596
rect 13112 25536 13176 25540
rect 13192 25596 13256 25600
rect 13192 25540 13196 25596
rect 13196 25540 13252 25596
rect 13252 25540 13256 25596
rect 13192 25536 13256 25540
rect 22952 25596 23016 25600
rect 22952 25540 22956 25596
rect 22956 25540 23012 25596
rect 23012 25540 23016 25596
rect 22952 25536 23016 25540
rect 23032 25596 23096 25600
rect 23032 25540 23036 25596
rect 23036 25540 23092 25596
rect 23092 25540 23096 25596
rect 23032 25536 23096 25540
rect 23112 25596 23176 25600
rect 23112 25540 23116 25596
rect 23116 25540 23172 25596
rect 23172 25540 23176 25596
rect 23112 25536 23176 25540
rect 23192 25596 23256 25600
rect 23192 25540 23196 25596
rect 23196 25540 23252 25596
rect 23252 25540 23256 25596
rect 23192 25536 23256 25540
rect 15332 25060 15396 25124
rect 7952 25052 8016 25056
rect 7952 24996 7956 25052
rect 7956 24996 8012 25052
rect 8012 24996 8016 25052
rect 7952 24992 8016 24996
rect 8032 25052 8096 25056
rect 8032 24996 8036 25052
rect 8036 24996 8092 25052
rect 8092 24996 8096 25052
rect 8032 24992 8096 24996
rect 8112 25052 8176 25056
rect 8112 24996 8116 25052
rect 8116 24996 8172 25052
rect 8172 24996 8176 25052
rect 8112 24992 8176 24996
rect 8192 25052 8256 25056
rect 8192 24996 8196 25052
rect 8196 24996 8252 25052
rect 8252 24996 8256 25052
rect 8192 24992 8256 24996
rect 17952 25052 18016 25056
rect 17952 24996 17956 25052
rect 17956 24996 18012 25052
rect 18012 24996 18016 25052
rect 17952 24992 18016 24996
rect 18032 25052 18096 25056
rect 18032 24996 18036 25052
rect 18036 24996 18092 25052
rect 18092 24996 18096 25052
rect 18032 24992 18096 24996
rect 18112 25052 18176 25056
rect 18112 24996 18116 25052
rect 18116 24996 18172 25052
rect 18172 24996 18176 25052
rect 18112 24992 18176 24996
rect 18192 25052 18256 25056
rect 18192 24996 18196 25052
rect 18196 24996 18252 25052
rect 18252 24996 18256 25052
rect 18192 24992 18256 24996
rect 19932 24984 19996 24988
rect 19932 24928 19946 24984
rect 19946 24928 19996 24984
rect 19932 24924 19996 24928
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 19012 23428 19076 23492
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 16804 22808 16868 22812
rect 16804 22752 16818 22808
rect 16818 22752 16868 22808
rect 16804 22748 16868 22752
rect 20484 22400 20548 22404
rect 20484 22344 20498 22400
rect 20498 22344 20548 22400
rect 20484 22340 20548 22344
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 22140 19756 22204 19820
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 17356 17988 17420 18052
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 12572 17444 12636 17508
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 17540 17308 17604 17372
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 17172 16688 17236 16692
rect 17172 16632 17186 16688
rect 17186 16632 17236 16688
rect 17172 16628 17236 16632
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 16804 16280 16868 16284
rect 16804 16224 16854 16280
rect 16854 16224 16868 16280
rect 16804 16220 16868 16224
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 16988 15268 17052 15332
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 13676 14180 13740 14244
rect 14780 14240 14844 14244
rect 14780 14184 14794 14240
rect 14794 14184 14844 14240
rect 14780 14180 14844 14184
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 17356 13560 17420 13564
rect 17356 13504 17406 13560
rect 17406 13504 17420 13560
rect 17356 13500 17420 13504
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 13676 11732 13740 11796
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 18460 10236 18524 10300
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 16804 8528 16868 8532
rect 16804 8472 16854 8528
rect 16854 8472 16868 8528
rect 16804 8468 16868 8472
rect 22324 8332 22388 8396
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 15332 7244 15396 7308
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 16804 6836 16868 6900
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 22324 4660 22388 4724
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 22140 4116 22204 4180
rect 18460 3844 18524 3908
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 12572 3572 12636 3636
rect 16988 3572 17052 3636
rect 19012 3436 19076 3500
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 17172 3028 17236 3092
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 14780 2484 14844 2548
rect 19932 2348 19996 2412
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 20484 1804 20548 1868
<< metal4 >>
rect 2944 53888 3264 54448
rect 2944 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3264 53888
rect 2944 52800 3264 53824
rect 2944 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3264 52800
rect 2944 51712 3264 52736
rect 2944 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3264 51712
rect 2944 50624 3264 51648
rect 2944 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3264 50624
rect 2944 49536 3264 50560
rect 2944 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3264 49536
rect 2944 48448 3264 49472
rect 2944 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3264 48448
rect 2944 47360 3264 48384
rect 2944 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3264 47360
rect 2944 46272 3264 47296
rect 2944 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3264 46272
rect 2944 45184 3264 46208
rect 2944 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3264 45184
rect 2944 44096 3264 45120
rect 2944 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3264 44096
rect 2944 43008 3264 44032
rect 2944 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3264 43008
rect 2944 41920 3264 42944
rect 2944 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3264 41920
rect 2944 40832 3264 41856
rect 2944 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3264 40832
rect 2944 39744 3264 40768
rect 2944 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3264 39744
rect 2944 38656 3264 39680
rect 2944 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3264 38656
rect 2944 37568 3264 38592
rect 2944 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3264 37568
rect 2944 36480 3264 37504
rect 2944 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3264 36480
rect 2944 35392 3264 36416
rect 2944 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3264 35392
rect 2944 34304 3264 35328
rect 2944 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3264 34304
rect 2944 33216 3264 34240
rect 2944 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3264 33216
rect 2944 32128 3264 33152
rect 2944 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3264 32128
rect 2944 31040 3264 32064
rect 2944 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3264 31040
rect 2944 29952 3264 30976
rect 2944 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3264 29952
rect 2944 28864 3264 29888
rect 2944 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3264 28864
rect 2944 27776 3264 28800
rect 2944 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3264 27776
rect 2944 26688 3264 27712
rect 2944 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3264 26688
rect 2944 25600 3264 26624
rect 2944 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3264 25600
rect 2944 24512 3264 25536
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 54432 8264 54448
rect 7944 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8264 54432
rect 7944 53344 8264 54368
rect 7944 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8264 53344
rect 7944 52256 8264 53280
rect 7944 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8264 52256
rect 7944 51168 8264 52192
rect 7944 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8264 51168
rect 7944 50080 8264 51104
rect 7944 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8264 50080
rect 7944 48992 8264 50016
rect 7944 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8264 48992
rect 7944 47904 8264 48928
rect 7944 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8264 47904
rect 7944 46816 8264 47840
rect 7944 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8264 46816
rect 7944 45728 8264 46752
rect 7944 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8264 45728
rect 7944 44640 8264 45664
rect 7944 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8264 44640
rect 7944 43552 8264 44576
rect 7944 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8264 43552
rect 7944 42464 8264 43488
rect 7944 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8264 42464
rect 7944 41376 8264 42400
rect 7944 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8264 41376
rect 7944 40288 8264 41312
rect 7944 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8264 40288
rect 7944 39200 8264 40224
rect 7944 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8264 39200
rect 7944 38112 8264 39136
rect 7944 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8264 38112
rect 7944 37024 8264 38048
rect 7944 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8264 37024
rect 7944 35936 8264 36960
rect 7944 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8264 35936
rect 7944 34848 8264 35872
rect 7944 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8264 34848
rect 7944 33760 8264 34784
rect 7944 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8264 33760
rect 7944 32672 8264 33696
rect 7944 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8264 32672
rect 7944 31584 8264 32608
rect 7944 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8264 31584
rect 7944 30496 8264 31520
rect 7944 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8264 30496
rect 7944 29408 8264 30432
rect 7944 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8264 29408
rect 7944 28320 8264 29344
rect 7944 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8264 28320
rect 7944 27232 8264 28256
rect 7944 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8264 27232
rect 7944 26144 8264 27168
rect 7944 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8264 26144
rect 7944 25056 8264 26080
rect 7944 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8264 25056
rect 7944 23968 8264 24992
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 12944 53888 13264 54448
rect 12944 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13264 53888
rect 12944 52800 13264 53824
rect 12944 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13264 52800
rect 12944 51712 13264 52736
rect 12944 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13264 51712
rect 12944 50624 13264 51648
rect 12944 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13264 50624
rect 12944 49536 13264 50560
rect 12944 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13264 49536
rect 12944 48448 13264 49472
rect 12944 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13264 48448
rect 12944 47360 13264 48384
rect 12944 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13264 47360
rect 12944 46272 13264 47296
rect 12944 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13264 46272
rect 12944 45184 13264 46208
rect 12944 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13264 45184
rect 12944 44096 13264 45120
rect 12944 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13264 44096
rect 12944 43008 13264 44032
rect 12944 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13264 43008
rect 12944 41920 13264 42944
rect 12944 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13264 41920
rect 12944 40832 13264 41856
rect 12944 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13264 40832
rect 12944 39744 13264 40768
rect 12944 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13264 39744
rect 12944 38656 13264 39680
rect 12944 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13264 38656
rect 12944 37568 13264 38592
rect 12944 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13264 37568
rect 12944 36480 13264 37504
rect 12944 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13264 36480
rect 12944 35392 13264 36416
rect 12944 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13264 35392
rect 12944 34304 13264 35328
rect 12944 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13264 34304
rect 12944 33216 13264 34240
rect 12944 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13264 33216
rect 12944 32128 13264 33152
rect 12944 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13264 32128
rect 12944 31040 13264 32064
rect 12944 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13264 31040
rect 12944 29952 13264 30976
rect 12944 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13264 29952
rect 12944 28864 13264 29888
rect 12944 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13264 28864
rect 12944 27776 13264 28800
rect 12944 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13264 27776
rect 12944 26688 13264 27712
rect 12944 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13264 26688
rect 12944 25600 13264 26624
rect 17944 54432 18264 54448
rect 17944 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18264 54432
rect 17944 53344 18264 54368
rect 17944 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18264 53344
rect 17944 52256 18264 53280
rect 17944 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18264 52256
rect 17944 51168 18264 52192
rect 17944 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18264 51168
rect 17944 50080 18264 51104
rect 17944 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18264 50080
rect 17944 48992 18264 50016
rect 17944 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18264 48992
rect 17944 47904 18264 48928
rect 17944 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18264 47904
rect 17944 46816 18264 47840
rect 17944 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18264 46816
rect 17944 45728 18264 46752
rect 17944 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18264 45728
rect 17944 44640 18264 45664
rect 17944 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18264 44640
rect 17944 43552 18264 44576
rect 17944 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18264 43552
rect 17944 42464 18264 43488
rect 17944 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18264 42464
rect 17944 41376 18264 42400
rect 17944 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18264 41376
rect 17944 40288 18264 41312
rect 17944 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18264 40288
rect 17944 39200 18264 40224
rect 17944 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18264 39200
rect 17944 38112 18264 39136
rect 17944 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18264 38112
rect 17944 37024 18264 38048
rect 17944 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18264 37024
rect 17944 35936 18264 36960
rect 17944 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18264 35936
rect 17944 34848 18264 35872
rect 17944 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18264 34848
rect 17944 33760 18264 34784
rect 17944 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18264 33760
rect 17944 32672 18264 33696
rect 17944 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18264 32672
rect 17944 31584 18264 32608
rect 17944 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18264 31584
rect 17944 30496 18264 31520
rect 17944 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18264 30496
rect 17944 29408 18264 30432
rect 17944 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18264 29408
rect 17944 28320 18264 29344
rect 17944 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18264 28320
rect 17944 27232 18264 28256
rect 17944 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18264 27232
rect 17944 26144 18264 27168
rect 17944 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18264 26144
rect 17539 25940 17605 25941
rect 17539 25876 17540 25940
rect 17604 25876 17605 25940
rect 17539 25875 17605 25876
rect 12944 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13264 25600
rect 12944 24512 13264 25536
rect 15331 25124 15397 25125
rect 15331 25060 15332 25124
rect 15396 25060 15397 25124
rect 15331 25059 15397 25060
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12571 17508 12637 17509
rect 12571 17444 12572 17508
rect 12636 17444 12637 17508
rect 12571 17443 12637 17444
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 12574 3637 12634 17443
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 13675 14244 13741 14245
rect 13675 14180 13676 14244
rect 13740 14180 13741 14244
rect 13675 14179 13741 14180
rect 14779 14244 14845 14245
rect 14779 14180 14780 14244
rect 14844 14180 14845 14244
rect 14779 14179 14845 14180
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 13678 11797 13738 14179
rect 13675 11796 13741 11797
rect 13675 11732 13676 11796
rect 13740 11732 13741 11796
rect 13675 11731 13741 11732
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12571 3636 12637 3637
rect 12571 3572 12572 3636
rect 12636 3572 12637 3636
rect 12571 3571 12637 3572
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 14782 2549 14842 14179
rect 15334 7309 15394 25059
rect 16803 22812 16869 22813
rect 16803 22748 16804 22812
rect 16868 22748 16869 22812
rect 16803 22747 16869 22748
rect 16806 16285 16866 22747
rect 17355 18052 17421 18053
rect 17355 17988 17356 18052
rect 17420 17988 17421 18052
rect 17355 17987 17421 17988
rect 17171 16692 17237 16693
rect 17171 16628 17172 16692
rect 17236 16628 17237 16692
rect 17171 16627 17237 16628
rect 16803 16284 16869 16285
rect 16803 16220 16804 16284
rect 16868 16220 16869 16284
rect 16803 16219 16869 16220
rect 16987 15332 17053 15333
rect 16987 15268 16988 15332
rect 17052 15268 17053 15332
rect 16987 15267 17053 15268
rect 16803 8532 16869 8533
rect 16803 8468 16804 8532
rect 16868 8468 16869 8532
rect 16803 8467 16869 8468
rect 15331 7308 15397 7309
rect 15331 7244 15332 7308
rect 15396 7244 15397 7308
rect 15331 7243 15397 7244
rect 16806 6901 16866 8467
rect 16803 6900 16869 6901
rect 16803 6836 16804 6900
rect 16868 6836 16869 6900
rect 16803 6835 16869 6836
rect 16990 3637 17050 15267
rect 16987 3636 17053 3637
rect 16987 3572 16988 3636
rect 17052 3572 17053 3636
rect 16987 3571 17053 3572
rect 17174 3093 17234 16627
rect 17358 13565 17418 17987
rect 17542 17373 17602 25875
rect 17944 25056 18264 26080
rect 17944 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18264 25056
rect 17944 23968 18264 24992
rect 22944 53888 23264 54448
rect 22944 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23264 53888
rect 22944 52800 23264 53824
rect 22944 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23264 52800
rect 22944 51712 23264 52736
rect 22944 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23264 51712
rect 22944 50624 23264 51648
rect 22944 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23264 50624
rect 22944 49536 23264 50560
rect 22944 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23264 49536
rect 22944 48448 23264 49472
rect 22944 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23264 48448
rect 22944 47360 23264 48384
rect 22944 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23264 47360
rect 22944 46272 23264 47296
rect 22944 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23264 46272
rect 22944 45184 23264 46208
rect 22944 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23264 45184
rect 22944 44096 23264 45120
rect 22944 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23264 44096
rect 22944 43008 23264 44032
rect 22944 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23264 43008
rect 22944 41920 23264 42944
rect 22944 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23264 41920
rect 22944 40832 23264 41856
rect 22944 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23264 40832
rect 22944 39744 23264 40768
rect 22944 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23264 39744
rect 22944 38656 23264 39680
rect 22944 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23264 38656
rect 22944 37568 23264 38592
rect 22944 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23264 37568
rect 22944 36480 23264 37504
rect 22944 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23264 36480
rect 22944 35392 23264 36416
rect 22944 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23264 35392
rect 22944 34304 23264 35328
rect 22944 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23264 34304
rect 22944 33216 23264 34240
rect 22944 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23264 33216
rect 22944 32128 23264 33152
rect 22944 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23264 32128
rect 22944 31040 23264 32064
rect 22944 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23264 31040
rect 22944 29952 23264 30976
rect 22944 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23264 29952
rect 22944 28864 23264 29888
rect 22944 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23264 28864
rect 22944 27776 23264 28800
rect 22944 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23264 27776
rect 22944 26688 23264 27712
rect 22944 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23264 26688
rect 22944 25600 23264 26624
rect 22944 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23264 25600
rect 19931 24988 19997 24989
rect 19931 24924 19932 24988
rect 19996 24924 19997 24988
rect 19931 24923 19997 24924
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 19011 23492 19077 23493
rect 19011 23428 19012 23492
rect 19076 23428 19077 23492
rect 19011 23427 19077 23428
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17539 17372 17605 17373
rect 17539 17308 17540 17372
rect 17604 17308 17605 17372
rect 17539 17307 17605 17308
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17355 13564 17421 13565
rect 17355 13500 17356 13564
rect 17420 13500 17421 13564
rect 17355 13499 17421 13500
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 18459 10300 18525 10301
rect 18459 10236 18460 10300
rect 18524 10236 18525 10300
rect 18459 10235 18525 10236
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 18462 3909 18522 10235
rect 18459 3908 18525 3909
rect 18459 3844 18460 3908
rect 18524 3844 18525 3908
rect 18459 3843 18525 3844
rect 19014 3501 19074 23427
rect 19011 3500 19077 3501
rect 19011 3436 19012 3500
rect 19076 3436 19077 3500
rect 19011 3435 19077 3436
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17171 3092 17237 3093
rect 17171 3028 17172 3092
rect 17236 3028 17237 3092
rect 17171 3027 17237 3028
rect 14779 2548 14845 2549
rect 14779 2484 14780 2548
rect 14844 2484 14845 2548
rect 14779 2483 14845 2484
rect 17944 2208 18264 3232
rect 19934 2413 19994 24923
rect 22944 24512 23264 25536
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 20483 22404 20549 22405
rect 20483 22340 20484 22404
rect 20548 22340 20549 22404
rect 20483 22339 20549 22340
rect 19931 2412 19997 2413
rect 19931 2348 19932 2412
rect 19996 2348 19997 2412
rect 19931 2347 19997 2348
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 20486 1869 20546 22339
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22139 19820 22205 19821
rect 22139 19756 22140 19820
rect 22204 19756 22205 19820
rect 22139 19755 22205 19756
rect 22142 16590 22202 19755
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22142 16530 22386 16590
rect 22326 12450 22386 16530
rect 22142 12390 22386 12450
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22142 4181 22202 12390
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22323 8396 22389 8397
rect 22323 8332 22324 8396
rect 22388 8332 22389 8396
rect 22323 8331 22389 8332
rect 22326 4725 22386 8331
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22323 4724 22389 4725
rect 22323 4660 22324 4724
rect 22388 4660 22389 4724
rect 22323 4659 22389 4660
rect 22139 4180 22205 4181
rect 22139 4116 22140 4180
rect 22204 4116 22205 4180
rect 22139 4115 22205 4116
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
rect 20483 1868 20549 1869
rect 20483 1804 20484 1868
rect 20548 1804 20549 1868
rect 20483 1803 20549 1804
use sky130_fd_sc_hd__clkbuf_2  _104_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _105_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14444 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _106_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12880 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _107_
timestamp 1676037725
transform 1 0 15456 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1676037725
transform 1 0 13524 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _109_
timestamp 1676037725
transform 1 0 21344 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1676037725
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _111_
timestamp 1676037725
transform 1 0 24472 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1676037725
transform -1 0 11224 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _114_
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1676037725
transform 1 0 24564 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1676037725
transform 1 0 24564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1676037725
transform 1 0 25024 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1676037725
transform 1 0 24840 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1676037725
transform 1 0 25024 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1676037725
transform 1 0 24564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1676037725
transform 1 0 21988 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1676037725
transform 1 0 24564 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1676037725
transform 1 0 21988 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 1676037725
transform 1 0 22724 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1676037725
transform 1 0 21988 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1676037725
transform 1 0 20792 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1676037725
transform 1 0 21620 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1676037725
transform 1 0 23736 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1676037725
transform 1 0 22172 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 1676037725
transform 1 0 20792 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1676037725
transform 1 0 21528 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1676037725
transform 1 0 19412 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1676037725
transform 1 0 19688 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1676037725
transform 1 0 16836 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _137_
timestamp 1676037725
transform 1 0 17112 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 1676037725
transform 1 0 13524 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1676037725
transform 1 0 13800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1676037725
transform 1 0 16744 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1676037725
transform 1 0 17480 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1676037725
transform 1 0 17756 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1676037725
transform 1 0 18492 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1676037725
transform 1 0 19228 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1676037725
transform 1 0 19412 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1676037725
transform 1 0 18584 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1676037725
transform 1 0 16008 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1676037725
transform 1 0 16376 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1676037725
transform 1 0 19964 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1676037725
transform 1 0 20792 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1676037725
transform 1 0 21896 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1676037725
transform 1 0 17480 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp 1676037725
transform 1 0 19412 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1676037725
transform 1 0 20976 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1676037725
transform 1 0 23092 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1676037725
transform 1 0 23828 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _159_
timestamp 1676037725
transform 1 0 20608 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1676037725
transform 1 0 18584 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _161_
timestamp 1676037725
transform 1 0 24564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _162_
timestamp 1676037725
transform 1 0 21988 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1676037725
transform 1 0 23552 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1676037725
transform 1 0 5152 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1676037725
transform 1 0 6532 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _166_
timestamp 1676037725
transform 1 0 7544 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp 1676037725
transform 1 0 9200 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1676037725
transform 1 0 8280 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _169_
timestamp 1676037725
transform 1 0 9384 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _170_
timestamp 1676037725
transform 1 0 10396 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _171_
timestamp 1676037725
transform 1 0 11408 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10948 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1676037725
transform 1 0 20240 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__A
timestamp 1676037725
transform 1 0 17388 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__A
timestamp 1676037725
transform 1 0 16744 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1676037725
transform 1 0 17388 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1676037725
transform 1 0 19044 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1676037725
transform 1 0 19964 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A
timestamp 1676037725
transform 1 0 21160 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A
timestamp 1676037725
transform 1 0 21344 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1676037725
transform 1 0 21988 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 7360 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 10304 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 8556 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 8556 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 10120 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 9292 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 8464 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 9568 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12052 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 10948 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 10028 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11868 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 10028 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 10948 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 16008 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 13432 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 16192 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 15272 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 9476 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 14168 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 9844 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 15732 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 14812 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 9660 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 17296 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11132 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8648 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1676037725
transform 1 0 18860 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1676037725
transform 1 0 12144 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1676037725
transform 1 0 13708 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1676037725
transform 1 0 16284 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1676037725
transform 1 0 20608 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1676037725
transform 1 0 16836 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1676037725
transform 1 0 15732 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1676037725
transform 1 0 15548 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1676037725
transform 1 0 15824 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1676037725
transform 1 0 19320 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1676037725
transform 1 0 19504 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1676037725
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1676037725
transform 1 0 24748 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1676037725
transform 1 0 24748 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1676037725
transform 1 0 25392 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1676037725
transform 1 0 24748 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1676037725
transform 1 0 25392 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1676037725
transform 1 0 24656 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1676037725
transform 1 0 25392 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1676037725
transform 1 0 24748 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1676037725
transform 1 0 25392 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1676037725
transform 1 0 24748 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1676037725
transform 1 0 25392 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1676037725
transform 1 0 25208 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1676037725
transform 1 0 24656 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1676037725
transform 1 0 25392 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1676037725
transform 1 0 24656 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1676037725
transform 1 0 25392 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1676037725
transform 1 0 24748 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1676037725
transform 1 0 25392 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1676037725
transform 1 0 24748 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1676037725
transform 1 0 25392 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1676037725
transform 1 0 24656 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1676037725
transform 1 0 25392 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1676037725
transform 1 0 24564 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1676037725
transform 1 0 22816 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1676037725
transform 1 0 25392 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1676037725
transform 1 0 25392 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1676037725
transform 1 0 24748 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1676037725
transform 1 0 24748 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1676037725
transform 1 0 24748 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1676037725
transform 1 0 2668 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1676037725
transform 1 0 6532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1676037725
transform 1 0 4140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1676037725
transform 1 0 6716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1676037725
transform 1 0 7728 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1676037725
transform 1 0 7544 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1676037725
transform 1 0 7636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1676037725
transform 1 0 8004 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1676037725
transform 1 0 7820 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1676037725
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1676037725
transform 1 0 9752 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1676037725
transform 1 0 9292 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1676037725
transform 1 0 8924 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1676037725
transform 1 0 9108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1676037725
transform 1 0 10580 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1676037725
transform 1 0 9292 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1676037725
transform 1 0 11224 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1676037725
transform 1 0 11684 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1676037725
transform 1 0 3956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1676037725
transform 1 0 3312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1676037725
transform 1 0 2852 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1676037725
transform 1 0 4600 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1676037725
transform 1 0 4508 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1676037725
transform 1 0 13800 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1676037725
transform 1 0 15364 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1676037725
transform 1 0 17296 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1676037725
transform 1 0 18124 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1676037725
transform 1 0 18952 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1676037725
transform 1 0 25392 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1676037725
transform 1 0 24472 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1676037725
transform 1 0 24472 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1676037725
transform 1 0 24472 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1676037725
transform 1 0 25392 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1676037725
transform 1 0 24104 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1676037725
transform 1 0 24380 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1676037725
transform 1 0 24656 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1676037725
transform 1 0 23368 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1676037725
transform 1 0 21252 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1676037725
transform 1 0 22540 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1676037725
transform 1 0 23736 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1676037725
transform 1 0 25116 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output124_A
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20608 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25392 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25392 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25300 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21436 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 23920 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25208 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25392 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24748 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25208 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25208 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21436 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 19964 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18952 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18860 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18768 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18768 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 19412 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21252 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22724 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24472 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25300 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24564 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24104 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24288 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23644 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21252 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21068 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23828 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25392 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22356 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 15456 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 11132 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13708 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12512 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13156 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13616 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 13432 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 15824 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 15272 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14996 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12880 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 11408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 10120 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 8372 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 10948 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 12696 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14352 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 15088 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14536 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14536 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 12236 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 10948 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 12052 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12788 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 15824 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16376 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16928 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 17204 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18124 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18676 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18400 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16928 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16008 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14352 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16100 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16928 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 20424 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22264 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 22448 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22632 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21252 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22264 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24012 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25024 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25024 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25116 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25116 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 19872 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 19320 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18860 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 20332 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 19136 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 25392 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 18860 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 22264 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 25024 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 25392 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_15.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 24012 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_19.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19964 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_29.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19688 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_31.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21436 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 22632 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_35.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 24472 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_45.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 22356 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_47.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21804 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_49.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 20332 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_51.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16744 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16560 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16008 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16192 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 16192 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 9016 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16192 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16376 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 16836 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 10304 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18032 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 17848 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 18676 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 18492 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 11132 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16192 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16376 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 17204 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 17020 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 15272 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15272 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 16836 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 16652 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_12.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 14260 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_12.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_14.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18032 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_14.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18216 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_16.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19044 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_16.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19228 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_18.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16192 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_20.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 13616 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_22.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 12880 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_24.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 12696 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_26.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14628 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_28.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18492 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_28.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18676 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_30.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_30.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19044 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_32.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18676 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_32.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18860 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_34.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 17848 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_34.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18032 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_36.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14352 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_38.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_40.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 17848 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_42.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_44.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 20424 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_44.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21252 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_46.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21160 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_46.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21344 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_48.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_48.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21436 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_50.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 22448 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_52.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 20148 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_54.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_56.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_58.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_58.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5060 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8188 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 6532 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7636 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9292 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 7268 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 6440 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7728 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9936 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 7728 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 6900 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7728 0 -1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9752 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 8004 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 9108 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 13892 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 14536 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 14996 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4_
timestamp 1676037725
transform 1 0 12604 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11592 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11408 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2_
timestamp 1676037725
transform 1 0 9016 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__194 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3_
timestamp 1676037725
transform 1 0 10396 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 10120 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l3_in_1_
timestamp 1676037725
transform 1 0 9108 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l4_in_0_
timestamp 1676037725
transform 1 0 8740 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15824 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 17112 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 15088 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3_
timestamp 1676037725
transform 1 0 15180 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4_
timestamp 1676037725
transform 1 0 14260 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12604 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2_
timestamp 1676037725
transform 1 0 9844 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__195
timestamp 1676037725
transform 1 0 11684 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3_
timestamp 1676037725
transform 1 0 12788 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 10212 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l3_in_1_
timestamp 1676037725
transform 1 0 9200 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l4_in_0_
timestamp 1676037725
transform 1 0 7820 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8924 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15916 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 13800 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3_
timestamp 1676037725
transform 1 0 11868 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4_
timestamp 1676037725
transform 1 0 13340 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12420 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2_
timestamp 1676037725
transform 1 0 10212 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__196
timestamp 1676037725
transform 1 0 15640 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3_
timestamp 1676037725
transform 1 0 14720 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 12696 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l3_in_1_
timestamp 1676037725
transform 1 0 10396 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l4_in_0_
timestamp 1676037725
transform 1 0 9108 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14260 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2_
timestamp 1676037725
transform 1 0 13064 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3_
timestamp 1676037725
transform 1 0 12604 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4_
timestamp 1676037725
transform 1 0 13800 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12144 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11592 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2_
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__197
timestamp 1676037725
transform 1 0 16008 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3_
timestamp 1676037725
transform 1 0 14812 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l3_in_1_
timestamp 1676037725
transform 1 0 10396 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l4_in_0_
timestamp 1676037725
transform 1 0 9476 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8648 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15640 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13248 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10580 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10212 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9384 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 14812 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 12512 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 10304 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 9568 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9384 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 13892 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 11592 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 9384 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 8924 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9108 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 12696 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 10304 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 7544 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 7912 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6624 0 -1 48960
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15916 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10212 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1676037725
transform 1 0 12604 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1676037725
transform 1 0 10212 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1676037725
transform 1 0 12420 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1676037725
transform 1 0 17296 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1676037725
transform 1 0 17204 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1676037725
transform 1 0 19228 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1676037725
transform 1 0 14076 0 -1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1676037725
transform 1 0 14352 0 1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1676037725
transform 1 0 14628 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1676037725
transform 1 0 15364 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1676037725
transform 1 0 20332 0 -1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1676037725
transform 1 0 22172 0 -1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1676037725
transform 1 0 19872 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1676037725
transform 1 0 22080 0 -1 32640
box -38 -48 1050 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35
timestamp 1676037725
transform 1 0 4324 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1676037725
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63
timestamp 1676037725
transform 1 0 6900 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77
timestamp 1676037725
transform 1 0 8188 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1676037725
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1676037725
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1676037725
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 1676037725
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1676037725
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_143
timestamp 1676037725
transform 1 0 14260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_161
timestamp 1676037725
transform 1 0 15916 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1676037725
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1676037725
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_215
timestamp 1676037725
transform 1 0 20884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_243
timestamp 1676037725
transform 1 0 23460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_258 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24840 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_21
timestamp 1676037725
transform 1 0 3036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_35
timestamp 1676037725
transform 1 0 4324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_41
timestamp 1676037725
transform 1 0 4876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1676037725
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 1676037725
transform 1 0 6808 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_83
timestamp 1676037725
transform 1 0 8740 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_91
timestamp 1676037725
transform 1 0 9476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1676037725
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_103
timestamp 1676037725
transform 1 0 10580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1676037725
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_145
timestamp 1676037725
transform 1 0 14444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1676037725
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1676037725
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_207
timestamp 1676037725
transform 1 0 20148 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_211
timestamp 1676037725
transform 1 0 20516 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1676037725
transform 1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1676037725
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_231
timestamp 1676037725
transform 1 0 22356 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_238
timestamp 1676037725
transform 1 0 23000 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_264
timestamp 1676037725
transform 1 0 25392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_22
timestamp 1676037725
transform 1 0 3128 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_33
timestamp 1676037725
transform 1 0 4140 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_37
timestamp 1676037725
transform 1 0 4508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_51
timestamp 1676037725
transform 1 0 5796 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_55
timestamp 1676037725
transform 1 0 6164 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_60
timestamp 1676037725
transform 1 0 6624 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_64
timestamp 1676037725
transform 1 0 6992 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_68
timestamp 1676037725
transform 1 0 7360 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_74
timestamp 1676037725
transform 1 0 7912 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_78
timestamp 1676037725
transform 1 0 8280 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1676037725
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_87
timestamp 1676037725
transform 1 0 9108 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_91
timestamp 1676037725
transform 1 0 9476 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_96
timestamp 1676037725
transform 1 0 9936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_100
timestamp 1676037725
transform 1 0 10304 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_104
timestamp 1676037725
transform 1 0 10672 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_118
timestamp 1676037725
transform 1 0 11960 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1676037725
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_159
timestamp 1676037725
transform 1 0 15732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_179
timestamp 1676037725
transform 1 0 17572 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_186
timestamp 1676037725
transform 1 0 18216 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1676037725
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1676037725
transform 1 0 20884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_235
timestamp 1676037725
transform 1 0 22724 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_242
timestamp 1676037725
transform 1 0 23368 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_246
timestamp 1676037725
transform 1 0 23736 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1676037725
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_262
timestamp 1676037725
transform 1 0 25208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_8
timestamp 1676037725
transform 1 0 1840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_21
timestamp 1676037725
transform 1 0 3036 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_36
timestamp 1676037725
transform 1 0 4416 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_40
timestamp 1676037725
transform 1 0 4784 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1676037725
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_92
timestamp 1676037725
transform 1 0 9568 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_96
timestamp 1676037725
transform 1 0 9936 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_102
timestamp 1676037725
transform 1 0 10488 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1676037725
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_117
timestamp 1676037725
transform 1 0 11868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_135
timestamp 1676037725
transform 1 0 13524 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_159
timestamp 1676037725
transform 1 0 15732 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1676037725
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_187
timestamp 1676037725
transform 1 0 18308 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_207
timestamp 1676037725
transform 1 0 20148 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_220
timestamp 1676037725
transform 1 0 21344 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_243
timestamp 1676037725
transform 1 0 23460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_263
timestamp 1676037725
transform 1 0 25300 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5
timestamp 1676037725
transform 1 0 1564 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_17
timestamp 1676037725
transform 1 0 2668 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1676037725
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_66
timestamp 1676037725
transform 1 0 7176 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_70
timestamp 1676037725
transform 1 0 7544 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1676037725
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_112
timestamp 1676037725
transform 1 0 11408 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_120
timestamp 1676037725
transform 1 0 12144 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_124
timestamp 1676037725
transform 1 0 12512 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1676037725
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_143
timestamp 1676037725
transform 1 0 14260 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1676037725
transform 1 0 14720 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_172
timestamp 1676037725
transform 1 0 16928 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_176
timestamp 1676037725
transform 1 0 17296 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 1676037725
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_220
timestamp 1676037725
transform 1 0 21344 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_240
timestamp 1676037725
transform 1 0 23184 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_248
timestamp 1676037725
transform 1 0 23920 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_259
timestamp 1676037725
transform 1 0 24932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_151
timestamp 1676037725
transform 1 0 14996 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_155
timestamp 1676037725
transform 1 0 15364 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1676037725
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_188
timestamp 1676037725
transform 1 0 18400 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_212
timestamp 1676037725
transform 1 0 20608 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_220
timestamp 1676037725
transform 1 0 21344 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_243
timestamp 1676037725
transform 1 0 23460 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_263
timestamp 1676037725
transform 1 0 25300 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_117
timestamp 1676037725
transform 1 0 11868 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1676037725
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_146
timestamp 1676037725
transform 1 0 14536 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_157
timestamp 1676037725
transform 1 0 15548 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_181
timestamp 1676037725
transform 1 0 17756 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1676037725
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1676037725
transform 1 0 20884 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_235
timestamp 1676037725
transform 1 0 22724 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_243
timestamp 1676037725
transform 1 0 23460 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1676037725
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_259
timestamp 1676037725
transform 1 0 24932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1676037725
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_124
timestamp 1676037725
transform 1 0 12512 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_130
timestamp 1676037725
transform 1 0 13064 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_142
timestamp 1676037725
transform 1 0 14168 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_146
timestamp 1676037725
transform 1 0 14536 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1676037725
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_174
timestamp 1676037725
transform 1 0 17112 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_182
timestamp 1676037725
transform 1 0 17848 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_202
timestamp 1676037725
transform 1 0 19688 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1676037725
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_247
timestamp 1676037725
transform 1 0 23828 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_254
timestamp 1676037725
transform 1 0 24472 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_261
timestamp 1676037725
transform 1 0 25116 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_265
timestamp 1676037725
transform 1 0 25484 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_125
timestamp 1676037725
transform 1 0 12604 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_129
timestamp 1676037725
transform 1 0 12972 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1676037725
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_147
timestamp 1676037725
transform 1 0 14628 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_160
timestamp 1676037725
transform 1 0 15824 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_164
timestamp 1676037725
transform 1 0 16192 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_170
timestamp 1676037725
transform 1 0 16744 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1676037725
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_208
timestamp 1676037725
transform 1 0 20240 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1676037725
transform 1 0 20608 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_230
timestamp 1676037725
transform 1 0 22264 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1676037725
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_264
timestamp 1676037725
transform 1 0 25392 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_85
timestamp 1676037725
transform 1 0 8924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_106
timestamp 1676037725
transform 1 0 10856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1676037725
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_9_130
timestamp 1676037725
transform 1 0 13064 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_136
timestamp 1676037725
transform 1 0 13616 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_157
timestamp 1676037725
transform 1 0 15548 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1676037725
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_171
timestamp 1676037725
transform 1 0 16836 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_174
timestamp 1676037725
transform 1 0 17112 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_185
timestamp 1676037725
transform 1 0 18124 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_209
timestamp 1676037725
transform 1 0 20332 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1676037725
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_244
timestamp 1676037725
transform 1 0 23552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1676037725
transform 1 0 25392 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_105
timestamp 1676037725
transform 1 0 10764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_117
timestamp 1676037725
transform 1 0 11868 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_125
timestamp 1676037725
transform 1 0 12604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1676037725
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_152
timestamp 1676037725
transform 1 0 15088 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_169
timestamp 1676037725
transform 1 0 16652 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1676037725
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_202
timestamp 1676037725
transform 1 0 19688 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_206
timestamp 1676037725
transform 1 0 20056 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_224
timestamp 1676037725
transform 1 0 21712 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_248
timestamp 1676037725
transform 1 0 23920 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_259
timestamp 1676037725
transform 1 0 24932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_118
timestamp 1676037725
transform 1 0 11960 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_130
timestamp 1676037725
transform 1 0 13064 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_134
timestamp 1676037725
transform 1 0 13432 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_142
timestamp 1676037725
transform 1 0 14168 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_148
timestamp 1676037725
transform 1 0 14720 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_159
timestamp 1676037725
transform 1 0 15732 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1676037725
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_180
timestamp 1676037725
transform 1 0 17664 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_184
timestamp 1676037725
transform 1 0 18032 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_202
timestamp 1676037725
transform 1 0 19688 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1676037725
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_244
timestamp 1676037725
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_264
timestamp 1676037725
transform 1 0 25392 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_107
timestamp 1676037725
transform 1 0 10948 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_111
timestamp 1676037725
transform 1 0 11316 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_123
timestamp 1676037725
transform 1 0 12420 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1676037725
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_152
timestamp 1676037725
transform 1 0 15088 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_160
timestamp 1676037725
transform 1 0 15824 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_170
timestamp 1676037725
transform 1 0 16744 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_183
timestamp 1676037725
transform 1 0 17940 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_189
timestamp 1676037725
transform 1 0 18492 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_228
timestamp 1676037725
transform 1 0 22080 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_232
timestamp 1676037725
transform 1 0 22448 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1676037725
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_258
timestamp 1676037725
transform 1 0 24840 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_109
timestamp 1676037725
transform 1 0 11132 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_135
timestamp 1676037725
transform 1 0 13524 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_148
timestamp 1676037725
transform 1 0 14720 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1676037725
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_175
timestamp 1676037725
transform 1 0 17204 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_196
timestamp 1676037725
transform 1 0 19136 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_200
timestamp 1676037725
transform 1 0 19504 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1676037725
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_230
timestamp 1676037725
transform 1 0 22264 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_254
timestamp 1676037725
transform 1 0 24472 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_261
timestamp 1676037725
transform 1 0 25116 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_265
timestamp 1676037725
transform 1 0 25484 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_110
timestamp 1676037725
transform 1 0 11224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_123
timestamp 1676037725
transform 1 0 12420 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_136
timestamp 1676037725
transform 1 0 13616 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 1676037725
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_155
timestamp 1676037725
transform 1 0 15364 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_166
timestamp 1676037725
transform 1 0 16376 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_174
timestamp 1676037725
transform 1 0 17112 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_182
timestamp 1676037725
transform 1 0 17848 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_192
timestamp 1676037725
transform 1 0 18768 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_203
timestamp 1676037725
transform 1 0 19780 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_209
timestamp 1676037725
transform 1 0 20332 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_231
timestamp 1676037725
transform 1 0 22356 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_235
timestamp 1676037725
transform 1 0 22724 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1676037725
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1676037725
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_258
timestamp 1676037725
transform 1 0 24840 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_98
timestamp 1676037725
transform 1 0 10120 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_102
timestamp 1676037725
transform 1 0 10488 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_106
timestamp 1676037725
transform 1 0 10856 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1676037725
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1676037725
transform 1 0 11960 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_131
timestamp 1676037725
transform 1 0 13156 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_137
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_147
timestamp 1676037725
transform 1 0 14628 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_155
timestamp 1676037725
transform 1 0 15364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_174
timestamp 1676037725
transform 1 0 17112 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_182
timestamp 1676037725
transform 1 0 17848 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_189
timestamp 1676037725
transform 1 0 18492 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_196
timestamp 1676037725
transform 1 0 19136 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_209
timestamp 1676037725
transform 1 0 20332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1676037725
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_230
timestamp 1676037725
transform 1 0 22264 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_234
timestamp 1676037725
transform 1 0 22632 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_238
timestamp 1676037725
transform 1 0 23000 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_259
timestamp 1676037725
transform 1 0 24932 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_263
timestamp 1676037725
transform 1 0 25300 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_107
timestamp 1676037725
transform 1 0 10948 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_111
timestamp 1676037725
transform 1 0 11316 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_134
timestamp 1676037725
transform 1 0 13432 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1676037725
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_146
timestamp 1676037725
transform 1 0 14536 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_170
timestamp 1676037725
transform 1 0 16744 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_174
timestamp 1676037725
transform 1 0 17112 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_182
timestamp 1676037725
transform 1 0 17848 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_199
timestamp 1676037725
transform 1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_210
timestamp 1676037725
transform 1 0 20424 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_218
timestamp 1676037725
transform 1 0 21160 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_225
timestamp 1676037725
transform 1 0 21804 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_229
timestamp 1676037725
transform 1 0 22172 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_233
timestamp 1676037725
transform 1 0 22540 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1676037725
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_259
timestamp 1676037725
transform 1 0 24932 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_263
timestamp 1676037725
transform 1 0 25300 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_65
timestamp 1676037725
transform 1 0 7084 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_87
timestamp 1676037725
transform 1 0 9108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_104
timestamp 1676037725
transform 1 0 10672 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_126
timestamp 1676037725
transform 1 0 12696 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_139
timestamp 1676037725
transform 1 0 13892 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_152
timestamp 1676037725
transform 1 0 15088 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1676037725
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_180
timestamp 1676037725
transform 1 0 17664 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_193
timestamp 1676037725
transform 1 0 18860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_201
timestamp 1676037725
transform 1 0 19596 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_209
timestamp 1676037725
transform 1 0 20332 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_216
timestamp 1676037725
transform 1 0 20976 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1676037725
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_244
timestamp 1676037725
transform 1 0 23552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_264
timestamp 1676037725
transform 1 0 25392 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_71
timestamp 1676037725
transform 1 0 7636 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1676037725
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_108
timestamp 1676037725
transform 1 0 11040 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_134
timestamp 1676037725
transform 1 0 13432 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_152
timestamp 1676037725
transform 1 0 15088 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_164
timestamp 1676037725
transform 1 0 16192 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_167
timestamp 1676037725
transform 1 0 16468 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_172
timestamp 1676037725
transform 1 0 16928 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_187
timestamp 1676037725
transform 1 0 18308 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_203
timestamp 1676037725
transform 1 0 19780 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_207
timestamp 1676037725
transform 1 0 20148 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_230
timestamp 1676037725
transform 1 0 22264 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_258
timestamp 1676037725
transform 1 0 24840 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_82
timestamp 1676037725
transform 1 0 8648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_95
timestamp 1676037725
transform 1 0 9844 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1676037725
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1676037725
transform 1 0 12420 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_134
timestamp 1676037725
transform 1 0 13432 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_147
timestamp 1676037725
transform 1 0 14628 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_160
timestamp 1676037725
transform 1 0 15824 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1676037725
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_180
timestamp 1676037725
transform 1 0 17664 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_187
timestamp 1676037725
transform 1 0 18308 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_191
timestamp 1676037725
transform 1 0 18676 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_201
timestamp 1676037725
transform 1 0 19596 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_208
timestamp 1676037725
transform 1 0 20240 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_212
timestamp 1676037725
transform 1 0 20608 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_230
timestamp 1676037725
transform 1 0 22264 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_236
timestamp 1676037725
transform 1 0 22816 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_259
timestamp 1676037725
transform 1 0 24932 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_263
timestamp 1676037725
transform 1 0 25300 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_79
timestamp 1676037725
transform 1 0 8372 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_121
timestamp 1676037725
transform 1 0 12236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_136
timestamp 1676037725
transform 1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_149
timestamp 1676037725
transform 1 0 14812 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_162
timestamp 1676037725
transform 1 0 16008 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_166
timestamp 1676037725
transform 1 0 16376 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_174
timestamp 1676037725
transform 1 0 17112 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_179
timestamp 1676037725
transform 1 0 17572 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_185
timestamp 1676037725
transform 1 0 18124 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1676037725
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_210
timestamp 1676037725
transform 1 0 20424 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_214
timestamp 1676037725
transform 1 0 20792 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_230
timestamp 1676037725
transform 1 0 22264 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_258
timestamp 1676037725
transform 1 0 24840 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_262
timestamp 1676037725
transform 1 0 25208 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1676037725
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1676037725
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1676037725
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_95
timestamp 1676037725
transform 1 0 9844 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1676037725
transform 1 0 11960 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_122
timestamp 1676037725
transform 1 0 12328 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_134
timestamp 1676037725
transform 1 0 13432 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_158
timestamp 1676037725
transform 1 0 15640 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_162
timestamp 1676037725
transform 1 0 16008 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_191
timestamp 1676037725
transform 1 0 18676 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_197
timestamp 1676037725
transform 1 0 19228 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_203
timestamp 1676037725
transform 1 0 19780 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_210
timestamp 1676037725
transform 1 0 20424 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_214
timestamp 1676037725
transform 1 0 20792 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_218
timestamp 1676037725
transform 1 0 21160 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_230
timestamp 1676037725
transform 1 0 22264 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_256
timestamp 1676037725
transform 1 0 24656 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_263
timestamp 1676037725
transform 1 0 25300 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_57
timestamp 1676037725
transform 1 0 6348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_78
timestamp 1676037725
transform 1 0 8280 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1676037725
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1676037725
transform 1 0 9476 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_94
timestamp 1676037725
transform 1 0 9752 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_119
timestamp 1676037725
transform 1 0 12052 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_132
timestamp 1676037725
transform 1 0 13248 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1676037725
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_152
timestamp 1676037725
transform 1 0 15088 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_156
timestamp 1676037725
transform 1 0 15456 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_164
timestamp 1676037725
transform 1 0 16192 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_176
timestamp 1676037725
transform 1 0 17296 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_183
timestamp 1676037725
transform 1 0 17940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1676037725
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_205
timestamp 1676037725
transform 1 0 19964 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_211
timestamp 1676037725
transform 1 0 20516 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_219
timestamp 1676037725
transform 1 0 21252 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_230
timestamp 1676037725
transform 1 0 22264 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_257
timestamp 1676037725
transform 1 0 24748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_261
timestamp 1676037725
transform 1 0 25116 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_265
timestamp 1676037725
transform 1 0 25484 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_94
timestamp 1676037725
transform 1 0 9752 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_107
timestamp 1676037725
transform 1 0 10948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1676037725
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_121
timestamp 1676037725
transform 1 0 12236 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_133
timestamp 1676037725
transform 1 0 13340 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_146
timestamp 1676037725
transform 1 0 14536 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_154
timestamp 1676037725
transform 1 0 15272 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_181
timestamp 1676037725
transform 1 0 17756 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_189
timestamp 1676037725
transform 1 0 18492 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_194
timestamp 1676037725
transform 1 0 18952 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_200
timestamp 1676037725
transform 1 0 19504 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_210
timestamp 1676037725
transform 1 0 20424 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_217
timestamp 1676037725
transform 1 0 21068 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_221
timestamp 1676037725
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_244
timestamp 1676037725
transform 1 0 23552 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_264
timestamp 1676037725
transform 1 0 25392 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_96
timestamp 1676037725
transform 1 0 9936 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_100
timestamp 1676037725
transform 1 0 10304 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_112
timestamp 1676037725
transform 1 0 11408 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_123
timestamp 1676037725
transform 1 0 12420 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_135
timestamp 1676037725
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1676037725
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_146
timestamp 1676037725
transform 1 0 14536 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_158
timestamp 1676037725
transform 1 0 15640 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_162
timestamp 1676037725
transform 1 0 16008 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_186
timestamp 1676037725
transform 1 0 18216 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_190
timestamp 1676037725
transform 1 0 18584 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_219
timestamp 1676037725
transform 1 0 21252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_226
timestamp 1676037725
transform 1 0 21896 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1676037725
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_258
timestamp 1676037725
transform 1 0 24840 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_262
timestamp 1676037725
transform 1 0 25208 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1676037725
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1676037725
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1676037725
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_79
timestamp 1676037725
transform 1 0 8372 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_83
timestamp 1676037725
transform 1 0 8740 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_95
timestamp 1676037725
transform 1 0 9844 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_107
timestamp 1676037725
transform 1 0 10948 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_119
timestamp 1676037725
transform 1 0 12052 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_129
timestamp 1676037725
transform 1 0 12972 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_142
timestamp 1676037725
transform 1 0 14168 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_155
timestamp 1676037725
transform 1 0 15364 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_162
timestamp 1676037725
transform 1 0 16008 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_172
timestamp 1676037725
transform 1 0 16928 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_178
timestamp 1676037725
transform 1 0 17480 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_185
timestamp 1676037725
transform 1 0 18124 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_192
timestamp 1676037725
transform 1 0 18768 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_196
timestamp 1676037725
transform 1 0 19136 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_208
timestamp 1676037725
transform 1 0 20240 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_212
timestamp 1676037725
transform 1 0 20608 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1676037725
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_247
timestamp 1676037725
transform 1 0 23828 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_251
timestamp 1676037725
transform 1 0 24196 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_264
timestamp 1676037725
transform 1 0 25392 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1676037725
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1676037725
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1676037725
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1676037725
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_108
timestamp 1676037725
transform 1 0 11040 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_136
timestamp 1676037725
transform 1 0 13616 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_144
timestamp 1676037725
transform 1 0 14352 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_155
timestamp 1676037725
transform 1 0 15364 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_168
timestamp 1676037725
transform 1 0 16560 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_173
timestamp 1676037725
transform 1 0 17020 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_186
timestamp 1676037725
transform 1 0 18216 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_190
timestamp 1676037725
transform 1 0 18584 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_199
timestamp 1676037725
transform 1 0 19412 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_204
timestamp 1676037725
transform 1 0 19872 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_228
timestamp 1676037725
transform 1 0 22080 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_232
timestamp 1676037725
transform 1 0 22448 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1676037725
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_258
timestamp 1676037725
transform 1 0 24840 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1676037725
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1676037725
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_80
timestamp 1676037725
transform 1 0 8464 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_95
timestamp 1676037725
transform 1 0 9844 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1676037725
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_115
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_119
timestamp 1676037725
transform 1 0 12052 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_136
timestamp 1676037725
transform 1 0 13616 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_144
timestamp 1676037725
transform 1 0 14352 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_175
timestamp 1676037725
transform 1 0 17204 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_179
timestamp 1676037725
transform 1 0 17572 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_186
timestamp 1676037725
transform 1 0 18216 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_210
timestamp 1676037725
transform 1 0 20424 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_214
timestamp 1676037725
transform 1 0 20792 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_218
timestamp 1676037725
transform 1 0 21160 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_229
timestamp 1676037725
transform 1 0 22172 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_239
timestamp 1676037725
transform 1 0 23092 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_264
timestamp 1676037725
transform 1 0 25392 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_69
timestamp 1676037725
transform 1 0 7452 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1676037725
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_90
timestamp 1676037725
transform 1 0 9384 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_117
timestamp 1676037725
transform 1 0 11868 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_130
timestamp 1676037725
transform 1 0 13064 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1676037725
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_153
timestamp 1676037725
transform 1 0 15180 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_162
timestamp 1676037725
transform 1 0 16008 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_168
timestamp 1676037725
transform 1 0 16560 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_181
timestamp 1676037725
transform 1 0 17756 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1676037725
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_201
timestamp 1676037725
transform 1 0 19596 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_206
timestamp 1676037725
transform 1 0 20056 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_217
timestamp 1676037725
transform 1 0 21068 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_225
timestamp 1676037725
transform 1 0 21804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_230
timestamp 1676037725
transform 1 0 22264 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_264
timestamp 1676037725
transform 1 0 25392 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1676037725
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1676037725
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1676037725
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_92
timestamp 1676037725
transform 1 0 9568 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_109
timestamp 1676037725
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_121
timestamp 1676037725
transform 1 0 12236 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_134
timestamp 1676037725
transform 1 0 13432 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_147
timestamp 1676037725
transform 1 0 14628 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_151
timestamp 1676037725
transform 1 0 14996 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1676037725
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_191
timestamp 1676037725
transform 1 0 18676 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_195
timestamp 1676037725
transform 1 0 19044 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_207
timestamp 1676037725
transform 1 0 20148 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_215
timestamp 1676037725
transform 1 0 20884 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1676037725
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_244
timestamp 1676037725
transform 1 0 23552 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_264
timestamp 1676037725
transform 1 0 25392 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1676037725
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_59
timestamp 1676037725
transform 1 0 6532 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_80
timestamp 1676037725
transform 1 0 8464 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_95
timestamp 1676037725
transform 1 0 9844 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_106
timestamp 1676037725
transform 1 0 10856 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_112
timestamp 1676037725
transform 1 0 11408 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_122
timestamp 1676037725
transform 1 0 12328 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_135
timestamp 1676037725
transform 1 0 13524 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_146
timestamp 1676037725
transform 1 0 14536 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_158
timestamp 1676037725
transform 1 0 15640 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_170
timestamp 1676037725
transform 1 0 16744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_180
timestamp 1676037725
transform 1 0 17664 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_186
timestamp 1676037725
transform 1 0 18216 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1676037725
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_209
timestamp 1676037725
transform 1 0 20332 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_217
timestamp 1676037725
transform 1 0 21068 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_222
timestamp 1676037725
transform 1 0 21528 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_226
timestamp 1676037725
transform 1 0 21896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_230
timestamp 1676037725
transform 1 0 22264 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_259
timestamp 1676037725
transform 1 0 24932 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_265
timestamp 1676037725
transform 1 0 25484 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1676037725
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1676037725
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1676037725
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_79
timestamp 1676037725
transform 1 0 8372 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_92
timestamp 1676037725
transform 1 0 9568 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_104
timestamp 1676037725
transform 1 0 10672 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1676037725
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_118
timestamp 1676037725
transform 1 0 11960 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_144
timestamp 1676037725
transform 1 0 14352 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_148
timestamp 1676037725
transform 1 0 14720 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_154
timestamp 1676037725
transform 1 0 15272 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_160
timestamp 1676037725
transform 1 0 15824 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1676037725
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_180
timestamp 1676037725
transform 1 0 17664 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_192
timestamp 1676037725
transform 1 0 18768 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_197
timestamp 1676037725
transform 1 0 19228 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_205
timestamp 1676037725
transform 1 0 19964 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1676037725
transform 1 0 20884 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_227
timestamp 1676037725
transform 1 0 21988 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_238
timestamp 1676037725
transform 1 0 23000 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_262
timestamp 1676037725
transform 1 0 25208 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1676037725
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1676037725
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1676037725
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_77
timestamp 1676037725
transform 1 0 8188 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_81
timestamp 1676037725
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_107
timestamp 1676037725
transform 1 0 10948 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_120
timestamp 1676037725
transform 1 0 12144 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_132
timestamp 1676037725
transform 1 0 13248 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_163
timestamp 1676037725
transform 1 0 16100 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_170
timestamp 1676037725
transform 1 0 16744 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_174
timestamp 1676037725
transform 1 0 17112 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_187
timestamp 1676037725
transform 1 0 18308 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1676037725
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_203
timestamp 1676037725
transform 1 0 19780 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_224
timestamp 1676037725
transform 1 0 21712 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_248
timestamp 1676037725
transform 1 0 23920 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_255
timestamp 1676037725
transform 1 0 24564 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_263
timestamp 1676037725
transform 1 0 25300 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1676037725
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1676037725
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1676037725
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1676037725
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_95
timestamp 1676037725
transform 1 0 9844 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_99
timestamp 1676037725
transform 1 0 10212 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1676037725
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_125
timestamp 1676037725
transform 1 0 12604 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_146
timestamp 1676037725
transform 1 0 14536 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_150
timestamp 1676037725
transform 1 0 14904 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_160
timestamp 1676037725
transform 1 0 15824 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_191
timestamp 1676037725
transform 1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_198
timestamp 1676037725
transform 1 0 19320 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_205
timestamp 1676037725
transform 1 0 19964 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_209
timestamp 1676037725
transform 1 0 20332 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_219
timestamp 1676037725
transform 1 0 21252 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1676037725
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_230
timestamp 1676037725
transform 1 0 22264 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_234
timestamp 1676037725
transform 1 0 22632 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_238
timestamp 1676037725
transform 1 0 23000 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_264
timestamp 1676037725
transform 1 0 25392 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1676037725
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1676037725
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1676037725
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1676037725
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1676037725
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1676037725
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_88
timestamp 1676037725
transform 1 0 9200 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_99
timestamp 1676037725
transform 1 0 10212 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_103
timestamp 1676037725
transform 1 0 10580 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_124
timestamp 1676037725
transform 1 0 12512 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_128
timestamp 1676037725
transform 1 0 12880 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_145
timestamp 1676037725
transform 1 0 14444 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_148
timestamp 1676037725
transform 1 0 14720 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_152
timestamp 1676037725
transform 1 0 15088 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_173
timestamp 1676037725
transform 1 0 17020 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1676037725
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_189
timestamp 1676037725
transform 1 0 18492 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_193
timestamp 1676037725
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_208
timestamp 1676037725
transform 1 0 20240 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_212
timestamp 1676037725
transform 1 0 20608 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_217
timestamp 1676037725
transform 1 0 21068 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_223
timestamp 1676037725
transform 1 0 21620 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_230
timestamp 1676037725
transform 1 0 22264 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1676037725
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_264
timestamp 1676037725
transform 1 0 25392 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1676037725
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1676037725
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1676037725
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1676037725
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_83
timestamp 1676037725
transform 1 0 8740 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_87
timestamp 1676037725
transform 1 0 9108 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_97
timestamp 1676037725
transform 1 0 10028 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1676037725
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_118
timestamp 1676037725
transform 1 0 11960 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_150
timestamp 1676037725
transform 1 0 14904 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_154
timestamp 1676037725
transform 1 0 15272 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1676037725
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1676037725
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_181
timestamp 1676037725
transform 1 0 17756 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_189
timestamp 1676037725
transform 1 0 18492 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_194
timestamp 1676037725
transform 1 0 18952 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_198
timestamp 1676037725
transform 1 0 19320 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_209
timestamp 1676037725
transform 1 0 20332 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_216
timestamp 1676037725
transform 1 0 20976 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_236
timestamp 1676037725
transform 1 0 22816 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_240
timestamp 1676037725
transform 1 0 23184 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_261
timestamp 1676037725
transform 1 0 25116 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_265
timestamp 1676037725
transform 1 0 25484 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1676037725
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1676037725
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1676037725
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1676037725
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1676037725
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_87
timestamp 1676037725
transform 1 0 9108 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_99
timestamp 1676037725
transform 1 0 10212 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_102
timestamp 1676037725
transform 1 0 10488 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_113
timestamp 1676037725
transform 1 0 11500 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_117
timestamp 1676037725
transform 1 0 11868 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_127
timestamp 1676037725
transform 1 0 12788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1676037725
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_158
timestamp 1676037725
transform 1 0 15640 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_162
timestamp 1676037725
transform 1 0 16008 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_183
timestamp 1676037725
transform 1 0 17940 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_187
timestamp 1676037725
transform 1 0 18308 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1676037725
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_201
timestamp 1676037725
transform 1 0 19596 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_211
timestamp 1676037725
transform 1 0 20516 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_218
timestamp 1676037725
transform 1 0 21160 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_242
timestamp 1676037725
transform 1 0 23368 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_249
timestamp 1676037725
transform 1 0 24012 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_264
timestamp 1676037725
transform 1 0 25392 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1676037725
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1676037725
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1676037725
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1676037725
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1676037725
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_69
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_75
timestamp 1676037725
transform 1 0 8004 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_96
timestamp 1676037725
transform 1 0 9936 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_100
timestamp 1676037725
transform 1 0 10304 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_121
timestamp 1676037725
transform 1 0 12236 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_142
timestamp 1676037725
transform 1 0 14168 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_146
timestamp 1676037725
transform 1 0 14536 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_158
timestamp 1676037725
transform 1 0 15640 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1676037725
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_174
timestamp 1676037725
transform 1 0 17112 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_186
timestamp 1676037725
transform 1 0 18216 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_190
timestamp 1676037725
transform 1 0 18584 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_195
timestamp 1676037725
transform 1 0 19044 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_201
timestamp 1676037725
transform 1 0 19596 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_205
timestamp 1676037725
transform 1 0 19964 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_211
timestamp 1676037725
transform 1 0 20516 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1676037725
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_244
timestamp 1676037725
transform 1 0 23552 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_264
timestamp 1676037725
transform 1 0 25392 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1676037725
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1676037725
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1676037725
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1676037725
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1676037725
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1676037725
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_96
timestamp 1676037725
transform 1 0 9936 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_108
timestamp 1676037725
transform 1 0 11040 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_119
timestamp 1676037725
transform 1 0 12052 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_127
timestamp 1676037725
transform 1 0 12788 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1676037725
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_145
timestamp 1676037725
transform 1 0 14444 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_157
timestamp 1676037725
transform 1 0 15548 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_161
timestamp 1676037725
transform 1 0 15916 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_173
timestamp 1676037725
transform 1 0 17020 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_181
timestamp 1676037725
transform 1 0 17756 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_191
timestamp 1676037725
transform 1 0 18676 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1676037725
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_209
timestamp 1676037725
transform 1 0 20332 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_216
timestamp 1676037725
transform 1 0 20976 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_222
timestamp 1676037725
transform 1 0 21528 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_226
timestamp 1676037725
transform 1 0 21896 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1676037725
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_264
timestamp 1676037725
transform 1 0 25392 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1676037725
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1676037725
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1676037725
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1676037725
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1676037725
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_69
timestamp 1676037725
transform 1 0 7452 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_95
timestamp 1676037725
transform 1 0 9844 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_99
timestamp 1676037725
transform 1 0 10212 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1676037725
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_125
timestamp 1676037725
transform 1 0 12604 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_131
timestamp 1676037725
transform 1 0 13156 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_141
timestamp 1676037725
transform 1 0 14076 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_154
timestamp 1676037725
transform 1 0 15272 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1676037725
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1676037725
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_180
timestamp 1676037725
transform 1 0 17664 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_187
timestamp 1676037725
transform 1 0 18308 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_195
timestamp 1676037725
transform 1 0 19044 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_206
timestamp 1676037725
transform 1 0 20056 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_219
timestamp 1676037725
transform 1 0 21252 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1676037725
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_232
timestamp 1676037725
transform 1 0 22448 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_260
timestamp 1676037725
transform 1 0 25024 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1676037725
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1676037725
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1676037725
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1676037725
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1676037725
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1676037725
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1676037725
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_107
timestamp 1676037725
transform 1 0 10948 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_114
timestamp 1676037725
transform 1 0 11592 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1676037725
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_143
timestamp 1676037725
transform 1 0 14260 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_155
timestamp 1676037725
transform 1 0 15364 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_181
timestamp 1676037725
transform 1 0 17756 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1676037725
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_219
timestamp 1676037725
transform 1 0 21252 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_224
timestamp 1676037725
transform 1 0 21712 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_246
timestamp 1676037725
transform 1 0 23736 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1676037725
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_258
timestamp 1676037725
transform 1 0 24840 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1676037725
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1676037725
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1676037725
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1676037725
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1676037725
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1676037725
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_81
timestamp 1676037725
transform 1 0 8556 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_89
timestamp 1676037725
transform 1 0 9292 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1676037725
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_124
timestamp 1676037725
transform 1 0 12512 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_128
timestamp 1676037725
transform 1 0 12880 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_149
timestamp 1676037725
transform 1 0 14812 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_153
timestamp 1676037725
transform 1 0 15180 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_156
timestamp 1676037725
transform 1 0 15456 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_180
timestamp 1676037725
transform 1 0 17664 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_193
timestamp 1676037725
transform 1 0 18860 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_199
timestamp 1676037725
transform 1 0 19412 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1676037725
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_237
timestamp 1676037725
transform 1 0 22908 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_243
timestamp 1676037725
transform 1 0 23460 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_264
timestamp 1676037725
transform 1 0 25392 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1676037725
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1676037725
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1676037725
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1676037725
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1676037725
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1676037725
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1676037725
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_97
timestamp 1676037725
transform 1 0 10028 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_105
timestamp 1676037725
transform 1 0 10764 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_126
timestamp 1676037725
transform 1 0 12696 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_130
timestamp 1676037725
transform 1 0 13064 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1676037725
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_152
timestamp 1676037725
transform 1 0 15088 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_156
timestamp 1676037725
transform 1 0 15456 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_168
timestamp 1676037725
transform 1 0 16560 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_175
timestamp 1676037725
transform 1 0 17204 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_182
timestamp 1676037725
transform 1 0 17848 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_188
timestamp 1676037725
transform 1 0 18400 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1676037725
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_199
timestamp 1676037725
transform 1 0 19412 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_206
timestamp 1676037725
transform 1 0 20056 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_210
timestamp 1676037725
transform 1 0 20424 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_217
timestamp 1676037725
transform 1 0 21068 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_221
timestamp 1676037725
transform 1 0 21436 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_225
timestamp 1676037725
transform 1 0 21804 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_233
timestamp 1676037725
transform 1 0 22540 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1676037725
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_259
timestamp 1676037725
transform 1 0 24932 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_264
timestamp 1676037725
transform 1 0 25392 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1676037725
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1676037725
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1676037725
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1676037725
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1676037725
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1676037725
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1676037725
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1676037725
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1676037725
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1676037725
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_119
timestamp 1676037725
transform 1 0 12052 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_129
timestamp 1676037725
transform 1 0 12972 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_144
timestamp 1676037725
transform 1 0 14352 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_148
timestamp 1676037725
transform 1 0 14720 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_158
timestamp 1676037725
transform 1 0 15640 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_165
timestamp 1676037725
transform 1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_174
timestamp 1676037725
transform 1 0 17112 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_178
timestamp 1676037725
transform 1 0 17480 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_190
timestamp 1676037725
transform 1 0 18584 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_194
timestamp 1676037725
transform 1 0 18952 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_197
timestamp 1676037725
transform 1 0 19228 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_209
timestamp 1676037725
transform 1 0 20332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_221
timestamp 1676037725
transform 1 0 21436 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_236
timestamp 1676037725
transform 1 0 22816 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_240
timestamp 1676037725
transform 1 0 23184 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_244
timestamp 1676037725
transform 1 0 23552 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_264
timestamp 1676037725
transform 1 0 25392 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1676037725
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1676037725
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1676037725
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1676037725
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1676037725
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1676037725
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1676037725
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_107
timestamp 1676037725
transform 1 0 10948 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_111
timestamp 1676037725
transform 1 0 11316 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_123
timestamp 1676037725
transform 1 0 12420 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_135
timestamp 1676037725
transform 1 0 13524 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1676037725
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_152
timestamp 1676037725
transform 1 0 15088 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_156
timestamp 1676037725
transform 1 0 15456 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_167
timestamp 1676037725
transform 1 0 16468 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_177
timestamp 1676037725
transform 1 0 17388 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_185
timestamp 1676037725
transform 1 0 18124 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1676037725
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1676037725
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_219
timestamp 1676037725
transform 1 0 21252 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_223
timestamp 1676037725
transform 1 0 21620 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_229
timestamp 1676037725
transform 1 0 22172 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_232
timestamp 1676037725
transform 1 0 22448 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_243
timestamp 1676037725
transform 1 0 23460 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1676037725
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_264
timestamp 1676037725
transform 1 0 25392 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1676037725
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1676037725
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1676037725
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1676037725
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1676037725
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1676037725
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_81
timestamp 1676037725
transform 1 0 8556 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_109
timestamp 1676037725
transform 1 0 11132 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_115
timestamp 1676037725
transform 1 0 11684 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_127
timestamp 1676037725
transform 1 0 12788 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_150
timestamp 1676037725
transform 1 0 14904 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_163
timestamp 1676037725
transform 1 0 16100 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1676037725
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_181
timestamp 1676037725
transform 1 0 17756 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_203
timestamp 1676037725
transform 1 0 19780 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_207
timestamp 1676037725
transform 1 0 20148 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_219
timestamp 1676037725
transform 1 0 21252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1676037725
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_227
timestamp 1676037725
transform 1 0 21988 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_240
timestamp 1676037725
transform 1 0 23184 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_264
timestamp 1676037725
transform 1 0 25392 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1676037725
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1676037725
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1676037725
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1676037725
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1676037725
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1676037725
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1676037725
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_97
timestamp 1676037725
transform 1 0 10028 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_101
timestamp 1676037725
transform 1 0 10396 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_122
timestamp 1676037725
transform 1 0 12328 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_126
timestamp 1676037725
transform 1 0 12696 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1676037725
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_162
timestamp 1676037725
transform 1 0 16008 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_168
timestamp 1676037725
transform 1 0 16560 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_176
timestamp 1676037725
transform 1 0 17296 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_187
timestamp 1676037725
transform 1 0 18308 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1676037725
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_203
timestamp 1676037725
transform 1 0 19780 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_224
timestamp 1676037725
transform 1 0 21712 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_248
timestamp 1676037725
transform 1 0 23920 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_264
timestamp 1676037725
transform 1 0 25392 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1676037725
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1676037725
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1676037725
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1676037725
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1676037725
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1676037725
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1676037725
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1676037725
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_105
timestamp 1676037725
transform 1 0 10764 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_109
timestamp 1676037725
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_135
timestamp 1676037725
transform 1 0 13524 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_139
timestamp 1676037725
transform 1 0 13892 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_151
timestamp 1676037725
transform 1 0 14996 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_162
timestamp 1676037725
transform 1 0 16008 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_180
timestamp 1676037725
transform 1 0 17664 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_187
timestamp 1676037725
transform 1 0 18308 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_193
timestamp 1676037725
transform 1 0 18860 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_196
timestamp 1676037725
transform 1 0 19136 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_200
timestamp 1676037725
transform 1 0 19504 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_205
timestamp 1676037725
transform 1 0 19964 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_220
timestamp 1676037725
transform 1 0 21344 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_236
timestamp 1676037725
transform 1 0 22816 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_260
timestamp 1676037725
transform 1 0 25024 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1676037725
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1676037725
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1676037725
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1676037725
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1676037725
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1676037725
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1676037725
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_107
timestamp 1676037725
transform 1 0 10948 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_111
timestamp 1676037725
transform 1 0 11316 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_132
timestamp 1676037725
transform 1 0 13248 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_136
timestamp 1676037725
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_158
timestamp 1676037725
transform 1 0 15640 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_166
timestamp 1676037725
transform 1 0 16376 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1676037725
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_208
timestamp 1676037725
transform 1 0 20240 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_232
timestamp 1676037725
transform 1 0 22448 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_245
timestamp 1676037725
transform 1 0 23644 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1676037725
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_264
timestamp 1676037725
transform 1 0 25392 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1676037725
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1676037725
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1676037725
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1676037725
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1676037725
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_81
timestamp 1676037725
transform 1 0 8556 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_89
timestamp 1676037725
transform 1 0 9292 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_100
timestamp 1676037725
transform 1 0 10304 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_119
timestamp 1676037725
transform 1 0 12052 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_129
timestamp 1676037725
transform 1 0 12972 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_153
timestamp 1676037725
transform 1 0 15180 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_166
timestamp 1676037725
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_180
timestamp 1676037725
transform 1 0 17664 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_186
timestamp 1676037725
transform 1 0 18216 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_201
timestamp 1676037725
transform 1 0 19596 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_207
timestamp 1676037725
transform 1 0 20148 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_219
timestamp 1676037725
transform 1 0 21252 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1676037725
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_227
timestamp 1676037725
transform 1 0 21988 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_240
timestamp 1676037725
transform 1 0 23184 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_253
timestamp 1676037725
transform 1 0 24380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_260
timestamp 1676037725
transform 1 0 25024 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1676037725
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1676037725
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1676037725
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1676037725
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1676037725
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1676037725
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1676037725
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1676037725
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_129
timestamp 1676037725
transform 1 0 12972 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_133
timestamp 1676037725
transform 1 0 13340 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1676037725
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_162
timestamp 1676037725
transform 1 0 16008 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_168
timestamp 1676037725
transform 1 0 16560 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_172
timestamp 1676037725
transform 1 0 16928 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_193
timestamp 1676037725
transform 1 0 18860 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_202
timestamp 1676037725
transform 1 0 19688 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_206
timestamp 1676037725
transform 1 0 20056 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_216
timestamp 1676037725
transform 1 0 20976 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_228
timestamp 1676037725
transform 1 0 22080 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_238
timestamp 1676037725
transform 1 0 23000 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_243
timestamp 1676037725
transform 1 0 23460 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_250
timestamp 1676037725
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_255
timestamp 1676037725
transform 1 0 24564 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_264
timestamp 1676037725
transform 1 0 25392 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1676037725
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1676037725
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1676037725
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1676037725
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1676037725
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1676037725
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_81
timestamp 1676037725
transform 1 0 8556 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_88
timestamp 1676037725
transform 1 0 9200 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_100
timestamp 1676037725
transform 1 0 10304 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_136
timestamp 1676037725
transform 1 0 13616 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_140
timestamp 1676037725
transform 1 0 13984 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_152
timestamp 1676037725
transform 1 0 15088 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_165
timestamp 1676037725
transform 1 0 16284 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_173
timestamp 1676037725
transform 1 0 17020 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_185
timestamp 1676037725
transform 1 0 18124 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_51_195
timestamp 1676037725
transform 1 0 19044 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_203
timestamp 1676037725
transform 1 0 19780 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_213
timestamp 1676037725
transform 1 0 20700 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1676037725
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_236
timestamp 1676037725
transform 1 0 22816 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_240
timestamp 1676037725
transform 1 0 23184 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_261
timestamp 1676037725
transform 1 0 25116 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_265
timestamp 1676037725
transform 1 0 25484 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1676037725
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1676037725
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1676037725
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1676037725
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1676037725
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1676037725
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1676037725
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_90
timestamp 1676037725
transform 1 0 9384 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_102
timestamp 1676037725
transform 1 0 10488 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_114
timestamp 1676037725
transform 1 0 11592 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_126
timestamp 1676037725
transform 1 0 12696 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1676037725
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_155
timestamp 1676037725
transform 1 0 15364 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_161
timestamp 1676037725
transform 1 0 15916 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_169
timestamp 1676037725
transform 1 0 16652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_190
timestamp 1676037725
transform 1 0 18584 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1676037725
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_205
timestamp 1676037725
transform 1 0 19964 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_209
timestamp 1676037725
transform 1 0 20332 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_233
timestamp 1676037725
transform 1 0 22540 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_237
timestamp 1676037725
transform 1 0 22908 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_249
timestamp 1676037725
transform 1 0 24012 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_258
timestamp 1676037725
transform 1 0 24840 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1676037725
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1676037725
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1676037725
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1676037725
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1676037725
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1676037725
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1676037725
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1676037725
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1676037725
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1676037725
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_125
timestamp 1676037725
transform 1 0 12604 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_154
timestamp 1676037725
transform 1 0 15272 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_158
timestamp 1676037725
transform 1 0 15640 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_53_171
timestamp 1676037725
transform 1 0 16836 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_197
timestamp 1676037725
transform 1 0 19228 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_201
timestamp 1676037725
transform 1 0 19596 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_204
timestamp 1676037725
transform 1 0 19872 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_215
timestamp 1676037725
transform 1 0 20884 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1676037725
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_231
timestamp 1676037725
transform 1 0 22356 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_252
timestamp 1676037725
transform 1 0 24288 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_256
timestamp 1676037725
transform 1 0 24656 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_260
timestamp 1676037725
transform 1 0 25024 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_264
timestamp 1676037725
transform 1 0 25392 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1676037725
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1676037725
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1676037725
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1676037725
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1676037725
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1676037725
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1676037725
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1676037725
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1676037725
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1676037725
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1676037725
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1676037725
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_153
timestamp 1676037725
transform 1 0 15180 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_166
timestamp 1676037725
transform 1 0 16376 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_190
timestamp 1676037725
transform 1 0 18584 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 1676037725
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_219
timestamp 1676037725
transform 1 0 21252 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_232
timestamp 1676037725
transform 1 0 22448 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_236
timestamp 1676037725
transform 1 0 22816 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_247
timestamp 1676037725
transform 1 0 23828 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1676037725
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_259
timestamp 1676037725
transform 1 0 24932 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_264
timestamp 1676037725
transform 1 0 25392 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1676037725
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1676037725
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1676037725
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1676037725
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1676037725
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1676037725
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1676037725
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1676037725
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1676037725
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1676037725
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1676037725
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1676037725
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_149
timestamp 1676037725
transform 1 0 14812 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1676037725
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_171
timestamp 1676037725
transform 1 0 16836 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_183
timestamp 1676037725
transform 1 0 17940 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_215
timestamp 1676037725
transform 1 0 20884 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_219
timestamp 1676037725
transform 1 0 21252 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_225
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_239
timestamp 1676037725
transform 1 0 23092 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_263
timestamp 1676037725
transform 1 0 25300 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1676037725
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1676037725
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1676037725
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1676037725
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1676037725
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1676037725
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1676037725
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1676037725
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1676037725
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1676037725
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1676037725
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_153
timestamp 1676037725
transform 1 0 15180 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_166
timestamp 1676037725
transform 1 0 16376 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_172
timestamp 1676037725
transform 1 0 16928 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_184
timestamp 1676037725
transform 1 0 18032 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_202
timestamp 1676037725
transform 1 0 19688 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_215
timestamp 1676037725
transform 1 0 20884 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_227
timestamp 1676037725
transform 1 0 21988 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1676037725
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_264
timestamp 1676037725
transform 1 0 25392 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1676037725
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1676037725
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1676037725
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1676037725
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1676037725
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1676037725
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1676037725
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1676037725
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1676037725
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1676037725
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1676037725
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1676037725
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1676037725
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1676037725
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1676037725
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1676037725
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_193
timestamp 1676037725
transform 1 0 18860 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_199
timestamp 1676037725
transform 1 0 19412 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_220
timestamp 1676037725
transform 1 0 21344 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_247
timestamp 1676037725
transform 1 0 23828 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_57_256
timestamp 1676037725
transform 1 0 24656 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_259
timestamp 1676037725
transform 1 0 24932 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_264
timestamp 1676037725
transform 1 0 25392 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1676037725
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1676037725
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1676037725
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1676037725
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1676037725
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1676037725
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1676037725
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1676037725
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1676037725
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_85
timestamp 1676037725
transform 1 0 8924 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_90
timestamp 1676037725
transform 1 0 9384 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_102
timestamp 1676037725
transform 1 0 10488 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_114
timestamp 1676037725
transform 1 0 11592 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_126
timestamp 1676037725
transform 1 0 12696 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_138
timestamp 1676037725
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_141
timestamp 1676037725
transform 1 0 14076 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_58_158
timestamp 1676037725
transform 1 0 15640 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_162
timestamp 1676037725
transform 1 0 16008 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_174
timestamp 1676037725
transform 1 0 17112 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_186
timestamp 1676037725
transform 1 0 18216 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_194
timestamp 1676037725
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_197
timestamp 1676037725
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_219
timestamp 1676037725
transform 1 0 21252 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_243
timestamp 1676037725
transform 1 0 23460 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_247
timestamp 1676037725
transform 1 0 23828 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1676037725
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_253
timestamp 1676037725
transform 1 0 24380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_259
timestamp 1676037725
transform 1 0 24932 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_264
timestamp 1676037725
transform 1 0 25392 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1676037725
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1676037725
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1676037725
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1676037725
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1676037725
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1676037725
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1676037725
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1676037725
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1676037725
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1676037725
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1676037725
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1676037725
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1676037725
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1676037725
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1676037725
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1676037725
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1676037725
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1676037725
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1676037725
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1676037725
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1676037725
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1676037725
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_217
timestamp 1676037725
transform 1 0 21068 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_221
timestamp 1676037725
transform 1 0 21436 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1676037725
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1676037725
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_249
timestamp 1676037725
transform 1 0 24012 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_259
timestamp 1676037725
transform 1 0 24932 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_264
timestamp 1676037725
transform 1 0 25392 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1676037725
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1676037725
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1676037725
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1676037725
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1676037725
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1676037725
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1676037725
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1676037725
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1676037725
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1676037725
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1676037725
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1676037725
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1676037725
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1676037725
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1676037725
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1676037725
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1676037725
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1676037725
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1676037725
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1676037725
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1676037725
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1676037725
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1676037725
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_221
timestamp 1676037725
transform 1 0 21436 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_227
timestamp 1676037725
transform 1 0 21988 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_233
timestamp 1676037725
transform 1 0 22540 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_244
timestamp 1676037725
transform 1 0 23552 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_253
timestamp 1676037725
transform 1 0 24380 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_264
timestamp 1676037725
transform 1 0 25392 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1676037725
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1676037725
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1676037725
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1676037725
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1676037725
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1676037725
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1676037725
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1676037725
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_81
timestamp 1676037725
transform 1 0 8556 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_89
timestamp 1676037725
transform 1 0 9292 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_110
timestamp 1676037725
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_115
timestamp 1676037725
transform 1 0 11684 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_127
timestamp 1676037725
transform 1 0 12788 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_139
timestamp 1676037725
transform 1 0 13892 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_151
timestamp 1676037725
transform 1 0 14996 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_163
timestamp 1676037725
transform 1 0 16100 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1676037725
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1676037725
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1676037725
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1676037725
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_205
timestamp 1676037725
transform 1 0 19964 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_211
timestamp 1676037725
transform 1 0 20516 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_222
timestamp 1676037725
transform 1 0 21528 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1676037725
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_236
timestamp 1676037725
transform 1 0 22816 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_248
timestamp 1676037725
transform 1 0 23920 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_260
timestamp 1676037725
transform 1 0 25024 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1676037725
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1676037725
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1676037725
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1676037725
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1676037725
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1676037725
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1676037725
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1676037725
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1676037725
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1676037725
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1676037725
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1676037725
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1676037725
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1676037725
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1676037725
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1676037725
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1676037725
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1676037725
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1676037725
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1676037725
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1676037725
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1676037725
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1676037725
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1676037725
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1676037725
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1676037725
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1676037725
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_253
timestamp 1676037725
transform 1 0 24380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_259
timestamp 1676037725
transform 1 0 24932 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_264
timestamp 1676037725
transform 1 0 25392 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1676037725
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1676037725
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1676037725
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1676037725
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1676037725
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1676037725
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1676037725
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1676037725
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1676037725
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1676037725
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1676037725
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1676037725
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1676037725
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1676037725
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1676037725
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1676037725
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1676037725
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1676037725
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1676037725
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1676037725
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1676037725
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1676037725
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1676037725
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1676037725
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1676037725
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1676037725
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_249
timestamp 1676037725
transform 1 0 24012 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_257
timestamp 1676037725
transform 1 0 24748 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_264
timestamp 1676037725
transform 1 0 25392 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1676037725
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1676037725
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1676037725
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1676037725
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1676037725
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1676037725
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1676037725
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1676037725
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1676037725
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1676037725
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1676037725
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1676037725
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1676037725
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1676037725
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1676037725
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1676037725
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1676037725
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1676037725
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1676037725
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1676037725
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1676037725
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1676037725
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1676037725
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1676037725
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1676037725
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1676037725
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1676037725
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_253
timestamp 1676037725
transform 1 0 24380 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_261
timestamp 1676037725
transform 1 0 25116 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1676037725
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1676037725
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1676037725
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1676037725
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1676037725
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1676037725
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1676037725
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1676037725
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_81
timestamp 1676037725
transform 1 0 8556 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_85
timestamp 1676037725
transform 1 0 8924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_97
timestamp 1676037725
transform 1 0 10028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_109
timestamp 1676037725
transform 1 0 11132 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1676037725
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1676037725
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1676037725
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1676037725
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1676037725
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1676037725
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1676037725
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1676037725
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1676037725
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1676037725
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1676037725
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1676037725
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1676037725
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1676037725
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_249
timestamp 1676037725
transform 1 0 24012 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_255
timestamp 1676037725
transform 1 0 24564 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_258
timestamp 1676037725
transform 1 0 24840 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_264
timestamp 1676037725
transform 1 0 25392 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1676037725
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1676037725
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1676037725
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1676037725
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1676037725
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1676037725
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1676037725
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1676037725
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1676037725
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1676037725
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1676037725
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1676037725
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1676037725
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1676037725
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1676037725
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1676037725
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1676037725
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1676037725
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1676037725
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1676037725
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1676037725
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1676037725
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1676037725
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1676037725
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1676037725
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1676037725
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1676037725
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_253
timestamp 1676037725
transform 1 0 24380 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_264
timestamp 1676037725
transform 1 0 25392 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1676037725
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1676037725
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1676037725
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1676037725
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1676037725
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1676037725
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1676037725
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1676037725
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1676037725
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1676037725
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1676037725
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1676037725
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1676037725
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1676037725
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1676037725
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1676037725
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1676037725
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1676037725
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1676037725
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1676037725
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1676037725
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1676037725
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1676037725
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1676037725
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1676037725
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1676037725
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1676037725
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_261
timestamp 1676037725
transform 1 0 25116 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1676037725
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1676037725
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1676037725
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1676037725
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1676037725
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1676037725
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1676037725
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1676037725
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1676037725
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1676037725
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1676037725
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1676037725
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1676037725
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1676037725
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1676037725
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1676037725
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1676037725
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1676037725
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1676037725
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1676037725
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1676037725
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1676037725
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1676037725
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1676037725
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1676037725
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1676037725
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1676037725
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_253
timestamp 1676037725
transform 1 0 24380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_259
timestamp 1676037725
transform 1 0 24932 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_264
timestamp 1676037725
transform 1 0 25392 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1676037725
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1676037725
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1676037725
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1676037725
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1676037725
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1676037725
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1676037725
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1676037725
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1676037725
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1676037725
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1676037725
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1676037725
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1676037725
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1676037725
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1676037725
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1676037725
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1676037725
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1676037725
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1676037725
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1676037725
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1676037725
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1676037725
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1676037725
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1676037725
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1676037725
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1676037725
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1676037725
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_264
timestamp 1676037725
transform 1 0 25392 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1676037725
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1676037725
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1676037725
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1676037725
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1676037725
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1676037725
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1676037725
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1676037725
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1676037725
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1676037725
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1676037725
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1676037725
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1676037725
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1676037725
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1676037725
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1676037725
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1676037725
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1676037725
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1676037725
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1676037725
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1676037725
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1676037725
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1676037725
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1676037725
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1676037725
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1676037725
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1676037725
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_253
timestamp 1676037725
transform 1 0 24380 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_261
timestamp 1676037725
transform 1 0 25116 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1676037725
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1676037725
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1676037725
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1676037725
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1676037725
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1676037725
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1676037725
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1676037725
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1676037725
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1676037725
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1676037725
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1676037725
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1676037725
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1676037725
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1676037725
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1676037725
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1676037725
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1676037725
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1676037725
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1676037725
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1676037725
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1676037725
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1676037725
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1676037725
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1676037725
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1676037725
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_249
timestamp 1676037725
transform 1 0 24012 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_259
timestamp 1676037725
transform 1 0 24932 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_264
timestamp 1676037725
transform 1 0 25392 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1676037725
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1676037725
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1676037725
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1676037725
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1676037725
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1676037725
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1676037725
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1676037725
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1676037725
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1676037725
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_97
timestamp 1676037725
transform 1 0 10028 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_107
timestamp 1676037725
transform 1 0 10948 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_119
timestamp 1676037725
transform 1 0 12052 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_131
timestamp 1676037725
transform 1 0 13156 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1676037725
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1676037725
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1676037725
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1676037725
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1676037725
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1676037725
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1676037725
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1676037725
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1676037725
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1676037725
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1676037725
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1676037725
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1676037725
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_253
timestamp 1676037725
transform 1 0 24380 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_259
timestamp 1676037725
transform 1 0 24932 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_264
timestamp 1676037725
transform 1 0 25392 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1676037725
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1676037725
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1676037725
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1676037725
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1676037725
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1676037725
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1676037725
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1676037725
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_81
timestamp 1676037725
transform 1 0 8556 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_89
timestamp 1676037725
transform 1 0 9292 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_110
timestamp 1676037725
transform 1 0 11224 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_115
timestamp 1676037725
transform 1 0 11684 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_127
timestamp 1676037725
transform 1 0 12788 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_139
timestamp 1676037725
transform 1 0 13892 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_151
timestamp 1676037725
transform 1 0 14996 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_163
timestamp 1676037725
transform 1 0 16100 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1676037725
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1676037725
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1676037725
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1676037725
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1676037725
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1676037725
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1676037725
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1676037725
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1676037725
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1676037725
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_261
timestamp 1676037725
transform 1 0 25116 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1676037725
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1676037725
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1676037725
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1676037725
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1676037725
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1676037725
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1676037725
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1676037725
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1676037725
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_85
timestamp 1676037725
transform 1 0 8924 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_91
timestamp 1676037725
transform 1 0 9476 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_100
timestamp 1676037725
transform 1 0 10304 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_112
timestamp 1676037725
transform 1 0 11408 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_124
timestamp 1676037725
transform 1 0 12512 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_136
timestamp 1676037725
transform 1 0 13616 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1676037725
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1676037725
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1676037725
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1676037725
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1676037725
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1676037725
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1676037725
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1676037725
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1676037725
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1676037725
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1676037725
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1676037725
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_74_253
timestamp 1676037725
transform 1 0 24380 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_258
timestamp 1676037725
transform 1 0 24840 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_264
timestamp 1676037725
transform 1 0 25392 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1676037725
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1676037725
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1676037725
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1676037725
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1676037725
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1676037725
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1676037725
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1676037725
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1676037725
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1676037725
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1676037725
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1676037725
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1676037725
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1676037725
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1676037725
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1676037725
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1676037725
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1676037725
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1676037725
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1676037725
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1676037725
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1676037725
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1676037725
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1676037725
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1676037725
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1676037725
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_249
timestamp 1676037725
transform 1 0 24012 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_257
timestamp 1676037725
transform 1 0 24748 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_264
timestamp 1676037725
transform 1 0 25392 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1676037725
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1676037725
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1676037725
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1676037725
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1676037725
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1676037725
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1676037725
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1676037725
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1676037725
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1676037725
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1676037725
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1676037725
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1676037725
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1676037725
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1676037725
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1676037725
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1676037725
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1676037725
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1676037725
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1676037725
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1676037725
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1676037725
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_229
timestamp 1676037725
transform 1 0 22172 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1676037725
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1676037725
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1676037725
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_253
timestamp 1676037725
transform 1 0 24380 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_261
timestamp 1676037725
transform 1 0 25116 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1676037725
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1676037725
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1676037725
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1676037725
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1676037725
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1676037725
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1676037725
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1676037725
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_81
timestamp 1676037725
transform 1 0 8556 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_93
timestamp 1676037725
transform 1 0 9660 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_101
timestamp 1676037725
transform 1 0 10396 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_77_109
timestamp 1676037725
transform 1 0 11132 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1676037725
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1676037725
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1676037725
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1676037725
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1676037725
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1676037725
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1676037725
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1676037725
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1676037725
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1676037725
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1676037725
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1676037725
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1676037725
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1676037725
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_249
timestamp 1676037725
transform 1 0 24012 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_255
timestamp 1676037725
transform 1 0 24564 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_258
timestamp 1676037725
transform 1 0 24840 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_264
timestamp 1676037725
transform 1 0 25392 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1676037725
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1676037725
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1676037725
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1676037725
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1676037725
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1676037725
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1676037725
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1676037725
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1676037725
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_85
timestamp 1676037725
transform 1 0 8924 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_107
timestamp 1676037725
transform 1 0 10948 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_111
timestamp 1676037725
transform 1 0 11316 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_123
timestamp 1676037725
transform 1 0 12420 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_135
timestamp 1676037725
transform 1 0 13524 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1676037725
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1676037725
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_153
timestamp 1676037725
transform 1 0 15180 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_157
timestamp 1676037725
transform 1 0 15548 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_179
timestamp 1676037725
transform 1 0 17572 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_191
timestamp 1676037725
transform 1 0 18676 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1676037725
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1676037725
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1676037725
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1676037725
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1676037725
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1676037725
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1676037725
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_253
timestamp 1676037725
transform 1 0 24380 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_264
timestamp 1676037725
transform 1 0 25392 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1676037725
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1676037725
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1676037725
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1676037725
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1676037725
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1676037725
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1676037725
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1676037725
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1676037725
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1676037725
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1676037725
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1676037725
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1676037725
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_125
timestamp 1676037725
transform 1 0 12604 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_147
timestamp 1676037725
transform 1 0 14628 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_159
timestamp 1676037725
transform 1 0 15732 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1676037725
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1676037725
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1676037725
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1676037725
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1676037725
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1676037725
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1676037725
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1676037725
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1676037725
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1676037725
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_261
timestamp 1676037725
transform 1 0 25116 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1676037725
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1676037725
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1676037725
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1676037725
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1676037725
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1676037725
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_65
timestamp 1676037725
transform 1 0 7084 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_73
timestamp 1676037725
transform 1 0 7820 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_82
timestamp 1676037725
transform 1 0 8648 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1676037725
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1676037725
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1676037725
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_121
timestamp 1676037725
transform 1 0 12236 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_129
timestamp 1676037725
transform 1 0 12972 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_135
timestamp 1676037725
transform 1 0 13524 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1676037725
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_141
timestamp 1676037725
transform 1 0 14076 0 1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_80_170
timestamp 1676037725
transform 1 0 16744 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_182
timestamp 1676037725
transform 1 0 17848 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_194
timestamp 1676037725
transform 1 0 18952 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1676037725
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1676037725
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1676037725
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1676037725
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1676037725
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1676037725
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_253
timestamp 1676037725
transform 1 0 24380 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_259
timestamp 1676037725
transform 1 0 24932 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_264
timestamp 1676037725
transform 1 0 25392 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1676037725
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1676037725
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1676037725
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1676037725
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1676037725
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1676037725
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1676037725
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1676037725
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1676037725
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_93
timestamp 1676037725
transform 1 0 9660 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_99
timestamp 1676037725
transform 1 0 10212 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_106
timestamp 1676037725
transform 1 0 10856 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_81_113
timestamp 1676037725
transform 1 0 11500 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_121
timestamp 1676037725
transform 1 0 12236 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_127
timestamp 1676037725
transform 1 0 12788 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_160
timestamp 1676037725
transform 1 0 15824 0 -1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1676037725
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1676037725
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1676037725
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1676037725
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1676037725
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1676037725
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1676037725
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1676037725
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1676037725
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_264
timestamp 1676037725
transform 1 0 25392 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1676037725
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1676037725
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1676037725
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1676037725
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1676037725
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1676037725
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1676037725
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1676037725
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1676037725
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1676037725
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1676037725
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_109
timestamp 1676037725
transform 1 0 11132 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_113
timestamp 1676037725
transform 1 0 11500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_117
timestamp 1676037725
transform 1 0 11868 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_129
timestamp 1676037725
transform 1 0 12972 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_137
timestamp 1676037725
transform 1 0 13708 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1676037725
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1676037725
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1676037725
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1676037725
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1676037725
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1676037725
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1676037725
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1676037725
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1676037725
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1676037725
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1676037725
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1676037725
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_253
timestamp 1676037725
transform 1 0 24380 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_261
timestamp 1676037725
transform 1 0 25116 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1676037725
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1676037725
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1676037725
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1676037725
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1676037725
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1676037725
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1676037725
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1676037725
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_81
timestamp 1676037725
transform 1 0 8556 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_89
timestamp 1676037725
transform 1 0 9292 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_96
timestamp 1676037725
transform 1 0 9936 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_108
timestamp 1676037725
transform 1 0 11040 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1676037725
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1676037725
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1676037725
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1676037725
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1676037725
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1676037725
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1676037725
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1676037725
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1676037725
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1676037725
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1676037725
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1676037725
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1676037725
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1676037725
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_249
timestamp 1676037725
transform 1 0 24012 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_259
timestamp 1676037725
transform 1 0 24932 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_264
timestamp 1676037725
transform 1 0 25392 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1676037725
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1676037725
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1676037725
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1676037725
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1676037725
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1676037725
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1676037725
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1676037725
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1676037725
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1676037725
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_97
timestamp 1676037725
transform 1 0 10028 0 1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_84_103
timestamp 1676037725
transform 1 0 10580 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_115
timestamp 1676037725
transform 1 0 11684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_127
timestamp 1676037725
transform 1 0 12788 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1676037725
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1676037725
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1676037725
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1676037725
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1676037725
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1676037725
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1676037725
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1676037725
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1676037725
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1676037725
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1676037725
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1676037725
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1676037725
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_84_253
timestamp 1676037725
transform 1 0 24380 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_259
timestamp 1676037725
transform 1 0 24932 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_264
timestamp 1676037725
transform 1 0 25392 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1676037725
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1676037725
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1676037725
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1676037725
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1676037725
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1676037725
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_85_57
timestamp 1676037725
transform 1 0 6348 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_85_80
timestamp 1676037725
transform 1 0 8464 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_84
timestamp 1676037725
transform 1 0 8832 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_96
timestamp 1676037725
transform 1 0 9936 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_108
timestamp 1676037725
transform 1 0 11040 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1676037725
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1676037725
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1676037725
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1676037725
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1676037725
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1676037725
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1676037725
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1676037725
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1676037725
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1676037725
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1676037725
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1676037725
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1676037725
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1676037725
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1676037725
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_261
timestamp 1676037725
transform 1 0 25116 0 -1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1676037725
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1676037725
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1676037725
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1676037725
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1676037725
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1676037725
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1676037725
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1676037725
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1676037725
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1676037725
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_97
timestamp 1676037725
transform 1 0 10028 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_105
timestamp 1676037725
transform 1 0 10764 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_111
timestamp 1676037725
transform 1 0 11316 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_116
timestamp 1676037725
transform 1 0 11776 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_128
timestamp 1676037725
transform 1 0 12880 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1676037725
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1676037725
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1676037725
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1676037725
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1676037725
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1676037725
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1676037725
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1676037725
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1676037725
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1676037725
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1676037725
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1676037725
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_86_253
timestamp 1676037725
transform 1 0 24380 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_86_258
timestamp 1676037725
transform 1 0 24840 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_264
timestamp 1676037725
transform 1 0 25392 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1676037725
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1676037725
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1676037725
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1676037725
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1676037725
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1676037725
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1676037725
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1676037725
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1676037725
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1676037725
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1676037725
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1676037725
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1676037725
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1676037725
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1676037725
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1676037725
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1676037725
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1676037725
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1676037725
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1676037725
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1676037725
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1676037725
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1676037725
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1676037725
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1676037725
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1676037725
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_249
timestamp 1676037725
transform 1 0 24012 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_253
timestamp 1676037725
transform 1 0 24380 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_264
timestamp 1676037725
transform 1 0 25392 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1676037725
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1676037725
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1676037725
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1676037725
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1676037725
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1676037725
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_65
timestamp 1676037725
transform 1 0 7084 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_69
timestamp 1676037725
transform 1 0 7452 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_76
timestamp 1676037725
transform 1 0 8096 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_88_85
timestamp 1676037725
transform 1 0 8924 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_89
timestamp 1676037725
transform 1 0 9292 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_94
timestamp 1676037725
transform 1 0 9752 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_106
timestamp 1676037725
transform 1 0 10856 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_118
timestamp 1676037725
transform 1 0 11960 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_130
timestamp 1676037725
transform 1 0 13064 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_138
timestamp 1676037725
transform 1 0 13800 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1676037725
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1676037725
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1676037725
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1676037725
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1676037725
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1676037725
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1676037725
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1676037725
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1676037725
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1676037725
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1676037725
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1676037725
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_253
timestamp 1676037725
transform 1 0 24380 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_88_261
timestamp 1676037725
transform 1 0 25116 0 1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1676037725
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1676037725
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1676037725
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1676037725
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1676037725
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1676037725
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1676037725
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1676037725
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1676037725
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1676037725
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1676037725
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1676037725
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1676037725
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1676037725
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1676037725
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1676037725
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1676037725
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1676037725
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1676037725
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1676037725
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1676037725
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1676037725
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1676037725
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1676037725
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1676037725
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1676037725
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_249
timestamp 1676037725
transform 1 0 24012 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_253
timestamp 1676037725
transform 1 0 24380 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_256
timestamp 1676037725
transform 1 0 24656 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_264
timestamp 1676037725
transform 1 0 25392 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1676037725
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1676037725
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1676037725
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1676037725
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1676037725
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1676037725
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_65
timestamp 1676037725
transform 1 0 7084 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_69
timestamp 1676037725
transform 1 0 7452 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_74
timestamp 1676037725
transform 1 0 7912 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_90_81
timestamp 1676037725
transform 1 0 8556 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_90_85
timestamp 1676037725
transform 1 0 8924 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_90_91
timestamp 1676037725
transform 1 0 9476 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_103
timestamp 1676037725
transform 1 0 10580 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_115
timestamp 1676037725
transform 1 0 11684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_127
timestamp 1676037725
transform 1 0 12788 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1676037725
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1676037725
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1676037725
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1676037725
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1676037725
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1676037725
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1676037725
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1676037725
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1676037725
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1676037725
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1676037725
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1676037725
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1676037725
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_90_253
timestamp 1676037725
transform 1 0 24380 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_256
timestamp 1676037725
transform 1 0 24656 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_264
timestamp 1676037725
transform 1 0 25392 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1676037725
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1676037725
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1676037725
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1676037725
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1676037725
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1676037725
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1676037725
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1676037725
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1676037725
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1676037725
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1676037725
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1676037725
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1676037725
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1676037725
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1676037725
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1676037725
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1676037725
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1676037725
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1676037725
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1676037725
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1676037725
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1676037725
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1676037725
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1676037725
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1676037725
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1676037725
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_249
timestamp 1676037725
transform 1 0 24012 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_91_259
timestamp 1676037725
transform 1 0 24932 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_264
timestamp 1676037725
transform 1 0 25392 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1676037725
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1676037725
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1676037725
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1676037725
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1676037725
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_53
timestamp 1676037725
transform 1 0 5980 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_62
timestamp 1676037725
transform 1 0 6808 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_74
timestamp 1676037725
transform 1 0 7912 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_82
timestamp 1676037725
transform 1 0 8648 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1676037725
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1676037725
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1676037725
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1676037725
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1676037725
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1676037725
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1676037725
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1676037725
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1676037725
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1676037725
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1676037725
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1676037725
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1676037725
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1676037725
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1676037725
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1676037725
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1676037725
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1676037725
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_92_253
timestamp 1676037725
transform 1 0 24380 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_256
timestamp 1676037725
transform 1 0 24656 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_264
timestamp 1676037725
transform 1 0 25392 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1676037725
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1676037725
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1676037725
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_39
timestamp 1676037725
transform 1 0 4692 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_43
timestamp 1676037725
transform 1 0 5060 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_47
timestamp 1676037725
transform 1 0 5428 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1676037725
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1676037725
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1676037725
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1676037725
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1676037725
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1676037725
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1676037725
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1676037725
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1676037725
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1676037725
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1676037725
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1676037725
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1676037725
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1676037725
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1676037725
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1676037725
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1676037725
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1676037725
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1676037725
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1676037725
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_237
timestamp 1676037725
transform 1 0 22908 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_241
timestamp 1676037725
transform 1 0 23276 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_244
timestamp 1676037725
transform 1 0 23552 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_93_256
timestamp 1676037725
transform 1 0 24656 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_264
timestamp 1676037725
transform 1 0 25392 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_3
timestamp 1676037725
transform 1 0 1380 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_21
timestamp 1676037725
transform 1 0 3036 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1676037725
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_29
timestamp 1676037725
transform 1 0 3772 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_47
timestamp 1676037725
transform 1 0 5428 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_59
timestamp 1676037725
transform 1 0 6532 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_76
timestamp 1676037725
transform 1 0 8096 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1676037725
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_97
timestamp 1676037725
transform 1 0 10028 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1676037725
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1676037725
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1676037725
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1676037725
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1676037725
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1676037725
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1676037725
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1676037725
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1676037725
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1676037725
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1676037725
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1676037725
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_233
timestamp 1676037725
transform 1 0 22540 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_237
timestamp 1676037725
transform 1 0 22908 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_242
timestamp 1676037725
transform 1 0 23368 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_250
timestamp 1676037725
transform 1 0 24104 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_94_255
timestamp 1676037725
transform 1 0 24564 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_258
timestamp 1676037725
transform 1 0 24840 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_264
timestamp 1676037725
transform 1 0 25392 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_3
timestamp 1676037725
transform 1 0 1380 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_9
timestamp 1676037725
transform 1 0 1932 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_26
timestamp 1676037725
transform 1 0 3496 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_29
timestamp 1676037725
transform 1 0 3772 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_37
timestamp 1676037725
transform 1 0 4508 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_54
timestamp 1676037725
transform 1 0 6072 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_57
timestamp 1676037725
transform 1 0 6348 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_65
timestamp 1676037725
transform 1 0 7084 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_82
timestamp 1676037725
transform 1 0 8648 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_85
timestamp 1676037725
transform 1 0 8924 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_89
timestamp 1676037725
transform 1 0 9292 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_95_106
timestamp 1676037725
transform 1 0 10856 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_95_113
timestamp 1676037725
transform 1 0 11500 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_119
timestamp 1676037725
transform 1 0 12052 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_136
timestamp 1676037725
transform 1 0 13616 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_141
timestamp 1676037725
transform 1 0 14076 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_146
timestamp 1676037725
transform 1 0 14536 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_153
timestamp 1676037725
transform 1 0 15180 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_157
timestamp 1676037725
transform 1 0 15548 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_95_165
timestamp 1676037725
transform 1 0 16284 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_169
timestamp 1676037725
transform 1 0 16652 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_174
timestamp 1676037725
transform 1 0 17112 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_178
timestamp 1676037725
transform 1 0 17480 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_183
timestamp 1676037725
transform 1 0 17940 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_187
timestamp 1676037725
transform 1 0 18308 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_193
timestamp 1676037725
transform 1 0 18860 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_197
timestamp 1676037725
transform 1 0 19228 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_209
timestamp 1676037725
transform 1 0 20332 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_217
timestamp 1676037725
transform 1 0 21068 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_221
timestamp 1676037725
transform 1 0 21436 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_225
timestamp 1676037725
transform 1 0 21804 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_231
timestamp 1676037725
transform 1 0 22356 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_235
timestamp 1676037725
transform 1 0 22724 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_239
timestamp 1676037725
transform 1 0 23092 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_244
timestamp 1676037725
transform 1 0 23552 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_248
timestamp 1676037725
transform 1 0 23920 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_253
timestamp 1676037725
transform 1 0 24380 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_259
timestamp 1676037725
transform 1 0 24932 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_263
timestamp 1676037725
transform 1 0 25300 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform 1 0 25116 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 1564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 23276 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1676037725
transform 1 0 25116 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1676037725
transform 1 0 25116 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 25116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1676037725
transform 1 0 25024 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1676037725
transform 1 0 25024 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1676037725
transform 1 0 25116 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1676037725
transform 1 0 25116 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1676037725
transform 1 0 25116 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1676037725
transform 1 0 25116 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1676037725
transform 1 0 25024 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1676037725
transform 1 0 25116 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1676037725
transform 1 0 25024 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1676037725
transform 1 0 25024 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1676037725
transform 1 0 25024 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1676037725
transform 1 0 25116 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1676037725
transform 1 0 25116 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1676037725
transform 1 0 25116 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1676037725
transform 1 0 25116 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1676037725
transform 1 0 25024 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1676037725
transform 1 0 25024 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1676037725
transform 1 0 24472 0 -1 50048
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1676037725
transform 1 0 23828 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1676037725
transform 1 0 23828 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1676037725
transform 1 0 23184 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1676037725
transform 1 0 25116 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1676037725
transform 1 0 25116 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1676037725
transform 1 0 25116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1676037725
transform 1 0 25116 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1676037725
transform 1 0 25116 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1676037725
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1676037725
transform 1 0 5152 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1676037725
transform 1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1676037725
transform 1 0 6348 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1676037725
transform 1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1676037725
transform 1 0 7176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1676037725
transform 1 0 7820 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1676037725
transform 1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1676037725
transform 1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1676037725
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1676037725
transform 1 0 2852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1676037725
transform 1 0 9292 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1676037725
transform 1 0 9660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1676037725
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1676037725
transform 1 0 10396 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1676037725
transform 1 0 10304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1676037725
transform 1 0 11684 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1676037725
transform 1 0 10948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1676037725
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1676037725
transform 1 0 11040 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input55
timestamp 1676037725
transform 1 0 2116 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1676037725
transform 1 0 2576 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1676037725
transform 1 0 3404 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1676037725
transform 1 0 1564 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1676037725
transform 1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1676037725
transform 1 0 4232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1676037725
transform 1 0 5152 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1676037725
transform 1 0 14260 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1676037725
transform 1 0 14904 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1676037725
transform 1 0 16836 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1676037725
transform 1 0 17664 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1676037725
transform 1 0 19412 0 -1 54400
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_16  input68
timestamp 1676037725
transform 1 0 23552 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  input69 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24840 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input70
timestamp 1676037725
transform 1 0 24840 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input71
timestamp 1676037725
transform 1 0 24840 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input72 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25024 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input73
timestamp 1676037725
transform 1 0 25024 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input74
timestamp 1676037725
transform 1 0 23736 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input75
timestamp 1676037725
transform 1 0 24288 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input76
timestamp 1676037725
transform 1 0 23000 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1676037725
transform 1 0 20700 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1676037725
transform 1 0 21988 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input79
timestamp 1676037725
transform 1 0 23184 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input80
timestamp 1676037725
transform 1 0 24564 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output81 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17480 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1676037725
transform 1 0 1564 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1676037725
transform 1 0 14904 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1676037725
transform 1 0 23920 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1676037725
transform 1 0 22632 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1676037725
transform 1 0 22080 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1676037725
transform 1 0 22632 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1676037725
transform 1 0 23920 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1676037725
transform 1 0 22632 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1676037725
transform 1 0 22632 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1676037725
transform 1 0 22080 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1676037725
transform 1 0 23920 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1676037725
transform 1 0 22632 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1676037725
transform 1 0 9752 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1676037725
transform 1 0 22632 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1676037725
transform 1 0 22080 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1676037725
transform 1 0 22632 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1676037725
transform 1 0 23920 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1676037725
transform 1 0 22632 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1676037725
transform 1 0 22080 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1676037725
transform 1 0 22632 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1676037725
transform 1 0 23920 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1676037725
transform 1 0 22632 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1676037725
transform 1 0 23920 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output105
timestamp 1676037725
transform 1 0 18216 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output106
timestamp 1676037725
transform 1 0 20056 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output107
timestamp 1676037725
transform 1 0 18216 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1676037725
transform 1 0 20792 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1676037725
transform 1 0 22632 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1676037725
transform 1 0 22080 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1676037725
transform 1 0 23920 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1676037725
transform 1 0 22632 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1676037725
transform 1 0 12328 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1676037725
transform 1 0 18676 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1676037725
transform 1 0 19412 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1676037725
transform 1 0 19412 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1676037725
transform 1 0 18676 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1676037725
transform 1 0 21988 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform 1 0 21252 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform 1 0 19412 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform 1 0 21988 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform 1 0 21712 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform 1 0 12328 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform 1 0 21988 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform 1 0 21252 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform 1 0 23828 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform 1 0 23828 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform 1 0 20056 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform 1 0 16928 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform 1 0 22080 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1676037725
transform 1 0 20240 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1676037725
transform 1 0 20056 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1676037725
transform 1 0 12052 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1676037725
transform 1 0 12972 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1676037725
transform 1 0 14260 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1676037725
transform 1 0 14444 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1676037725
transform 1 0 16836 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1676037725
transform 1 0 16100 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1676037725
transform 1 0 16836 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1676037725
transform 1 0 16836 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1676037725
transform 1 0 2024 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1676037725
transform 1 0 3956 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1676037725
transform 1 0 4600 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1676037725
transform 1 0 6624 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1676037725
transform 1 0 7176 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1676037725
transform 1 0 9384 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1676037725
transform 1 0 10764 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1676037725
transform 1 0 12144 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 25852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 25852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 25852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 25852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 25852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 25852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 25852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 25852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 25852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 25852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 25852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 25852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 25852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 25852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 25852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 25852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 25852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 25852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 25852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 25852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 25852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 25852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 25852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1676037725
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1676037725
transform -1 0 25852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1676037725
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1676037725
transform -1 0 25852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1676037725
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1676037725
transform -1 0 25852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1676037725
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1676037725
transform -1 0 25852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1676037725
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1676037725
transform -1 0 25852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1676037725
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1676037725
transform -1 0 25852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1676037725
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1676037725
transform -1 0 25852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1676037725
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1676037725
transform -1 0 25852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1676037725
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1676037725
transform -1 0 25852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1676037725
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1676037725
transform -1 0 25852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1676037725
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1676037725
transform -1 0 25852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1676037725
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1676037725
transform -1 0 25852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1676037725
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1676037725
transform -1 0 25852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1676037725
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1676037725
transform -1 0 25852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1676037725
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1676037725
transform -1 0 25852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1676037725
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1676037725
transform -1 0 25852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1676037725
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1676037725
transform -1 0 25852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1676037725
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1676037725
transform -1 0 25852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1676037725
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1676037725
transform -1 0 25852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1676037725
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1676037725
transform -1 0 25852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1676037725
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1676037725
transform -1 0 25852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1676037725
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1676037725
transform -1 0 25852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1676037725
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1676037725
transform -1 0 25852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1676037725
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1676037725
transform -1 0 25852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1676037725
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1676037725
transform -1 0 25852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1676037725
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1676037725
transform -1 0 25852 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1676037725
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1676037725
transform -1 0 25852 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1676037725
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1676037725
transform -1 0 25852 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1676037725
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1676037725
transform -1 0 25852 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1676037725
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1676037725
transform -1 0 25852 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1676037725
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1676037725
transform -1 0 25852 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1676037725
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1676037725
transform -1 0 25852 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1676037725
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1676037725
transform -1 0 25852 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1676037725
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1676037725
transform -1 0 25852 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1676037725
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1676037725
transform -1 0 25852 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1676037725
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1676037725
transform -1 0 25852 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1676037725
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1676037725
transform -1 0 25852 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1676037725
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1676037725
transform -1 0 25852 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18584 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19872 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22080 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23368 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23552 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23276 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21528 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19688 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21896 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23184 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23552 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23552 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23184 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22080 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19872 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17940 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17020 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16744 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16744 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17388 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20700 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22448 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23276 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23460 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21620 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19504 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19044 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20608 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23460 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20332 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13340 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 9108 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11684 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10488 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 9292 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11132 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11776 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 11408 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13340 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13064 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 11960 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12972 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10856 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 9108 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9384 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 8096 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 6532 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6624 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9108 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10672 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12328 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13064 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12696 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12512 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11776 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10396 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9108 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9108 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9016 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10764 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11684 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13800 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15180 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16100 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16376 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14904 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13156 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13892 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 15088 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15916 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17112 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19596 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20516 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20424 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20240 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22816 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23092 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23092 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22632 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22080 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19504 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18768 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 18492 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17296 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_1.mux_l1_in_1__198
timestamp 1676037725
transform 1 0 20700 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19504 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20056 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18584 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_3.mux_l2_in_0__153
timestamp 1676037725
transform 1 0 24564 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21988 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_5.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_5.mux_l2_in_0__160
timestamp 1676037725
transform 1 0 21252 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_5.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22172 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20884 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_7.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_7.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19228 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_7.mux_l1_in_1__162
timestamp 1676037725
transform 1 0 19688 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_7.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19504 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17848 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_9.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22632 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_9.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_9.mux_l2_in_0__163
timestamp 1676037725
transform 1 0 21988 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20240 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_11.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_11.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_11.mux_l2_in_0__199
timestamp 1676037725
transform 1 0 20884 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20792 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_13.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_13.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22080 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_13.mux_l2_in_0__200
timestamp 1676037725
transform 1 0 24564 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19596 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_15.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22816 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_15.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20424 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_15.mux_l2_in_0__201
timestamp 1676037725
transform 1 0 20700 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18492 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_17.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_17.mux_l2_in_0__202
timestamp 1676037725
transform 1 0 18676 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_17.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17848 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_19.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20148 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_19.mux_l2_in_0__151
timestamp 1676037725
transform 1 0 18216 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_19.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17756 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16100 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_29.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20056 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_29.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17480 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_29.mux_l2_in_0__152
timestamp 1676037725
transform 1 0 18032 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15916 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_31.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21620 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_31.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_31.mux_l2_in_0__154
timestamp 1676037725
transform 1 0 19688 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18676 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_33.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23000 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_33.mux_l2_in_0__155
timestamp 1676037725
transform 1 0 24564 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_33.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22356 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21068 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_35.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_35.mux_l2_in_0__156
timestamp 1676037725
transform 1 0 24748 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_35.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21252 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_45.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22724 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_45.mux_l2_in_0__157
timestamp 1676037725
transform 1 0 21252 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_45.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19688 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_47.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_47.mux_l2_in_0__158
timestamp 1676037725
transform 1 0 20056 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_47.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19872 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19044 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_49.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_49.mux_l2_in_0__159
timestamp 1676037725
transform 1 0 19412 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_49.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18768 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15548 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_51.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23552 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_51.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22264 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_51.mux_l2_in_0__161
timestamp 1676037725
transform 1 0 21252 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19964 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15548 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15548 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12144 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_0.mux_l2_in_1__164
timestamp 1676037725
transform 1 0 7176 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 7636 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16928 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14812 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15180 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 9200 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_2.mux_l2_in_1__170
timestamp 1676037725
transform 1 0 9936 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 12144 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16836 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15180 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15456 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 10672 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_4.mux_l2_in_1__181
timestamp 1676037725
transform 1 0 11684 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 13524 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17572 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 16836 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15272 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11316 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_6.mux_l2_in_1__192
timestamp 1676037725
transform 1 0 11684 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 14444 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18032 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15180 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15640 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13248 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_8.mux_l2_in_1__193
timestamp 1676037725
transform 1 0 9108 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l2_in_1_
timestamp 1676037725
transform 1 0 9016 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l3_in_0_
timestamp 1676037725
transform 1 0 11960 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16836 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14260 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11224 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 6624 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_10.mux_l2_in_1__165
timestamp 1676037725
transform 1 0 7360 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 9936 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14996 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_12.mux_l1_in_1_
timestamp 1676037725
transform 1 0 7820 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_12.mux_l1_in_1__166
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11500 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16468 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15732 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_14.mux_l1_in_1__167
timestamp 1676037725
transform 1 0 14260 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_14.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12236 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14812 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18676 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_16.mux_l1_in_1__168
timestamp 1676037725
transform 1 0 13432 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_16.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12788 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14996 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18952 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14536 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14536 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_18.mux_l2_in_0__169
timestamp 1676037725
transform 1 0 15732 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18676 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11408 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_20.mux_l2_in_0__171
timestamp 1676037725
transform 1 0 14260 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12328 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18032 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_22.mux_l1_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_22.mux_l2_in_0__172
timestamp 1676037725
transform 1 0 12328 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_22.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12236 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_24.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_24.mux_l2_in_0__173
timestamp 1676037725
transform 1 0 16100 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_24.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18216 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_26.mux_l1_in_0_
timestamp 1676037725
transform 1 0 13800 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_26.mux_l2_in_0__174
timestamp 1676037725
transform 1 0 17664 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_26.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16468 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20148 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_28.mux_l1_in_1__175
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_28.mux_l1_in_1_
timestamp 1676037725
transform 1 0 13708 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19780 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18032 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_30.mux_l1_in_1__176
timestamp 1676037725
transform 1 0 15732 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_30.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15732 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17480 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20792 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17848 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_32.mux_l1_in_1__177
timestamp 1676037725
transform 1 0 15732 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_32.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21620 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_34.mux_l1_in_1__178
timestamp 1676037725
transform 1 0 13156 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_34.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12972 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21528 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 13340 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_36.mux_l2_in_0__179
timestamp 1676037725
transform 1 0 16836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14720 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14352 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_38.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14996 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_38.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_38.mux_l2_in_0__180
timestamp 1676037725
transform 1 0 16100 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_40.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_40.mux_l2_in_0__182
timestamp 1676037725
transform 1 0 16100 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_40.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23092 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_42.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_42.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_42.mux_l2_in_0__183
timestamp 1676037725
transform 1 0 21988 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_44.mux_l1_in_1__184
timestamp 1676037725
transform 1 0 16652 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_44.mux_l1_in_1_
timestamp 1676037725
transform 1 0 18032 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19596 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19688 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_46.mux_l1_in_1_
timestamp 1676037725
transform 1 0 18768 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_46.mux_l1_in_1__185
timestamp 1676037725
transform 1 0 18676 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20424 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_48.mux_l1_in_1__186
timestamp 1676037725
transform 1 0 20700 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_48.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19596 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21436 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22816 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_50.mux_l2_in_0__187
timestamp 1676037725
transform 1 0 24196 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_52.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19504 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_52.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_52.mux_l2_in_0__188
timestamp 1676037725
transform 1 0 22724 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_54.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_54.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20516 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_54.mux_l2_in_0__189
timestamp 1676037725
transform 1 0 21252 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_56.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17940 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_56.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17296 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_56.mux_l2_in_0__190
timestamp 1676037725
transform 1 0 23828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_58.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16928 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_58.mux_l1_in_1__191
timestamp 1676037725
transform 1 0 11684 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_58.mux_l1_in_1_
timestamp 1676037725
transform 1 0 11040 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_58.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21804 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 3680 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 8832 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 13984 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 19136 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 24288 0 -1 54400
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 25870 56200 25926 57000 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 1490 0 1546 800 0 FreeSans 224 90 0 0 ccff_head_0
port 3 nsew signal input
flabel metal3 s 26200 688 27000 808 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 1030 56200 1086 57000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 26200 25984 27000 26104 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 6 nsew signal input
flabel metal3 s 26200 34144 27000 34264 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 7 nsew signal input
flabel metal3 s 26200 34960 27000 35080 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 8 nsew signal input
flabel metal3 s 26200 35776 27000 35896 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 9 nsew signal input
flabel metal3 s 26200 36592 27000 36712 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 10 nsew signal input
flabel metal3 s 26200 37408 27000 37528 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 11 nsew signal input
flabel metal3 s 26200 38224 27000 38344 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 12 nsew signal input
flabel metal3 s 26200 39040 27000 39160 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 13 nsew signal input
flabel metal3 s 26200 39856 27000 39976 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 14 nsew signal input
flabel metal3 s 26200 40672 27000 40792 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 15 nsew signal input
flabel metal3 s 26200 41488 27000 41608 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 16 nsew signal input
flabel metal3 s 26200 26800 27000 26920 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 17 nsew signal input
flabel metal3 s 26200 42304 27000 42424 0 FreeSans 480 0 0 0 chanx_right_in[20]
port 18 nsew signal input
flabel metal3 s 26200 43120 27000 43240 0 FreeSans 480 0 0 0 chanx_right_in[21]
port 19 nsew signal input
flabel metal3 s 26200 43936 27000 44056 0 FreeSans 480 0 0 0 chanx_right_in[22]
port 20 nsew signal input
flabel metal3 s 26200 44752 27000 44872 0 FreeSans 480 0 0 0 chanx_right_in[23]
port 21 nsew signal input
flabel metal3 s 26200 45568 27000 45688 0 FreeSans 480 0 0 0 chanx_right_in[24]
port 22 nsew signal input
flabel metal3 s 26200 46384 27000 46504 0 FreeSans 480 0 0 0 chanx_right_in[25]
port 23 nsew signal input
flabel metal3 s 26200 47200 27000 47320 0 FreeSans 480 0 0 0 chanx_right_in[26]
port 24 nsew signal input
flabel metal3 s 26200 48016 27000 48136 0 FreeSans 480 0 0 0 chanx_right_in[27]
port 25 nsew signal input
flabel metal3 s 26200 48832 27000 48952 0 FreeSans 480 0 0 0 chanx_right_in[28]
port 26 nsew signal input
flabel metal3 s 26200 49648 27000 49768 0 FreeSans 480 0 0 0 chanx_right_in[29]
port 27 nsew signal input
flabel metal3 s 26200 27616 27000 27736 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 28 nsew signal input
flabel metal3 s 26200 28432 27000 28552 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 29 nsew signal input
flabel metal3 s 26200 29248 27000 29368 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 30 nsew signal input
flabel metal3 s 26200 30064 27000 30184 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 31 nsew signal input
flabel metal3 s 26200 30880 27000 31000 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 32 nsew signal input
flabel metal3 s 26200 31696 27000 31816 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 33 nsew signal input
flabel metal3 s 26200 32512 27000 32632 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 34 nsew signal input
flabel metal3 s 26200 33328 27000 33448 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 35 nsew signal input
flabel metal3 s 26200 1504 27000 1624 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 36 nsew signal tristate
flabel metal3 s 26200 9664 27000 9784 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 37 nsew signal tristate
flabel metal3 s 26200 10480 27000 10600 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 38 nsew signal tristate
flabel metal3 s 26200 11296 27000 11416 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 39 nsew signal tristate
flabel metal3 s 26200 12112 27000 12232 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 40 nsew signal tristate
flabel metal3 s 26200 12928 27000 13048 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 41 nsew signal tristate
flabel metal3 s 26200 13744 27000 13864 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 42 nsew signal tristate
flabel metal3 s 26200 14560 27000 14680 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 43 nsew signal tristate
flabel metal3 s 26200 15376 27000 15496 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 44 nsew signal tristate
flabel metal3 s 26200 16192 27000 16312 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 45 nsew signal tristate
flabel metal3 s 26200 17008 27000 17128 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 46 nsew signal tristate
flabel metal3 s 26200 2320 27000 2440 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 47 nsew signal tristate
flabel metal3 s 26200 17824 27000 17944 0 FreeSans 480 0 0 0 chanx_right_out[20]
port 48 nsew signal tristate
flabel metal3 s 26200 18640 27000 18760 0 FreeSans 480 0 0 0 chanx_right_out[21]
port 49 nsew signal tristate
flabel metal3 s 26200 19456 27000 19576 0 FreeSans 480 0 0 0 chanx_right_out[22]
port 50 nsew signal tristate
flabel metal3 s 26200 20272 27000 20392 0 FreeSans 480 0 0 0 chanx_right_out[23]
port 51 nsew signal tristate
flabel metal3 s 26200 21088 27000 21208 0 FreeSans 480 0 0 0 chanx_right_out[24]
port 52 nsew signal tristate
flabel metal3 s 26200 21904 27000 22024 0 FreeSans 480 0 0 0 chanx_right_out[25]
port 53 nsew signal tristate
flabel metal3 s 26200 22720 27000 22840 0 FreeSans 480 0 0 0 chanx_right_out[26]
port 54 nsew signal tristate
flabel metal3 s 26200 23536 27000 23656 0 FreeSans 480 0 0 0 chanx_right_out[27]
port 55 nsew signal tristate
flabel metal3 s 26200 24352 27000 24472 0 FreeSans 480 0 0 0 chanx_right_out[28]
port 56 nsew signal tristate
flabel metal3 s 26200 25168 27000 25288 0 FreeSans 480 0 0 0 chanx_right_out[29]
port 57 nsew signal tristate
flabel metal3 s 26200 3136 27000 3256 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 58 nsew signal tristate
flabel metal3 s 26200 3952 27000 4072 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 59 nsew signal tristate
flabel metal3 s 26200 4768 27000 4888 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 60 nsew signal tristate
flabel metal3 s 26200 5584 27000 5704 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 61 nsew signal tristate
flabel metal3 s 26200 6400 27000 6520 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 62 nsew signal tristate
flabel metal3 s 26200 7216 27000 7336 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 63 nsew signal tristate
flabel metal3 s 26200 8032 27000 8152 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 64 nsew signal tristate
flabel metal3 s 26200 8848 27000 8968 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 65 nsew signal tristate
flabel metal2 s 1858 0 1914 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[0]
port 66 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[10]
port 67 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[11]
port 68 nsew signal input
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[12]
port 69 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[13]
port 70 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[14]
port 71 nsew signal input
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[15]
port 72 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[16]
port 73 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[17]
port 74 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[18]
port 75 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[19]
port 76 nsew signal input
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[1]
port 77 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[20]
port 78 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[21]
port 79 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[22]
port 80 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[23]
port 81 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[24]
port 82 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[25]
port 83 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[26]
port 84 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[27]
port 85 nsew signal input
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[28]
port 86 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[29]
port 87 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[2]
port 88 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[3]
port 89 nsew signal input
flabel metal2 s 3330 0 3386 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[4]
port 90 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[5]
port 91 nsew signal input
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[6]
port 92 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[7]
port 93 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[8]
port 94 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[9]
port 95 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[0]
port 96 nsew signal tristate
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[10]
port 97 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[11]
port 98 nsew signal tristate
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[12]
port 99 nsew signal tristate
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[13]
port 100 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[14]
port 101 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[15]
port 102 nsew signal tristate
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[16]
port 103 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[17]
port 104 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[18]
port 105 nsew signal tristate
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[19]
port 106 nsew signal tristate
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[1]
port 107 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[20]
port 108 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[21]
port 109 nsew signal tristate
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[22]
port 110 nsew signal tristate
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[23]
port 111 nsew signal tristate
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[24]
port 112 nsew signal tristate
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[25]
port 113 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[26]
port 114 nsew signal tristate
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[27]
port 115 nsew signal tristate
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[28]
port 116 nsew signal tristate
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[29]
port 117 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[2]
port 118 nsew signal tristate
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[3]
port 119 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[4]
port 120 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[5]
port 121 nsew signal tristate
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[6]
port 122 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[7]
port 123 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[8]
port 124 nsew signal tristate
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[9]
port 125 nsew signal tristate
flabel metal2 s 2410 56200 2466 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[0]
port 126 nsew signal tristate
flabel metal2 s 3790 56200 3846 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[1]
port 127 nsew signal tristate
flabel metal2 s 5170 56200 5226 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[2]
port 128 nsew signal tristate
flabel metal2 s 6550 56200 6606 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[3]
port 129 nsew signal tristate
flabel metal2 s 13450 56200 13506 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[0]
port 130 nsew signal input
flabel metal2 s 14830 56200 14886 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[1]
port 131 nsew signal input
flabel metal2 s 16210 56200 16266 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[2]
port 132 nsew signal input
flabel metal2 s 17590 56200 17646 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[3]
port 133 nsew signal input
flabel metal2 s 7930 56200 7986 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[0]
port 134 nsew signal tristate
flabel metal2 s 9310 56200 9366 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[1]
port 135 nsew signal tristate
flabel metal2 s 10690 56200 10746 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[2]
port 136 nsew signal tristate
flabel metal2 s 12070 56200 12126 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[3]
port 137 nsew signal tristate
flabel metal2 s 18970 56200 19026 57000 0 FreeSans 224 90 0 0 isol_n
port 138 nsew signal input
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 prog_clk
port 139 nsew signal input
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 prog_reset
port 140 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 reset
port 141 nsew signal input
flabel metal3 s 26200 50464 27000 50584 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 142 nsew signal input
flabel metal3 s 26200 51280 27000 51400 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
port 143 nsew signal input
flabel metal3 s 26200 52096 27000 52216 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 144 nsew signal input
flabel metal3 s 26200 52912 27000 53032 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
port 145 nsew signal input
flabel metal3 s 26200 53728 27000 53848 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 146 nsew signal input
flabel metal3 s 26200 54544 27000 54664 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
port 147 nsew signal input
flabel metal3 s 26200 55360 27000 55480 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
port 148 nsew signal input
flabel metal3 s 26200 56176 27000 56296 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
port 149 nsew signal input
flabel metal2 s 20350 56200 20406 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 150 nsew signal input
flabel metal2 s 21730 56200 21786 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
port 151 nsew signal input
flabel metal2 s 23110 56200 23166 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
port 152 nsew signal input
flabel metal2 s 24490 56200 24546 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
port 153 nsew signal input
flabel metal3 s 0 1776 800 1896 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_0__pin_inpad_0_
port 154 nsew signal tristate
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_1__pin_inpad_0_
port 155 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_2__pin_inpad_0_
port 156 nsew signal tristate
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_3__pin_inpad_0_
port 157 nsew signal tristate
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 test_enable
port 158 nsew signal input
rlabel metal1 13478 54400 13478 54400 0 VGND
rlabel metal1 13478 53856 13478 53856 0 VPWR
rlabel metal1 9890 29070 9890 29070 0 cby_0__8_.cby_0__1_.ccff_tail
rlabel metal1 9752 41582 9752 41582 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 9292 42670 9292 42670 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 9016 44302 9016 44302 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 8280 37978 8280 37978 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 8464 16218 8464 16218 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.ccff_tail
rlabel metal1 15364 12750 15364 12750 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
rlabel metal1 9752 12750 9752 12750 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
rlabel metal1 9660 15538 9660 15538 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
rlabel metal1 8050 14586 8050 14586 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.ccff_tail
rlabel metal1 14858 14484 14858 14484 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
rlabel metal1 13524 10098 13524 10098 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
rlabel metal1 9798 13396 9798 13396 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
rlabel metal1 9200 23154 9200 23154 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.ccff_tail
rlabel metal1 16376 10574 16376 10574 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
rlabel metal1 13294 14450 13294 14450 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
rlabel metal1 10994 20400 10994 20400 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
rlabel metal2 13386 15793 13386 15793 0 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
rlabel metal1 9016 23630 9016 23630 0 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
rlabel metal1 10994 23698 10994 23698 0 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
rlabel metal1 13570 9146 13570 9146 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9200 15674 9200 15674 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 9062 30702 9062 30702 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13846 9418 13846 9418 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14582 10676 14582 10676 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal3 12627 12444 12627 12444 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 12650 13294 12650 13294 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11086 15062 11086 15062 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 10994 14994 10994 14994 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9154 12954 9154 12954 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 10258 12954 10258 12954 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 10166 17238 10166 17238 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 15042 8058 15042 8058 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9062 13498 9062 13498 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 8832 30226 8832 30226 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 15272 8874 15272 8874 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 15134 10234 15134 10234 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13570 11118 13570 11118 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 14398 14246 14398 14246 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12834 9078 12834 9078 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 10626 11696 10626 11696 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9798 11866 9798 11866 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 11546 13158 11546 13158 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 8050 17510 8050 17510 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 13340 12818 13340 12818 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9982 23018 9982 23018 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 9200 23290 9200 23290 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13524 12886 13524 12886 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13616 10506 13616 10506 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 12834 13056 12834 13056 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 12282 16150 12282 16150 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12558 12614 12558 12614 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 12558 14586 12558 14586 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 10258 18394 10258 18394 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 13708 23222 13708 23222 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 9706 22950 9706 22950 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 14352 15436 14352 15436 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10396 23834 10396 23834 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 9200 29274 9200 29274 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13386 16218 13386 16218 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 13110 12104 13110 12104 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12604 12410 12604 12410 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 10534 18496 10534 18496 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11638 16218 11638 16218 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 11592 15674 11592 15674 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 10488 23630 10488 23630 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 13846 24922 13846 24922 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 10120 29138 10120 29138 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 9752 42126 9752 42126 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 11040 44166 11040 44166 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 11224 49130 11224 49130 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel metal1 15502 44778 15502 44778 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 9568 44778 9568 44778 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal2 10810 48994 10810 48994 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal1 10396 49130 10396 49130 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel metal2 15042 46172 15042 46172 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 10166 45050 10166 45050 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal1 9200 44370 9200 44370 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal1 9568 50286 9568 50286 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel metal1 13938 46614 13938 46614 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 7912 50422 7912 50422 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal2 8510 48756 8510 48756 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel metal1 12788 45526 12788 45526 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 25622 51986 25622 51986 0 ccff_head
rlabel metal1 1656 4114 1656 4114 0 ccff_head_0
rlabel metal3 25860 748 25860 748 0 ccff_tail
rlabel metal1 1564 53618 1564 53618 0 ccff_tail_0
rlabel metal1 24702 25466 24702 25466 0 chanx_right_in[0]
rlabel metal2 25346 34391 25346 34391 0 chanx_right_in[10]
rlabel via2 25346 35037 25346 35037 0 chanx_right_in[11]
rlabel metal2 25346 35989 25346 35989 0 chanx_right_in[12]
rlabel metal2 25530 36873 25530 36873 0 chanx_right_in[13]
rlabel metal2 25162 37655 25162 37655 0 chanx_right_in[14]
rlabel via2 25346 38301 25346 38301 0 chanx_right_in[15]
rlabel metal2 25346 39253 25346 39253 0 chanx_right_in[16]
rlabel metal2 25530 40137 25530 40137 0 chanx_right_in[17]
rlabel metal2 25346 40919 25346 40919 0 chanx_right_in[18]
rlabel via2 25162 41565 25162 41565 0 chanx_right_in[19]
rlabel metal2 25346 26061 25346 26061 0 chanx_right_in[1]
rlabel metal2 25162 42483 25162 42483 0 chanx_right_in[20]
rlabel metal2 25530 43401 25530 43401 0 chanx_right_in[21]
rlabel metal2 24794 44183 24794 44183 0 chanx_right_in[22]
rlabel via2 25346 44829 25346 44829 0 chanx_right_in[23]
rlabel metal2 25346 45781 25346 45781 0 chanx_right_in[24]
rlabel metal2 25346 46495 25346 46495 0 chanx_right_in[25]
rlabel metal2 25346 47447 25346 47447 0 chanx_right_in[26]
rlabel via2 25162 48093 25162 48093 0 chanx_right_in[27]
rlabel metal2 25162 49011 25162 49011 0 chanx_right_in[28]
rlabel metal2 25530 49929 25530 49929 0 chanx_right_in[29]
rlabel metal2 24058 27013 24058 27013 0 chanx_right_in[2]
rlabel metal2 24518 28985 24518 28985 0 chanx_right_in[3]
rlabel metal1 23414 29580 23414 29580 0 chanx_right_in[4]
rlabel metal2 25346 29869 25346 29869 0 chanx_right_in[5]
rlabel via2 25530 30923 25530 30923 0 chanx_right_in[6]
rlabel via2 25346 31773 25346 31773 0 chanx_right_in[7]
rlabel metal1 25438 33490 25438 33490 0 chanx_right_in[8]
rlabel metal2 25346 33677 25346 33677 0 chanx_right_in[9]
rlabel metal2 22310 2057 22310 2057 0 chanx_right_out[0]
rlabel metal2 24794 9061 24794 9061 0 chanx_right_out[10]
rlabel metal3 25124 10540 25124 10540 0 chanx_right_out[11]
rlabel metal1 24104 11798 24104 11798 0 chanx_right_out[12]
rlabel metal3 25676 12172 25676 12172 0 chanx_right_out[13]
rlabel metal3 25584 12988 25584 12988 0 chanx_right_out[14]
rlabel metal2 23874 13583 23874 13583 0 chanx_right_out[15]
rlabel metal1 24380 14450 24380 14450 0 chanx_right_out[16]
rlabel metal2 23322 15249 23322 15249 0 chanx_right_out[17]
rlabel metal2 24794 15589 24794 15589 0 chanx_right_out[18]
rlabel metal3 25124 17068 25124 17068 0 chanx_right_out[19]
rlabel metal2 22126 2091 22126 2091 0 chanx_right_out[1]
rlabel metal1 24426 17714 24426 17714 0 chanx_right_out[20]
rlabel metal1 24104 18326 24104 18326 0 chanx_right_out[21]
rlabel metal2 23874 19159 23874 19159 0 chanx_right_out[22]
rlabel metal2 24702 19261 24702 19261 0 chanx_right_out[23]
rlabel metal1 24380 20978 24380 20978 0 chanx_right_out[24]
rlabel metal3 24894 21964 24894 21964 0 chanx_right_out[25]
rlabel metal3 25630 22780 25630 22780 0 chanx_right_out[26]
rlabel metal2 24794 23069 24794 23069 0 chanx_right_out[27]
rlabel metal3 25124 24412 25124 24412 0 chanx_right_out[28]
rlabel metal2 25162 25517 25162 25517 0 chanx_right_out[29]
rlabel metal2 21574 4012 21574 4012 0 chanx_right_out[2]
rlabel metal2 22494 9078 22494 9078 0 chanx_right_out[3]
rlabel metal2 22034 5627 22034 5627 0 chanx_right_out[4]
rlabel metal2 22862 6171 22862 6171 0 chanx_right_out[5]
rlabel metal3 25676 6460 25676 6460 0 chanx_right_out[6]
rlabel metal1 24104 7310 24104 7310 0 chanx_right_out[7]
rlabel metal2 25162 7769 25162 7769 0 chanx_right_out[8]
rlabel metal3 25676 8908 25676 8908 0 chanx_right_out[9]
rlabel metal1 2162 4114 2162 4114 0 chany_bottom_in_0[0]
rlabel metal1 5382 2414 5382 2414 0 chany_bottom_in_0[10]
rlabel metal1 4738 2380 4738 2380 0 chany_bottom_in_0[11]
rlabel metal1 6348 3502 6348 3502 0 chany_bottom_in_0[12]
rlabel metal1 6716 2278 6716 2278 0 chany_bottom_in_0[13]
rlabel metal1 7176 3502 7176 3502 0 chany_bottom_in_0[14]
rlabel metal2 7406 3196 7406 3196 0 chany_bottom_in_0[15]
rlabel metal2 7774 1520 7774 1520 0 chany_bottom_in_0[16]
rlabel metal1 7958 2414 7958 2414 0 chany_bottom_in_0[17]
rlabel metal1 8786 3502 8786 3502 0 chany_bottom_in_0[18]
rlabel metal1 8418 2346 8418 2346 0 chany_bottom_in_0[19]
rlabel metal2 2254 2132 2254 2132 0 chany_bottom_in_0[1]
rlabel metal1 9384 4114 9384 4114 0 chany_bottom_in_0[20]
rlabel metal1 9660 3502 9660 3502 0 chany_bottom_in_0[21]
rlabel metal1 9338 2380 9338 2380 0 chany_bottom_in_0[22]
rlabel metal1 9568 3026 9568 3026 0 chany_bottom_in_0[23]
rlabel metal2 10718 1761 10718 1761 0 chany_bottom_in_0[24]
rlabel metal1 10534 3060 10534 3060 0 chany_bottom_in_0[25]
rlabel metal2 11454 1761 11454 1761 0 chany_bottom_in_0[26]
rlabel metal2 11178 3740 11178 3740 0 chany_bottom_in_0[27]
rlabel metal1 11914 2448 11914 2448 0 chany_bottom_in_0[28]
rlabel metal2 12558 3740 12558 3740 0 chany_bottom_in_0[29]
rlabel metal1 2392 3026 2392 3026 0 chany_bottom_in_0[2]
rlabel metal1 2806 2414 2806 2414 0 chany_bottom_in_0[3]
rlabel metal2 3358 1761 3358 1761 0 chany_bottom_in_0[4]
rlabel metal2 2898 3740 2898 3740 0 chany_bottom_in_0[5]
rlabel metal1 4232 4114 4232 4114 0 chany_bottom_in_0[6]
rlabel metal1 4508 3162 4508 3162 0 chany_bottom_in_0[7]
rlabel metal2 4830 1761 4830 1761 0 chany_bottom_in_0[8]
rlabel metal1 5796 2278 5796 2278 0 chany_bottom_in_0[9]
rlabel metal2 12926 1231 12926 1231 0 chany_bottom_out_0[0]
rlabel metal1 17894 3094 17894 3094 0 chany_bottom_out_0[10]
rlabel metal1 18676 2890 18676 2890 0 chany_bottom_out_0[11]
rlabel metal2 17342 1503 17342 1503 0 chany_bottom_out_0[12]
rlabel metal1 18814 3570 18814 3570 0 chany_bottom_out_0[13]
rlabel metal2 18078 823 18078 823 0 chany_bottom_out_0[14]
rlabel metal1 22356 2482 22356 2482 0 chany_bottom_out_0[15]
rlabel metal2 18814 1231 18814 1231 0 chany_bottom_out_0[16]
rlabel metal2 19182 1761 19182 1761 0 chany_bottom_out_0[17]
rlabel metal2 19550 2438 19550 2438 0 chany_bottom_out_0[18]
rlabel metal2 19918 1095 19918 1095 0 chany_bottom_out_0[19]
rlabel metal2 13294 1554 13294 1554 0 chany_bottom_out_0[1]
rlabel metal2 20378 5372 20378 5372 0 chany_bottom_out_0[20]
rlabel metal2 20654 1761 20654 1761 0 chany_bottom_out_0[21]
rlabel metal2 21022 2370 21022 2370 0 chany_bottom_out_0[22]
rlabel metal2 21390 2948 21390 2948 0 chany_bottom_out_0[23]
rlabel metal1 21528 6222 21528 6222 0 chany_bottom_out_0[24]
rlabel metal2 22126 823 22126 823 0 chany_bottom_out_0[25]
rlabel metal1 22540 8398 22540 8398 0 chany_bottom_out_0[26]
rlabel metal2 21482 5576 21482 5576 0 chany_bottom_out_0[27]
rlabel metal2 23230 1010 23230 1010 0 chany_bottom_out_0[28]
rlabel metal2 23598 1299 23598 1299 0 chany_bottom_out_0[29]
rlabel metal2 13662 1860 13662 1860 0 chany_bottom_out_0[2]
rlabel metal1 14398 3570 14398 3570 0 chany_bottom_out_0[3]
rlabel metal2 14398 1622 14398 1622 0 chany_bottom_out_0[4]
rlabel metal1 15042 2958 15042 2958 0 chany_bottom_out_0[5]
rlabel metal1 16238 2822 16238 2822 0 chany_bottom_out_0[6]
rlabel metal1 16054 3570 16054 3570 0 chany_bottom_out_0[7]
rlabel metal1 16606 2958 16606 2958 0 chany_bottom_out_0[8]
rlabel metal1 16790 4046 16790 4046 0 chany_bottom_out_0[9]
rlabel metal1 21758 32198 21758 32198 0 clknet_0_prog_clk
rlabel metal1 9798 14382 9798 14382 0 clknet_4_0_0_prog_clk
rlabel metal1 6670 48586 6670 48586 0 clknet_4_10_0_prog_clk
rlabel metal2 16790 32062 16790 32062 0 clknet_4_11_0_prog_clk
rlabel metal1 18170 20570 18170 20570 0 clknet_4_12_0_prog_clk
rlabel metal1 23322 21556 23322 21556 0 clknet_4_13_0_prog_clk
rlabel metal2 19458 31994 19458 31994 0 clknet_4_14_0_prog_clk
rlabel metal1 19964 43758 19964 43758 0 clknet_4_15_0_prog_clk
rlabel metal1 13662 13362 13662 13362 0 clknet_4_1_0_prog_clk
rlabel metal1 7958 23698 7958 23698 0 clknet_4_2_0_prog_clk
rlabel metal1 11546 24242 11546 24242 0 clknet_4_3_0_prog_clk
rlabel metal2 16882 13129 16882 13129 0 clknet_4_4_0_prog_clk
rlabel metal1 22908 12750 22908 12750 0 clknet_4_5_0_prog_clk
rlabel metal1 15916 20978 15916 20978 0 clknet_4_6_0_prog_clk
rlabel metal1 23414 19380 23414 19380 0 clknet_4_7_0_prog_clk
rlabel metal2 11454 29138 11454 29138 0 clknet_4_8_0_prog_clk
rlabel metal1 10281 26214 10281 26214 0 clknet_4_9_0_prog_clk
rlabel metal1 2484 54094 2484 54094 0 gfpga_pad_io_soc_dir[0]
rlabel metal1 4140 53618 4140 53618 0 gfpga_pad_io_soc_dir[1]
rlabel metal2 5198 55158 5198 55158 0 gfpga_pad_io_soc_dir[2]
rlabel metal2 6578 54920 6578 54920 0 gfpga_pad_io_soc_dir[3]
rlabel metal2 13662 56236 13662 56236 0 gfpga_pad_io_soc_in[0]
rlabel metal1 14996 54162 14996 54162 0 gfpga_pad_io_soc_in[1]
rlabel metal1 16836 54162 16836 54162 0 gfpga_pad_io_soc_in[2]
rlabel metal1 17756 54162 17756 54162 0 gfpga_pad_io_soc_in[3]
rlabel metal2 7958 55711 7958 55711 0 gfpga_pad_io_soc_out[0]
rlabel metal1 9614 54094 9614 54094 0 gfpga_pad_io_soc_out[1]
rlabel metal1 10718 53652 10718 53652 0 gfpga_pad_io_soc_out[2]
rlabel metal2 12282 56236 12282 56236 0 gfpga_pad_io_soc_out[3]
rlabel metal1 19228 54162 19228 54162 0 isol_n
rlabel metal1 25024 51782 25024 51782 0 net1
rlabel metal2 21942 35564 21942 35564 0 net10
rlabel metal2 22126 22780 22126 22780 0 net100
rlabel metal2 23782 22644 23782 22644 0 net101
rlabel metal1 23414 22610 23414 22610 0 net102
rlabel metal1 21482 25432 21482 25432 0 net103
rlabel metal2 23966 25670 23966 25670 0 net104
rlabel metal1 13524 4658 13524 4658 0 net105
rlabel metal1 15778 5236 15778 5236 0 net106
rlabel metal1 18262 6324 18262 6324 0 net107
rlabel metal1 21275 13430 21275 13430 0 net108
rlabel metal1 23644 2550 23644 2550 0 net109
rlabel metal1 23598 31790 23598 31790 0 net11
rlabel metal2 23828 13940 23828 13940 0 net110
rlabel metal1 15502 4216 15502 4216 0 net111
rlabel via2 12282 4709 12282 4709 0 net112
rlabel metal1 19826 13838 19826 13838 0 net113
rlabel metal1 18952 3026 18952 3026 0 net114
rlabel metal1 19688 2414 19688 2414 0 net115
rlabel metal1 17618 4556 17618 4556 0 net116
rlabel metal2 19458 6188 19458 6188 0 net117
rlabel metal2 18814 5780 18814 5780 0 net118
rlabel metal1 18676 2346 18676 2346 0 net119
rlabel metal1 25346 32878 25346 32878 0 net12
rlabel metal1 21068 3502 21068 3502 0 net120
rlabel metal2 19642 8364 19642 8364 0 net121
rlabel metal1 25162 18666 25162 18666 0 net122
rlabel metal1 22402 4624 22402 4624 0 net123
rlabel metal1 15364 2346 15364 2346 0 net124
rlabel metal2 22126 5644 22126 5644 0 net125
rlabel metal1 21206 5678 21206 5678 0 net126
rlabel metal1 21689 5066 21689 5066 0 net127
rlabel metal1 23828 5202 23828 5202 0 net128
rlabel metal2 20286 6086 20286 6086 0 net129
rlabel via2 13570 14229 13570 14229 0 net13
rlabel metal1 20562 3162 20562 3162 0 net130
rlabel metal2 22126 3910 22126 3910 0 net131
rlabel metal1 20470 7922 20470 7922 0 net132
rlabel metal2 20102 5712 20102 5712 0 net133
rlabel metal2 12282 4335 12282 4335 0 net134
rlabel via3 17181 16660 17181 16660 0 net135
rlabel metal3 17181 15300 17181 15300 0 net136
rlabel metal1 14858 2414 14858 2414 0 net137
rlabel metal1 14490 3026 14490 3026 0 net138
rlabel metal1 16836 2414 16836 2414 0 net139
rlabel metal2 25162 23936 25162 23936 0 net14
rlabel metal1 16698 3502 16698 3502 0 net140
rlabel metal1 18354 13362 18354 13362 0 net141
rlabel metal1 18906 13226 18906 13226 0 net142
rlabel metal1 4646 53210 4646 53210 0 net143
rlabel metal1 5382 52666 5382 52666 0 net144
rlabel metal2 4830 52768 4830 52768 0 net145
rlabel metal1 8556 51510 8556 51510 0 net146
rlabel metal1 7866 51578 7866 51578 0 net147
rlabel metal2 9614 52326 9614 52326 0 net148
rlabel metal2 10718 51442 10718 51442 0 net149
rlabel metal2 20148 13260 20148 13260 0 net15
rlabel metal2 11730 51748 11730 51748 0 net150
rlabel metal1 18262 26010 18262 26010 0 net151
rlabel metal1 17940 27438 17940 27438 0 net152
rlabel metal1 24840 17510 24840 17510 0 net153
rlabel metal2 19734 28288 19734 28288 0 net154
rlabel metal1 22862 26962 22862 26962 0 net155
rlabel metal2 24978 28798 24978 28798 0 net156
rlabel metal1 21850 30226 21850 30226 0 net157
rlabel metal1 20194 30362 20194 30362 0 net158
rlabel metal2 19182 29376 19182 29376 0 net159
rlabel metal1 19044 14042 19044 14042 0 net16
rlabel metal1 21942 19346 21942 19346 0 net160
rlabel metal1 21988 17170 21988 17170 0 net161
rlabel metal1 19688 22746 19688 22746 0 net162
rlabel metal2 22034 21250 22034 21250 0 net163
rlabel metal1 7636 17306 7636 17306 0 net164
rlabel metal1 7222 12274 7222 12274 0 net165
rlabel metal2 8234 12546 8234 12546 0 net166
rlabel metal1 13478 17646 13478 17646 0 net167
rlabel metal2 13202 17408 13202 17408 0 net168
rlabel metal1 15640 16218 15640 16218 0 net169
rlabel metal1 15916 18394 15916 18394 0 net17
rlabel metal2 9982 21250 9982 21250 0 net170
rlabel metal1 13524 10778 13524 10778 0 net171
rlabel metal2 12650 7616 12650 7616 0 net172
rlabel metal1 15410 7854 15410 7854 0 net173
rlabel metal1 17296 14314 17296 14314 0 net174
rlabel metal1 14214 15130 14214 15130 0 net175
rlabel metal1 15962 16558 15962 16558 0 net176
rlabel metal1 15870 15130 15870 15130 0 net177
rlabel metal2 13386 8126 13386 8126 0 net178
rlabel metal1 16008 5542 16008 5542 0 net179
rlabel metal1 24104 35054 24104 35054 0 net18
rlabel metal1 17250 4250 17250 4250 0 net180
rlabel metal1 11408 21658 11408 21658 0 net181
rlabel metal1 21068 7446 21068 7446 0 net182
rlabel metal1 21574 9690 21574 9690 0 net183
rlabel metal2 18446 11968 18446 11968 0 net184
rlabel metal1 18952 12274 18952 12274 0 net185
rlabel metal2 20010 11390 20010 11390 0 net186
rlabel metal2 24242 8126 24242 8126 0 net187
rlabel metal1 23736 3162 23736 3162 0 net188
rlabel metal1 21114 3162 21114 3162 0 net189
rlabel metal1 23690 35802 23690 35802 0 net19
rlabel metal1 23920 3570 23920 3570 0 net190
rlabel metal1 11592 7854 11592 7854 0 net191
rlabel metal2 11730 19584 11730 19584 0 net192
rlabel metal2 9430 17408 9430 17408 0 net193
rlabel metal1 10948 12954 10948 12954 0 net194
rlabel metal2 12098 10302 12098 10302 0 net195
rlabel metal1 15410 23086 15410 23086 0 net196
rlabel metal1 15640 25874 15640 25874 0 net197
rlabel metal1 20332 21522 20332 21522 0 net198
rlabel metal1 24058 21930 24058 21930 0 net199
rlabel metal1 1610 4012 1610 4012 0 net2
rlabel metal1 23322 35734 23322 35734 0 net20
rlabel metal1 24380 24242 24380 24242 0 net200
rlabel metal1 20792 23154 20792 23154 0 net201
rlabel metal2 18538 24650 18538 24650 0 net202
rlabel metal1 25254 29206 25254 29206 0 net21
rlabel via2 16882 16235 16882 16235 0 net22
rlabel via2 17434 17323 17434 17323 0 net23
rlabel metal1 20102 25194 20102 25194 0 net24
rlabel metal1 25024 20978 25024 20978 0 net25
rlabel metal1 24702 23154 24702 23154 0 net26
rlabel metal1 22586 26010 22586 26010 0 net27
rlabel metal1 23230 26350 23230 26350 0 net28
rlabel metal1 25116 26282 25116 26282 0 net29
rlabel metal2 22724 21148 22724 21148 0 net3
rlabel metal1 25116 31926 25116 31926 0 net30
rlabel metal1 25300 33286 25300 33286 0 net31
rlabel metal1 25714 33830 25714 33830 0 net32
rlabel metal2 2254 5848 2254 5848 0 net33
rlabel via2 5474 2499 5474 2499 0 net34
rlabel metal1 8234 2618 8234 2618 0 net35
rlabel metal2 6394 4964 6394 4964 0 net36
rlabel metal1 8602 3162 8602 3162 0 net37
rlabel metal1 13984 12818 13984 12818 0 net38
rlabel metal2 7222 7072 7222 7072 0 net39
rlabel metal1 20700 29546 20700 29546 0 net4
rlabel metal1 15778 13294 15778 13294 0 net40
rlabel metal2 8418 2108 8418 2108 0 net41
rlabel metal1 9660 3706 9660 3706 0 net42
rlabel metal1 7176 2278 7176 2278 0 net43
rlabel metal1 5750 17102 5750 17102 0 net44
rlabel metal1 14122 6698 14122 6698 0 net45
rlabel metal2 14260 7548 14260 7548 0 net46
rlabel metal1 10396 2278 10396 2278 0 net47
rlabel metal1 15226 9894 15226 9894 0 net48
rlabel metal1 16698 12886 16698 12886 0 net49
rlabel metal1 24334 17578 24334 17578 0 net5
rlabel metal1 17664 8806 17664 8806 0 net50
rlabel metal3 14766 12444 14766 12444 0 net51
rlabel metal1 19596 10642 19596 10642 0 net52
rlabel metal1 16277 7854 16277 7854 0 net53
rlabel metal1 14720 8806 14720 8806 0 net54
rlabel metal1 2438 2924 2438 2924 0 net55
rlabel metal1 2898 2516 2898 2516 0 net56
rlabel metal2 11270 16133 11270 16133 0 net57
rlabel metal1 1886 3468 1886 3468 0 net58
rlabel metal1 7038 12750 7038 12750 0 net59
rlabel metal1 25668 18734 25668 18734 0 net6
rlabel metal1 8004 12750 8004 12750 0 net60
rlabel via2 12742 17493 12742 17493 0 net61
rlabel via1 13846 15997 13846 15997 0 net62
rlabel metal1 13524 53958 13524 53958 0 net63
rlabel metal2 13938 50286 13938 50286 0 net64
rlabel metal2 15686 50014 15686 50014 0 net65
rlabel metal1 15916 44914 15916 44914 0 net66
rlabel metal1 18262 54162 18262 54162 0 net67
rlabel metal1 22717 19754 22717 19754 0 net68
rlabel metal1 13432 11254 13432 11254 0 net69
rlabel metal2 16146 13124 16146 13124 0 net7
rlabel metal1 26128 51306 26128 51306 0 net70
rlabel metal2 17986 31756 17986 31756 0 net71
rlabel metal2 15640 45540 15640 45540 0 net72
rlabel metal1 25898 53414 25898 53414 0 net73
rlabel metal2 20102 21760 20102 21760 0 net74
rlabel metal2 24518 52768 24518 52768 0 net75
rlabel metal1 23046 53414 23046 53414 0 net76
rlabel metal1 16974 33082 16974 33082 0 net77
rlabel metal1 19504 22066 19504 22066 0 net78
rlabel metal1 23046 53958 23046 53958 0 net79
rlabel metal2 16330 12801 16330 12801 0 net8
rlabel metal2 16882 32878 16882 32878 0 net80
rlabel metal1 23276 17102 23276 17102 0 net81
rlabel metal1 1794 53516 1794 53516 0 net82
rlabel metal1 15870 6290 15870 6290 0 net83
rlabel metal1 15134 8500 15134 8500 0 net84
rlabel metal1 23184 11118 23184 11118 0 net85
rlabel metal1 24288 9146 24288 9146 0 net86
rlabel metal1 23966 11322 23966 11322 0 net87
rlabel metal1 24564 11730 24564 11730 0 net88
rlabel metal1 23184 13294 23184 13294 0 net89
rlabel metal2 25116 34918 25116 34918 0 net9
rlabel metal1 24564 13498 24564 13498 0 net90
rlabel metal2 22862 13022 22862 13022 0 net91
rlabel metal1 24380 12410 24380 12410 0 net92
rlabel metal2 22402 15198 22402 15198 0 net93
rlabel metal1 9890 2482 9890 2482 0 net94
rlabel metal2 24610 17204 24610 17204 0 net95
rlabel metal2 22126 18428 22126 18428 0 net96
rlabel metal2 22770 19482 22770 19482 0 net97
rlabel metal1 23828 18258 23828 18258 0 net98
rlabel metal1 22402 20910 22402 20910 0 net99
rlabel metal2 18906 23970 18906 23970 0 prog_clk
rlabel metal1 24518 2618 24518 2618 0 prog_reset
rlabel metal2 24978 50711 24978 50711 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel via2 24978 51323 24978 51323 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
rlabel metal2 24978 52275 24978 52275 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel metal2 25070 53023 25070 53023 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 25070 53669 25070 53669 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal1 24564 53754 24564 53754 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
rlabel metal3 25584 55420 25584 55420 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
rlabel via2 23437 56100 23437 56100 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
rlabel metal2 20562 56236 20562 56236 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 21896 54162 21896 54162 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 23184 54162 23184 54162 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 24564 54162 24564 54162 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 18768 44778 18768 44778 0 right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 23782 19890 23782 19890 0 right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 21114 35564 21114 35564 0 right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 18446 21318 18446 21318 0 right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 18630 15640 18630 15640 0 sb_0__8_.mem_bottom_track_1.ccff_head
rlabel metal2 21666 19482 21666 19482 0 sb_0__8_.mem_bottom_track_1.ccff_tail
rlabel metal2 20194 18530 20194 18530 0 sb_0__8_.mem_bottom_track_1.mem_out\[0\]
rlabel metal1 23138 21318 23138 21318 0 sb_0__8_.mem_bottom_track_11.ccff_head
rlabel metal1 25438 24718 25438 24718 0 sb_0__8_.mem_bottom_track_11.ccff_tail
rlabel metal1 25116 23834 25116 23834 0 sb_0__8_.mem_bottom_track_11.mem_out\[0\]
rlabel metal2 22402 27608 22402 27608 0 sb_0__8_.mem_bottom_track_13.ccff_tail
rlabel metal1 25162 27540 25162 27540 0 sb_0__8_.mem_bottom_track_13.mem_out\[0\]
rlabel metal1 20700 26418 20700 26418 0 sb_0__8_.mem_bottom_track_15.ccff_tail
rlabel metal1 23506 28594 23506 28594 0 sb_0__8_.mem_bottom_track_15.mem_out\[0\]
rlabel metal1 19366 26758 19366 26758 0 sb_0__8_.mem_bottom_track_17.ccff_tail
rlabel metal2 22586 27438 22586 27438 0 sb_0__8_.mem_bottom_track_17.mem_out\[0\]
rlabel metal1 18768 29818 18768 29818 0 sb_0__8_.mem_bottom_track_19.ccff_tail
rlabel metal2 18906 29172 18906 29172 0 sb_0__8_.mem_bottom_track_19.mem_out\[0\]
rlabel metal1 18124 31858 18124 31858 0 sb_0__8_.mem_bottom_track_29.ccff_tail
rlabel metal1 17795 31994 17795 31994 0 sb_0__8_.mem_bottom_track_29.mem_out\[0\]
rlabel metal2 25162 19924 25162 19924 0 sb_0__8_.mem_bottom_track_3.ccff_tail
rlabel metal1 23920 20026 23920 20026 0 sb_0__8_.mem_bottom_track_3.mem_out\[0\]
rlabel metal2 21022 29614 21022 29614 0 sb_0__8_.mem_bottom_track_31.ccff_tail
rlabel metal1 20240 31858 20240 31858 0 sb_0__8_.mem_bottom_track_31.mem_out\[0\]
rlabel metal1 23644 30158 23644 30158 0 sb_0__8_.mem_bottom_track_33.ccff_tail
rlabel metal1 23046 31824 23046 31824 0 sb_0__8_.mem_bottom_track_33.mem_out\[0\]
rlabel metal1 25162 32538 25162 32538 0 sb_0__8_.mem_bottom_track_35.ccff_tail
rlabel metal1 24380 32334 24380 32334 0 sb_0__8_.mem_bottom_track_35.mem_out\[0\]
rlabel metal1 22011 33898 22011 33898 0 sb_0__8_.mem_bottom_track_45.ccff_tail
rlabel metal1 22356 33422 22356 33422 0 sb_0__8_.mem_bottom_track_45.mem_out\[0\]
rlabel via1 20562 33422 20562 33422 0 sb_0__8_.mem_bottom_track_47.ccff_tail
rlabel metal1 19826 33592 19826 33592 0 sb_0__8_.mem_bottom_track_47.mem_out\[0\]
rlabel metal1 20884 32198 20884 32198 0 sb_0__8_.mem_bottom_track_49.ccff_tail
rlabel metal2 21206 33082 21206 33082 0 sb_0__8_.mem_bottom_track_49.mem_out\[0\]
rlabel metal1 24196 21658 24196 21658 0 sb_0__8_.mem_bottom_track_5.ccff_tail
rlabel metal1 24472 21454 24472 21454 0 sb_0__8_.mem_bottom_track_5.mem_out\[0\]
rlabel metal1 24012 17102 24012 17102 0 sb_0__8_.mem_bottom_track_51.mem_out\[0\]
rlabel metal1 20838 24378 20838 24378 0 sb_0__8_.mem_bottom_track_7.ccff_tail
rlabel metal1 23092 22066 23092 22066 0 sb_0__8_.mem_bottom_track_7.mem_out\[0\]
rlabel metal2 22402 25568 22402 25568 0 sb_0__8_.mem_bottom_track_9.mem_out\[0\]
rlabel metal1 11454 26554 11454 26554 0 sb_0__8_.mem_right_track_0.ccff_tail
rlabel metal2 16146 32402 16146 32402 0 sb_0__8_.mem_right_track_0.mem_out\[0\]
rlabel metal2 12374 30090 12374 30090 0 sb_0__8_.mem_right_track_0.mem_out\[1\]
rlabel metal1 10994 24038 10994 24038 0 sb_0__8_.mem_right_track_10.ccff_head
rlabel metal1 8372 19142 8372 19142 0 sb_0__8_.mem_right_track_10.ccff_tail
rlabel metal1 11178 24616 11178 24616 0 sb_0__8_.mem_right_track_10.mem_out\[0\]
rlabel metal1 8418 22406 8418 22406 0 sb_0__8_.mem_right_track_10.mem_out\[1\]
rlabel metal2 10902 19244 10902 19244 0 sb_0__8_.mem_right_track_12.ccff_tail
rlabel metal1 10672 23222 10672 23222 0 sb_0__8_.mem_right_track_12.mem_out\[0\]
rlabel metal1 13754 21658 13754 21658 0 sb_0__8_.mem_right_track_14.ccff_tail
rlabel metal1 12926 21046 12926 21046 0 sb_0__8_.mem_right_track_14.mem_out\[0\]
rlabel metal2 14490 19754 14490 19754 0 sb_0__8_.mem_right_track_16.ccff_tail
rlabel metal1 13248 20366 13248 20366 0 sb_0__8_.mem_right_track_16.mem_out\[0\]
rlabel metal1 13616 16422 13616 16422 0 sb_0__8_.mem_right_track_18.ccff_tail
rlabel metal1 15134 15980 15134 15980 0 sb_0__8_.mem_right_track_18.mem_out\[0\]
rlabel metal2 11086 28322 11086 28322 0 sb_0__8_.mem_right_track_2.ccff_tail
rlabel metal1 11822 27880 11822 27880 0 sb_0__8_.mem_right_track_2.mem_out\[0\]
rlabel metal2 9614 27166 9614 27166 0 sb_0__8_.mem_right_track_2.mem_out\[1\]
rlabel metal1 12650 10574 12650 10574 0 sb_0__8_.mem_right_track_20.ccff_tail
rlabel metal2 12190 12789 12190 12789 0 sb_0__8_.mem_right_track_20.mem_out\[0\]
rlabel metal1 12834 7276 12834 7276 0 sb_0__8_.mem_right_track_22.ccff_tail
rlabel metal2 10994 7514 10994 7514 0 sb_0__8_.mem_right_track_22.mem_out\[0\]
rlabel metal2 12558 8160 12558 8160 0 sb_0__8_.mem_right_track_24.ccff_tail
rlabel metal1 11592 5882 11592 5882 0 sb_0__8_.mem_right_track_24.mem_out\[0\]
rlabel metal1 15226 14042 15226 14042 0 sb_0__8_.mem_right_track_26.ccff_tail
rlabel metal1 14352 12750 14352 12750 0 sb_0__8_.mem_right_track_26.mem_out\[0\]
rlabel metal1 15916 20026 15916 20026 0 sb_0__8_.mem_right_track_28.ccff_tail
rlabel metal1 15870 16966 15870 16966 0 sb_0__8_.mem_right_track_28.mem_out\[0\]
rlabel metal2 17158 21182 17158 21182 0 sb_0__8_.mem_right_track_30.ccff_tail
rlabel metal1 16698 20774 16698 20774 0 sb_0__8_.mem_right_track_30.mem_out\[0\]
rlabel metal1 18538 17714 18538 17714 0 sb_0__8_.mem_right_track_32.ccff_tail
rlabel metal1 17112 18326 17112 18326 0 sb_0__8_.mem_right_track_32.mem_out\[0\]
rlabel metal2 16698 9282 16698 9282 0 sb_0__8_.mem_right_track_34.ccff_tail
rlabel metal1 18032 15674 18032 15674 0 sb_0__8_.mem_right_track_34.mem_out\[0\]
rlabel metal1 14582 4998 14582 4998 0 sb_0__8_.mem_right_track_36.ccff_tail
rlabel metal1 13938 6188 13938 6188 0 sb_0__8_.mem_right_track_36.mem_out\[0\]
rlabel metal1 16737 5882 16737 5882 0 sb_0__8_.mem_right_track_38.ccff_tail
rlabel metal2 15410 5678 15410 5678 0 sb_0__8_.mem_right_track_38.mem_out\[0\]
rlabel metal1 13662 28594 13662 28594 0 sb_0__8_.mem_right_track_4.ccff_tail
rlabel metal2 12098 29988 12098 29988 0 sb_0__8_.mem_right_track_4.mem_out\[0\]
rlabel metal1 11546 28458 11546 28458 0 sb_0__8_.mem_right_track_4.mem_out\[1\]
rlabel metal1 21298 7276 21298 7276 0 sb_0__8_.mem_right_track_40.ccff_tail
rlabel metal1 17572 5882 17572 5882 0 sb_0__8_.mem_right_track_40.mem_out\[0\]
rlabel metal2 21298 11424 21298 11424 0 sb_0__8_.mem_right_track_42.ccff_tail
rlabel metal2 20838 10608 20838 10608 0 sb_0__8_.mem_right_track_42.mem_out\[0\]
rlabel metal1 20884 15334 20884 15334 0 sb_0__8_.mem_right_track_44.ccff_tail
rlabel metal2 19734 18190 19734 18190 0 sb_0__8_.mem_right_track_44.mem_out\[0\]
rlabel metal1 23184 15538 23184 15538 0 sb_0__8_.mem_right_track_46.ccff_tail
rlabel metal1 22540 16014 22540 16014 0 sb_0__8_.mem_right_track_46.mem_out\[0\]
rlabel metal2 23414 13668 23414 13668 0 sb_0__8_.mem_right_track_48.ccff_tail
rlabel metal2 23414 18463 23414 18463 0 sb_0__8_.mem_right_track_48.mem_out\[0\]
rlabel metal2 23414 10268 23414 10268 0 sb_0__8_.mem_right_track_50.ccff_tail
rlabel metal1 24058 12614 24058 12614 0 sb_0__8_.mem_right_track_50.mem_out\[0\]
rlabel metal2 23874 7004 23874 7004 0 sb_0__8_.mem_right_track_52.ccff_tail
rlabel metal3 21298 9996 21298 9996 0 sb_0__8_.mem_right_track_52.mem_out\[0\]
rlabel metal1 21252 4794 21252 4794 0 sb_0__8_.mem_right_track_54.ccff_tail
rlabel metal1 21942 6834 21942 6834 0 sb_0__8_.mem_right_track_54.mem_out\[0\]
rlabel metal1 17756 7310 17756 7310 0 sb_0__8_.mem_right_track_56.ccff_tail
rlabel metal1 18860 7310 18860 7310 0 sb_0__8_.mem_right_track_56.mem_out\[0\]
rlabel metal1 17335 13702 17335 13702 0 sb_0__8_.mem_right_track_58.mem_out\[0\]
rlabel metal1 13846 24038 13846 24038 0 sb_0__8_.mem_right_track_6.ccff_tail
rlabel metal1 13432 27030 13432 27030 0 sb_0__8_.mem_right_track_6.mem_out\[0\]
rlabel metal1 12144 24106 12144 24106 0 sb_0__8_.mem_right_track_6.mem_out\[1\]
rlabel metal2 14766 25024 14766 25024 0 sb_0__8_.mem_right_track_8.mem_out\[0\]
rlabel metal1 9384 24106 9384 24106 0 sb_0__8_.mem_right_track_8.mem_out\[1\]
rlabel metal2 14674 10336 14674 10336 0 sb_0__8_.mux_bottom_track_1.out
rlabel metal1 20654 19482 20654 19482 0 sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 20470 20400 20470 20400 0 sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18998 15062 18998 15062 0 sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18170 10642 18170 10642 0 sb_0__8_.mux_bottom_track_11.out
rlabel metal1 24840 26486 24840 26486 0 sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24334 21862 24334 21862 0 sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 19596 11186 19596 11186 0 sb_0__8_.mux_bottom_track_13.out
rlabel metal1 23046 24786 23046 24786 0 sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22264 18156 22264 18156 0 sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16698 9622 16698 9622 0 sb_0__8_.mux_bottom_track_15.out
rlabel metal2 20930 25092 20930 25092 0 sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 20608 19890 20608 19890 0 sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 19826 9010 19826 9010 0 sb_0__8_.mux_bottom_track_17.out
rlabel metal1 19688 24038 19688 24038 0 sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18262 16082 18262 16082 0 sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17572 13532 17572 13532 0 sb_0__8_.mux_bottom_track_19.out
rlabel metal1 18354 25942 18354 25942 0 sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17066 26010 17066 26010 0 sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15640 19482 15640 19482 0 sb_0__8_.mux_bottom_track_29.out
rlabel metal1 17802 27302 17802 27302 0 sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16330 19346 16330 19346 0 sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 22034 6664 22034 6664 0 sb_0__8_.mux_bottom_track_3.out
rlabel metal1 25070 17748 25070 17748 0 sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24104 17510 24104 17510 0 sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 18492 15980 18492 15980 0 sb_0__8_.mux_bottom_track_31.out
rlabel metal2 21666 30022 21666 30022 0 sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19274 19822 19274 19822 0 sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21344 18054 21344 18054 0 sb_0__8_.mux_bottom_track_33.out
rlabel metal1 22908 31926 22908 31926 0 sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22172 19924 22172 19924 0 sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21344 18598 21344 18598 0 sb_0__8_.mux_bottom_track_35.out
rlabel metal1 24840 28458 24840 28458 0 sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21482 18802 21482 18802 0 sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19642 20230 19642 20230 0 sb_0__8_.mux_bottom_track_45.out
rlabel metal1 22678 34918 22678 34918 0 sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21436 20434 21436 20434 0 sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17986 9962 17986 9962 0 sb_0__8_.mux_bottom_track_47.out
rlabel metal2 22034 33601 22034 33601 0 sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19412 20434 19412 20434 0 sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 15732 13260 15732 13260 0 sb_0__8_.mux_bottom_track_49.out
rlabel metal1 20056 35530 20056 35530 0 sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17388 21454 17388 21454 0 sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21942 13515 21942 13515 0 sb_0__8_.mux_bottom_track_5.out
rlabel metal1 22632 19482 22632 19482 0 sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22356 19482 22356 19482 0 sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13386 9894 13386 9894 0 sb_0__8_.mux_bottom_track_51.out
rlabel metal1 23598 17306 23598 17306 0 sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22448 16966 22448 16966 0 sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14996 14756 14996 14756 0 sb_0__8_.mux_bottom_track_7.out
rlabel metal2 20010 24446 20010 24446 0 sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19596 23086 19596 23086 0 sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 19136 20434 19136 20434 0 sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 17526 8704 17526 8704 0 sb_0__8_.mux_bottom_track_9.out
rlabel metal1 22586 26486 22586 26486 0 sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21114 14382 21114 14382 0 sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21758 25296 21758 25296 0 sb_0__8_.mux_right_track_0.out
rlabel metal1 14122 32742 14122 32742 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14076 31926 14076 31926 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12236 24786 12236 24786 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 11684 24854 11684 24854 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 14582 24684 14582 24684 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 15180 19210 15180 19210 0 sb_0__8_.mux_right_track_10.out
rlabel metal2 11730 24310 11730 24310 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11730 23018 11730 23018 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10902 22950 10902 22950 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 6854 12954 6854 12954 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 15226 19414 15226 19414 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 22218 20230 22218 20230 0 sb_0__8_.mux_right_track_12.out
rlabel metal1 12604 22950 12604 22950 0 sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9614 12682 9614 12682 0 sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 15870 19380 15870 19380 0 sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22954 20468 22954 20468 0 sb_0__8_.mux_right_track_14.out
rlabel metal1 15548 22134 15548 22134 0 sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15226 19856 15226 19856 0 sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14858 21726 14858 21726 0 sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 21574 19074 21574 19074 0 sb_0__8_.mux_right_track_16.out
rlabel metal1 16192 24582 16192 24582 0 sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13248 17034 13248 17034 0 sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 19182 19822 19182 19822 0 sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 24794 16524 24794 16524 0 sb_0__8_.mux_right_track_18.out
rlabel metal1 14812 16218 14812 16218 0 sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18538 16558 18538 16558 0 sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21022 25296 21022 25296 0 sb_0__8_.mux_right_track_2.out
rlabel metal1 14168 27438 14168 27438 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13616 27370 13616 27370 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12650 26656 12650 26656 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 12558 23596 12558 23596 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 12305 25738 12305 25738 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 22310 13396 22310 13396 0 sb_0__8_.mux_right_track_20.out
rlabel metal2 12834 10982 12834 10982 0 sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16514 12750 16514 12750 0 sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 16882 10336 16882 10336 0 sb_0__8_.mux_right_track_22.out
rlabel metal1 10948 6426 10948 6426 0 sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14352 7446 14352 7446 0 sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20378 11662 20378 11662 0 sb_0__8_.mux_right_track_24.out
rlabel metal2 13386 7072 13386 7072 0 sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14674 7718 14674 7718 0 sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24196 13294 24196 13294 0 sb_0__8_.mux_right_track_26.out
rlabel metal1 15226 12614 15226 12614 0 sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 20378 14212 20378 14212 0 sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 24426 14110 24426 14110 0 sb_0__8_.mux_right_track_28.out
rlabel metal1 17112 23494 17112 23494 0 sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15226 14858 15226 14858 0 sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19688 17646 19688 17646 0 sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 24702 14518 24702 14518 0 sb_0__8_.mux_right_track_30.out
rlabel metal2 17940 19890 17940 19890 0 sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15870 16422 15870 16422 0 sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21022 17680 21022 17680 0 sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 24610 15402 24610 15402 0 sb_0__8_.mux_right_track_32.out
rlabel metal1 18676 17578 18676 17578 0 sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15594 16354 15594 16354 0 sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21850 16660 21850 16660 0 sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 23782 10098 23782 10098 0 sb_0__8_.mux_right_track_34.out
rlabel metal1 16836 18598 16836 18598 0 sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13294 8058 13294 8058 0 sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21758 11356 21758 11356 0 sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 14398 6528 14398 6528 0 sb_0__8_.mux_right_track_36.out
rlabel metal1 14306 5746 14306 5746 0 sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14766 6324 14766 6324 0 sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14858 6069 14858 6069 0 sb_0__8_.mux_right_track_38.out
rlabel metal1 18124 5678 18124 5678 0 sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20562 5712 20562 5712 0 sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 19182 24514 19182 24514 0 sb_0__8_.mux_right_track_4.out
rlabel metal1 15640 29274 15640 29274 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15962 29614 15962 29614 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14030 27421 14030 27421 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13202 21352 13202 21352 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17710 25262 17710 25262 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 17342 4369 17342 4369 0 sb_0__8_.mux_right_track_40.out
rlabel metal1 20240 7310 20240 7310 0 sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22586 5338 22586 5338 0 sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 15732 3944 15732 3944 0 sb_0__8_.mux_right_track_42.out
rlabel metal1 21298 10710 21298 10710 0 sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19090 10676 19090 10676 0 sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24564 16014 24564 16014 0 sb_0__8_.mux_right_track_44.out
rlabel metal2 20102 18088 20102 18088 0 sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19734 14994 19734 14994 0 sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24058 14824 24058 14824 0 sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 24886 2414 24886 2414 0 sb_0__8_.mux_right_track_46.out
rlabel metal1 19826 21862 19826 21862 0 sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19458 12614 19458 12614 0 sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21482 15776 21482 15776 0 sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21390 13260 21390 13260 0 sb_0__8_.mux_right_track_48.out
rlabel metal1 21620 14450 21620 14450 0 sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21850 13333 21850 13333 0 sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23276 14586 23276 14586 0 sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 23874 2142 23874 2142 0 sb_0__8_.mux_right_track_50.out
rlabel metal1 21344 12614 21344 12614 0 sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23092 9962 23092 9962 0 sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17986 3927 17986 3927 0 sb_0__8_.mux_right_track_52.out
rlabel metal2 21390 8534 21390 8534 0 sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 19274 4930 19274 4930 0 sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16974 2618 16974 2618 0 sb_0__8_.mux_right_track_54.out
rlabel metal2 21022 5406 21022 5406 0 sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18906 2448 18906 2448 0 sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20470 2618 20470 2618 0 sb_0__8_.mux_right_track_56.out
rlabel metal1 18170 10166 18170 10166 0 sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19642 2278 19642 2278 0 sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21965 8806 21965 8806 0 sb_0__8_.mux_right_track_58.out
rlabel metal1 17296 12954 17296 12954 0 sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 17250 10540 17250 10540 0 sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17158 12614 17158 12614 0 sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23046 23528 23046 23528 0 sb_0__8_.mux_right_track_6.out
rlabel metal2 15778 28016 15778 28016 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16284 27098 16284 27098 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14950 25296 14950 25296 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14444 23698 14444 23698 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 18262 23732 18262 23732 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 16882 22882 16882 22882 0 sb_0__8_.mux_right_track_8.out
rlabel metal2 13754 25534 13754 25534 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13662 25126 13662 25126 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12880 23494 12880 23494 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 9062 17272 9062 17272 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 12052 22134 12052 22134 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X
<< properties >>
string FIXED_BBOX 0 0 27000 57000
<< end >>
