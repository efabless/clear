magic
tech sky130A
magscale 1 2
timestamp 1656248018
<< viali >>
rect 6377 17289 6411 17323
rect 6745 17289 6779 17323
rect 7113 17289 7147 17323
rect 7481 17289 7515 17323
rect 7849 17289 7883 17323
rect 8217 17289 8251 17323
rect 8585 17289 8619 17323
rect 9045 17289 9079 17323
rect 9413 17289 9447 17323
rect 15577 17289 15611 17323
rect 5733 17221 5767 17255
rect 10057 17221 10091 17255
rect 15025 17221 15059 17255
rect 1777 17153 1811 17187
rect 2145 17153 2179 17187
rect 2513 17153 2547 17187
rect 2881 17153 2915 17187
rect 2973 17153 3007 17187
rect 3341 17153 3375 17187
rect 3801 17153 3835 17187
rect 4169 17153 4203 17187
rect 4537 17153 4571 17187
rect 5181 17153 5215 17187
rect 5641 17153 5675 17187
rect 6561 17153 6595 17187
rect 6929 17153 6963 17187
rect 7297 17153 7331 17187
rect 7665 17153 7699 17187
rect 8033 17153 8067 17187
rect 8401 17153 8435 17187
rect 8769 17153 8803 17187
rect 9229 17153 9263 17187
rect 9597 17153 9631 17187
rect 11345 17153 11379 17187
rect 13277 17153 13311 17187
rect 13553 17153 13587 17187
rect 13737 17153 13771 17187
rect 15485 17153 15519 17187
rect 5917 17085 5951 17119
rect 9781 17085 9815 17119
rect 9965 17085 9999 17119
rect 11069 17085 11103 17119
rect 11529 17085 11563 17119
rect 11805 17085 11839 17119
rect 13001 17085 13035 17119
rect 14105 17085 14139 17119
rect 14381 17085 14415 17119
rect 1593 17017 1627 17051
rect 3157 17017 3191 17051
rect 3525 17017 3559 17051
rect 3985 17017 4019 17051
rect 4353 17017 4387 17051
rect 4721 17017 4755 17051
rect 1961 16949 1995 16983
rect 2329 16949 2363 16983
rect 2697 16949 2731 16983
rect 4997 16949 5031 16983
rect 5273 16949 5307 16983
rect 6101 16949 6135 16983
rect 10425 16949 10459 16983
rect 13461 16949 13495 16983
rect 13921 16949 13955 16983
rect 15301 16949 15335 16983
rect 6837 16745 6871 16779
rect 7665 16745 7699 16779
rect 9137 16745 9171 16779
rect 10241 16745 10275 16779
rect 11437 16745 11471 16779
rect 13737 16745 13771 16779
rect 15669 16745 15703 16779
rect 3341 16677 3375 16711
rect 4077 16677 4111 16711
rect 4353 16677 4387 16711
rect 10425 16677 10459 16711
rect 15301 16677 15335 16711
rect 7481 16609 7515 16643
rect 8493 16609 8527 16643
rect 9965 16609 9999 16643
rect 10977 16609 11011 16643
rect 12173 16609 12207 16643
rect 12449 16609 12483 16643
rect 13369 16609 13403 16643
rect 14105 16609 14139 16643
rect 14381 16609 14415 16643
rect 1501 16541 1535 16575
rect 1777 16541 1811 16575
rect 2329 16541 2363 16575
rect 2421 16541 2455 16575
rect 3065 16541 3099 16575
rect 3157 16541 3191 16575
rect 3433 16541 3467 16575
rect 3893 16541 3927 16575
rect 4169 16541 4203 16575
rect 4445 16541 4479 16575
rect 4997 16541 5031 16575
rect 5365 16541 5399 16575
rect 5632 16541 5666 16575
rect 7205 16541 7239 16575
rect 7849 16541 7883 16575
rect 8401 16541 8435 16575
rect 9321 16541 9355 16575
rect 10885 16541 10919 16575
rect 13093 16541 13127 16575
rect 13461 16541 13495 16575
rect 13921 16541 13955 16575
rect 15209 16541 15243 16575
rect 15485 16541 15519 16575
rect 7297 16473 7331 16507
rect 10793 16473 10827 16507
rect 11345 16473 11379 16507
rect 2145 16405 2179 16439
rect 2605 16405 2639 16439
rect 2881 16405 2915 16439
rect 3617 16405 3651 16439
rect 4629 16405 4663 16439
rect 4813 16405 4847 16439
rect 5181 16405 5215 16439
rect 6745 16405 6779 16439
rect 7941 16405 7975 16439
rect 8309 16405 8343 16439
rect 9045 16405 9079 16439
rect 9413 16405 9447 16439
rect 9781 16405 9815 16439
rect 9873 16405 9907 16439
rect 13645 16405 13679 16439
rect 15025 16405 15059 16439
rect 1501 16201 1535 16235
rect 1869 16201 1903 16235
rect 2329 16201 2363 16235
rect 2605 16201 2639 16235
rect 3249 16201 3283 16235
rect 3801 16201 3835 16235
rect 5457 16201 5491 16235
rect 6009 16201 6043 16235
rect 6745 16201 6779 16235
rect 7205 16201 7239 16235
rect 7573 16201 7607 16235
rect 8033 16201 8067 16235
rect 8493 16201 8527 16235
rect 12357 16201 12391 16235
rect 5733 16133 5767 16167
rect 9882 16133 9916 16167
rect 1685 16065 1719 16099
rect 2053 16065 2087 16099
rect 2145 16065 2179 16099
rect 2789 16065 2823 16099
rect 3065 16065 3099 16099
rect 3525 16065 3559 16099
rect 3617 16065 3651 16099
rect 5006 16065 5040 16099
rect 5273 16065 5307 16099
rect 5641 16065 5675 16099
rect 6193 16065 6227 16099
rect 6561 16065 6595 16099
rect 6929 16065 6963 16099
rect 7389 16065 7423 16099
rect 7757 16065 7791 16099
rect 8217 16065 8251 16099
rect 8677 16065 8711 16099
rect 10241 16065 10275 16099
rect 10977 16065 11011 16099
rect 11897 16065 11931 16099
rect 12541 16065 12575 16099
rect 13645 16065 13679 16099
rect 14565 16065 14599 16099
rect 15485 16065 15519 16099
rect 7113 15997 7147 16031
rect 10149 15997 10183 16031
rect 11069 15997 11103 16031
rect 11161 15997 11195 16031
rect 11989 15997 12023 16031
rect 12081 15997 12115 16031
rect 13277 15997 13311 16031
rect 13553 15997 13587 16031
rect 13921 15997 13955 16031
rect 3341 15929 3375 15963
rect 6377 15929 6411 15963
rect 8401 15929 8435 15963
rect 10609 15929 10643 15963
rect 2421 15861 2455 15895
rect 2973 15861 3007 15895
rect 3893 15861 3927 15895
rect 7849 15861 7883 15895
rect 8769 15861 8803 15895
rect 10425 15861 10459 15895
rect 11529 15861 11563 15895
rect 14795 15861 14829 15895
rect 15669 15861 15703 15895
rect 7389 15657 7423 15691
rect 10977 15657 11011 15691
rect 13737 15657 13771 15691
rect 14197 15657 14231 15691
rect 1777 15589 1811 15623
rect 7297 15589 7331 15623
rect 9321 15589 9355 15623
rect 13461 15589 13495 15623
rect 14473 15589 14507 15623
rect 11437 15521 11471 15555
rect 11529 15521 11563 15555
rect 12357 15521 12391 15555
rect 13185 15521 13219 15555
rect 14749 15521 14783 15555
rect 1685 15453 1719 15487
rect 1961 15453 1995 15487
rect 2145 15453 2179 15487
rect 3617 15453 3651 15487
rect 5273 15453 5307 15487
rect 5457 15453 5491 15487
rect 8769 15453 8803 15487
rect 9137 15453 9171 15487
rect 10434 15453 10468 15487
rect 10701 15453 10735 15487
rect 13645 15453 13679 15487
rect 14381 15453 14415 15487
rect 14657 15453 14691 15487
rect 15025 15453 15059 15487
rect 3372 15385 3406 15419
rect 5006 15385 5040 15419
rect 5702 15385 5736 15419
rect 8524 15385 8558 15419
rect 9045 15385 9079 15419
rect 1501 15317 1535 15351
rect 2237 15317 2271 15351
rect 3893 15317 3927 15351
rect 6837 15317 6871 15351
rect 7113 15317 7147 15351
rect 10793 15317 10827 15351
rect 11345 15317 11379 15351
rect 11805 15317 11839 15351
rect 12173 15317 12207 15351
rect 12265 15317 12299 15351
rect 12633 15317 12667 15351
rect 13001 15317 13035 15351
rect 13093 15317 13127 15351
rect 1777 15113 1811 15147
rect 2513 15113 2547 15147
rect 7021 15113 7055 15147
rect 8953 15113 8987 15147
rect 11529 15113 11563 15147
rect 12909 15113 12943 15147
rect 13369 15113 13403 15147
rect 13645 15113 13679 15147
rect 14381 15113 14415 15147
rect 7380 15045 7414 15079
rect 13001 15045 13035 15079
rect 2421 14977 2455 15011
rect 2697 14977 2731 15011
rect 2789 14977 2823 15011
rect 3056 14977 3090 15011
rect 10250 14977 10284 15011
rect 10977 14977 11011 15011
rect 11897 14977 11931 15011
rect 13737 14977 13771 15011
rect 14841 14977 14875 15011
rect 1501 14909 1535 14943
rect 1685 14909 1719 14943
rect 4445 14909 4479 14943
rect 5273 14909 5307 14943
rect 7113 14909 7147 14943
rect 10517 14909 10551 14943
rect 10701 14909 10735 14943
rect 10885 14909 10919 14943
rect 11989 14909 12023 14943
rect 12081 14909 12115 14943
rect 12449 14909 12483 14943
rect 13093 14909 13127 14943
rect 14105 14909 14139 14943
rect 14289 14909 14323 14943
rect 2237 14841 2271 14875
rect 4169 14841 4203 14875
rect 8493 14841 8527 14875
rect 11345 14841 11379 14875
rect 2145 14773 2179 14807
rect 4537 14773 4571 14807
rect 4813 14773 4847 14807
rect 5733 14773 5767 14807
rect 9137 14773 9171 14807
rect 12541 14773 12575 14807
rect 14749 14773 14783 14807
rect 15071 14773 15105 14807
rect 1777 14569 1811 14603
rect 3433 14569 3467 14603
rect 10425 14569 10459 14603
rect 12357 14569 12391 14603
rect 13185 14569 13219 14603
rect 14105 14569 14139 14603
rect 14381 14569 14415 14603
rect 3985 14501 4019 14535
rect 2881 14433 2915 14467
rect 3157 14433 3191 14467
rect 3893 14433 3927 14467
rect 4905 14433 4939 14467
rect 10793 14433 10827 14467
rect 11621 14433 11655 14467
rect 12817 14433 12851 14467
rect 12909 14433 12943 14467
rect 13829 14433 13863 14467
rect 15669 14433 15703 14467
rect 1685 14365 1719 14399
rect 1961 14365 1995 14399
rect 2237 14365 2271 14399
rect 6469 14365 6503 14399
rect 7941 14365 7975 14399
rect 10977 14365 11011 14399
rect 11805 14365 11839 14399
rect 11897 14365 11931 14399
rect 14473 14365 14507 14399
rect 15393 14365 15427 14399
rect 6224 14297 6258 14331
rect 7674 14297 7708 14331
rect 12725 14297 12759 14331
rect 13553 14297 13587 14331
rect 1501 14229 1535 14263
rect 3525 14229 3559 14263
rect 4169 14229 4203 14263
rect 5089 14229 5123 14263
rect 6561 14229 6595 14263
rect 10609 14229 10643 14263
rect 11069 14229 11103 14263
rect 11437 14229 11471 14263
rect 12265 14229 12299 14263
rect 13645 14229 13679 14263
rect 1409 14025 1443 14059
rect 2237 14025 2271 14059
rect 2513 14025 2547 14059
rect 2881 14025 2915 14059
rect 3157 14025 3191 14059
rect 4629 14025 4663 14059
rect 5641 14025 5675 14059
rect 6377 14025 6411 14059
rect 6929 14025 6963 14059
rect 9413 14025 9447 14059
rect 11069 14025 11103 14059
rect 11345 14025 11379 14059
rect 12725 14025 12759 14059
rect 13185 14025 13219 14059
rect 13461 14025 13495 14059
rect 13829 14025 13863 14059
rect 15117 14025 15151 14059
rect 15485 14025 15519 14059
rect 15669 14025 15703 14059
rect 5549 13957 5583 13991
rect 9321 13957 9355 13991
rect 14197 13957 14231 13991
rect 1777 13889 1811 13923
rect 2421 13889 2455 13923
rect 2697 13889 2731 13923
rect 3249 13889 3283 13923
rect 3505 13889 3539 13923
rect 7113 13889 7147 13923
rect 7369 13889 7403 13923
rect 10526 13889 10560 13923
rect 10793 13889 10827 13923
rect 11897 13889 11931 13923
rect 12817 13889 12851 13923
rect 1869 13821 1903 13855
rect 2053 13821 2087 13855
rect 11621 13821 11655 13855
rect 11805 13821 11839 13855
rect 12909 13821 12943 13855
rect 13737 13821 13771 13855
rect 14289 13821 14323 13855
rect 14473 13821 14507 13855
rect 14933 13821 14967 13855
rect 15025 13821 15059 13855
rect 8493 13753 8527 13787
rect 12265 13753 12299 13787
rect 12357 13685 12391 13719
rect 1869 13481 1903 13515
rect 4169 13481 4203 13515
rect 10425 13481 10459 13515
rect 11897 13481 11931 13515
rect 13553 13481 13587 13515
rect 13737 13481 13771 13515
rect 14105 13481 14139 13515
rect 14565 13481 14599 13515
rect 14657 13481 14691 13515
rect 7389 13413 7423 13447
rect 12725 13413 12759 13447
rect 5733 13345 5767 13379
rect 5825 13345 5859 13379
rect 11621 13345 11655 13379
rect 12449 13345 12483 13379
rect 13277 13345 13311 13379
rect 15209 13345 15243 13379
rect 1685 13277 1719 13311
rect 8769 13277 8803 13311
rect 9045 13277 9079 13311
rect 15117 13277 15151 13311
rect 15669 13277 15703 13311
rect 5488 13209 5522 13243
rect 6092 13209 6126 13243
rect 8502 13209 8536 13243
rect 9312 13209 9346 13243
rect 12265 13209 12299 13243
rect 12357 13209 12391 13243
rect 13093 13209 13127 13243
rect 1501 13141 1535 13175
rect 4353 13141 4387 13175
rect 7205 13141 7239 13175
rect 11069 13141 11103 13175
rect 11437 13141 11471 13175
rect 11529 13141 11563 13175
rect 13185 13141 13219 13175
rect 14289 13141 14323 13175
rect 15025 13141 15059 13175
rect 15485 13141 15519 13175
rect 2789 12937 2823 12971
rect 4445 12937 4479 12971
rect 7021 12937 7055 12971
rect 7205 12937 7239 12971
rect 8953 12937 8987 12971
rect 9321 12937 9355 12971
rect 11713 12937 11747 12971
rect 13369 12937 13403 12971
rect 13737 12937 13771 12971
rect 14657 12937 14691 12971
rect 15577 12937 15611 12971
rect 7564 12869 7598 12903
rect 12357 12869 12391 12903
rect 12817 12869 12851 12903
rect 12909 12869 12943 12903
rect 15117 12869 15151 12903
rect 1685 12801 1719 12835
rect 1961 12801 1995 12835
rect 2881 12801 2915 12835
rect 3148 12801 3182 12835
rect 5558 12801 5592 12835
rect 5825 12801 5859 12835
rect 7297 12801 7331 12835
rect 10629 12801 10663 12835
rect 14565 12801 14599 12835
rect 15485 12801 15519 12835
rect 10885 12733 10919 12767
rect 12633 12733 12667 12767
rect 13829 12733 13863 12767
rect 14013 12733 14047 12767
rect 14749 12733 14783 12767
rect 14197 12665 14231 12699
rect 15301 12665 15335 12699
rect 1501 12597 1535 12631
rect 1777 12597 1811 12631
rect 4261 12597 4295 12631
rect 8677 12597 8711 12631
rect 9505 12597 9539 12631
rect 13277 12597 13311 12631
rect 2145 12393 2179 12427
rect 4905 12393 4939 12427
rect 8769 12393 8803 12427
rect 13553 12393 13587 12427
rect 14105 12393 14139 12427
rect 3801 12325 3835 12359
rect 4261 12325 4295 12359
rect 13829 12325 13863 12359
rect 1593 12257 1627 12291
rect 2237 12257 2271 12291
rect 4629 12257 4663 12291
rect 12633 12257 12667 12291
rect 12909 12257 12943 12291
rect 14657 12257 14691 12291
rect 15025 12257 15059 12291
rect 1777 12189 1811 12223
rect 6285 12189 6319 12223
rect 7205 12189 7239 12223
rect 7389 12189 7423 12223
rect 7656 12189 7690 12223
rect 14565 12189 14599 12223
rect 15301 12189 15335 12223
rect 2482 12121 2516 12155
rect 6018 12121 6052 12155
rect 13093 12121 13127 12155
rect 13185 12121 13219 12155
rect 13737 12121 13771 12155
rect 1685 12053 1719 12087
rect 3617 12053 3651 12087
rect 4445 12053 4479 12087
rect 14473 12053 14507 12087
rect 15209 12053 15243 12087
rect 15669 12053 15703 12087
rect 6101 11849 6135 11883
rect 7941 11849 7975 11883
rect 11529 11849 11563 11883
rect 11989 11849 12023 11883
rect 14197 11849 14231 11883
rect 15485 11849 15519 11883
rect 15669 11849 15703 11883
rect 6644 11781 6678 11815
rect 9505 11781 9539 11815
rect 10710 11781 10744 11815
rect 14841 11781 14875 11815
rect 1685 11713 1719 11747
rect 2964 11713 2998 11747
rect 4528 11713 4562 11747
rect 6377 11713 6411 11747
rect 10977 11713 11011 11747
rect 11897 11713 11931 11747
rect 12817 11713 12851 11747
rect 14105 11713 14139 11747
rect 14933 11713 14967 11747
rect 2697 11645 2731 11679
rect 4261 11645 4295 11679
rect 12081 11645 12115 11679
rect 12357 11645 12391 11679
rect 13093 11645 13127 11679
rect 14289 11645 14323 11679
rect 14749 11645 14783 11679
rect 1501 11509 1535 11543
rect 4077 11509 4111 11543
rect 5641 11509 5675 11543
rect 7757 11509 7791 11543
rect 9597 11509 9631 11543
rect 13737 11509 13771 11543
rect 15301 11509 15335 11543
rect 1501 11305 1535 11339
rect 4077 11305 4111 11339
rect 4261 11305 4295 11339
rect 4445 11305 4479 11339
rect 5641 11305 5675 11339
rect 7205 11305 7239 11339
rect 11253 11305 11287 11339
rect 13185 11305 13219 11339
rect 14841 11305 14875 11339
rect 3525 11237 3559 11271
rect 9045 11237 9079 11271
rect 9229 11237 9263 11271
rect 13093 11237 13127 11271
rect 2145 11169 2179 11203
rect 5825 11169 5859 11203
rect 10701 11169 10735 11203
rect 11897 11169 11931 11203
rect 12449 11169 12483 11203
rect 13645 11169 13679 11203
rect 13737 11169 13771 11203
rect 15393 11169 15427 11203
rect 1685 11101 1719 11135
rect 3985 11101 4019 11135
rect 6092 11101 6126 11135
rect 7389 11101 7423 11135
rect 11621 11101 11655 11135
rect 12725 11101 12759 11135
rect 13553 11101 13587 11135
rect 14381 11101 14415 11135
rect 15209 11101 15243 11135
rect 2412 11033 2446 11067
rect 7656 11033 7690 11067
rect 10456 11033 10490 11067
rect 12633 11033 12667 11067
rect 15301 11033 15335 11067
rect 8769 10965 8803 10999
rect 9321 10965 9355 10999
rect 11713 10965 11747 10999
rect 12173 10965 12207 10999
rect 1777 10761 1811 10795
rect 2237 10761 2271 10795
rect 3157 10761 3191 10795
rect 3801 10761 3835 10795
rect 7021 10761 7055 10795
rect 13461 10761 13495 10795
rect 14841 10761 14875 10795
rect 15209 10761 15243 10795
rect 9505 10693 9539 10727
rect 14473 10693 14507 10727
rect 1685 10625 1719 10659
rect 2605 10625 2639 10659
rect 3893 10625 3927 10659
rect 4160 10625 4194 10659
rect 7113 10625 7147 10659
rect 7380 10625 7414 10659
rect 10710 10625 10744 10659
rect 10977 10625 11011 10659
rect 13369 10625 13403 10659
rect 14381 10625 14415 10659
rect 1593 10557 1627 10591
rect 2697 10557 2731 10591
rect 2881 10557 2915 10591
rect 12909 10557 12943 10591
rect 13553 10557 13587 10591
rect 14565 10557 14599 10591
rect 15301 10557 15335 10591
rect 15393 10557 15427 10591
rect 2145 10489 2179 10523
rect 13001 10489 13035 10523
rect 14013 10489 14047 10523
rect 5273 10421 5307 10455
rect 8493 10421 8527 10455
rect 9597 10421 9631 10455
rect 1501 10217 1535 10251
rect 6929 10217 6963 10251
rect 10609 10217 10643 10251
rect 14105 10217 14139 10251
rect 14933 10217 14967 10251
rect 7389 10149 7423 10183
rect 10517 10081 10551 10115
rect 12541 10081 12575 10115
rect 12725 10081 12759 10115
rect 13001 10081 13035 10115
rect 13185 10081 13219 10115
rect 13829 10081 13863 10115
rect 14749 10081 14783 10115
rect 15393 10081 15427 10115
rect 15485 10081 15519 10115
rect 1685 10013 1719 10047
rect 5549 10013 5583 10047
rect 5816 10013 5850 10047
rect 7297 10013 7331 10047
rect 8769 10013 8803 10047
rect 10250 10013 10284 10047
rect 11989 10013 12023 10047
rect 12449 10013 12483 10047
rect 15301 10013 15335 10047
rect 4445 9945 4479 9979
rect 5365 9945 5399 9979
rect 8502 9945 8536 9979
rect 11722 9945 11756 9979
rect 14565 9945 14599 9979
rect 9137 9877 9171 9911
rect 12081 9877 12115 9911
rect 13277 9877 13311 9911
rect 13645 9877 13679 9911
rect 14473 9877 14507 9911
rect 1777 9673 1811 9707
rect 10701 9673 10735 9707
rect 13185 9673 13219 9707
rect 14841 9673 14875 9707
rect 6193 9605 6227 9639
rect 8769 9605 8803 9639
rect 8953 9605 8987 9639
rect 10250 9605 10284 9639
rect 14105 9605 14139 9639
rect 15209 9605 15243 9639
rect 1685 9537 1719 9571
rect 1961 9537 1995 9571
rect 3240 9537 3274 9571
rect 5661 9537 5695 9571
rect 5917 9537 5951 9571
rect 7490 9537 7524 9571
rect 10517 9537 10551 9571
rect 11989 9537 12023 9571
rect 14013 9537 14047 9571
rect 14565 9537 14599 9571
rect 2973 9469 3007 9503
rect 7757 9469 7791 9503
rect 12081 9469 12115 9503
rect 12173 9469 12207 9503
rect 13277 9469 13311 9503
rect 13369 9469 13403 9503
rect 14197 9469 14231 9503
rect 15301 9469 15335 9503
rect 15485 9469 15519 9503
rect 1501 9401 1535 9435
rect 4353 9401 4387 9435
rect 11621 9401 11655 9435
rect 12541 9401 12575 9435
rect 12817 9401 12851 9435
rect 2881 9333 2915 9367
rect 4537 9333 4571 9367
rect 6377 9333 6411 9367
rect 9137 9333 9171 9367
rect 12633 9333 12667 9367
rect 13645 9333 13679 9367
rect 14749 9333 14783 9367
rect 1777 9129 1811 9163
rect 3985 9129 4019 9163
rect 9229 9129 9263 9163
rect 9413 9129 9447 9163
rect 11805 9129 11839 9163
rect 12541 9061 12575 9095
rect 14933 9061 14967 9095
rect 15577 9061 15611 9095
rect 2237 8993 2271 9027
rect 5457 8993 5491 9027
rect 8769 8993 8803 9027
rect 13553 8993 13587 9027
rect 15301 8993 15335 9027
rect 1685 8925 1719 8959
rect 1961 8925 1995 8959
rect 3893 8925 3927 8959
rect 5365 8925 5399 8959
rect 7297 8925 7331 8959
rect 10793 8925 10827 8959
rect 13277 8925 13311 8959
rect 13829 8925 13863 8959
rect 14657 8925 14691 8959
rect 15393 8925 15427 8959
rect 2482 8857 2516 8891
rect 5098 8857 5132 8891
rect 8502 8857 8536 8891
rect 10526 8857 10560 8891
rect 11989 8857 12023 8891
rect 12817 8857 12851 8891
rect 13369 8857 13403 8891
rect 1501 8789 1535 8823
rect 3617 8789 3651 8823
rect 7389 8789 7423 8823
rect 12173 8789 12207 8823
rect 12449 8789 12483 8823
rect 12909 8789 12943 8823
rect 14105 8789 14139 8823
rect 14473 8789 14507 8823
rect 1869 8585 1903 8619
rect 2237 8585 2271 8619
rect 7757 8585 7791 8619
rect 9045 8585 9079 8619
rect 10609 8585 10643 8619
rect 13553 8585 13587 8619
rect 14197 8585 14231 8619
rect 14565 8585 14599 8619
rect 15577 8585 15611 8619
rect 1777 8517 1811 8551
rect 9474 8517 9508 8551
rect 12725 8517 12759 8551
rect 3718 8449 3752 8483
rect 3985 8449 4019 8483
rect 4077 8449 4111 8483
rect 4344 8449 4378 8483
rect 6644 8449 6678 8483
rect 9229 8449 9263 8483
rect 11897 8449 11931 8483
rect 14105 8449 14139 8483
rect 1685 8381 1719 8415
rect 6377 8381 6411 8415
rect 11345 8381 11379 8415
rect 11989 8381 12023 8415
rect 12081 8381 12115 8415
rect 12817 8381 12851 8415
rect 12909 8381 12943 8415
rect 13369 8381 13403 8415
rect 13461 8381 13495 8415
rect 14657 8381 14691 8415
rect 14749 8381 14783 8415
rect 15117 8381 15151 8415
rect 12357 8313 12391 8347
rect 15485 8313 15519 8347
rect 2605 8245 2639 8279
rect 5457 8245 5491 8279
rect 6193 8245 6227 8279
rect 11529 8245 11563 8279
rect 13921 8245 13955 8279
rect 2145 8041 2179 8075
rect 9229 8041 9263 8075
rect 12541 8041 12575 8075
rect 13921 8041 13955 8075
rect 15577 8041 15611 8075
rect 3617 7973 3651 8007
rect 6285 7973 6319 8007
rect 12081 7973 12115 8007
rect 14289 7973 14323 8007
rect 1593 7905 1627 7939
rect 2237 7905 2271 7939
rect 7665 7905 7699 7939
rect 10793 7905 10827 7939
rect 11621 7905 11655 7939
rect 12173 7905 12207 7939
rect 13001 7905 13035 7939
rect 13185 7905 13219 7939
rect 13737 7905 13771 7939
rect 15301 7905 15335 7939
rect 2504 7837 2538 7871
rect 3985 7837 4019 7871
rect 4169 7837 4203 7871
rect 4353 7837 4387 7871
rect 4629 7837 4663 7871
rect 4813 7837 4847 7871
rect 10537 7837 10571 7871
rect 11345 7837 11379 7871
rect 15117 7837 15151 7871
rect 1777 7769 1811 7803
rect 5080 7769 5114 7803
rect 7398 7769 7432 7803
rect 12909 7769 12943 7803
rect 15209 7769 15243 7803
rect 1685 7701 1719 7735
rect 6193 7701 6227 7735
rect 8585 7701 8619 7735
rect 9413 7701 9447 7735
rect 10977 7701 11011 7735
rect 11437 7701 11471 7735
rect 11805 7701 11839 7735
rect 12449 7701 12483 7735
rect 13461 7701 13495 7735
rect 14105 7701 14139 7735
rect 14565 7701 14599 7735
rect 14749 7701 14783 7735
rect 1501 7497 1535 7531
rect 1777 7497 1811 7531
rect 6193 7497 6227 7531
rect 7481 7497 7515 7531
rect 9229 7497 9263 7531
rect 9321 7497 9355 7531
rect 11161 7497 11195 7531
rect 11897 7497 11931 7531
rect 15485 7497 15519 7531
rect 3065 7429 3099 7463
rect 5742 7429 5776 7463
rect 10434 7429 10468 7463
rect 12909 7429 12943 7463
rect 1685 7361 1719 7395
rect 1961 7361 1995 7395
rect 4270 7361 4304 7395
rect 4537 7361 4571 7395
rect 6009 7361 6043 7395
rect 8789 7361 8823 7395
rect 9045 7361 9079 7395
rect 10701 7361 10735 7395
rect 11989 7361 12023 7395
rect 12541 7361 12575 7395
rect 13461 7361 13495 7395
rect 13921 7361 13955 7395
rect 14013 7361 14047 7395
rect 14565 7365 14599 7399
rect 15025 7361 15059 7395
rect 15117 7361 15151 7395
rect 15669 7361 15703 7395
rect 10977 7293 11011 7327
rect 12081 7293 12115 7327
rect 14105 7293 14139 7327
rect 15209 7293 15243 7327
rect 4629 7225 4663 7259
rect 7665 7225 7699 7259
rect 12725 7225 12759 7259
rect 13277 7225 13311 7259
rect 3157 7157 3191 7191
rect 11345 7157 11379 7191
rect 11529 7157 11563 7191
rect 13093 7157 13127 7191
rect 13553 7157 13587 7191
rect 14381 7157 14415 7191
rect 14657 7157 14691 7191
rect 4537 6953 4571 6987
rect 6469 6953 6503 6987
rect 8033 6953 8067 6987
rect 8401 6953 8435 6987
rect 11161 6953 11195 6987
rect 8493 6885 8527 6919
rect 8769 6885 8803 6919
rect 10885 6885 10919 6919
rect 1961 6817 1995 6851
rect 6561 6817 6595 6851
rect 9505 6817 9539 6851
rect 9873 6817 9907 6851
rect 11713 6817 11747 6851
rect 12541 6817 12575 6851
rect 13369 6817 13403 6851
rect 14473 6817 14507 6851
rect 14841 6817 14875 6851
rect 1685 6749 1719 6783
rect 6817 6749 6851 6783
rect 8217 6725 8251 6759
rect 9413 6749 9447 6783
rect 10793 6749 10827 6783
rect 11529 6749 11563 6783
rect 13277 6749 13311 6783
rect 13921 6749 13955 6783
rect 14565 6749 14599 6783
rect 15117 6749 15151 6783
rect 2237 6681 2271 6715
rect 12357 6681 12391 6715
rect 13185 6681 13219 6715
rect 1501 6613 1535 6647
rect 2145 6613 2179 6647
rect 2605 6613 2639 6647
rect 7941 6613 7975 6647
rect 8953 6613 8987 6647
rect 9321 6613 9355 6647
rect 10149 6613 10183 6647
rect 10333 6613 10367 6647
rect 10609 6613 10643 6647
rect 11621 6613 11655 6647
rect 11989 6613 12023 6647
rect 12449 6613 12483 6647
rect 12817 6613 12851 6647
rect 13737 6613 13771 6647
rect 14105 6613 14139 6647
rect 14749 6613 14783 6647
rect 1593 6409 1627 6443
rect 1961 6409 1995 6443
rect 2973 6409 3007 6443
rect 3341 6409 3375 6443
rect 3893 6409 3927 6443
rect 5641 6409 5675 6443
rect 6193 6409 6227 6443
rect 7021 6409 7055 6443
rect 10609 6409 10643 6443
rect 10977 6409 11011 6443
rect 11161 6409 11195 6443
rect 12265 6409 12299 6443
rect 12633 6409 12667 6443
rect 13461 6409 13495 6443
rect 13829 6409 13863 6443
rect 13921 6409 13955 6443
rect 14473 6409 14507 6443
rect 14933 6409 14967 6443
rect 15301 6409 15335 6443
rect 4997 6341 5031 6375
rect 7665 6341 7699 6375
rect 7849 6341 7883 6375
rect 8208 6341 8242 6375
rect 9781 6341 9815 6375
rect 9873 6341 9907 6375
rect 3433 6273 3467 6307
rect 5549 6273 5583 6307
rect 6469 6273 6503 6307
rect 7113 6273 7147 6307
rect 7941 6273 7975 6307
rect 10517 6273 10551 6307
rect 12173 6273 12207 6307
rect 13001 6273 13035 6307
rect 14289 6273 14323 6307
rect 15577 6273 15611 6307
rect 2053 6205 2087 6239
rect 2237 6205 2271 6239
rect 3617 6205 3651 6239
rect 5825 6205 5859 6239
rect 6837 6205 6871 6239
rect 9965 6205 9999 6239
rect 10425 6205 10459 6239
rect 11713 6205 11747 6239
rect 12449 6205 12483 6239
rect 13093 6205 13127 6239
rect 13185 6205 13219 6239
rect 14013 6205 14047 6239
rect 14657 6205 14691 6239
rect 14841 6205 14875 6239
rect 9321 6137 9355 6171
rect 9413 6137 9447 6171
rect 1409 6069 1443 6103
rect 3985 6069 4019 6103
rect 4629 6069 4663 6103
rect 5181 6069 5215 6103
rect 6653 6069 6687 6103
rect 7481 6069 7515 6103
rect 11253 6069 11287 6103
rect 11805 6069 11839 6103
rect 15393 6069 15427 6103
rect 1777 5865 1811 5899
rect 2329 5865 2363 5899
rect 4629 5865 4663 5899
rect 14289 5865 14323 5899
rect 3433 5797 3467 5831
rect 3801 5797 3835 5831
rect 7941 5797 7975 5831
rect 9229 5797 9263 5831
rect 9413 5797 9447 5831
rect 10517 5797 10551 5831
rect 2881 5729 2915 5763
rect 4445 5729 4479 5763
rect 5273 5729 5307 5763
rect 6745 5729 6779 5763
rect 7113 5729 7147 5763
rect 7297 5729 7331 5763
rect 8585 5729 8619 5763
rect 9689 5729 9723 5763
rect 11345 5729 11379 5763
rect 12357 5729 12391 5763
rect 12449 5729 12483 5763
rect 13369 5729 13403 5763
rect 15117 5729 15151 5763
rect 1685 5661 1719 5695
rect 1961 5661 1995 5695
rect 3617 5661 3651 5695
rect 4169 5661 4203 5695
rect 4813 5661 4847 5695
rect 5181 5661 5215 5695
rect 5549 5661 5583 5695
rect 6561 5661 6595 5695
rect 7573 5661 7607 5695
rect 9045 5661 9079 5695
rect 10333 5661 10367 5695
rect 11161 5661 11195 5695
rect 11621 5661 11655 5695
rect 12265 5661 12299 5695
rect 14105 5661 14139 5695
rect 14565 5661 14599 5695
rect 14841 5661 14875 5695
rect 2237 5593 2271 5627
rect 2697 5593 2731 5627
rect 2789 5593 2823 5627
rect 6653 5593 6687 5627
rect 8401 5593 8435 5627
rect 9873 5593 9907 5627
rect 11069 5593 11103 5627
rect 13093 5593 13127 5627
rect 13553 5593 13587 5627
rect 13921 5593 13955 5627
rect 1501 5525 1535 5559
rect 3157 5525 3191 5559
rect 4261 5525 4295 5559
rect 4997 5525 5031 5559
rect 6193 5525 6227 5559
rect 7481 5525 7515 5559
rect 8033 5525 8067 5559
rect 8493 5525 8527 5559
rect 9781 5525 9815 5559
rect 10241 5525 10275 5559
rect 10701 5525 10735 5559
rect 11805 5525 11839 5559
rect 11897 5525 11931 5559
rect 12725 5525 12759 5559
rect 13185 5525 13219 5559
rect 14381 5525 14415 5559
rect 14749 5525 14783 5559
rect 2605 5321 2639 5355
rect 3065 5321 3099 5355
rect 3617 5321 3651 5355
rect 5549 5321 5583 5355
rect 7297 5321 7331 5355
rect 8585 5321 8619 5355
rect 8953 5321 8987 5355
rect 10057 5321 10091 5355
rect 10517 5321 10551 5355
rect 10885 5321 10919 5355
rect 10977 5321 11011 5355
rect 11805 5321 11839 5355
rect 12265 5321 12299 5355
rect 13369 5321 13403 5355
rect 14105 5321 14139 5355
rect 14657 5321 14691 5355
rect 15117 5321 15151 5355
rect 15485 5321 15519 5355
rect 2145 5253 2179 5287
rect 3157 5253 3191 5287
rect 5917 5253 5951 5287
rect 6653 5253 6687 5287
rect 6837 5253 6871 5287
rect 8125 5253 8159 5287
rect 9413 5253 9447 5287
rect 13553 5253 13587 5287
rect 15025 5253 15059 5287
rect 1685 5185 1719 5219
rect 2237 5185 2271 5219
rect 3985 5185 4019 5219
rect 5457 5185 5491 5219
rect 9045 5185 9079 5219
rect 10149 5185 10183 5219
rect 11897 5185 11931 5219
rect 12725 5185 12759 5219
rect 13185 5185 13219 5219
rect 14013 5185 14047 5219
rect 15669 5185 15703 5219
rect 1961 5117 1995 5151
rect 3341 5117 3375 5151
rect 4077 5117 4111 5151
rect 4261 5117 4295 5151
rect 4537 5117 4571 5151
rect 5641 5117 5675 5151
rect 7389 5117 7423 5151
rect 7573 5117 7607 5151
rect 7849 5117 7883 5151
rect 8033 5117 8067 5151
rect 9137 5117 9171 5151
rect 9873 5117 9907 5151
rect 10701 5117 10735 5151
rect 11621 5117 11655 5151
rect 12817 5117 12851 5151
rect 13001 5117 13035 5151
rect 14289 5117 14323 5151
rect 15209 5117 15243 5151
rect 5089 5049 5123 5083
rect 6193 5049 6227 5083
rect 13645 5049 13679 5083
rect 1501 4981 1535 5015
rect 2697 4981 2731 5015
rect 4721 4981 4755 5015
rect 4905 4981 4939 5015
rect 6377 4981 6411 5015
rect 6929 4981 6963 5015
rect 8493 4981 8527 5015
rect 11345 4981 11379 5015
rect 12357 4981 12391 5015
rect 14473 4981 14507 5015
rect 1685 4777 1719 4811
rect 2421 4777 2455 4811
rect 3801 4777 3835 4811
rect 5549 4777 5583 4811
rect 6653 4777 6687 4811
rect 8309 4777 8343 4811
rect 9413 4777 9447 4811
rect 9689 4777 9723 4811
rect 10517 4777 10551 4811
rect 12725 4777 12759 4811
rect 13921 4777 13955 4811
rect 14565 4777 14599 4811
rect 1593 4709 1627 4743
rect 3433 4709 3467 4743
rect 11437 4709 11471 4743
rect 3249 4641 3283 4675
rect 4445 4641 4479 4675
rect 4997 4641 5031 4675
rect 5089 4641 5123 4675
rect 6285 4641 6319 4675
rect 6469 4641 6503 4675
rect 7113 4641 7147 4675
rect 7297 4641 7331 4675
rect 7941 4641 7975 4675
rect 8033 4641 8067 4675
rect 9873 4641 9907 4675
rect 10057 4641 10091 4675
rect 11161 4641 11195 4675
rect 11989 4641 12023 4675
rect 12541 4641 12575 4675
rect 13369 4641 13403 4675
rect 14289 4641 14323 4675
rect 15025 4641 15059 4675
rect 15117 4641 15151 4675
rect 1409 4573 1443 4607
rect 1869 4573 1903 4607
rect 2145 4573 2179 4607
rect 2237 4573 2271 4607
rect 4261 4573 4295 4607
rect 6193 4573 6227 4607
rect 7021 4573 7055 4607
rect 7849 4573 7883 4607
rect 8469 4573 8503 4607
rect 8585 4549 8619 4583
rect 9321 4573 9355 4607
rect 10977 4573 11011 4607
rect 11805 4573 11839 4607
rect 12449 4573 12483 4607
rect 15393 4573 15427 4607
rect 2605 4505 2639 4539
rect 2789 4505 2823 4539
rect 4721 4505 4755 4539
rect 5641 4505 5675 4539
rect 10149 4505 10183 4539
rect 11069 4505 11103 4539
rect 13093 4505 13127 4539
rect 13553 4505 13587 4539
rect 14197 4505 14231 4539
rect 14933 4505 14967 4539
rect 1961 4437 1995 4471
rect 3065 4437 3099 4471
rect 3617 4437 3651 4471
rect 4169 4437 4203 4471
rect 5181 4437 5215 4471
rect 5825 4437 5859 4471
rect 7481 4437 7515 4471
rect 8769 4437 8803 4471
rect 9045 4437 9079 4471
rect 10609 4437 10643 4471
rect 11897 4437 11931 4471
rect 12265 4437 12299 4471
rect 13185 4437 13219 4471
rect 15577 4437 15611 4471
rect 1869 4233 1903 4267
rect 10149 4233 10183 4267
rect 10517 4233 10551 4267
rect 11897 4233 11931 4267
rect 13185 4233 13219 4267
rect 14933 4233 14967 4267
rect 1501 4165 1535 4199
rect 5641 4165 5675 4199
rect 6745 4165 6779 4199
rect 8953 4165 8987 4199
rect 12817 4165 12851 4199
rect 1961 4097 1995 4131
rect 2605 4097 2639 4131
rect 2881 4097 2915 4131
rect 3157 4097 3191 4131
rect 3433 4097 3467 4131
rect 3893 4097 3927 4131
rect 4721 4097 4755 4131
rect 4813 4097 4847 4131
rect 5549 4097 5583 4131
rect 6185 4097 6219 4131
rect 7389 4097 7423 4131
rect 7665 4097 7699 4131
rect 8125 4097 8159 4131
rect 9505 4097 9539 4131
rect 10057 4097 10091 4131
rect 10977 4097 11011 4131
rect 12725 4097 12759 4131
rect 13553 4097 13587 4131
rect 14013 4097 14047 4131
rect 14473 4097 14507 4131
rect 15393 4097 15427 4131
rect 1777 4029 1811 4063
rect 3617 4029 3651 4063
rect 3801 4029 3835 4063
rect 4997 4029 5031 4063
rect 5825 4029 5859 4063
rect 6837 4029 6871 4063
rect 6929 4029 6963 4063
rect 7849 4029 7883 4063
rect 8033 4029 8067 4063
rect 9045 4029 9079 4063
rect 9137 4029 9171 4063
rect 9965 4029 9999 4063
rect 11069 4029 11103 4063
rect 11253 4029 11287 4063
rect 11989 4029 12023 4063
rect 12173 4029 12207 4063
rect 12909 4029 12943 4063
rect 13645 4029 13679 4063
rect 13737 4029 13771 4063
rect 14657 4029 14691 4063
rect 14841 4029 14875 4063
rect 2329 3961 2363 3995
rect 2973 3961 3007 3995
rect 4261 3961 4295 3995
rect 8493 3961 8527 3995
rect 9689 3961 9723 3995
rect 12357 3961 12391 3995
rect 14197 3961 14231 3995
rect 2421 3893 2455 3927
rect 2697 3893 2731 3927
rect 3249 3893 3283 3927
rect 4353 3893 4387 3927
rect 5181 3893 5215 3927
rect 6009 3893 6043 3927
rect 6377 3893 6411 3927
rect 7205 3893 7239 3927
rect 7481 3893 7515 3927
rect 8585 3893 8619 3927
rect 10609 3893 10643 3927
rect 11529 3893 11563 3927
rect 14289 3893 14323 3927
rect 15301 3893 15335 3927
rect 15577 3893 15611 3927
rect 1501 3689 1535 3723
rect 6285 3689 6319 3723
rect 6837 3689 6871 3723
rect 7849 3689 7883 3723
rect 8953 3689 8987 3723
rect 9965 3689 9999 3723
rect 11069 3689 11103 3723
rect 14933 3689 14967 3723
rect 3341 3621 3375 3655
rect 3801 3621 3835 3655
rect 5457 3621 5491 3655
rect 9137 3621 9171 3655
rect 4261 3553 4295 3587
rect 4353 3553 4387 3587
rect 6009 3553 6043 3587
rect 7297 3553 7331 3587
rect 7481 3553 7515 3587
rect 8585 3553 8619 3587
rect 9597 3553 9631 3587
rect 9689 3553 9723 3587
rect 10517 3553 10551 3587
rect 11253 3553 11287 3587
rect 12081 3553 12115 3587
rect 12357 3553 12391 3587
rect 12449 3553 12483 3587
rect 12725 3553 12759 3587
rect 14289 3553 14323 3587
rect 15393 3553 15427 3587
rect 15485 3553 15519 3587
rect 1685 3485 1719 3519
rect 2053 3485 2087 3519
rect 2329 3485 2363 3519
rect 2605 3485 2639 3519
rect 2881 3485 2915 3519
rect 3157 3485 3191 3519
rect 3525 3485 3559 3519
rect 3985 3485 4019 3519
rect 4445 3485 4479 3519
rect 5181 3485 5215 3519
rect 5825 3485 5859 3519
rect 6469 3485 6503 3519
rect 6561 3461 6595 3495
rect 7205 3485 7239 3519
rect 7941 3485 7975 3519
rect 8309 3485 8343 3519
rect 10333 3485 10367 3519
rect 13553 3485 13587 3519
rect 13645 3485 13679 3519
rect 15301 3485 15335 3519
rect 5917 3417 5951 3451
rect 8125 3417 8159 3451
rect 1869 3349 1903 3383
rect 2145 3349 2179 3383
rect 2421 3349 2455 3383
rect 2697 3349 2731 3383
rect 2973 3349 3007 3383
rect 4813 3349 4847 3383
rect 4997 3349 5031 3383
rect 5365 3349 5399 3383
rect 6745 3349 6779 3383
rect 8493 3349 8527 3383
rect 9505 3349 9539 3383
rect 10425 3349 10459 3383
rect 10793 3349 10827 3383
rect 13369 3349 13403 3383
rect 13829 3349 13863 3383
rect 14381 3349 14415 3383
rect 14473 3349 14507 3383
rect 14841 3349 14875 3383
rect 3801 3145 3835 3179
rect 4905 3145 4939 3179
rect 4997 3145 5031 3179
rect 5457 3145 5491 3179
rect 5917 3145 5951 3179
rect 7665 3145 7699 3179
rect 10057 3145 10091 3179
rect 10425 3145 10459 3179
rect 10977 3145 11011 3179
rect 2605 3077 2639 3111
rect 4169 3077 4203 3111
rect 5825 3077 5859 3111
rect 8033 3077 8067 3111
rect 15393 3077 15427 3111
rect 1685 3009 1719 3043
rect 2053 3009 2087 3043
rect 2421 3009 2455 3043
rect 2973 3009 3007 3043
rect 3341 3009 3375 3043
rect 3702 3009 3736 3043
rect 6646 3009 6680 3043
rect 7113 3009 7147 3043
rect 7205 3009 7239 3043
rect 8125 3009 8159 3043
rect 8493 3009 8527 3043
rect 9505 3009 9539 3043
rect 9965 3009 9999 3043
rect 11069 3009 11103 3043
rect 11529 3009 11563 3043
rect 12449 3009 12483 3043
rect 12725 3009 12759 3043
rect 13645 3009 13679 3043
rect 14657 3009 14691 3043
rect 14749 3009 14783 3043
rect 15117 3009 15151 3043
rect 4261 2941 4295 2975
rect 4445 2941 4479 2975
rect 4813 2941 4847 2975
rect 6101 2941 6135 2975
rect 7389 2941 7423 2975
rect 8217 2941 8251 2975
rect 8769 2941 8803 2975
rect 10517 2941 10551 2975
rect 10609 2941 10643 2975
rect 11805 2941 11839 2975
rect 13369 2941 13403 2975
rect 14841 2941 14875 2975
rect 3157 2873 3191 2907
rect 5365 2873 5399 2907
rect 6745 2873 6779 2907
rect 9689 2873 9723 2907
rect 14289 2873 14323 2907
rect 1501 2805 1535 2839
rect 1869 2805 1903 2839
rect 2237 2805 2271 2839
rect 2789 2805 2823 2839
rect 3525 2805 3559 2839
rect 6469 2805 6503 2839
rect 9781 2805 9815 2839
rect 11253 2805 11287 2839
rect 2329 2601 2363 2635
rect 4537 2601 4571 2635
rect 6561 2601 6595 2635
rect 9321 2601 9355 2635
rect 1961 2533 1995 2567
rect 2697 2533 2731 2567
rect 4261 2533 4295 2567
rect 7389 2533 7423 2567
rect 8125 2533 8159 2567
rect 13645 2533 13679 2567
rect 15577 2533 15611 2567
rect 5089 2465 5123 2499
rect 10793 2465 10827 2499
rect 11529 2465 11563 2499
rect 11805 2465 11839 2499
rect 14105 2465 14139 2499
rect 14381 2465 14415 2499
rect 1777 2397 1811 2431
rect 2145 2397 2179 2431
rect 2513 2397 2547 2431
rect 2881 2397 2915 2431
rect 3249 2397 3283 2431
rect 3617 2397 3651 2431
rect 4077 2397 4111 2431
rect 4445 2397 4479 2431
rect 4905 2397 4939 2431
rect 4997 2397 5031 2431
rect 5825 2397 5859 2431
rect 6193 2397 6227 2431
rect 6377 2397 6411 2431
rect 6929 2397 6963 2431
rect 7297 2397 7331 2431
rect 8309 2397 8343 2431
rect 9137 2397 9171 2431
rect 9413 2397 9447 2431
rect 9597 2397 9631 2431
rect 9873 2397 9907 2431
rect 10517 2397 10551 2431
rect 12449 2397 12483 2431
rect 12725 2397 12759 2431
rect 13461 2397 13495 2431
rect 13921 2397 13955 2431
rect 15025 2397 15059 2431
rect 15393 2397 15427 2431
rect 7573 2329 7607 2363
rect 7849 2329 7883 2363
rect 8493 2329 8527 2363
rect 8677 2329 8711 2363
rect 1593 2261 1627 2295
rect 3065 2261 3099 2295
rect 3433 2261 3467 2295
rect 3893 2261 3927 2295
rect 5457 2261 5491 2295
rect 5641 2261 5675 2295
rect 6009 2261 6043 2295
rect 6745 2261 6779 2295
rect 7113 2261 7147 2295
rect 7941 2261 7975 2295
rect 8953 2261 8987 2295
rect 13737 2261 13771 2295
rect 15209 2261 15243 2295
<< metal1 >>
rect 11698 17892 11704 17944
rect 11756 17932 11762 17944
rect 13078 17932 13084 17944
rect 11756 17904 13084 17932
rect 11756 17892 11762 17904
rect 13078 17892 13084 17904
rect 13136 17892 13142 17944
rect 9674 17824 9680 17876
rect 9732 17864 9738 17876
rect 10226 17864 10232 17876
rect 9732 17836 10232 17864
rect 9732 17824 9738 17836
rect 10226 17824 10232 17836
rect 10284 17864 10290 17876
rect 13722 17864 13728 17876
rect 10284 17836 13728 17864
rect 10284 17824 10290 17836
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 12434 17756 12440 17808
rect 12492 17796 12498 17808
rect 13354 17796 13360 17808
rect 12492 17768 13360 17796
rect 12492 17756 12498 17768
rect 13354 17756 13360 17768
rect 13412 17756 13418 17808
rect 9214 17688 9220 17740
rect 9272 17728 9278 17740
rect 13446 17728 13452 17740
rect 9272 17700 13452 17728
rect 9272 17688 9278 17700
rect 13446 17688 13452 17700
rect 13504 17688 13510 17740
rect 12618 17620 12624 17672
rect 12676 17660 12682 17672
rect 15654 17660 15660 17672
rect 12676 17632 15660 17660
rect 12676 17620 12682 17632
rect 15654 17620 15660 17632
rect 15712 17660 15718 17672
rect 16114 17660 16120 17672
rect 15712 17632 16120 17660
rect 15712 17620 15718 17632
rect 16114 17620 16120 17632
rect 16172 17620 16178 17672
rect 11330 17552 11336 17604
rect 11388 17592 11394 17604
rect 16482 17592 16488 17604
rect 11388 17564 16488 17592
rect 11388 17552 11394 17564
rect 16482 17552 16488 17564
rect 16540 17552 16546 17604
rect 12802 17484 12808 17536
rect 12860 17524 12866 17536
rect 13630 17524 13636 17536
rect 12860 17496 13636 17524
rect 12860 17484 12866 17496
rect 13630 17484 13636 17496
rect 13688 17484 13694 17536
rect 1104 17434 16008 17456
rect 1104 17382 4698 17434
rect 4750 17382 4762 17434
rect 4814 17382 4826 17434
rect 4878 17382 4890 17434
rect 4942 17382 4954 17434
rect 5006 17382 8446 17434
rect 8498 17382 8510 17434
rect 8562 17382 8574 17434
rect 8626 17382 8638 17434
rect 8690 17382 8702 17434
rect 8754 17382 12194 17434
rect 12246 17382 12258 17434
rect 12310 17382 12322 17434
rect 12374 17382 12386 17434
rect 12438 17382 12450 17434
rect 12502 17382 16008 17434
rect 1104 17360 16008 17382
rect 1394 17280 1400 17332
rect 1452 17320 1458 17332
rect 6365 17323 6423 17329
rect 6365 17320 6377 17323
rect 1452 17292 6377 17320
rect 1452 17280 1458 17292
rect 6365 17289 6377 17292
rect 6411 17289 6423 17323
rect 6365 17283 6423 17289
rect 6733 17323 6791 17329
rect 6733 17289 6745 17323
rect 6779 17320 6791 17323
rect 6914 17320 6920 17332
rect 6779 17292 6920 17320
rect 6779 17289 6791 17292
rect 6733 17283 6791 17289
rect 6914 17280 6920 17292
rect 6972 17280 6978 17332
rect 7101 17323 7159 17329
rect 7101 17289 7113 17323
rect 7147 17320 7159 17323
rect 7282 17320 7288 17332
rect 7147 17292 7288 17320
rect 7147 17289 7159 17292
rect 7101 17283 7159 17289
rect 7282 17280 7288 17292
rect 7340 17280 7346 17332
rect 7469 17323 7527 17329
rect 7469 17289 7481 17323
rect 7515 17320 7527 17323
rect 7650 17320 7656 17332
rect 7515 17292 7656 17320
rect 7515 17289 7527 17292
rect 7469 17283 7527 17289
rect 7650 17280 7656 17292
rect 7708 17280 7714 17332
rect 7837 17323 7895 17329
rect 7837 17289 7849 17323
rect 7883 17320 7895 17323
rect 8018 17320 8024 17332
rect 7883 17292 8024 17320
rect 7883 17289 7895 17292
rect 7837 17283 7895 17289
rect 8018 17280 8024 17292
rect 8076 17280 8082 17332
rect 8205 17323 8263 17329
rect 8205 17289 8217 17323
rect 8251 17320 8263 17323
rect 8294 17320 8300 17332
rect 8251 17292 8300 17320
rect 8251 17289 8263 17292
rect 8205 17283 8263 17289
rect 8294 17280 8300 17292
rect 8352 17280 8358 17332
rect 8573 17323 8631 17329
rect 8573 17289 8585 17323
rect 8619 17320 8631 17323
rect 8846 17320 8852 17332
rect 8619 17292 8852 17320
rect 8619 17289 8631 17292
rect 8573 17283 8631 17289
rect 8846 17280 8852 17292
rect 8904 17280 8910 17332
rect 9033 17323 9091 17329
rect 9033 17289 9045 17323
rect 9079 17320 9091 17323
rect 9122 17320 9128 17332
rect 9079 17292 9128 17320
rect 9079 17289 9091 17292
rect 9033 17283 9091 17289
rect 9122 17280 9128 17292
rect 9180 17280 9186 17332
rect 9401 17323 9459 17329
rect 9401 17289 9413 17323
rect 9447 17320 9459 17323
rect 9490 17320 9496 17332
rect 9447 17292 9496 17320
rect 9447 17289 9459 17292
rect 9401 17283 9459 17289
rect 9490 17280 9496 17292
rect 9548 17280 9554 17332
rect 11146 17320 11152 17332
rect 9646 17292 11152 17320
rect 2314 17212 2320 17264
rect 2372 17252 2378 17264
rect 5442 17252 5448 17264
rect 2372 17224 3004 17252
rect 2372 17212 2378 17224
rect 1765 17187 1823 17193
rect 1765 17153 1777 17187
rect 1811 17184 1823 17187
rect 2038 17184 2044 17196
rect 1811 17156 2044 17184
rect 1811 17153 1823 17156
rect 1765 17147 1823 17153
rect 2038 17144 2044 17156
rect 2096 17144 2102 17196
rect 2133 17187 2191 17193
rect 2133 17153 2145 17187
rect 2179 17153 2191 17187
rect 2498 17184 2504 17196
rect 2459 17156 2504 17184
rect 2133 17147 2191 17153
rect 2148 17116 2176 17147
rect 2498 17144 2504 17156
rect 2556 17144 2562 17196
rect 2976 17193 3004 17224
rect 4724 17224 5448 17252
rect 2869 17187 2927 17193
rect 2869 17153 2881 17187
rect 2915 17153 2927 17187
rect 2869 17147 2927 17153
rect 2961 17187 3019 17193
rect 2961 17153 2973 17187
rect 3007 17153 3019 17187
rect 3326 17184 3332 17196
rect 3287 17156 3332 17184
rect 2961 17147 3019 17153
rect 2590 17116 2596 17128
rect 2148 17088 2596 17116
rect 2590 17076 2596 17088
rect 2648 17076 2654 17128
rect 2884 17116 2912 17147
rect 3326 17144 3332 17156
rect 3384 17144 3390 17196
rect 3786 17184 3792 17196
rect 3747 17156 3792 17184
rect 3786 17144 3792 17156
rect 3844 17144 3850 17196
rect 3878 17144 3884 17196
rect 3936 17184 3942 17196
rect 4157 17187 4215 17193
rect 4157 17184 4169 17187
rect 3936 17156 4169 17184
rect 3936 17144 3942 17156
rect 4157 17153 4169 17156
rect 4203 17153 4215 17187
rect 4157 17147 4215 17153
rect 4338 17144 4344 17196
rect 4396 17184 4402 17196
rect 4525 17187 4583 17193
rect 4525 17184 4537 17187
rect 4396 17156 4537 17184
rect 4396 17144 4402 17156
rect 4525 17153 4537 17156
rect 4571 17153 4583 17187
rect 4525 17147 4583 17153
rect 3418 17116 3424 17128
rect 2884 17088 3424 17116
rect 3418 17076 3424 17088
rect 3476 17076 3482 17128
rect 1581 17051 1639 17057
rect 1581 17017 1593 17051
rect 1627 17048 1639 17051
rect 1670 17048 1676 17060
rect 1627 17020 1676 17048
rect 1627 17017 1639 17020
rect 1581 17011 1639 17017
rect 1670 17008 1676 17020
rect 1728 17008 1734 17060
rect 3145 17051 3203 17057
rect 3145 17017 3157 17051
rect 3191 17048 3203 17051
rect 3234 17048 3240 17060
rect 3191 17020 3240 17048
rect 3191 17017 3203 17020
rect 3145 17011 3203 17017
rect 3234 17008 3240 17020
rect 3292 17008 3298 17060
rect 3513 17051 3571 17057
rect 3513 17017 3525 17051
rect 3559 17048 3571 17051
rect 3602 17048 3608 17060
rect 3559 17020 3608 17048
rect 3559 17017 3571 17020
rect 3513 17011 3571 17017
rect 3602 17008 3608 17020
rect 3660 17008 3666 17060
rect 3970 17048 3976 17060
rect 3931 17020 3976 17048
rect 3970 17008 3976 17020
rect 4028 17008 4034 17060
rect 4341 17051 4399 17057
rect 4341 17017 4353 17051
rect 4387 17048 4399 17051
rect 4614 17048 4620 17060
rect 4387 17020 4620 17048
rect 4387 17017 4399 17020
rect 4341 17011 4399 17017
rect 4614 17008 4620 17020
rect 4672 17008 4678 17060
rect 4724 17057 4752 17224
rect 5442 17212 5448 17224
rect 5500 17212 5506 17264
rect 5721 17255 5779 17261
rect 5721 17221 5733 17255
rect 5767 17252 5779 17255
rect 6270 17252 6276 17264
rect 5767 17224 6276 17252
rect 5767 17221 5779 17224
rect 5721 17215 5779 17221
rect 6270 17212 6276 17224
rect 6328 17212 6334 17264
rect 9306 17212 9312 17264
rect 9364 17252 9370 17264
rect 9646 17252 9674 17292
rect 11146 17280 11152 17292
rect 11204 17280 11210 17332
rect 11514 17280 11520 17332
rect 11572 17320 11578 17332
rect 15565 17323 15623 17329
rect 15565 17320 15577 17323
rect 11572 17292 15577 17320
rect 11572 17280 11578 17292
rect 15565 17289 15577 17292
rect 15611 17289 15623 17323
rect 15565 17283 15623 17289
rect 9364 17224 9674 17252
rect 10045 17255 10103 17261
rect 9364 17212 9370 17224
rect 10045 17221 10057 17255
rect 10091 17252 10103 17255
rect 15013 17255 15071 17261
rect 15013 17252 15025 17255
rect 10091 17224 15025 17252
rect 10091 17221 10103 17224
rect 10045 17215 10103 17221
rect 15013 17221 15025 17224
rect 15059 17221 15071 17255
rect 15013 17215 15071 17221
rect 5166 17184 5172 17196
rect 5127 17156 5172 17184
rect 5166 17144 5172 17156
rect 5224 17144 5230 17196
rect 5626 17184 5632 17196
rect 5587 17156 5632 17184
rect 5626 17144 5632 17156
rect 5684 17144 5690 17196
rect 5994 17144 6000 17196
rect 6052 17184 6058 17196
rect 6549 17187 6607 17193
rect 6549 17184 6561 17187
rect 6052 17156 6561 17184
rect 6052 17144 6058 17156
rect 6549 17153 6561 17156
rect 6595 17153 6607 17187
rect 6549 17147 6607 17153
rect 6917 17187 6975 17193
rect 6917 17153 6929 17187
rect 6963 17153 6975 17187
rect 7282 17184 7288 17196
rect 7243 17156 7288 17184
rect 6917 17147 6975 17153
rect 5905 17119 5963 17125
rect 5000 17088 5580 17116
rect 4709 17051 4767 17057
rect 4709 17017 4721 17051
rect 4755 17017 4767 17051
rect 4709 17011 4767 17017
rect 1949 16983 2007 16989
rect 1949 16949 1961 16983
rect 1995 16980 2007 16983
rect 2130 16980 2136 16992
rect 1995 16952 2136 16980
rect 1995 16949 2007 16952
rect 1949 16943 2007 16949
rect 2130 16940 2136 16952
rect 2188 16940 2194 16992
rect 2317 16983 2375 16989
rect 2317 16949 2329 16983
rect 2363 16980 2375 16983
rect 2406 16980 2412 16992
rect 2363 16952 2412 16980
rect 2363 16949 2375 16952
rect 2317 16943 2375 16949
rect 2406 16940 2412 16952
rect 2464 16940 2470 16992
rect 2685 16983 2743 16989
rect 2685 16949 2697 16983
rect 2731 16980 2743 16983
rect 2866 16980 2872 16992
rect 2731 16952 2872 16980
rect 2731 16949 2743 16952
rect 2685 16943 2743 16949
rect 2866 16940 2872 16952
rect 2924 16940 2930 16992
rect 5000 16989 5028 17088
rect 5552 17048 5580 17088
rect 5905 17085 5917 17119
rect 5951 17116 5963 17119
rect 6932 17116 6960 17147
rect 7282 17144 7288 17156
rect 7340 17144 7346 17196
rect 7650 17184 7656 17196
rect 7611 17156 7656 17184
rect 7650 17144 7656 17156
rect 7708 17144 7714 17196
rect 8021 17187 8079 17193
rect 8021 17153 8033 17187
rect 8067 17153 8079 17187
rect 8386 17184 8392 17196
rect 8347 17156 8392 17184
rect 8021 17147 8079 17153
rect 7558 17116 7564 17128
rect 5951 17088 6868 17116
rect 6932 17088 7564 17116
rect 5951 17085 5963 17088
rect 5905 17079 5963 17085
rect 6178 17048 6184 17060
rect 5552 17020 6184 17048
rect 6178 17008 6184 17020
rect 6236 17008 6242 17060
rect 4985 16983 5043 16989
rect 4985 16949 4997 16983
rect 5031 16949 5043 16983
rect 5258 16980 5264 16992
rect 5219 16952 5264 16980
rect 4985 16943 5043 16949
rect 5258 16940 5264 16952
rect 5316 16940 5322 16992
rect 5534 16940 5540 16992
rect 5592 16980 5598 16992
rect 6089 16983 6147 16989
rect 6089 16980 6101 16983
rect 5592 16952 6101 16980
rect 5592 16940 5598 16952
rect 6089 16949 6101 16952
rect 6135 16949 6147 16983
rect 6840 16980 6868 17088
rect 7558 17076 7564 17088
rect 7616 17076 7622 17128
rect 8036 17116 8064 17147
rect 8386 17144 8392 17156
rect 8444 17144 8450 17196
rect 8757 17187 8815 17193
rect 8757 17153 8769 17187
rect 8803 17153 8815 17187
rect 9214 17184 9220 17196
rect 9175 17156 9220 17184
rect 8757 17147 8815 17153
rect 8294 17116 8300 17128
rect 8036 17088 8300 17116
rect 8294 17076 8300 17088
rect 8352 17076 8358 17128
rect 8772 17048 8800 17147
rect 9214 17144 9220 17156
rect 9272 17144 9278 17196
rect 9585 17187 9643 17193
rect 9585 17153 9597 17187
rect 9631 17184 9643 17187
rect 11330 17184 11336 17196
rect 9631 17156 11192 17184
rect 11291 17156 11336 17184
rect 9631 17153 9643 17156
rect 9585 17147 9643 17153
rect 9766 17116 9772 17128
rect 9727 17088 9772 17116
rect 9766 17076 9772 17088
rect 9824 17076 9830 17128
rect 9950 17076 9956 17128
rect 10008 17116 10014 17128
rect 10778 17116 10784 17128
rect 10008 17088 10784 17116
rect 10008 17076 10014 17088
rect 10778 17076 10784 17088
rect 10836 17076 10842 17128
rect 11057 17119 11115 17125
rect 11057 17085 11069 17119
rect 11103 17085 11115 17119
rect 11164 17116 11192 17156
rect 11330 17144 11336 17156
rect 11388 17144 11394 17196
rect 11440 17156 11928 17184
rect 11440 17116 11468 17156
rect 11164 17088 11468 17116
rect 11057 17079 11115 17085
rect 11072 17048 11100 17079
rect 11514 17076 11520 17128
rect 11572 17116 11578 17128
rect 11790 17116 11796 17128
rect 11572 17088 11617 17116
rect 11751 17088 11796 17116
rect 11572 17076 11578 17088
rect 11790 17076 11796 17088
rect 11848 17076 11854 17128
rect 11900 17116 11928 17156
rect 12066 17144 12072 17196
rect 12124 17184 12130 17196
rect 13262 17184 13268 17196
rect 12124 17156 13268 17184
rect 12124 17144 12130 17156
rect 13262 17144 13268 17156
rect 13320 17144 13326 17196
rect 13541 17187 13599 17193
rect 13541 17153 13553 17187
rect 13587 17153 13599 17187
rect 13722 17184 13728 17196
rect 13683 17156 13728 17184
rect 13541 17147 13599 17153
rect 12894 17116 12900 17128
rect 11900 17088 12900 17116
rect 12894 17076 12900 17088
rect 12952 17076 12958 17128
rect 12986 17076 12992 17128
rect 13044 17116 13050 17128
rect 13044 17088 13089 17116
rect 13044 17076 13050 17088
rect 12710 17048 12716 17060
rect 8772 17020 11008 17048
rect 11072 17020 12716 17048
rect 9214 16980 9220 16992
rect 6840 16952 9220 16980
rect 6089 16943 6147 16949
rect 9214 16940 9220 16952
rect 9272 16940 9278 16992
rect 10134 16940 10140 16992
rect 10192 16980 10198 16992
rect 10413 16983 10471 16989
rect 10413 16980 10425 16983
rect 10192 16952 10425 16980
rect 10192 16940 10198 16952
rect 10413 16949 10425 16952
rect 10459 16949 10471 16983
rect 10980 16980 11008 17020
rect 12710 17008 12716 17020
rect 12768 17008 12774 17060
rect 13078 17008 13084 17060
rect 13136 17048 13142 17060
rect 13556 17048 13584 17147
rect 13722 17144 13728 17156
rect 13780 17144 13786 17196
rect 13906 17144 13912 17196
rect 13964 17184 13970 17196
rect 15473 17187 15531 17193
rect 15473 17184 15485 17187
rect 13964 17156 15485 17184
rect 13964 17144 13970 17156
rect 15473 17153 15485 17156
rect 15519 17184 15531 17187
rect 16022 17184 16028 17196
rect 15519 17156 16028 17184
rect 15519 17153 15531 17156
rect 15473 17147 15531 17153
rect 16022 17144 16028 17156
rect 16080 17144 16086 17196
rect 13630 17076 13636 17128
rect 13688 17116 13694 17128
rect 14093 17119 14151 17125
rect 14093 17116 14105 17119
rect 13688 17088 14105 17116
rect 13688 17076 13694 17088
rect 14093 17085 14105 17088
rect 14139 17085 14151 17119
rect 14093 17079 14151 17085
rect 14369 17119 14427 17125
rect 14369 17085 14381 17119
rect 14415 17116 14427 17119
rect 16574 17116 16580 17128
rect 14415 17088 16580 17116
rect 14415 17085 14427 17088
rect 14369 17079 14427 17085
rect 16574 17076 16580 17088
rect 16632 17076 16638 17128
rect 13136 17020 13584 17048
rect 13136 17008 13142 17020
rect 12250 16980 12256 16992
rect 10980 16952 12256 16980
rect 10413 16943 10471 16949
rect 12250 16940 12256 16952
rect 12308 16940 12314 16992
rect 13449 16983 13507 16989
rect 13449 16949 13461 16983
rect 13495 16980 13507 16983
rect 13722 16980 13728 16992
rect 13495 16952 13728 16980
rect 13495 16949 13507 16952
rect 13449 16943 13507 16949
rect 13722 16940 13728 16952
rect 13780 16940 13786 16992
rect 13909 16983 13967 16989
rect 13909 16949 13921 16983
rect 13955 16980 13967 16983
rect 15194 16980 15200 16992
rect 13955 16952 15200 16980
rect 13955 16949 13967 16952
rect 13909 16943 13967 16949
rect 15194 16940 15200 16952
rect 15252 16940 15258 16992
rect 15289 16983 15347 16989
rect 15289 16949 15301 16983
rect 15335 16980 15347 16983
rect 16390 16980 16396 16992
rect 15335 16952 16396 16980
rect 15335 16949 15347 16952
rect 15289 16943 15347 16949
rect 16390 16940 16396 16952
rect 16448 16940 16454 16992
rect 1104 16890 16008 16912
rect 1104 16838 2824 16890
rect 2876 16838 2888 16890
rect 2940 16838 2952 16890
rect 3004 16838 3016 16890
rect 3068 16838 3080 16890
rect 3132 16838 6572 16890
rect 6624 16838 6636 16890
rect 6688 16838 6700 16890
rect 6752 16838 6764 16890
rect 6816 16838 6828 16890
rect 6880 16838 10320 16890
rect 10372 16838 10384 16890
rect 10436 16838 10448 16890
rect 10500 16838 10512 16890
rect 10564 16838 10576 16890
rect 10628 16838 14068 16890
rect 14120 16838 14132 16890
rect 14184 16838 14196 16890
rect 14248 16838 14260 16890
rect 14312 16838 14324 16890
rect 14376 16838 16008 16890
rect 1104 16816 16008 16838
rect 5994 16776 6000 16788
rect 2746 16748 6000 16776
rect 1762 16668 1768 16720
rect 1820 16708 1826 16720
rect 2746 16708 2774 16748
rect 5994 16736 6000 16748
rect 6052 16736 6058 16788
rect 6270 16736 6276 16788
rect 6328 16776 6334 16788
rect 6825 16779 6883 16785
rect 6825 16776 6837 16779
rect 6328 16748 6837 16776
rect 6328 16736 6334 16748
rect 6825 16745 6837 16748
rect 6871 16745 6883 16779
rect 6825 16739 6883 16745
rect 7282 16736 7288 16788
rect 7340 16776 7346 16788
rect 7653 16779 7711 16785
rect 7653 16776 7665 16779
rect 7340 16748 7665 16776
rect 7340 16736 7346 16748
rect 7653 16745 7665 16748
rect 7699 16745 7711 16779
rect 7653 16739 7711 16745
rect 8386 16736 8392 16788
rect 8444 16776 8450 16788
rect 9125 16779 9183 16785
rect 9125 16776 9137 16779
rect 8444 16748 9137 16776
rect 8444 16736 8450 16748
rect 9125 16745 9137 16748
rect 9171 16745 9183 16779
rect 9858 16776 9864 16788
rect 9125 16739 9183 16745
rect 9232 16748 9864 16776
rect 1820 16680 2774 16708
rect 3329 16711 3387 16717
rect 1820 16668 1826 16680
rect 3329 16677 3341 16711
rect 3375 16708 3387 16711
rect 3786 16708 3792 16720
rect 3375 16680 3792 16708
rect 3375 16677 3387 16680
rect 3329 16671 3387 16677
rect 3786 16668 3792 16680
rect 3844 16668 3850 16720
rect 4065 16711 4123 16717
rect 4065 16677 4077 16711
rect 4111 16677 4123 16711
rect 4338 16708 4344 16720
rect 4299 16680 4344 16708
rect 4065 16671 4123 16677
rect 4080 16640 4108 16671
rect 4338 16668 4344 16680
rect 4396 16668 4402 16720
rect 7926 16668 7932 16720
rect 7984 16708 7990 16720
rect 9232 16708 9260 16748
rect 9858 16736 9864 16748
rect 9916 16736 9922 16788
rect 10226 16776 10232 16788
rect 10187 16748 10232 16776
rect 10226 16736 10232 16748
rect 10284 16736 10290 16788
rect 10318 16736 10324 16788
rect 10376 16776 10382 16788
rect 11425 16779 11483 16785
rect 11425 16776 11437 16779
rect 10376 16748 11437 16776
rect 10376 16736 10382 16748
rect 11425 16745 11437 16748
rect 11471 16745 11483 16779
rect 12434 16776 12440 16788
rect 11425 16739 11483 16745
rect 12176 16748 12440 16776
rect 10413 16711 10471 16717
rect 10413 16708 10425 16711
rect 7984 16680 9260 16708
rect 9324 16680 9674 16708
rect 7984 16668 7990 16680
rect 7466 16640 7472 16652
rect 1412 16612 1900 16640
rect 4080 16612 4568 16640
rect 7427 16612 7472 16640
rect 290 16532 296 16584
rect 348 16572 354 16584
rect 1412 16572 1440 16612
rect 348 16544 1440 16572
rect 348 16532 354 16544
rect 1486 16532 1492 16584
rect 1544 16572 1550 16584
rect 1762 16572 1768 16584
rect 1544 16544 1637 16572
rect 1723 16544 1768 16572
rect 1544 16532 1550 16544
rect 1762 16532 1768 16544
rect 1820 16532 1826 16584
rect 1872 16572 1900 16612
rect 2317 16575 2375 16581
rect 1872 16544 2268 16572
rect 1504 16504 1532 16532
rect 2038 16504 2044 16516
rect 1504 16476 2044 16504
rect 2038 16464 2044 16476
rect 2096 16464 2102 16516
rect 1578 16396 1584 16448
rect 1636 16436 1642 16448
rect 2133 16439 2191 16445
rect 2133 16436 2145 16439
rect 1636 16408 2145 16436
rect 1636 16396 1642 16408
rect 2133 16405 2145 16408
rect 2179 16405 2191 16439
rect 2240 16436 2268 16544
rect 2317 16541 2329 16575
rect 2363 16541 2375 16575
rect 2317 16535 2375 16541
rect 2332 16504 2360 16535
rect 2406 16532 2412 16584
rect 2464 16572 2470 16584
rect 3050 16572 3056 16584
rect 2464 16544 2509 16572
rect 3011 16544 3056 16572
rect 2464 16532 2470 16544
rect 3050 16532 3056 16544
rect 3108 16532 3114 16584
rect 3142 16532 3148 16584
rect 3200 16572 3206 16584
rect 3421 16575 3479 16581
rect 3200 16544 3245 16572
rect 3200 16532 3206 16544
rect 3421 16541 3433 16575
rect 3467 16572 3479 16575
rect 3786 16572 3792 16584
rect 3467 16544 3792 16572
rect 3467 16541 3479 16544
rect 3421 16535 3479 16541
rect 3786 16532 3792 16544
rect 3844 16532 3850 16584
rect 3881 16575 3939 16581
rect 3881 16541 3893 16575
rect 3927 16572 3939 16575
rect 4062 16572 4068 16584
rect 3927 16544 4068 16572
rect 3927 16541 3939 16544
rect 3881 16535 3939 16541
rect 4062 16532 4068 16544
rect 4120 16532 4126 16584
rect 4157 16575 4215 16581
rect 4157 16541 4169 16575
rect 4203 16541 4215 16575
rect 4157 16535 4215 16541
rect 2682 16504 2688 16516
rect 2332 16476 2688 16504
rect 2682 16464 2688 16476
rect 2740 16464 2746 16516
rect 2593 16439 2651 16445
rect 2593 16436 2605 16439
rect 2240 16408 2605 16436
rect 2133 16399 2191 16405
rect 2593 16405 2605 16408
rect 2639 16405 2651 16439
rect 2866 16436 2872 16448
rect 2827 16408 2872 16436
rect 2593 16399 2651 16405
rect 2866 16396 2872 16408
rect 2924 16396 2930 16448
rect 3605 16439 3663 16445
rect 3605 16405 3617 16439
rect 3651 16436 3663 16439
rect 3878 16436 3884 16448
rect 3651 16408 3884 16436
rect 3651 16405 3663 16408
rect 3605 16399 3663 16405
rect 3878 16396 3884 16408
rect 3936 16396 3942 16448
rect 4172 16436 4200 16535
rect 4246 16532 4252 16584
rect 4304 16572 4310 16584
rect 4433 16575 4491 16581
rect 4433 16572 4445 16575
rect 4304 16544 4445 16572
rect 4304 16532 4310 16544
rect 4433 16541 4445 16544
rect 4479 16541 4491 16575
rect 4540 16572 4568 16612
rect 7466 16600 7472 16612
rect 7524 16600 7530 16652
rect 8496 16649 8524 16680
rect 8481 16643 8539 16649
rect 7668 16612 7972 16640
rect 5626 16581 5632 16584
rect 4985 16575 5043 16581
rect 4985 16572 4997 16575
rect 4540 16544 4997 16572
rect 4433 16535 4491 16541
rect 4985 16541 4997 16544
rect 5031 16541 5043 16575
rect 4985 16535 5043 16541
rect 5353 16575 5411 16581
rect 5353 16541 5365 16575
rect 5399 16541 5411 16575
rect 5620 16572 5632 16581
rect 5587 16544 5632 16572
rect 5353 16535 5411 16541
rect 5620 16535 5632 16544
rect 5368 16504 5396 16535
rect 5626 16532 5632 16535
rect 5684 16532 5690 16584
rect 7193 16575 7251 16581
rect 7193 16541 7205 16575
rect 7239 16572 7251 16575
rect 7668 16572 7696 16612
rect 7834 16572 7840 16584
rect 7239 16544 7696 16572
rect 7795 16544 7840 16572
rect 7239 16541 7251 16544
rect 7193 16535 7251 16541
rect 7834 16532 7840 16544
rect 7892 16532 7898 16584
rect 7944 16572 7972 16612
rect 8481 16609 8493 16643
rect 8527 16609 8539 16643
rect 9324 16640 9352 16680
rect 8481 16603 8539 16609
rect 9232 16612 9352 16640
rect 9646 16640 9674 16680
rect 9784 16680 10425 16708
rect 9784 16640 9812 16680
rect 10413 16677 10425 16680
rect 10459 16677 10471 16711
rect 10413 16671 10471 16677
rect 10502 16668 10508 16720
rect 10560 16708 10566 16720
rect 11790 16708 11796 16720
rect 10560 16680 11796 16708
rect 10560 16668 10566 16680
rect 11790 16668 11796 16680
rect 11848 16668 11854 16720
rect 9646 16612 9812 16640
rect 8389 16575 8447 16581
rect 7944 16544 8340 16572
rect 4816 16476 5396 16504
rect 7285 16507 7343 16513
rect 4338 16436 4344 16448
rect 4172 16408 4344 16436
rect 4338 16396 4344 16408
rect 4396 16396 4402 16448
rect 4430 16396 4436 16448
rect 4488 16436 4494 16448
rect 4617 16439 4675 16445
rect 4617 16436 4629 16439
rect 4488 16408 4629 16436
rect 4488 16396 4494 16408
rect 4617 16405 4629 16408
rect 4663 16405 4675 16439
rect 4617 16399 4675 16405
rect 4706 16396 4712 16448
rect 4764 16436 4770 16448
rect 4816 16445 4844 16476
rect 7285 16473 7297 16507
rect 7331 16504 7343 16507
rect 8312 16504 8340 16544
rect 8389 16541 8401 16575
rect 8435 16572 8447 16575
rect 9232 16572 9260 16612
rect 9858 16600 9864 16652
rect 9916 16640 9922 16652
rect 9953 16643 10011 16649
rect 9953 16640 9965 16643
rect 9916 16612 9965 16640
rect 9916 16600 9922 16612
rect 9953 16609 9965 16612
rect 9999 16609 10011 16643
rect 10965 16643 11023 16649
rect 10965 16640 10977 16643
rect 9953 16603 10011 16609
rect 10253 16612 10977 16640
rect 8435 16544 9260 16572
rect 9309 16575 9367 16581
rect 8435 16541 8447 16544
rect 8389 16535 8447 16541
rect 9309 16541 9321 16575
rect 9355 16572 9367 16575
rect 10042 16572 10048 16584
rect 9355 16544 10048 16572
rect 9355 16541 9367 16544
rect 9309 16535 9367 16541
rect 10042 16532 10048 16544
rect 10100 16532 10106 16584
rect 7331 16476 7972 16504
rect 8312 16476 9444 16504
rect 7331 16473 7343 16476
rect 7285 16467 7343 16473
rect 4801 16439 4859 16445
rect 4801 16436 4813 16439
rect 4764 16408 4813 16436
rect 4764 16396 4770 16408
rect 4801 16405 4813 16408
rect 4847 16405 4859 16439
rect 4801 16399 4859 16405
rect 5074 16396 5080 16448
rect 5132 16436 5138 16448
rect 5169 16439 5227 16445
rect 5169 16436 5181 16439
rect 5132 16408 5181 16436
rect 5132 16396 5138 16408
rect 5169 16405 5181 16408
rect 5215 16405 5227 16439
rect 5169 16399 5227 16405
rect 6733 16439 6791 16445
rect 6733 16405 6745 16439
rect 6779 16436 6791 16439
rect 7006 16436 7012 16448
rect 6779 16408 7012 16436
rect 6779 16405 6791 16408
rect 6733 16399 6791 16405
rect 7006 16396 7012 16408
rect 7064 16396 7070 16448
rect 7944 16445 7972 16476
rect 7929 16439 7987 16445
rect 7929 16405 7941 16439
rect 7975 16405 7987 16439
rect 7929 16399 7987 16405
rect 8297 16439 8355 16445
rect 8297 16405 8309 16439
rect 8343 16436 8355 16439
rect 8386 16436 8392 16448
rect 8343 16408 8392 16436
rect 8343 16405 8355 16408
rect 8297 16399 8355 16405
rect 8386 16396 8392 16408
rect 8444 16396 8450 16448
rect 9033 16439 9091 16445
rect 9033 16405 9045 16439
rect 9079 16436 9091 16439
rect 9306 16436 9312 16448
rect 9079 16408 9312 16436
rect 9079 16405 9091 16408
rect 9033 16399 9091 16405
rect 9306 16396 9312 16408
rect 9364 16396 9370 16448
rect 9416 16445 9444 16476
rect 9490 16464 9496 16516
rect 9548 16504 9554 16516
rect 10253 16504 10281 16612
rect 10965 16609 10977 16612
rect 11011 16609 11023 16643
rect 10965 16603 11023 16609
rect 11146 16600 11152 16652
rect 11204 16600 11210 16652
rect 12176 16649 12204 16748
rect 12434 16736 12440 16748
rect 12492 16736 12498 16788
rect 12894 16736 12900 16788
rect 12952 16776 12958 16788
rect 13725 16779 13783 16785
rect 13725 16776 13737 16779
rect 12952 16748 13737 16776
rect 12952 16736 12958 16748
rect 13725 16745 13737 16748
rect 13771 16745 13783 16779
rect 13725 16739 13783 16745
rect 15657 16779 15715 16785
rect 15657 16745 15669 16779
rect 15703 16776 15715 16779
rect 16482 16776 16488 16788
rect 15703 16748 16488 16776
rect 15703 16745 15715 16748
rect 15657 16739 15715 16745
rect 16482 16736 16488 16748
rect 16540 16736 16546 16788
rect 12250 16668 12256 16720
rect 12308 16708 12314 16720
rect 15289 16711 15347 16717
rect 15289 16708 15301 16711
rect 12308 16680 15301 16708
rect 12308 16668 12314 16680
rect 15289 16677 15301 16680
rect 15335 16677 15347 16711
rect 15289 16671 15347 16677
rect 12161 16643 12219 16649
rect 12161 16609 12173 16643
rect 12207 16609 12219 16643
rect 12161 16603 12219 16609
rect 12437 16643 12495 16649
rect 12437 16609 12449 16643
rect 12483 16609 12495 16643
rect 12437 16603 12495 16609
rect 10873 16575 10931 16581
rect 10873 16541 10885 16575
rect 10919 16572 10931 16575
rect 10919 16568 11054 16572
rect 11164 16568 11192 16600
rect 10919 16544 11192 16568
rect 10919 16541 10931 16544
rect 10873 16535 10931 16541
rect 11026 16540 11192 16544
rect 11238 16532 11244 16584
rect 11296 16572 11302 16584
rect 12452 16572 12480 16603
rect 13354 16600 13360 16652
rect 13412 16640 13418 16652
rect 14090 16640 14096 16652
rect 13412 16612 13457 16640
rect 14051 16612 14096 16640
rect 13412 16600 13418 16612
rect 14090 16600 14096 16612
rect 14148 16600 14154 16652
rect 14369 16643 14427 16649
rect 14369 16609 14381 16643
rect 14415 16640 14427 16643
rect 14826 16640 14832 16652
rect 14415 16612 14832 16640
rect 14415 16609 14427 16612
rect 14369 16603 14427 16609
rect 14826 16600 14832 16612
rect 14884 16600 14890 16652
rect 12618 16572 12624 16584
rect 11296 16544 11744 16572
rect 12452 16544 12624 16572
rect 11296 16532 11302 16544
rect 9548 16476 10281 16504
rect 9548 16464 9554 16476
rect 10410 16464 10416 16516
rect 10468 16504 10474 16516
rect 10781 16507 10839 16513
rect 10781 16504 10793 16507
rect 10468 16476 10793 16504
rect 10468 16464 10474 16476
rect 10781 16473 10793 16476
rect 10827 16504 10839 16507
rect 11333 16507 11391 16513
rect 11333 16504 11345 16507
rect 10827 16476 11345 16504
rect 10827 16473 10839 16476
rect 10781 16467 10839 16473
rect 11333 16473 11345 16476
rect 11379 16473 11391 16507
rect 11716 16504 11744 16544
rect 12618 16532 12624 16544
rect 12676 16532 12682 16584
rect 12710 16532 12716 16584
rect 12768 16572 12774 16584
rect 12986 16572 12992 16584
rect 12768 16544 12992 16572
rect 12768 16532 12774 16544
rect 12986 16532 12992 16544
rect 13044 16532 13050 16584
rect 13078 16532 13084 16584
rect 13136 16572 13142 16584
rect 13449 16575 13507 16581
rect 13136 16544 13181 16572
rect 13136 16532 13142 16544
rect 13449 16541 13461 16575
rect 13495 16572 13507 16575
rect 13630 16572 13636 16584
rect 13495 16544 13636 16572
rect 13495 16541 13507 16544
rect 13449 16535 13507 16541
rect 13630 16532 13636 16544
rect 13688 16532 13694 16584
rect 13909 16575 13967 16581
rect 13909 16541 13921 16575
rect 13955 16572 13967 16575
rect 15197 16575 15255 16581
rect 13955 16544 15148 16572
rect 13955 16541 13967 16544
rect 13909 16535 13967 16541
rect 12894 16504 12900 16516
rect 11716 16476 12900 16504
rect 11333 16467 11391 16473
rect 12894 16464 12900 16476
rect 12952 16464 12958 16516
rect 13262 16464 13268 16516
rect 13320 16504 13326 16516
rect 13814 16504 13820 16516
rect 13320 16476 13820 16504
rect 13320 16464 13326 16476
rect 13814 16464 13820 16476
rect 13872 16464 13878 16516
rect 9401 16439 9459 16445
rect 9401 16405 9413 16439
rect 9447 16405 9459 16439
rect 9401 16399 9459 16405
rect 9582 16396 9588 16448
rect 9640 16436 9646 16448
rect 9769 16439 9827 16445
rect 9769 16436 9781 16439
rect 9640 16408 9781 16436
rect 9640 16396 9646 16408
rect 9769 16405 9781 16408
rect 9815 16405 9827 16439
rect 9769 16399 9827 16405
rect 9861 16439 9919 16445
rect 9861 16405 9873 16439
rect 9907 16436 9919 16439
rect 11146 16436 11152 16448
rect 9907 16408 11152 16436
rect 9907 16405 9919 16408
rect 9861 16399 9919 16405
rect 11146 16396 11152 16408
rect 11204 16436 11210 16448
rect 12066 16436 12072 16448
rect 11204 16408 12072 16436
rect 11204 16396 11210 16408
rect 12066 16396 12072 16408
rect 12124 16396 12130 16448
rect 12618 16396 12624 16448
rect 12676 16436 12682 16448
rect 13633 16439 13691 16445
rect 13633 16436 13645 16439
rect 12676 16408 13645 16436
rect 12676 16396 12682 16408
rect 13633 16405 13645 16408
rect 13679 16405 13691 16439
rect 15010 16436 15016 16448
rect 14971 16408 15016 16436
rect 13633 16399 13691 16405
rect 15010 16396 15016 16408
rect 15068 16396 15074 16448
rect 15120 16436 15148 16544
rect 15197 16541 15209 16575
rect 15243 16541 15255 16575
rect 15197 16535 15255 16541
rect 15473 16575 15531 16581
rect 15473 16541 15485 16575
rect 15519 16572 15531 16575
rect 15838 16572 15844 16584
rect 15519 16544 15844 16572
rect 15519 16541 15531 16544
rect 15473 16535 15531 16541
rect 15212 16504 15240 16535
rect 15838 16532 15844 16544
rect 15896 16532 15902 16584
rect 16574 16504 16580 16516
rect 15212 16476 16580 16504
rect 16574 16464 16580 16476
rect 16632 16464 16638 16516
rect 15562 16436 15568 16448
rect 15120 16408 15568 16436
rect 15562 16396 15568 16408
rect 15620 16396 15626 16448
rect 1104 16346 16008 16368
rect 1104 16294 4698 16346
rect 4750 16294 4762 16346
rect 4814 16294 4826 16346
rect 4878 16294 4890 16346
rect 4942 16294 4954 16346
rect 5006 16294 8446 16346
rect 8498 16294 8510 16346
rect 8562 16294 8574 16346
rect 8626 16294 8638 16346
rect 8690 16294 8702 16346
rect 8754 16294 12194 16346
rect 12246 16294 12258 16346
rect 12310 16294 12322 16346
rect 12374 16294 12386 16346
rect 12438 16294 12450 16346
rect 12502 16294 16008 16346
rect 1104 16272 16008 16294
rect 1486 16232 1492 16244
rect 1447 16204 1492 16232
rect 1486 16192 1492 16204
rect 1544 16192 1550 16244
rect 1854 16232 1860 16244
rect 1815 16204 1860 16232
rect 1854 16192 1860 16204
rect 1912 16192 1918 16244
rect 2314 16232 2320 16244
rect 2275 16204 2320 16232
rect 2314 16192 2320 16204
rect 2372 16192 2378 16244
rect 2593 16235 2651 16241
rect 2593 16201 2605 16235
rect 2639 16201 2651 16235
rect 2593 16195 2651 16201
rect 3237 16235 3295 16241
rect 3237 16201 3249 16235
rect 3283 16232 3295 16235
rect 3326 16232 3332 16244
rect 3283 16204 3332 16232
rect 3283 16201 3295 16204
rect 3237 16195 3295 16201
rect 2608 16164 2636 16195
rect 3326 16192 3332 16204
rect 3384 16192 3390 16244
rect 3789 16235 3847 16241
rect 3789 16201 3801 16235
rect 3835 16232 3847 16235
rect 4246 16232 4252 16244
rect 3835 16204 4252 16232
rect 3835 16201 3847 16204
rect 3789 16195 3847 16201
rect 4246 16192 4252 16204
rect 4304 16192 4310 16244
rect 5166 16192 5172 16244
rect 5224 16232 5230 16244
rect 5445 16235 5503 16241
rect 5445 16232 5457 16235
rect 5224 16204 5457 16232
rect 5224 16192 5230 16204
rect 5445 16201 5457 16204
rect 5491 16201 5503 16235
rect 5445 16195 5503 16201
rect 5810 16192 5816 16244
rect 5868 16232 5874 16244
rect 5997 16235 6055 16241
rect 5997 16232 6009 16235
rect 5868 16204 6009 16232
rect 5868 16192 5874 16204
rect 5997 16201 6009 16204
rect 6043 16201 6055 16235
rect 5997 16195 6055 16201
rect 6454 16192 6460 16244
rect 6512 16232 6518 16244
rect 6733 16235 6791 16241
rect 6733 16232 6745 16235
rect 6512 16204 6745 16232
rect 6512 16192 6518 16204
rect 6733 16201 6745 16204
rect 6779 16201 6791 16235
rect 6733 16195 6791 16201
rect 7193 16235 7251 16241
rect 7193 16201 7205 16235
rect 7239 16201 7251 16235
rect 7558 16232 7564 16244
rect 7519 16204 7564 16232
rect 7193 16195 7251 16201
rect 4062 16164 4068 16176
rect 2056 16136 2636 16164
rect 2792 16136 4068 16164
rect 1673 16099 1731 16105
rect 1673 16065 1685 16099
rect 1719 16096 1731 16099
rect 1762 16096 1768 16108
rect 1719 16068 1768 16096
rect 1719 16065 1731 16068
rect 1673 16059 1731 16065
rect 1762 16056 1768 16068
rect 1820 16056 1826 16108
rect 2056 16105 2084 16136
rect 2041 16099 2099 16105
rect 2041 16065 2053 16099
rect 2087 16065 2099 16099
rect 2041 16059 2099 16065
rect 2130 16056 2136 16108
rect 2188 16096 2194 16108
rect 2792 16105 2820 16136
rect 4062 16124 4068 16136
rect 4120 16124 4126 16176
rect 4614 16124 4620 16176
rect 4672 16164 4678 16176
rect 5721 16167 5779 16173
rect 4672 16136 5304 16164
rect 4672 16124 4678 16136
rect 2777 16099 2835 16105
rect 2188 16068 2233 16096
rect 2188 16056 2194 16068
rect 2777 16065 2789 16099
rect 2823 16065 2835 16099
rect 2777 16059 2835 16065
rect 3053 16099 3111 16105
rect 3053 16065 3065 16099
rect 3099 16096 3111 16099
rect 3234 16096 3240 16108
rect 3099 16068 3240 16096
rect 3099 16065 3111 16068
rect 3053 16059 3111 16065
rect 3234 16056 3240 16068
rect 3292 16056 3298 16108
rect 3513 16099 3571 16105
rect 3513 16065 3525 16099
rect 3559 16065 3571 16099
rect 3513 16059 3571 16065
rect 658 15988 664 16040
rect 716 16028 722 16040
rect 2866 16028 2872 16040
rect 716 16000 2872 16028
rect 716 15988 722 16000
rect 2866 15988 2872 16000
rect 2924 15988 2930 16040
rect 3528 16028 3556 16059
rect 3602 16056 3608 16108
rect 3660 16096 3666 16108
rect 3660 16068 3705 16096
rect 3660 16056 3666 16068
rect 4522 16056 4528 16108
rect 4580 16096 4586 16108
rect 5276 16105 5304 16136
rect 5721 16133 5733 16167
rect 5767 16164 5779 16167
rect 7098 16164 7104 16176
rect 5767 16136 7104 16164
rect 5767 16133 5779 16136
rect 5721 16127 5779 16133
rect 4994 16099 5052 16105
rect 4994 16096 5006 16099
rect 4580 16068 5006 16096
rect 4580 16056 4586 16068
rect 4994 16065 5006 16068
rect 5040 16065 5052 16099
rect 4994 16059 5052 16065
rect 5261 16099 5319 16105
rect 5261 16065 5273 16099
rect 5307 16065 5319 16099
rect 5626 16096 5632 16108
rect 5587 16068 5632 16096
rect 5261 16059 5319 16065
rect 5626 16056 5632 16068
rect 5684 16056 5690 16108
rect 6564 16105 6592 16136
rect 7098 16124 7104 16136
rect 7156 16124 7162 16176
rect 6181 16099 6239 16105
rect 6181 16065 6193 16099
rect 6227 16096 6239 16099
rect 6549 16099 6607 16105
rect 6227 16068 6408 16096
rect 6227 16065 6239 16068
rect 6181 16059 6239 16065
rect 3694 16028 3700 16040
rect 3528 16000 3700 16028
rect 3694 15988 3700 16000
rect 3752 15988 3758 16040
rect 3329 15963 3387 15969
rect 3329 15929 3341 15963
rect 3375 15960 3387 15963
rect 3418 15960 3424 15972
rect 3375 15932 3424 15960
rect 3375 15929 3387 15932
rect 3329 15923 3387 15929
rect 3418 15920 3424 15932
rect 3476 15920 3482 15972
rect 6380 15969 6408 16068
rect 6549 16065 6561 16099
rect 6595 16065 6607 16099
rect 6549 16059 6607 16065
rect 6917 16099 6975 16105
rect 6917 16065 6929 16099
rect 6963 16096 6975 16099
rect 7208 16096 7236 16195
rect 7558 16192 7564 16204
rect 7616 16192 7622 16244
rect 7650 16192 7656 16244
rect 7708 16232 7714 16244
rect 8021 16235 8079 16241
rect 8021 16232 8033 16235
rect 7708 16204 8033 16232
rect 7708 16192 7714 16204
rect 8021 16201 8033 16204
rect 8067 16201 8079 16235
rect 8021 16195 8079 16201
rect 8294 16192 8300 16244
rect 8352 16232 8358 16244
rect 8481 16235 8539 16241
rect 8481 16232 8493 16235
rect 8352 16204 8493 16232
rect 8352 16192 8358 16204
rect 8481 16201 8493 16204
rect 8527 16201 8539 16235
rect 8481 16195 8539 16201
rect 8570 16192 8576 16244
rect 8628 16232 8634 16244
rect 9582 16232 9588 16244
rect 8628 16204 9588 16232
rect 8628 16192 8634 16204
rect 9582 16192 9588 16204
rect 9640 16232 9646 16244
rect 9766 16232 9772 16244
rect 9640 16204 9772 16232
rect 9640 16192 9646 16204
rect 9766 16192 9772 16204
rect 9824 16192 9830 16244
rect 12066 16192 12072 16244
rect 12124 16232 12130 16244
rect 12345 16235 12403 16241
rect 12345 16232 12357 16235
rect 12124 16204 12357 16232
rect 12124 16192 12130 16204
rect 12345 16201 12357 16204
rect 12391 16201 12403 16235
rect 12345 16195 12403 16201
rect 13170 16192 13176 16244
rect 13228 16232 13234 16244
rect 14090 16232 14096 16244
rect 13228 16204 14096 16232
rect 13228 16192 13234 16204
rect 14090 16192 14096 16204
rect 14148 16192 14154 16244
rect 9122 16124 9128 16176
rect 9180 16164 9186 16176
rect 9870 16167 9928 16173
rect 9870 16164 9882 16167
rect 9180 16136 9882 16164
rect 9180 16124 9186 16136
rect 9870 16133 9882 16136
rect 9916 16133 9928 16167
rect 9870 16127 9928 16133
rect 10042 16124 10048 16176
rect 10100 16164 10106 16176
rect 10318 16164 10324 16176
rect 10100 16136 10324 16164
rect 10100 16124 10106 16136
rect 10318 16124 10324 16136
rect 10376 16124 10382 16176
rect 10686 16124 10692 16176
rect 10744 16164 10750 16176
rect 10744 16136 12434 16164
rect 10744 16124 10750 16136
rect 6963 16068 7236 16096
rect 7377 16099 7435 16105
rect 6963 16065 6975 16068
rect 6917 16059 6975 16065
rect 7377 16065 7389 16099
rect 7423 16096 7435 16099
rect 7650 16096 7656 16108
rect 7423 16068 7656 16096
rect 7423 16065 7435 16068
rect 7377 16059 7435 16065
rect 7101 16031 7159 16037
rect 7101 15997 7113 16031
rect 7147 16028 7159 16031
rect 7392 16028 7420 16059
rect 7650 16056 7656 16068
rect 7708 16056 7714 16108
rect 7745 16099 7803 16105
rect 7745 16065 7757 16099
rect 7791 16065 7803 16099
rect 7745 16059 7803 16065
rect 7147 16000 7420 16028
rect 7147 15997 7159 16000
rect 7101 15991 7159 15997
rect 7558 15988 7564 16040
rect 7616 16028 7622 16040
rect 7760 16028 7788 16059
rect 8202 16056 8208 16108
rect 8260 16096 8266 16108
rect 8665 16099 8723 16105
rect 8260 16068 8305 16096
rect 8260 16056 8266 16068
rect 8665 16065 8677 16099
rect 8711 16096 8723 16099
rect 9582 16096 9588 16108
rect 8711 16068 9588 16096
rect 8711 16065 8723 16068
rect 8665 16059 8723 16065
rect 9582 16056 9588 16068
rect 9640 16056 9646 16108
rect 10226 16096 10232 16108
rect 10187 16068 10232 16096
rect 10226 16056 10232 16068
rect 10284 16056 10290 16108
rect 10962 16096 10968 16108
rect 10923 16068 10968 16096
rect 10962 16056 10968 16068
rect 11020 16056 11026 16108
rect 11882 16096 11888 16108
rect 11795 16068 11888 16096
rect 11882 16056 11888 16068
rect 11940 16096 11946 16108
rect 12158 16096 12164 16108
rect 11940 16068 12164 16096
rect 11940 16056 11946 16068
rect 12158 16056 12164 16068
rect 12216 16056 12222 16108
rect 12406 16096 12434 16136
rect 13538 16124 13544 16176
rect 13596 16164 13602 16176
rect 14734 16164 14740 16176
rect 13596 16136 13676 16164
rect 13596 16124 13602 16136
rect 12526 16096 12532 16108
rect 12406 16068 12532 16096
rect 12526 16056 12532 16068
rect 12584 16056 12590 16108
rect 12894 16056 12900 16108
rect 12952 16096 12958 16108
rect 13648 16105 13676 16136
rect 13832 16136 14740 16164
rect 13633 16099 13691 16105
rect 12952 16068 13400 16096
rect 12952 16056 12958 16068
rect 7616 16000 7788 16028
rect 7616 15988 7622 16000
rect 8110 15988 8116 16040
rect 8168 16028 8174 16040
rect 10137 16031 10195 16037
rect 8168 16000 9168 16028
rect 8168 15988 8174 16000
rect 6365 15963 6423 15969
rect 6365 15929 6377 15963
rect 6411 15929 6423 15963
rect 6365 15923 6423 15929
rect 7650 15920 7656 15972
rect 7708 15960 7714 15972
rect 8389 15963 8447 15969
rect 8389 15960 8401 15963
rect 7708 15932 8401 15960
rect 7708 15920 7714 15932
rect 8389 15929 8401 15932
rect 8435 15960 8447 15963
rect 8938 15960 8944 15972
rect 8435 15932 8944 15960
rect 8435 15929 8447 15932
rect 8389 15923 8447 15929
rect 8938 15920 8944 15932
rect 8996 15920 9002 15972
rect 2314 15852 2320 15904
rect 2372 15892 2378 15904
rect 2409 15895 2467 15901
rect 2409 15892 2421 15895
rect 2372 15864 2421 15892
rect 2372 15852 2378 15864
rect 2409 15861 2421 15864
rect 2455 15861 2467 15895
rect 2409 15855 2467 15861
rect 2961 15895 3019 15901
rect 2961 15861 2973 15895
rect 3007 15892 3019 15895
rect 3602 15892 3608 15904
rect 3007 15864 3608 15892
rect 3007 15861 3019 15864
rect 2961 15855 3019 15861
rect 3602 15852 3608 15864
rect 3660 15852 3666 15904
rect 3878 15892 3884 15904
rect 3839 15864 3884 15892
rect 3878 15852 3884 15864
rect 3936 15852 3942 15904
rect 7098 15852 7104 15904
rect 7156 15892 7162 15904
rect 7837 15895 7895 15901
rect 7837 15892 7849 15895
rect 7156 15864 7849 15892
rect 7156 15852 7162 15864
rect 7837 15861 7849 15864
rect 7883 15892 7895 15895
rect 8202 15892 8208 15904
rect 7883 15864 8208 15892
rect 7883 15861 7895 15864
rect 7837 15855 7895 15861
rect 8202 15852 8208 15864
rect 8260 15852 8266 15904
rect 8294 15852 8300 15904
rect 8352 15892 8358 15904
rect 8757 15895 8815 15901
rect 8757 15892 8769 15895
rect 8352 15864 8769 15892
rect 8352 15852 8358 15864
rect 8757 15861 8769 15864
rect 8803 15861 8815 15895
rect 9140 15892 9168 16000
rect 10137 15997 10149 16031
rect 10183 16028 10195 16031
rect 10686 16028 10692 16040
rect 10183 16000 10692 16028
rect 10183 15997 10195 16000
rect 10137 15991 10195 15997
rect 10686 15988 10692 16000
rect 10744 15988 10750 16040
rect 10870 15988 10876 16040
rect 10928 16028 10934 16040
rect 11057 16031 11115 16037
rect 11057 16028 11069 16031
rect 10928 16000 11069 16028
rect 10928 15988 10934 16000
rect 11057 15997 11069 16000
rect 11103 15997 11115 16031
rect 11057 15991 11115 15997
rect 11149 16031 11207 16037
rect 11149 15997 11161 16031
rect 11195 15997 11207 16031
rect 11974 16028 11980 16040
rect 11935 16000 11980 16028
rect 11149 15991 11207 15997
rect 10226 15920 10232 15972
rect 10284 15960 10290 15972
rect 10597 15963 10655 15969
rect 10597 15960 10609 15963
rect 10284 15932 10609 15960
rect 10284 15920 10290 15932
rect 10597 15929 10609 15932
rect 10643 15929 10655 15963
rect 10597 15923 10655 15929
rect 10778 15920 10784 15972
rect 10836 15960 10842 15972
rect 11164 15960 11192 15991
rect 11974 15988 11980 16000
rect 12032 15988 12038 16040
rect 12066 15988 12072 16040
rect 12124 16028 12130 16040
rect 12124 16000 12169 16028
rect 12124 15988 12130 16000
rect 12710 15988 12716 16040
rect 12768 16028 12774 16040
rect 13265 16031 13323 16037
rect 13265 16028 13277 16031
rect 12768 16000 13277 16028
rect 12768 15988 12774 16000
rect 13265 15997 13277 16000
rect 13311 15997 13323 16031
rect 13265 15991 13323 15997
rect 10836 15932 11192 15960
rect 10836 15920 10842 15932
rect 11330 15920 11336 15972
rect 11388 15960 11394 15972
rect 12894 15960 12900 15972
rect 11388 15932 12900 15960
rect 11388 15920 11394 15932
rect 12894 15920 12900 15932
rect 12952 15920 12958 15972
rect 13372 15960 13400 16068
rect 13633 16065 13645 16099
rect 13679 16065 13691 16099
rect 13633 16059 13691 16065
rect 13541 16031 13599 16037
rect 13541 15997 13553 16031
rect 13587 16028 13599 16031
rect 13832 16028 13860 16136
rect 14734 16124 14740 16136
rect 14792 16164 14798 16176
rect 15746 16164 15752 16176
rect 14792 16136 15752 16164
rect 14792 16124 14798 16136
rect 15746 16124 15752 16136
rect 15804 16124 15810 16176
rect 14458 16056 14464 16108
rect 14516 16096 14522 16108
rect 14553 16099 14611 16105
rect 14553 16096 14565 16099
rect 14516 16068 14565 16096
rect 14516 16056 14522 16068
rect 14553 16065 14565 16068
rect 14599 16065 14611 16099
rect 14553 16059 14611 16065
rect 15378 16056 15384 16108
rect 15436 16096 15442 16108
rect 15473 16099 15531 16105
rect 15473 16096 15485 16099
rect 15436 16068 15485 16096
rect 15436 16056 15442 16068
rect 15473 16065 15485 16068
rect 15519 16065 15531 16099
rect 15473 16059 15531 16065
rect 13587 16000 13860 16028
rect 13909 16031 13967 16037
rect 13587 15997 13599 16000
rect 13541 15991 13599 15997
rect 13909 15997 13921 16031
rect 13955 16028 13967 16031
rect 13998 16028 14004 16040
rect 13955 16000 14004 16028
rect 13955 15997 13967 16000
rect 13909 15991 13967 15997
rect 13998 15988 14004 16000
rect 14056 15988 14062 16040
rect 13630 15960 13636 15972
rect 13372 15932 13636 15960
rect 13630 15920 13636 15932
rect 13688 15920 13694 15972
rect 10410 15892 10416 15904
rect 9140 15864 10416 15892
rect 8757 15855 8815 15861
rect 10410 15852 10416 15864
rect 10468 15852 10474 15904
rect 11422 15852 11428 15904
rect 11480 15892 11486 15904
rect 11517 15895 11575 15901
rect 11517 15892 11529 15895
rect 11480 15864 11529 15892
rect 11480 15852 11486 15864
rect 11517 15861 11529 15864
rect 11563 15861 11575 15895
rect 11517 15855 11575 15861
rect 13262 15852 13268 15904
rect 13320 15892 13326 15904
rect 14783 15895 14841 15901
rect 14783 15892 14795 15895
rect 13320 15864 14795 15892
rect 13320 15852 13326 15864
rect 14783 15861 14795 15864
rect 14829 15861 14841 15895
rect 14783 15855 14841 15861
rect 15286 15852 15292 15904
rect 15344 15892 15350 15904
rect 15657 15895 15715 15901
rect 15657 15892 15669 15895
rect 15344 15864 15669 15892
rect 15344 15852 15350 15864
rect 15657 15861 15669 15864
rect 15703 15861 15715 15895
rect 15657 15855 15715 15861
rect 1104 15802 16008 15824
rect 1104 15750 2824 15802
rect 2876 15750 2888 15802
rect 2940 15750 2952 15802
rect 3004 15750 3016 15802
rect 3068 15750 3080 15802
rect 3132 15750 6572 15802
rect 6624 15750 6636 15802
rect 6688 15750 6700 15802
rect 6752 15750 6764 15802
rect 6816 15750 6828 15802
rect 6880 15750 10320 15802
rect 10372 15750 10384 15802
rect 10436 15750 10448 15802
rect 10500 15750 10512 15802
rect 10564 15750 10576 15802
rect 10628 15750 14068 15802
rect 14120 15750 14132 15802
rect 14184 15750 14196 15802
rect 14248 15750 14260 15802
rect 14312 15750 14324 15802
rect 14376 15750 16008 15802
rect 1104 15728 16008 15750
rect 5258 15688 5264 15700
rect 1964 15660 5264 15688
rect 1765 15623 1823 15629
rect 1765 15589 1777 15623
rect 1811 15589 1823 15623
rect 1765 15583 1823 15589
rect 1673 15487 1731 15493
rect 1673 15453 1685 15487
rect 1719 15484 1731 15487
rect 1780 15484 1808 15583
rect 1964 15493 1992 15660
rect 5258 15648 5264 15660
rect 5316 15648 5322 15700
rect 7374 15688 7380 15700
rect 7287 15660 7380 15688
rect 7374 15648 7380 15660
rect 7432 15688 7438 15700
rect 10962 15688 10968 15700
rect 7432 15660 10732 15688
rect 10923 15660 10968 15688
rect 7432 15648 7438 15660
rect 7285 15623 7343 15629
rect 7285 15589 7297 15623
rect 7331 15620 7343 15623
rect 7650 15620 7656 15632
rect 7331 15592 7656 15620
rect 7331 15589 7343 15592
rect 7285 15583 7343 15589
rect 7650 15580 7656 15592
rect 7708 15580 7714 15632
rect 8754 15580 8760 15632
rect 8812 15620 8818 15632
rect 9030 15620 9036 15632
rect 8812 15592 9036 15620
rect 8812 15580 8818 15592
rect 9030 15580 9036 15592
rect 9088 15580 9094 15632
rect 9214 15580 9220 15632
rect 9272 15620 9278 15632
rect 9309 15623 9367 15629
rect 9309 15620 9321 15623
rect 9272 15592 9321 15620
rect 9272 15580 9278 15592
rect 9309 15589 9321 15592
rect 9355 15589 9367 15623
rect 10704 15620 10732 15660
rect 10962 15648 10968 15660
rect 11020 15648 11026 15700
rect 12526 15648 12532 15700
rect 12584 15688 12590 15700
rect 13725 15691 13783 15697
rect 13725 15688 13737 15691
rect 12584 15660 13737 15688
rect 12584 15648 12590 15660
rect 13725 15657 13737 15660
rect 13771 15657 13783 15691
rect 13725 15651 13783 15657
rect 13906 15648 13912 15700
rect 13964 15688 13970 15700
rect 14185 15691 14243 15697
rect 14185 15688 14197 15691
rect 13964 15660 14197 15688
rect 13964 15648 13970 15660
rect 14185 15657 14197 15660
rect 14231 15657 14243 15691
rect 14185 15651 14243 15657
rect 11330 15620 11336 15632
rect 10704 15592 11336 15620
rect 9309 15583 9367 15589
rect 11330 15580 11336 15592
rect 11388 15580 11394 15632
rect 11606 15580 11612 15632
rect 11664 15620 11670 15632
rect 13078 15620 13084 15632
rect 11664 15592 13084 15620
rect 11664 15580 11670 15592
rect 13078 15580 13084 15592
rect 13136 15580 13142 15632
rect 13446 15620 13452 15632
rect 13407 15592 13452 15620
rect 13446 15580 13452 15592
rect 13504 15580 13510 15632
rect 14458 15620 14464 15632
rect 14419 15592 14464 15620
rect 14458 15580 14464 15592
rect 14516 15580 14522 15632
rect 14642 15580 14648 15632
rect 14700 15620 14706 15632
rect 14700 15592 14780 15620
rect 14700 15580 14706 15592
rect 3970 15552 3976 15564
rect 3528 15524 3976 15552
rect 1719 15456 1808 15484
rect 1949 15487 2007 15493
rect 1719 15453 1731 15456
rect 1673 15447 1731 15453
rect 1949 15453 1961 15487
rect 1995 15453 2007 15487
rect 1949 15447 2007 15453
rect 2133 15487 2191 15493
rect 2133 15453 2145 15487
rect 2179 15484 2191 15487
rect 3528 15484 3556 15524
rect 3970 15512 3976 15524
rect 4028 15512 4034 15564
rect 11422 15552 11428 15564
rect 8680 15524 9260 15552
rect 11383 15524 11428 15552
rect 2179 15456 3556 15484
rect 3605 15487 3663 15493
rect 2179 15453 2191 15456
rect 2133 15447 2191 15453
rect 3160 15428 3188 15456
rect 3605 15453 3617 15487
rect 3651 15453 3663 15487
rect 3605 15447 3663 15453
rect 2314 15376 2320 15428
rect 2372 15416 2378 15428
rect 2774 15416 2780 15428
rect 2372 15388 2780 15416
rect 2372 15376 2378 15388
rect 2774 15376 2780 15388
rect 2832 15376 2838 15428
rect 3142 15376 3148 15428
rect 3200 15376 3206 15428
rect 3360 15419 3418 15425
rect 3360 15385 3372 15419
rect 3406 15416 3418 15419
rect 3510 15416 3516 15428
rect 3406 15388 3516 15416
rect 3406 15385 3418 15388
rect 3360 15379 3418 15385
rect 3510 15376 3516 15388
rect 3568 15376 3574 15428
rect 1486 15348 1492 15360
rect 1447 15320 1492 15348
rect 1486 15308 1492 15320
rect 1544 15308 1550 15360
rect 2222 15348 2228 15360
rect 2183 15320 2228 15348
rect 2222 15308 2228 15320
rect 2280 15308 2286 15360
rect 2792 15348 2820 15376
rect 3620 15348 3648 15447
rect 4614 15444 4620 15496
rect 4672 15484 4678 15496
rect 5261 15487 5319 15493
rect 5261 15484 5273 15487
rect 4672 15456 5273 15484
rect 4672 15444 4678 15456
rect 5261 15453 5273 15456
rect 5307 15484 5319 15487
rect 5445 15487 5503 15493
rect 5445 15484 5457 15487
rect 5307 15456 5457 15484
rect 5307 15453 5319 15456
rect 5261 15447 5319 15453
rect 5445 15453 5457 15456
rect 5491 15453 5503 15487
rect 5445 15447 5503 15453
rect 7466 15444 7472 15496
rect 7524 15484 7530 15496
rect 8680 15484 8708 15524
rect 7524 15456 8708 15484
rect 8757 15487 8815 15493
rect 7524 15444 7530 15456
rect 8757 15453 8769 15487
rect 8803 15484 8815 15487
rect 8938 15484 8944 15496
rect 8803 15456 8944 15484
rect 8803 15453 8815 15456
rect 8757 15447 8815 15453
rect 8938 15444 8944 15456
rect 8996 15484 9002 15496
rect 9125 15487 9183 15493
rect 9125 15484 9137 15487
rect 8996 15456 9137 15484
rect 8996 15444 9002 15456
rect 9125 15453 9137 15456
rect 9171 15453 9183 15487
rect 9232 15484 9260 15524
rect 11422 15512 11428 15524
rect 11480 15512 11486 15564
rect 11514 15512 11520 15564
rect 11572 15552 11578 15564
rect 11572 15524 11617 15552
rect 11572 15512 11578 15524
rect 12066 15512 12072 15564
rect 12124 15552 12130 15564
rect 12345 15555 12403 15561
rect 12345 15552 12357 15555
rect 12124 15524 12357 15552
rect 12124 15512 12130 15524
rect 12345 15521 12357 15524
rect 12391 15521 12403 15555
rect 12345 15515 12403 15521
rect 12894 15512 12900 15564
rect 12952 15552 12958 15564
rect 13173 15555 13231 15561
rect 13173 15552 13185 15555
rect 12952 15524 13185 15552
rect 12952 15512 12958 15524
rect 13173 15521 13185 15524
rect 13219 15521 13231 15555
rect 13173 15515 13231 15521
rect 13906 15512 13912 15564
rect 13964 15552 13970 15564
rect 14752 15561 14780 15592
rect 14737 15555 14795 15561
rect 14737 15552 14749 15555
rect 13964 15524 14749 15552
rect 13964 15512 13970 15524
rect 14737 15521 14749 15524
rect 14783 15521 14795 15555
rect 14737 15515 14795 15521
rect 10422 15487 10480 15493
rect 10422 15484 10434 15487
rect 9232 15456 10434 15484
rect 9125 15447 9183 15453
rect 10422 15453 10434 15456
rect 10468 15453 10480 15487
rect 10422 15447 10480 15453
rect 10594 15444 10600 15496
rect 10652 15484 10658 15496
rect 10689 15487 10747 15493
rect 10689 15484 10701 15487
rect 10652 15456 10701 15484
rect 10652 15444 10658 15456
rect 10689 15453 10701 15456
rect 10735 15453 10747 15487
rect 10689 15447 10747 15453
rect 12158 15444 12164 15496
rect 12216 15484 12222 15496
rect 12216 15456 12940 15484
rect 12216 15444 12222 15456
rect 4994 15419 5052 15425
rect 4994 15385 5006 15419
rect 5040 15416 5052 15419
rect 5040 15388 5120 15416
rect 5040 15385 5052 15388
rect 4994 15379 5052 15385
rect 3878 15348 3884 15360
rect 2792 15320 3648 15348
rect 3839 15320 3884 15348
rect 3878 15308 3884 15320
rect 3936 15308 3942 15360
rect 5092 15348 5120 15388
rect 5166 15376 5172 15428
rect 5224 15416 5230 15428
rect 5690 15419 5748 15425
rect 5690 15416 5702 15419
rect 5224 15388 5702 15416
rect 5224 15376 5230 15388
rect 5690 15385 5702 15388
rect 5736 15385 5748 15419
rect 5690 15379 5748 15385
rect 6914 15376 6920 15428
rect 6972 15416 6978 15428
rect 8110 15416 8116 15428
rect 6972 15388 8116 15416
rect 6972 15376 6978 15388
rect 8110 15376 8116 15388
rect 8168 15376 8174 15428
rect 8512 15419 8570 15425
rect 8512 15385 8524 15419
rect 8558 15416 8570 15419
rect 8662 15416 8668 15428
rect 8558 15388 8668 15416
rect 8558 15385 8570 15388
rect 8512 15379 8570 15385
rect 8662 15376 8668 15388
rect 8720 15376 8726 15428
rect 9033 15419 9091 15425
rect 9033 15385 9045 15419
rect 9079 15416 9091 15419
rect 9950 15416 9956 15428
rect 9079 15388 9956 15416
rect 9079 15385 9091 15388
rect 9033 15379 9091 15385
rect 9950 15376 9956 15388
rect 10008 15376 10014 15428
rect 10962 15376 10968 15428
rect 11020 15416 11026 15428
rect 12802 15416 12808 15428
rect 11020 15388 12808 15416
rect 11020 15376 11026 15388
rect 12802 15376 12808 15388
rect 12860 15376 12866 15428
rect 12912 15416 12940 15456
rect 13262 15444 13268 15496
rect 13320 15484 13326 15496
rect 13633 15487 13691 15493
rect 13633 15484 13645 15487
rect 13320 15456 13645 15484
rect 13320 15444 13326 15456
rect 13633 15453 13645 15456
rect 13679 15453 13691 15487
rect 13633 15447 13691 15453
rect 14369 15487 14427 15493
rect 14369 15453 14381 15487
rect 14415 15453 14427 15487
rect 14642 15484 14648 15496
rect 14603 15456 14648 15484
rect 14369 15447 14427 15453
rect 12912 15388 13768 15416
rect 5902 15348 5908 15360
rect 5092 15320 5908 15348
rect 5902 15308 5908 15320
rect 5960 15308 5966 15360
rect 6822 15348 6828 15360
rect 6783 15320 6828 15348
rect 6822 15308 6828 15320
rect 6880 15308 6886 15360
rect 7101 15351 7159 15357
rect 7101 15317 7113 15351
rect 7147 15348 7159 15351
rect 7834 15348 7840 15360
rect 7147 15320 7840 15348
rect 7147 15317 7159 15320
rect 7101 15311 7159 15317
rect 7834 15308 7840 15320
rect 7892 15348 7898 15360
rect 8846 15348 8852 15360
rect 7892 15320 8852 15348
rect 7892 15308 7898 15320
rect 8846 15308 8852 15320
rect 8904 15308 8910 15360
rect 9766 15308 9772 15360
rect 9824 15348 9830 15360
rect 10781 15351 10839 15357
rect 10781 15348 10793 15351
rect 9824 15320 10793 15348
rect 9824 15308 9830 15320
rect 10781 15317 10793 15320
rect 10827 15317 10839 15351
rect 11330 15348 11336 15360
rect 11291 15320 11336 15348
rect 10781 15311 10839 15317
rect 11330 15308 11336 15320
rect 11388 15308 11394 15360
rect 11790 15348 11796 15360
rect 11751 15320 11796 15348
rect 11790 15308 11796 15320
rect 11848 15308 11854 15360
rect 11974 15308 11980 15360
rect 12032 15348 12038 15360
rect 12161 15351 12219 15357
rect 12161 15348 12173 15351
rect 12032 15320 12173 15348
rect 12032 15308 12038 15320
rect 12161 15317 12173 15320
rect 12207 15317 12219 15351
rect 12161 15311 12219 15317
rect 12253 15351 12311 15357
rect 12253 15317 12265 15351
rect 12299 15348 12311 15351
rect 12621 15351 12679 15357
rect 12621 15348 12633 15351
rect 12299 15320 12633 15348
rect 12299 15317 12311 15320
rect 12253 15311 12311 15317
rect 12621 15317 12633 15320
rect 12667 15317 12679 15351
rect 12986 15348 12992 15360
rect 12947 15320 12992 15348
rect 12621 15311 12679 15317
rect 12986 15308 12992 15320
rect 13044 15308 13050 15360
rect 13078 15308 13084 15360
rect 13136 15348 13142 15360
rect 13136 15320 13181 15348
rect 13136 15308 13142 15320
rect 13446 15308 13452 15360
rect 13504 15348 13510 15360
rect 13630 15348 13636 15360
rect 13504 15320 13636 15348
rect 13504 15308 13510 15320
rect 13630 15308 13636 15320
rect 13688 15308 13694 15360
rect 13740 15348 13768 15388
rect 13814 15376 13820 15428
rect 13872 15416 13878 15428
rect 13998 15416 14004 15428
rect 13872 15388 14004 15416
rect 13872 15376 13878 15388
rect 13998 15376 14004 15388
rect 14056 15376 14062 15428
rect 14384 15416 14412 15447
rect 14642 15444 14648 15456
rect 14700 15444 14706 15496
rect 15013 15487 15071 15493
rect 15013 15453 15025 15487
rect 15059 15484 15071 15487
rect 16206 15484 16212 15496
rect 15059 15456 16212 15484
rect 15059 15453 15071 15456
rect 15013 15447 15071 15453
rect 16206 15444 16212 15456
rect 16264 15444 16270 15496
rect 15930 15416 15936 15428
rect 14384 15388 15936 15416
rect 15930 15376 15936 15388
rect 15988 15376 15994 15428
rect 16666 15348 16672 15360
rect 13740 15320 16672 15348
rect 16666 15308 16672 15320
rect 16724 15308 16730 15360
rect 1104 15258 16008 15280
rect 1104 15206 4698 15258
rect 4750 15206 4762 15258
rect 4814 15206 4826 15258
rect 4878 15206 4890 15258
rect 4942 15206 4954 15258
rect 5006 15206 8446 15258
rect 8498 15206 8510 15258
rect 8562 15206 8574 15258
rect 8626 15206 8638 15258
rect 8690 15206 8702 15258
rect 8754 15206 12194 15258
rect 12246 15206 12258 15258
rect 12310 15206 12322 15258
rect 12374 15206 12386 15258
rect 12438 15206 12450 15258
rect 12502 15206 16008 15258
rect 1104 15184 16008 15206
rect 1765 15147 1823 15153
rect 1765 15113 1777 15147
rect 1811 15144 1823 15147
rect 2130 15144 2136 15156
rect 1811 15116 2136 15144
rect 1811 15113 1823 15116
rect 1765 15107 1823 15113
rect 2130 15104 2136 15116
rect 2188 15104 2194 15156
rect 2498 15144 2504 15156
rect 2459 15116 2504 15144
rect 2498 15104 2504 15116
rect 2556 15104 2562 15156
rect 7009 15147 7067 15153
rect 7009 15113 7021 15147
rect 7055 15144 7067 15147
rect 7650 15144 7656 15156
rect 7055 15116 7656 15144
rect 7055 15113 7067 15116
rect 7009 15107 7067 15113
rect 4154 15036 4160 15088
rect 4212 15076 4218 15088
rect 4798 15076 4804 15088
rect 4212 15048 4804 15076
rect 4212 15036 4218 15048
rect 4798 15036 4804 15048
rect 4856 15036 4862 15088
rect 2406 15008 2412 15020
rect 2367 14980 2412 15008
rect 2406 14968 2412 14980
rect 2464 14968 2470 15020
rect 2498 14968 2504 15020
rect 2556 15008 2562 15020
rect 2685 15011 2743 15017
rect 2685 15008 2697 15011
rect 2556 14980 2697 15008
rect 2556 14968 2562 14980
rect 2685 14977 2697 14980
rect 2731 14977 2743 15011
rect 2685 14971 2743 14977
rect 2774 14968 2780 15020
rect 2832 15008 2838 15020
rect 3044 15011 3102 15017
rect 2832 14980 2877 15008
rect 2832 14968 2838 14980
rect 3044 14977 3056 15011
rect 3090 15008 3102 15011
rect 4246 15008 4252 15020
rect 3090 14980 4252 15008
rect 3090 14977 3102 14980
rect 3044 14971 3102 14977
rect 4246 14968 4252 14980
rect 4304 14968 4310 15020
rect 6086 14968 6092 15020
rect 6144 15008 6150 15020
rect 6914 15008 6920 15020
rect 6144 14980 6920 15008
rect 6144 14968 6150 14980
rect 6914 14968 6920 14980
rect 6972 14968 6978 15020
rect 1394 14900 1400 14952
rect 1452 14940 1458 14952
rect 1489 14943 1547 14949
rect 1489 14940 1501 14943
rect 1452 14912 1501 14940
rect 1452 14900 1458 14912
rect 1489 14909 1501 14912
rect 1535 14909 1547 14943
rect 1670 14940 1676 14952
rect 1631 14912 1676 14940
rect 1489 14903 1547 14909
rect 1670 14900 1676 14912
rect 1728 14900 1734 14952
rect 4433 14943 4491 14949
rect 4433 14909 4445 14943
rect 4479 14940 4491 14943
rect 4614 14940 4620 14952
rect 4479 14912 4620 14940
rect 4479 14909 4491 14912
rect 4433 14903 4491 14909
rect 4614 14900 4620 14912
rect 4672 14940 4678 14952
rect 5261 14943 5319 14949
rect 5261 14940 5273 14943
rect 4672 14912 5273 14940
rect 4672 14900 4678 14912
rect 5261 14909 5273 14912
rect 5307 14909 5319 14943
rect 7024 14940 7052 15107
rect 7650 15104 7656 15116
rect 7708 15104 7714 15156
rect 8938 15144 8944 15156
rect 8899 15116 8944 15144
rect 8938 15104 8944 15116
rect 8996 15104 9002 15156
rect 9646 15116 10732 15144
rect 7374 15085 7380 15088
rect 7368 15076 7380 15085
rect 7335 15048 7380 15076
rect 7368 15039 7380 15048
rect 7374 15036 7380 15039
rect 7432 15036 7438 15088
rect 7558 15036 7564 15088
rect 7616 15076 7622 15088
rect 9646 15076 9674 15116
rect 7616 15048 9674 15076
rect 7616 15036 7622 15048
rect 10134 15036 10140 15088
rect 10192 15076 10198 15088
rect 10704 15076 10732 15116
rect 10870 15104 10876 15156
rect 10928 15144 10934 15156
rect 11517 15147 11575 15153
rect 11517 15144 11529 15147
rect 10928 15116 11529 15144
rect 10928 15104 10934 15116
rect 11517 15113 11529 15116
rect 11563 15113 11575 15147
rect 11517 15107 11575 15113
rect 11882 15104 11888 15156
rect 11940 15144 11946 15156
rect 12158 15144 12164 15156
rect 11940 15116 12164 15144
rect 11940 15104 11946 15116
rect 12158 15104 12164 15116
rect 12216 15104 12222 15156
rect 12897 15147 12955 15153
rect 12897 15144 12909 15147
rect 12406 15116 12909 15144
rect 11054 15076 11060 15088
rect 10192 15048 10660 15076
rect 10704 15048 11060 15076
rect 10192 15036 10198 15048
rect 9858 14968 9864 15020
rect 9916 15008 9922 15020
rect 10238 15011 10296 15017
rect 10238 15008 10250 15011
rect 9916 14980 10250 15008
rect 9916 14968 9922 14980
rect 10238 14977 10250 14980
rect 10284 14977 10296 15011
rect 10632 15008 10660 15048
rect 11054 15036 11060 15048
rect 11112 15036 11118 15088
rect 12406 15076 12434 15116
rect 12897 15113 12909 15116
rect 12943 15113 12955 15147
rect 13354 15144 13360 15156
rect 13315 15116 13360 15144
rect 12897 15107 12955 15113
rect 13354 15104 13360 15116
rect 13412 15104 13418 15156
rect 13633 15147 13691 15153
rect 13633 15113 13645 15147
rect 13679 15144 13691 15147
rect 14369 15147 14427 15153
rect 13679 15116 14044 15144
rect 13679 15113 13691 15116
rect 13633 15107 13691 15113
rect 11808 15048 12434 15076
rect 12989 15079 13047 15085
rect 10965 15011 11023 15017
rect 10965 15008 10977 15011
rect 10632 14980 10977 15008
rect 10238 14971 10296 14977
rect 10965 14977 10977 14980
rect 11011 14977 11023 15011
rect 10965 14971 11023 14977
rect 7101 14943 7159 14949
rect 7101 14940 7113 14943
rect 5261 14903 5319 14909
rect 6886 14912 7113 14940
rect 1854 14832 1860 14884
rect 1912 14872 1918 14884
rect 2225 14875 2283 14881
rect 2225 14872 2237 14875
rect 1912 14844 2237 14872
rect 1912 14832 1918 14844
rect 2225 14841 2237 14844
rect 2271 14841 2283 14875
rect 2225 14835 2283 14841
rect 4157 14875 4215 14881
rect 4157 14841 4169 14875
rect 4203 14872 4215 14875
rect 5994 14872 6000 14884
rect 4203 14844 6000 14872
rect 4203 14841 4215 14844
rect 4157 14835 4215 14841
rect 5994 14832 6000 14844
rect 6052 14832 6058 14884
rect 2038 14764 2044 14816
rect 2096 14804 2102 14816
rect 2133 14807 2191 14813
rect 2133 14804 2145 14807
rect 2096 14776 2145 14804
rect 2096 14764 2102 14776
rect 2133 14773 2145 14776
rect 2179 14773 2191 14807
rect 2133 14767 2191 14773
rect 3418 14764 3424 14816
rect 3476 14804 3482 14816
rect 4338 14804 4344 14816
rect 3476 14776 4344 14804
rect 3476 14764 3482 14776
rect 4338 14764 4344 14776
rect 4396 14804 4402 14816
rect 4525 14807 4583 14813
rect 4525 14804 4537 14807
rect 4396 14776 4537 14804
rect 4396 14764 4402 14776
rect 4525 14773 4537 14776
rect 4571 14773 4583 14807
rect 4798 14804 4804 14816
rect 4711 14776 4804 14804
rect 4525 14767 4583 14773
rect 4798 14764 4804 14776
rect 4856 14804 4862 14816
rect 5350 14804 5356 14816
rect 4856 14776 5356 14804
rect 4856 14764 4862 14776
rect 5350 14764 5356 14776
rect 5408 14764 5414 14816
rect 5626 14764 5632 14816
rect 5684 14804 5690 14816
rect 5721 14807 5779 14813
rect 5721 14804 5733 14807
rect 5684 14776 5733 14804
rect 5684 14764 5690 14776
rect 5721 14773 5733 14776
rect 5767 14773 5779 14807
rect 5721 14767 5779 14773
rect 6454 14764 6460 14816
rect 6512 14804 6518 14816
rect 6886 14804 6914 14912
rect 7101 14909 7113 14912
rect 7147 14909 7159 14943
rect 7101 14903 7159 14909
rect 8110 14900 8116 14952
rect 8168 14940 8174 14952
rect 9122 14940 9128 14952
rect 8168 14912 9128 14940
rect 8168 14900 8174 14912
rect 9122 14900 9128 14912
rect 9180 14900 9186 14952
rect 10505 14943 10563 14949
rect 10505 14909 10517 14943
rect 10551 14940 10563 14943
rect 10594 14940 10600 14952
rect 10551 14912 10600 14940
rect 10551 14909 10563 14912
rect 10505 14903 10563 14909
rect 10594 14900 10600 14912
rect 10652 14900 10658 14952
rect 10689 14943 10747 14949
rect 10689 14909 10701 14943
rect 10735 14909 10747 14943
rect 10689 14903 10747 14909
rect 10873 14943 10931 14949
rect 10873 14909 10885 14943
rect 10919 14940 10931 14943
rect 11238 14940 11244 14952
rect 10919 14912 11244 14940
rect 10919 14909 10931 14912
rect 10873 14903 10931 14909
rect 8481 14875 8539 14881
rect 8481 14841 8493 14875
rect 8527 14872 8539 14875
rect 9490 14872 9496 14884
rect 8527 14844 9496 14872
rect 8527 14841 8539 14844
rect 8481 14835 8539 14841
rect 9490 14832 9496 14844
rect 9548 14832 9554 14884
rect 10704 14872 10732 14903
rect 11238 14900 11244 14912
rect 11296 14900 11302 14952
rect 10612 14844 10732 14872
rect 11333 14875 11391 14881
rect 9122 14804 9128 14816
rect 6512 14776 6914 14804
rect 9083 14776 9128 14804
rect 6512 14764 6518 14776
rect 9122 14764 9128 14776
rect 9180 14764 9186 14816
rect 10134 14764 10140 14816
rect 10192 14804 10198 14816
rect 10612 14804 10640 14844
rect 11333 14841 11345 14875
rect 11379 14872 11391 14875
rect 11808 14872 11836 15048
rect 12989 15045 13001 15079
rect 13035 15076 13047 15079
rect 13814 15076 13820 15088
rect 13035 15048 13820 15076
rect 13035 15045 13047 15048
rect 12989 15039 13047 15045
rect 13814 15036 13820 15048
rect 13872 15036 13878 15088
rect 14016 15076 14044 15116
rect 14369 15113 14381 15147
rect 14415 15144 14427 15147
rect 15194 15144 15200 15156
rect 14415 15116 15200 15144
rect 14415 15113 14427 15116
rect 14369 15107 14427 15113
rect 15194 15104 15200 15116
rect 15252 15104 15258 15156
rect 14918 15076 14924 15088
rect 14016 15048 14412 15076
rect 11885 15011 11943 15017
rect 11885 14977 11897 15011
rect 11931 15008 11943 15011
rect 13725 15011 13783 15017
rect 11931 14980 12204 15008
rect 11931 14977 11943 14980
rect 11885 14971 11943 14977
rect 11977 14943 12035 14949
rect 11977 14940 11989 14943
rect 11900 14912 11989 14940
rect 11900 14884 11928 14912
rect 11977 14909 11989 14912
rect 12023 14909 12035 14943
rect 11977 14903 12035 14909
rect 12069 14943 12127 14949
rect 12069 14909 12081 14943
rect 12115 14909 12127 14943
rect 12069 14903 12127 14909
rect 11379 14844 11836 14872
rect 11379 14841 11391 14844
rect 11333 14835 11391 14841
rect 11882 14832 11888 14884
rect 11940 14832 11946 14884
rect 12084 14872 12112 14903
rect 11992 14844 12112 14872
rect 10192 14776 10640 14804
rect 10192 14764 10198 14776
rect 11146 14764 11152 14816
rect 11204 14804 11210 14816
rect 11514 14804 11520 14816
rect 11204 14776 11520 14804
rect 11204 14764 11210 14776
rect 11514 14764 11520 14776
rect 11572 14804 11578 14816
rect 11992 14804 12020 14844
rect 11572 14776 12020 14804
rect 11572 14764 11578 14776
rect 12066 14764 12072 14816
rect 12124 14804 12130 14816
rect 12176 14804 12204 14980
rect 13725 14977 13737 15011
rect 13771 15008 13783 15011
rect 13998 15008 14004 15020
rect 13771 14980 14004 15008
rect 13771 14977 13783 14980
rect 13725 14971 13783 14977
rect 13998 14968 14004 14980
rect 14056 14968 14062 15020
rect 12437 14943 12495 14949
rect 12437 14909 12449 14943
rect 12483 14940 12495 14943
rect 12710 14940 12716 14952
rect 12483 14912 12716 14940
rect 12483 14909 12495 14912
rect 12437 14903 12495 14909
rect 12710 14900 12716 14912
rect 12768 14900 12774 14952
rect 13081 14943 13139 14949
rect 13081 14909 13093 14943
rect 13127 14909 13139 14943
rect 13081 14903 13139 14909
rect 12250 14832 12256 14884
rect 12308 14872 12314 14884
rect 13096 14872 13124 14903
rect 13354 14900 13360 14952
rect 13412 14940 13418 14952
rect 14093 14943 14151 14949
rect 14093 14940 14105 14943
rect 13412 14912 14105 14940
rect 13412 14900 13418 14912
rect 14093 14909 14105 14912
rect 14139 14909 14151 14943
rect 14093 14903 14151 14909
rect 14277 14943 14335 14949
rect 14277 14909 14289 14943
rect 14323 14909 14335 14943
rect 14384 14940 14412 15048
rect 14844 15048 14924 15076
rect 14844 15017 14872 15048
rect 14918 15036 14924 15048
rect 14976 15036 14982 15088
rect 14829 15011 14887 15017
rect 14829 14977 14841 15011
rect 14875 14977 14887 15011
rect 15654 15008 15660 15020
rect 14829 14971 14887 14977
rect 14936 14980 15660 15008
rect 14936 14940 14964 14980
rect 15654 14968 15660 14980
rect 15712 14968 15718 15020
rect 14384 14912 14964 14940
rect 14277 14903 14335 14909
rect 12308 14844 13124 14872
rect 14292 14872 14320 14903
rect 15838 14872 15844 14884
rect 14292 14844 15844 14872
rect 12308 14832 12314 14844
rect 15838 14832 15844 14844
rect 15896 14832 15902 14884
rect 12124 14776 12204 14804
rect 12124 14764 12130 14776
rect 12526 14764 12532 14816
rect 12584 14804 12590 14816
rect 12584 14776 12629 14804
rect 12584 14764 12590 14776
rect 12986 14764 12992 14816
rect 13044 14804 13050 14816
rect 13538 14804 13544 14816
rect 13044 14776 13544 14804
rect 13044 14764 13050 14776
rect 13538 14764 13544 14776
rect 13596 14764 13602 14816
rect 14734 14804 14740 14816
rect 14695 14776 14740 14804
rect 14734 14764 14740 14776
rect 14792 14764 14798 14816
rect 14918 14764 14924 14816
rect 14976 14804 14982 14816
rect 15059 14807 15117 14813
rect 15059 14804 15071 14807
rect 14976 14776 15071 14804
rect 14976 14764 14982 14776
rect 15059 14773 15071 14776
rect 15105 14773 15117 14807
rect 15059 14767 15117 14773
rect 1104 14714 16008 14736
rect 1104 14662 2824 14714
rect 2876 14662 2888 14714
rect 2940 14662 2952 14714
rect 3004 14662 3016 14714
rect 3068 14662 3080 14714
rect 3132 14662 6572 14714
rect 6624 14662 6636 14714
rect 6688 14662 6700 14714
rect 6752 14662 6764 14714
rect 6816 14662 6828 14714
rect 6880 14662 10320 14714
rect 10372 14662 10384 14714
rect 10436 14662 10448 14714
rect 10500 14662 10512 14714
rect 10564 14662 10576 14714
rect 10628 14662 14068 14714
rect 14120 14662 14132 14714
rect 14184 14662 14196 14714
rect 14248 14662 14260 14714
rect 14312 14662 14324 14714
rect 14376 14662 16008 14714
rect 1104 14640 16008 14662
rect 1762 14600 1768 14612
rect 1723 14572 1768 14600
rect 1762 14560 1768 14572
rect 1820 14560 1826 14612
rect 3421 14603 3479 14609
rect 3421 14600 3433 14603
rect 2746 14572 3433 14600
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14396 1731 14399
rect 1762 14396 1768 14408
rect 1719 14368 1768 14396
rect 1719 14365 1731 14368
rect 1673 14359 1731 14365
rect 1762 14356 1768 14368
rect 1820 14356 1826 14408
rect 1946 14396 1952 14408
rect 1907 14368 1952 14396
rect 1946 14356 1952 14368
rect 2004 14356 2010 14408
rect 2222 14396 2228 14408
rect 2135 14368 2228 14396
rect 2222 14356 2228 14368
rect 2280 14396 2286 14408
rect 2746 14396 2774 14572
rect 3421 14569 3433 14572
rect 3467 14600 3479 14603
rect 9582 14600 9588 14612
rect 3467 14572 9588 14600
rect 3467 14569 3479 14572
rect 3421 14563 3479 14569
rect 9582 14560 9588 14572
rect 9640 14560 9646 14612
rect 10413 14603 10471 14609
rect 10413 14569 10425 14603
rect 10459 14600 10471 14603
rect 10962 14600 10968 14612
rect 10459 14572 10968 14600
rect 10459 14569 10471 14572
rect 10413 14563 10471 14569
rect 10962 14560 10968 14572
rect 11020 14560 11026 14612
rect 11330 14560 11336 14612
rect 11388 14600 11394 14612
rect 12345 14603 12403 14609
rect 12345 14600 12357 14603
rect 11388 14572 12357 14600
rect 11388 14560 11394 14572
rect 12345 14569 12357 14572
rect 12391 14569 12403 14603
rect 13173 14603 13231 14609
rect 12345 14563 12403 14569
rect 12544 14572 13124 14600
rect 3786 14492 3792 14544
rect 3844 14532 3850 14544
rect 3973 14535 4031 14541
rect 3973 14532 3985 14535
rect 3844 14504 3985 14532
rect 3844 14492 3850 14504
rect 3973 14501 3985 14504
rect 4019 14501 4031 14535
rect 3973 14495 4031 14501
rect 11514 14492 11520 14544
rect 11572 14532 11578 14544
rect 12158 14532 12164 14544
rect 11572 14504 12164 14532
rect 11572 14492 11578 14504
rect 12158 14492 12164 14504
rect 12216 14492 12222 14544
rect 2866 14424 2872 14476
rect 2924 14464 2930 14476
rect 3142 14464 3148 14476
rect 2924 14436 3148 14464
rect 2924 14424 2930 14436
rect 3142 14424 3148 14436
rect 3200 14464 3206 14476
rect 3881 14467 3939 14473
rect 3881 14464 3893 14467
rect 3200 14436 3893 14464
rect 3200 14424 3206 14436
rect 3881 14433 3893 14436
rect 3927 14464 3939 14467
rect 4154 14464 4160 14476
rect 3927 14436 4160 14464
rect 3927 14433 3939 14436
rect 3881 14427 3939 14433
rect 4154 14424 4160 14436
rect 4212 14464 4218 14476
rect 4614 14464 4620 14476
rect 4212 14436 4620 14464
rect 4212 14424 4218 14436
rect 4614 14424 4620 14436
rect 4672 14464 4678 14476
rect 4893 14467 4951 14473
rect 4893 14464 4905 14467
rect 4672 14436 4905 14464
rect 4672 14424 4678 14436
rect 4893 14433 4905 14436
rect 4939 14464 4951 14467
rect 5442 14464 5448 14476
rect 4939 14436 5448 14464
rect 4939 14433 4951 14436
rect 4893 14427 4951 14433
rect 5442 14424 5448 14436
rect 5500 14424 5506 14476
rect 10781 14467 10839 14473
rect 10781 14433 10793 14467
rect 10827 14433 10839 14467
rect 10781 14427 10839 14433
rect 11609 14467 11667 14473
rect 11609 14433 11621 14467
rect 11655 14464 11667 14467
rect 12544 14464 12572 14572
rect 12618 14492 12624 14544
rect 12676 14532 12682 14544
rect 13096 14532 13124 14572
rect 13173 14569 13185 14603
rect 13219 14600 13231 14603
rect 13538 14600 13544 14612
rect 13219 14572 13544 14600
rect 13219 14569 13231 14572
rect 13173 14563 13231 14569
rect 13538 14560 13544 14572
rect 13596 14560 13602 14612
rect 13630 14560 13636 14612
rect 13688 14600 13694 14612
rect 14093 14603 14151 14609
rect 14093 14600 14105 14603
rect 13688 14572 14105 14600
rect 13688 14560 13694 14572
rect 14093 14569 14105 14572
rect 14139 14569 14151 14603
rect 14093 14563 14151 14569
rect 14369 14603 14427 14609
rect 14369 14569 14381 14603
rect 14415 14600 14427 14603
rect 14642 14600 14648 14612
rect 14415 14572 14648 14600
rect 14415 14569 14427 14572
rect 14369 14563 14427 14569
rect 14642 14560 14648 14572
rect 14700 14560 14706 14612
rect 12676 14504 12940 14532
rect 13096 14504 13860 14532
rect 12676 14492 12682 14504
rect 12802 14464 12808 14476
rect 11655 14436 12572 14464
rect 12763 14436 12808 14464
rect 11655 14433 11667 14436
rect 11609 14427 11667 14433
rect 6454 14396 6460 14408
rect 2280 14368 2774 14396
rect 6415 14368 6460 14396
rect 2280 14356 2286 14368
rect 6454 14356 6460 14368
rect 6512 14396 6518 14408
rect 7929 14399 7987 14405
rect 7929 14396 7941 14399
rect 6512 14368 7941 14396
rect 6512 14356 6518 14368
rect 7929 14365 7941 14368
rect 7975 14365 7987 14399
rect 7929 14359 7987 14365
rect 8202 14356 8208 14408
rect 8260 14396 8266 14408
rect 9950 14396 9956 14408
rect 8260 14368 9956 14396
rect 8260 14356 8266 14368
rect 9950 14356 9956 14368
rect 10008 14396 10014 14408
rect 10796 14396 10824 14427
rect 10962 14396 10968 14408
rect 10008 14368 10824 14396
rect 10923 14368 10968 14396
rect 10008 14356 10014 14368
rect 10962 14356 10968 14368
rect 11020 14356 11026 14408
rect 2774 14288 2780 14340
rect 2832 14328 2838 14340
rect 6086 14328 6092 14340
rect 2832 14300 6092 14328
rect 2832 14288 2838 14300
rect 6086 14288 6092 14300
rect 6144 14288 6150 14340
rect 6212 14331 6270 14337
rect 6212 14297 6224 14331
rect 6258 14328 6270 14331
rect 6362 14328 6368 14340
rect 6258 14300 6368 14328
rect 6258 14297 6270 14300
rect 6212 14291 6270 14297
rect 6362 14288 6368 14300
rect 6420 14328 6426 14340
rect 6638 14328 6644 14340
rect 6420 14300 6644 14328
rect 6420 14288 6426 14300
rect 6638 14288 6644 14300
rect 6696 14288 6702 14340
rect 7650 14288 7656 14340
rect 7708 14337 7714 14340
rect 7708 14328 7720 14337
rect 8294 14328 8300 14340
rect 7708 14300 8300 14328
rect 7708 14291 7720 14300
rect 7708 14288 7714 14291
rect 8294 14288 8300 14300
rect 8352 14288 8358 14340
rect 9030 14288 9036 14340
rect 9088 14328 9094 14340
rect 11624 14328 11652 14427
rect 12802 14424 12808 14436
rect 12860 14424 12866 14476
rect 12912 14473 12940 14504
rect 12897 14467 12955 14473
rect 12897 14433 12909 14467
rect 12943 14433 12955 14467
rect 12897 14427 12955 14433
rect 12986 14424 12992 14476
rect 13044 14464 13050 14476
rect 13170 14464 13176 14476
rect 13044 14436 13176 14464
rect 13044 14424 13050 14436
rect 13170 14424 13176 14436
rect 13228 14424 13234 14476
rect 13832 14473 13860 14504
rect 13817 14467 13875 14473
rect 13817 14433 13829 14467
rect 13863 14464 13875 14467
rect 13998 14464 14004 14476
rect 13863 14436 14004 14464
rect 13863 14433 13875 14436
rect 13817 14427 13875 14433
rect 13998 14424 14004 14436
rect 14056 14424 14062 14476
rect 15654 14464 15660 14476
rect 15567 14436 15660 14464
rect 15654 14424 15660 14436
rect 15712 14464 15718 14476
rect 16850 14464 16856 14476
rect 15712 14436 16856 14464
rect 15712 14424 15718 14436
rect 16850 14424 16856 14436
rect 16908 14424 16914 14476
rect 11698 14356 11704 14408
rect 11756 14396 11762 14408
rect 11793 14399 11851 14405
rect 11793 14396 11805 14399
rect 11756 14368 11805 14396
rect 11756 14356 11762 14368
rect 11793 14365 11805 14368
rect 11839 14365 11851 14399
rect 11793 14359 11851 14365
rect 11885 14399 11943 14405
rect 11885 14365 11897 14399
rect 11931 14396 11943 14399
rect 14461 14399 14519 14405
rect 14461 14396 14473 14399
rect 11931 14368 14473 14396
rect 11931 14365 11943 14368
rect 11885 14359 11943 14365
rect 14461 14365 14473 14368
rect 14507 14365 14519 14399
rect 15378 14396 15384 14408
rect 15291 14368 15384 14396
rect 14461 14359 14519 14365
rect 15378 14356 15384 14368
rect 15436 14396 15442 14408
rect 16758 14396 16764 14408
rect 15436 14368 16764 14396
rect 15436 14356 15442 14368
rect 16758 14356 16764 14368
rect 16816 14356 16822 14408
rect 9088 14300 11652 14328
rect 12713 14331 12771 14337
rect 9088 14288 9094 14300
rect 12713 14297 12725 14331
rect 12759 14328 12771 14331
rect 13170 14328 13176 14340
rect 12759 14300 13176 14328
rect 12759 14297 12771 14300
rect 12713 14291 12771 14297
rect 13170 14288 13176 14300
rect 13228 14288 13234 14340
rect 13538 14328 13544 14340
rect 13499 14300 13544 14328
rect 13538 14288 13544 14300
rect 13596 14288 13602 14340
rect 1486 14260 1492 14272
rect 1447 14232 1492 14260
rect 1486 14220 1492 14232
rect 1544 14220 1550 14272
rect 3234 14220 3240 14272
rect 3292 14260 3298 14272
rect 3513 14263 3571 14269
rect 3513 14260 3525 14263
rect 3292 14232 3525 14260
rect 3292 14220 3298 14232
rect 3513 14229 3525 14232
rect 3559 14229 3571 14263
rect 3513 14223 3571 14229
rect 4062 14220 4068 14272
rect 4120 14260 4126 14272
rect 4157 14263 4215 14269
rect 4157 14260 4169 14263
rect 4120 14232 4169 14260
rect 4120 14220 4126 14232
rect 4157 14229 4169 14232
rect 4203 14229 4215 14263
rect 4157 14223 4215 14229
rect 5077 14263 5135 14269
rect 5077 14229 5089 14263
rect 5123 14260 5135 14263
rect 5166 14260 5172 14272
rect 5123 14232 5172 14260
rect 5123 14229 5135 14232
rect 5077 14223 5135 14229
rect 5166 14220 5172 14232
rect 5224 14220 5230 14272
rect 5810 14220 5816 14272
rect 5868 14260 5874 14272
rect 6549 14263 6607 14269
rect 6549 14260 6561 14263
rect 5868 14232 6561 14260
rect 5868 14220 5874 14232
rect 6549 14229 6561 14232
rect 6595 14229 6607 14263
rect 6549 14223 6607 14229
rect 7190 14220 7196 14272
rect 7248 14260 7254 14272
rect 10597 14263 10655 14269
rect 10597 14260 10609 14263
rect 7248 14232 10609 14260
rect 7248 14220 7254 14232
rect 10597 14229 10609 14232
rect 10643 14260 10655 14263
rect 10686 14260 10692 14272
rect 10643 14232 10692 14260
rect 10643 14229 10655 14232
rect 10597 14223 10655 14229
rect 10686 14220 10692 14232
rect 10744 14260 10750 14272
rect 11057 14263 11115 14269
rect 11057 14260 11069 14263
rect 10744 14232 11069 14260
rect 10744 14220 10750 14232
rect 11057 14229 11069 14232
rect 11103 14229 11115 14263
rect 11422 14260 11428 14272
rect 11383 14232 11428 14260
rect 11057 14223 11115 14229
rect 11422 14220 11428 14232
rect 11480 14220 11486 14272
rect 11514 14220 11520 14272
rect 11572 14260 11578 14272
rect 11698 14260 11704 14272
rect 11572 14232 11704 14260
rect 11572 14220 11578 14232
rect 11698 14220 11704 14232
rect 11756 14220 11762 14272
rect 12250 14220 12256 14272
rect 12308 14260 12314 14272
rect 12308 14232 12353 14260
rect 12308 14220 12314 14232
rect 12434 14220 12440 14272
rect 12492 14260 12498 14272
rect 12618 14260 12624 14272
rect 12492 14232 12624 14260
rect 12492 14220 12498 14232
rect 12618 14220 12624 14232
rect 12676 14220 12682 14272
rect 13633 14263 13691 14269
rect 13633 14229 13645 14263
rect 13679 14260 13691 14263
rect 14090 14260 14096 14272
rect 13679 14232 14096 14260
rect 13679 14229 13691 14232
rect 13633 14223 13691 14229
rect 14090 14220 14096 14232
rect 14148 14220 14154 14272
rect 1104 14170 16008 14192
rect 1104 14118 4698 14170
rect 4750 14118 4762 14170
rect 4814 14118 4826 14170
rect 4878 14118 4890 14170
rect 4942 14118 4954 14170
rect 5006 14118 8446 14170
rect 8498 14118 8510 14170
rect 8562 14118 8574 14170
rect 8626 14118 8638 14170
rect 8690 14118 8702 14170
rect 8754 14118 12194 14170
rect 12246 14118 12258 14170
rect 12310 14118 12322 14170
rect 12374 14118 12386 14170
rect 12438 14118 12450 14170
rect 12502 14118 16008 14170
rect 1104 14096 16008 14118
rect 1397 14059 1455 14065
rect 1397 14025 1409 14059
rect 1443 14056 1455 14059
rect 1670 14056 1676 14068
rect 1443 14028 1676 14056
rect 1443 14025 1455 14028
rect 1397 14019 1455 14025
rect 1670 14016 1676 14028
rect 1728 14016 1734 14068
rect 1762 14016 1768 14068
rect 1820 14056 1826 14068
rect 2225 14059 2283 14065
rect 2225 14056 2237 14059
rect 1820 14028 2237 14056
rect 1820 14016 1826 14028
rect 2225 14025 2237 14028
rect 2271 14025 2283 14059
rect 2225 14019 2283 14025
rect 2501 14059 2559 14065
rect 2501 14025 2513 14059
rect 2547 14056 2559 14059
rect 2590 14056 2596 14068
rect 2547 14028 2596 14056
rect 2547 14025 2559 14028
rect 2501 14019 2559 14025
rect 2590 14016 2596 14028
rect 2648 14016 2654 14068
rect 2866 14056 2872 14068
rect 2827 14028 2872 14056
rect 2866 14016 2872 14028
rect 2924 14016 2930 14068
rect 3142 14056 3148 14068
rect 3103 14028 3148 14056
rect 3142 14016 3148 14028
rect 3200 14016 3206 14068
rect 4614 14056 4620 14068
rect 4575 14028 4620 14056
rect 4614 14016 4620 14028
rect 4672 14016 4678 14068
rect 5442 14016 5448 14068
rect 5500 14056 5506 14068
rect 5629 14059 5687 14065
rect 5629 14056 5641 14059
rect 5500 14028 5641 14056
rect 5500 14016 5506 14028
rect 5629 14025 5641 14028
rect 5675 14056 5687 14059
rect 5718 14056 5724 14068
rect 5675 14028 5724 14056
rect 5675 14025 5687 14028
rect 5629 14019 5687 14025
rect 5718 14016 5724 14028
rect 5776 14056 5782 14068
rect 6365 14059 6423 14065
rect 6365 14056 6377 14059
rect 5776 14028 6377 14056
rect 5776 14016 5782 14028
rect 6365 14025 6377 14028
rect 6411 14056 6423 14059
rect 6454 14056 6460 14068
rect 6411 14028 6460 14056
rect 6411 14025 6423 14028
rect 6365 14019 6423 14025
rect 6454 14016 6460 14028
rect 6512 14056 6518 14068
rect 6914 14056 6920 14068
rect 6512 14028 6920 14056
rect 6512 14016 6518 14028
rect 6914 14016 6920 14028
rect 6972 14056 6978 14068
rect 6972 14028 7065 14056
rect 6972 14016 6978 14028
rect 7282 14016 7288 14068
rect 7340 14056 7346 14068
rect 8018 14056 8024 14068
rect 7340 14028 8024 14056
rect 7340 14016 7346 14028
rect 8018 14016 8024 14028
rect 8076 14016 8082 14068
rect 9401 14059 9459 14065
rect 9401 14056 9413 14059
rect 8588 14028 9413 14056
rect 2314 13948 2320 14000
rect 2372 13988 2378 14000
rect 2372 13960 3004 13988
rect 2372 13948 2378 13960
rect 1765 13923 1823 13929
rect 1765 13889 1777 13923
rect 1811 13920 1823 13923
rect 2406 13920 2412 13932
rect 1811 13892 2268 13920
rect 2367 13892 2412 13920
rect 1811 13889 1823 13892
rect 1765 13883 1823 13889
rect 1857 13855 1915 13861
rect 1857 13821 1869 13855
rect 1903 13821 1915 13855
rect 1857 13815 1915 13821
rect 2041 13855 2099 13861
rect 2041 13821 2053 13855
rect 2087 13821 2099 13855
rect 2240 13852 2268 13892
rect 2406 13880 2412 13892
rect 2464 13880 2470 13932
rect 2685 13923 2743 13929
rect 2685 13889 2697 13923
rect 2731 13920 2743 13923
rect 2866 13920 2872 13932
rect 2731 13892 2872 13920
rect 2731 13889 2743 13892
rect 2685 13883 2743 13889
rect 2866 13880 2872 13892
rect 2924 13880 2930 13932
rect 2774 13852 2780 13864
rect 2240 13824 2780 13852
rect 2041 13815 2099 13821
rect 1872 13716 1900 13815
rect 2056 13784 2084 13815
rect 2774 13812 2780 13824
rect 2832 13812 2838 13864
rect 2976 13852 3004 13960
rect 3160 13920 3188 14016
rect 3878 13948 3884 14000
rect 3936 13988 3942 14000
rect 5537 13991 5595 13997
rect 5537 13988 5549 13991
rect 3936 13960 5549 13988
rect 3936 13948 3942 13960
rect 5537 13957 5549 13960
rect 5583 13988 5595 13991
rect 6086 13988 6092 14000
rect 5583 13960 6092 13988
rect 5583 13957 5595 13960
rect 5537 13951 5595 13957
rect 6086 13948 6092 13960
rect 6144 13948 6150 14000
rect 8588 13988 8616 14028
rect 9401 14025 9413 14028
rect 9447 14025 9459 14059
rect 9401 14019 9459 14025
rect 9674 14016 9680 14068
rect 9732 14056 9738 14068
rect 11057 14059 11115 14065
rect 11057 14056 11069 14059
rect 9732 14028 11069 14056
rect 9732 14016 9738 14028
rect 11057 14025 11069 14028
rect 11103 14025 11115 14059
rect 11057 14019 11115 14025
rect 11333 14059 11391 14065
rect 11333 14025 11345 14059
rect 11379 14056 11391 14059
rect 11606 14056 11612 14068
rect 11379 14028 11612 14056
rect 11379 14025 11391 14028
rect 11333 14019 11391 14025
rect 11606 14016 11612 14028
rect 11664 14016 11670 14068
rect 12618 14016 12624 14068
rect 12676 14056 12682 14068
rect 12713 14059 12771 14065
rect 12713 14056 12725 14059
rect 12676 14028 12725 14056
rect 12676 14016 12682 14028
rect 12713 14025 12725 14028
rect 12759 14025 12771 14059
rect 13170 14056 13176 14068
rect 13131 14028 13176 14056
rect 12713 14019 12771 14025
rect 13170 14016 13176 14028
rect 13228 14016 13234 14068
rect 13446 14056 13452 14068
rect 13407 14028 13452 14056
rect 13446 14016 13452 14028
rect 13504 14016 13510 14068
rect 13814 14056 13820 14068
rect 13775 14028 13820 14056
rect 13814 14016 13820 14028
rect 13872 14016 13878 14068
rect 15105 14059 15163 14065
rect 15105 14025 15117 14059
rect 15151 14056 15163 14059
rect 15194 14056 15200 14068
rect 15151 14028 15200 14056
rect 15151 14025 15163 14028
rect 15105 14019 15163 14025
rect 15194 14016 15200 14028
rect 15252 14016 15258 14068
rect 15378 14016 15384 14068
rect 15436 14056 15442 14068
rect 15473 14059 15531 14065
rect 15473 14056 15485 14059
rect 15436 14028 15485 14056
rect 15436 14016 15442 14028
rect 15473 14025 15485 14028
rect 15519 14025 15531 14059
rect 15654 14056 15660 14068
rect 15615 14028 15660 14056
rect 15473 14019 15531 14025
rect 15654 14016 15660 14028
rect 15712 14016 15718 14068
rect 6840 13960 8616 13988
rect 9309 13991 9367 13997
rect 3237 13923 3295 13929
rect 3237 13920 3249 13923
rect 3160 13892 3249 13920
rect 3237 13889 3249 13892
rect 3283 13889 3295 13923
rect 3493 13923 3551 13929
rect 3493 13920 3505 13923
rect 3237 13883 3295 13889
rect 3344 13892 3505 13920
rect 3344 13852 3372 13892
rect 3493 13889 3505 13892
rect 3539 13889 3551 13923
rect 3493 13883 3551 13889
rect 3970 13880 3976 13932
rect 4028 13920 4034 13932
rect 4028 13892 4292 13920
rect 4028 13880 4034 13892
rect 2976 13824 3372 13852
rect 4264 13852 4292 13892
rect 5902 13880 5908 13932
rect 5960 13920 5966 13932
rect 6840 13920 6868 13960
rect 9309 13957 9321 13991
rect 9355 13988 9367 13991
rect 10594 13988 10600 14000
rect 9355 13960 10600 13988
rect 9355 13957 9367 13960
rect 9309 13951 9367 13957
rect 10594 13948 10600 13960
rect 10652 13948 10658 14000
rect 12434 13948 12440 14000
rect 12492 13988 12498 14000
rect 14185 13991 14243 13997
rect 14185 13988 14197 13991
rect 12492 13960 14197 13988
rect 12492 13948 12498 13960
rect 14185 13957 14197 13960
rect 14231 13957 14243 13991
rect 14185 13951 14243 13957
rect 5960 13892 6868 13920
rect 5960 13880 5966 13892
rect 6914 13880 6920 13932
rect 6972 13920 6978 13932
rect 7101 13923 7159 13929
rect 7101 13920 7113 13923
rect 6972 13892 7113 13920
rect 6972 13880 6978 13892
rect 7101 13889 7113 13892
rect 7147 13889 7159 13923
rect 7101 13883 7159 13889
rect 7190 13880 7196 13932
rect 7248 13920 7254 13932
rect 7357 13923 7415 13929
rect 7357 13920 7369 13923
rect 7248 13892 7369 13920
rect 7248 13880 7254 13892
rect 7357 13889 7369 13892
rect 7403 13889 7415 13923
rect 7357 13883 7415 13889
rect 8294 13880 8300 13932
rect 8352 13920 8358 13932
rect 9030 13920 9036 13932
rect 8352 13892 9036 13920
rect 8352 13880 8358 13892
rect 9030 13880 9036 13892
rect 9088 13880 9094 13932
rect 10226 13880 10232 13932
rect 10284 13920 10290 13932
rect 10514 13923 10572 13929
rect 10514 13920 10526 13923
rect 10284 13892 10526 13920
rect 10284 13880 10290 13892
rect 10514 13889 10526 13892
rect 10560 13889 10572 13923
rect 10612 13920 10640 13948
rect 10781 13923 10839 13929
rect 10781 13920 10793 13923
rect 10612 13892 10793 13920
rect 10514 13883 10572 13889
rect 10781 13889 10793 13892
rect 10827 13889 10839 13923
rect 10781 13883 10839 13889
rect 11054 13880 11060 13932
rect 11112 13920 11118 13932
rect 11514 13920 11520 13932
rect 11112 13892 11520 13920
rect 11112 13880 11118 13892
rect 11514 13880 11520 13892
rect 11572 13920 11578 13932
rect 11885 13923 11943 13929
rect 11885 13920 11897 13923
rect 11572 13892 11897 13920
rect 11572 13880 11578 13892
rect 11885 13889 11897 13892
rect 11931 13889 11943 13923
rect 11885 13883 11943 13889
rect 12805 13923 12863 13929
rect 12805 13889 12817 13923
rect 12851 13920 12863 13923
rect 14642 13920 14648 13932
rect 12851 13892 14648 13920
rect 12851 13889 12863 13892
rect 12805 13883 12863 13889
rect 14642 13880 14648 13892
rect 14700 13880 14706 13932
rect 6454 13852 6460 13864
rect 4264 13824 6460 13852
rect 6454 13812 6460 13824
rect 6512 13812 6518 13864
rect 11609 13855 11667 13861
rect 11609 13821 11621 13855
rect 11655 13821 11667 13855
rect 11790 13852 11796 13864
rect 11751 13824 11796 13852
rect 11609 13815 11667 13821
rect 2056 13756 2774 13784
rect 2314 13716 2320 13728
rect 1872 13688 2320 13716
rect 2314 13676 2320 13688
rect 2372 13676 2378 13728
rect 2746 13716 2774 13756
rect 4706 13744 4712 13796
rect 4764 13784 4770 13796
rect 4764 13756 6316 13784
rect 4764 13744 4770 13756
rect 6178 13716 6184 13728
rect 2746 13688 6184 13716
rect 6178 13676 6184 13688
rect 6236 13676 6242 13728
rect 6288 13716 6316 13756
rect 8110 13744 8116 13796
rect 8168 13784 8174 13796
rect 8481 13787 8539 13793
rect 8481 13784 8493 13787
rect 8168 13756 8493 13784
rect 8168 13744 8174 13756
rect 8481 13753 8493 13756
rect 8527 13753 8539 13787
rect 11624 13784 11652 13815
rect 11790 13812 11796 13824
rect 11848 13812 11854 13864
rect 12894 13852 12900 13864
rect 12855 13824 12900 13852
rect 12894 13812 12900 13824
rect 12952 13812 12958 13864
rect 13725 13855 13783 13861
rect 13725 13821 13737 13855
rect 13771 13852 13783 13855
rect 13814 13852 13820 13864
rect 13771 13824 13820 13852
rect 13771 13821 13783 13824
rect 13725 13815 13783 13821
rect 13814 13812 13820 13824
rect 13872 13812 13878 13864
rect 13906 13812 13912 13864
rect 13964 13852 13970 13864
rect 14277 13855 14335 13861
rect 14277 13852 14289 13855
rect 13964 13824 14289 13852
rect 13964 13812 13970 13824
rect 14277 13821 14289 13824
rect 14323 13821 14335 13855
rect 14277 13815 14335 13821
rect 14461 13855 14519 13861
rect 14461 13821 14473 13855
rect 14507 13821 14519 13855
rect 14461 13815 14519 13821
rect 14921 13855 14979 13861
rect 14921 13821 14933 13855
rect 14967 13821 14979 13855
rect 14921 13815 14979 13821
rect 15013 13855 15071 13861
rect 15013 13821 15025 13855
rect 15059 13852 15071 13855
rect 15838 13852 15844 13864
rect 15059 13824 15844 13852
rect 15059 13821 15071 13824
rect 15013 13815 15071 13821
rect 11698 13784 11704 13796
rect 11624 13756 11704 13784
rect 8481 13747 8539 13753
rect 11698 13744 11704 13756
rect 11756 13744 11762 13796
rect 12066 13744 12072 13796
rect 12124 13784 12130 13796
rect 12253 13787 12311 13793
rect 12253 13784 12265 13787
rect 12124 13756 12265 13784
rect 12124 13744 12130 13756
rect 12253 13753 12265 13756
rect 12299 13753 12311 13787
rect 12253 13747 12311 13753
rect 13446 13744 13452 13796
rect 13504 13784 13510 13796
rect 13998 13784 14004 13796
rect 13504 13756 14004 13784
rect 13504 13744 13510 13756
rect 13998 13744 14004 13756
rect 14056 13744 14062 13796
rect 14476 13728 14504 13815
rect 14936 13784 14964 13815
rect 15838 13812 15844 13824
rect 15896 13812 15902 13864
rect 15102 13784 15108 13796
rect 14936 13756 15108 13784
rect 15102 13744 15108 13756
rect 15160 13744 15166 13796
rect 11606 13716 11612 13728
rect 6288 13688 11612 13716
rect 11606 13676 11612 13688
rect 11664 13676 11670 13728
rect 11974 13676 11980 13728
rect 12032 13716 12038 13728
rect 12345 13719 12403 13725
rect 12345 13716 12357 13719
rect 12032 13688 12357 13716
rect 12032 13676 12038 13688
rect 12345 13685 12357 13688
rect 12391 13685 12403 13719
rect 12345 13679 12403 13685
rect 13630 13676 13636 13728
rect 13688 13716 13694 13728
rect 14090 13716 14096 13728
rect 13688 13688 14096 13716
rect 13688 13676 13694 13688
rect 14090 13676 14096 13688
rect 14148 13676 14154 13728
rect 14458 13676 14464 13728
rect 14516 13676 14522 13728
rect 1104 13626 16008 13648
rect 1104 13574 2824 13626
rect 2876 13574 2888 13626
rect 2940 13574 2952 13626
rect 3004 13574 3016 13626
rect 3068 13574 3080 13626
rect 3132 13574 6572 13626
rect 6624 13574 6636 13626
rect 6688 13574 6700 13626
rect 6752 13574 6764 13626
rect 6816 13574 6828 13626
rect 6880 13574 10320 13626
rect 10372 13574 10384 13626
rect 10436 13574 10448 13626
rect 10500 13574 10512 13626
rect 10564 13574 10576 13626
rect 10628 13574 14068 13626
rect 14120 13574 14132 13626
rect 14184 13574 14196 13626
rect 14248 13574 14260 13626
rect 14312 13574 14324 13626
rect 14376 13574 16008 13626
rect 1104 13552 16008 13574
rect 1857 13515 1915 13521
rect 1857 13481 1869 13515
rect 1903 13512 1915 13515
rect 2222 13512 2228 13524
rect 1903 13484 2228 13512
rect 1903 13481 1915 13484
rect 1857 13475 1915 13481
rect 2222 13472 2228 13484
rect 2280 13472 2286 13524
rect 4154 13512 4160 13524
rect 4115 13484 4160 13512
rect 4154 13472 4160 13484
rect 4212 13472 4218 13524
rect 6178 13472 6184 13524
rect 6236 13512 6242 13524
rect 9306 13512 9312 13524
rect 6236 13484 9312 13512
rect 6236 13472 6242 13484
rect 9306 13472 9312 13484
rect 9364 13472 9370 13524
rect 10134 13472 10140 13524
rect 10192 13512 10198 13524
rect 10413 13515 10471 13521
rect 10413 13512 10425 13515
rect 10192 13484 10425 13512
rect 10192 13472 10198 13484
rect 10413 13481 10425 13484
rect 10459 13512 10471 13515
rect 10870 13512 10876 13524
rect 10459 13484 10876 13512
rect 10459 13481 10471 13484
rect 10413 13475 10471 13481
rect 10870 13472 10876 13484
rect 10928 13472 10934 13524
rect 11606 13472 11612 13524
rect 11664 13512 11670 13524
rect 11664 13484 11753 13512
rect 11664 13472 11670 13484
rect 7377 13447 7435 13453
rect 7377 13413 7389 13447
rect 7423 13413 7435 13447
rect 7377 13407 7435 13413
rect 10980 13416 11652 13444
rect 3602 13336 3608 13388
rect 3660 13376 3666 13388
rect 4154 13376 4160 13388
rect 3660 13348 4160 13376
rect 3660 13336 3666 13348
rect 4154 13336 4160 13348
rect 4212 13376 4218 13388
rect 4706 13376 4712 13388
rect 4212 13348 4712 13376
rect 4212 13336 4218 13348
rect 4706 13336 4712 13348
rect 4764 13336 4770 13388
rect 5718 13376 5724 13388
rect 5679 13348 5724 13376
rect 5718 13336 5724 13348
rect 5776 13376 5782 13388
rect 5813 13379 5871 13385
rect 5813 13376 5825 13379
rect 5776 13348 5825 13376
rect 5776 13336 5782 13348
rect 5813 13345 5825 13348
rect 5859 13345 5871 13379
rect 5813 13339 5871 13345
rect 1673 13311 1731 13317
rect 1673 13277 1685 13311
rect 1719 13308 1731 13311
rect 1854 13308 1860 13320
rect 1719 13280 1860 13308
rect 1719 13277 1731 13280
rect 1673 13271 1731 13277
rect 1854 13268 1860 13280
rect 1912 13268 1918 13320
rect 7392 13308 7420 13407
rect 6021 13280 7420 13308
rect 8757 13311 8815 13317
rect 5442 13240 5448 13252
rect 5500 13249 5506 13252
rect 5500 13243 5534 13249
rect 5386 13212 5448 13240
rect 5442 13200 5448 13212
rect 5522 13240 5534 13243
rect 6021 13240 6049 13280
rect 8757 13277 8769 13311
rect 8803 13308 8815 13311
rect 9030 13308 9036 13320
rect 8803 13280 9036 13308
rect 8803 13277 8815 13280
rect 8757 13271 8815 13277
rect 9030 13268 9036 13280
rect 9088 13268 9094 13320
rect 10980 13308 11008 13416
rect 11624 13385 11652 13416
rect 11609 13379 11667 13385
rect 11609 13345 11621 13379
rect 11655 13345 11667 13379
rect 11725 13376 11753 13484
rect 11790 13472 11796 13524
rect 11848 13512 11854 13524
rect 11885 13515 11943 13521
rect 11885 13512 11897 13515
rect 11848 13484 11897 13512
rect 11848 13472 11854 13484
rect 11885 13481 11897 13484
rect 11931 13481 11943 13515
rect 11885 13475 11943 13481
rect 12250 13472 12256 13524
rect 12308 13512 12314 13524
rect 13538 13512 13544 13524
rect 12308 13484 13544 13512
rect 12308 13472 12314 13484
rect 13004 13456 13032 13484
rect 13538 13472 13544 13484
rect 13596 13472 13602 13524
rect 13722 13512 13728 13524
rect 13683 13484 13728 13512
rect 13722 13472 13728 13484
rect 13780 13472 13786 13524
rect 13814 13472 13820 13524
rect 13872 13512 13878 13524
rect 14093 13515 14151 13521
rect 14093 13512 14105 13515
rect 13872 13484 14105 13512
rect 13872 13472 13878 13484
rect 14093 13481 14105 13484
rect 14139 13481 14151 13515
rect 14550 13512 14556 13524
rect 14511 13484 14556 13512
rect 14093 13475 14151 13481
rect 14550 13472 14556 13484
rect 14608 13472 14614 13524
rect 14642 13472 14648 13524
rect 14700 13512 14706 13524
rect 14700 13484 14745 13512
rect 14700 13472 14706 13484
rect 15194 13472 15200 13524
rect 15252 13512 15258 13524
rect 15252 13484 15700 13512
rect 15252 13472 15258 13484
rect 11974 13404 11980 13456
rect 12032 13444 12038 13456
rect 12713 13447 12771 13453
rect 12713 13444 12725 13447
rect 12032 13416 12725 13444
rect 12032 13404 12038 13416
rect 12713 13413 12725 13416
rect 12759 13413 12771 13447
rect 12713 13407 12771 13413
rect 12986 13404 12992 13456
rect 13044 13404 13050 13456
rect 13170 13404 13176 13456
rect 13228 13444 13234 13456
rect 13740 13444 13768 13472
rect 15102 13444 15108 13456
rect 13228 13416 13768 13444
rect 14568 13416 15108 13444
rect 13228 13404 13234 13416
rect 14568 13388 14596 13416
rect 15102 13404 15108 13416
rect 15160 13404 15166 13456
rect 15562 13404 15568 13456
rect 15620 13404 15626 13456
rect 11790 13376 11796 13388
rect 11725 13348 11796 13376
rect 11609 13339 11667 13345
rect 11790 13336 11796 13348
rect 11848 13336 11854 13388
rect 12066 13336 12072 13388
rect 12124 13376 12130 13388
rect 12437 13379 12495 13385
rect 12437 13376 12449 13379
rect 12124 13348 12449 13376
rect 12124 13336 12130 13348
rect 12437 13345 12449 13348
rect 12483 13345 12495 13379
rect 12437 13339 12495 13345
rect 12802 13336 12808 13388
rect 12860 13376 12866 13388
rect 13265 13379 13323 13385
rect 13265 13376 13277 13379
rect 12860 13348 13277 13376
rect 12860 13336 12866 13348
rect 13265 13345 13277 13348
rect 13311 13345 13323 13379
rect 13265 13339 13323 13345
rect 14550 13336 14556 13388
rect 14608 13336 14614 13388
rect 15197 13379 15255 13385
rect 15197 13376 15209 13379
rect 14660 13348 15209 13376
rect 9232 13280 11008 13308
rect 11256 13280 12388 13308
rect 6086 13249 6092 13252
rect 5522 13212 6049 13240
rect 5522 13209 5534 13212
rect 5500 13203 5534 13209
rect 6080 13203 6092 13249
rect 6144 13240 6150 13252
rect 6144 13212 6180 13240
rect 5500 13200 5506 13203
rect 6086 13200 6092 13203
rect 6144 13200 6150 13212
rect 6362 13200 6368 13252
rect 6420 13240 6426 13252
rect 8490 13243 8548 13249
rect 8490 13240 8502 13243
rect 6420 13212 8502 13240
rect 6420 13200 6426 13212
rect 8490 13209 8502 13212
rect 8536 13240 8548 13243
rect 9232 13240 9260 13280
rect 8536 13212 9260 13240
rect 9300 13243 9358 13249
rect 8536 13209 8548 13212
rect 8490 13203 8548 13209
rect 9300 13209 9312 13243
rect 9346 13240 9358 13243
rect 9674 13240 9680 13252
rect 9346 13212 9680 13240
rect 9346 13209 9358 13212
rect 9300 13203 9358 13209
rect 1486 13172 1492 13184
rect 1447 13144 1492 13172
rect 1486 13132 1492 13144
rect 1544 13132 1550 13184
rect 4246 13132 4252 13184
rect 4304 13172 4310 13184
rect 4341 13175 4399 13181
rect 4341 13172 4353 13175
rect 4304 13144 4353 13172
rect 4304 13132 4310 13144
rect 4341 13141 4353 13144
rect 4387 13172 4399 13175
rect 5074 13172 5080 13184
rect 4387 13144 5080 13172
rect 4387 13141 4399 13144
rect 4341 13135 4399 13141
rect 5074 13132 5080 13144
rect 5132 13132 5138 13184
rect 5902 13132 5908 13184
rect 5960 13172 5966 13184
rect 6178 13172 6184 13184
rect 5960 13144 6184 13172
rect 5960 13132 5966 13144
rect 6178 13132 6184 13144
rect 6236 13132 6242 13184
rect 7193 13175 7251 13181
rect 7193 13141 7205 13175
rect 7239 13172 7251 13175
rect 7282 13172 7288 13184
rect 7239 13144 7288 13172
rect 7239 13141 7251 13144
rect 7193 13135 7251 13141
rect 7282 13132 7288 13144
rect 7340 13132 7346 13184
rect 8938 13132 8944 13184
rect 8996 13172 9002 13184
rect 9324 13172 9352 13203
rect 9674 13200 9680 13212
rect 9732 13200 9738 13252
rect 10778 13200 10784 13252
rect 10836 13240 10842 13252
rect 11256 13240 11284 13280
rect 12250 13240 12256 13252
rect 10836 13212 11284 13240
rect 12211 13212 12256 13240
rect 10836 13200 10842 13212
rect 12250 13200 12256 13212
rect 12308 13200 12314 13252
rect 12360 13249 12388 13280
rect 12345 13243 12403 13249
rect 12345 13209 12357 13243
rect 12391 13209 12403 13243
rect 12345 13203 12403 13209
rect 13081 13243 13139 13249
rect 13081 13209 13093 13243
rect 13127 13240 13139 13243
rect 13262 13240 13268 13252
rect 13127 13212 13268 13240
rect 13127 13209 13139 13212
rect 13081 13203 13139 13209
rect 13262 13200 13268 13212
rect 13320 13200 13326 13252
rect 13814 13240 13820 13252
rect 13372 13212 13820 13240
rect 11054 13172 11060 13184
rect 8996 13144 9352 13172
rect 11015 13144 11060 13172
rect 8996 13132 9002 13144
rect 11054 13132 11060 13144
rect 11112 13132 11118 13184
rect 11422 13172 11428 13184
rect 11383 13144 11428 13172
rect 11422 13132 11428 13144
rect 11480 13132 11486 13184
rect 11517 13175 11575 13181
rect 11517 13141 11529 13175
rect 11563 13172 11575 13175
rect 11606 13172 11612 13184
rect 11563 13144 11612 13172
rect 11563 13141 11575 13144
rect 11517 13135 11575 13141
rect 11606 13132 11612 13144
rect 11664 13132 11670 13184
rect 13173 13175 13231 13181
rect 13173 13141 13185 13175
rect 13219 13172 13231 13175
rect 13372 13172 13400 13212
rect 13814 13200 13820 13212
rect 13872 13200 13878 13252
rect 14660 13240 14688 13348
rect 15197 13345 15209 13348
rect 15243 13345 15255 13379
rect 15580 13376 15608 13404
rect 15197 13339 15255 13345
rect 15304 13348 15608 13376
rect 15105 13311 15163 13317
rect 15105 13277 15117 13311
rect 15151 13308 15163 13311
rect 15151 13280 15240 13308
rect 15151 13277 15163 13280
rect 15105 13271 15163 13277
rect 15212 13252 15240 13280
rect 14016 13212 14688 13240
rect 14016 13184 14044 13212
rect 15194 13200 15200 13252
rect 15252 13200 15258 13252
rect 15304 13184 15332 13348
rect 15672 13317 15700 13484
rect 15657 13311 15715 13317
rect 15657 13277 15669 13311
rect 15703 13277 15715 13311
rect 15657 13271 15715 13277
rect 13219 13144 13400 13172
rect 13219 13141 13231 13144
rect 13173 13135 13231 13141
rect 13446 13132 13452 13184
rect 13504 13172 13510 13184
rect 13998 13172 14004 13184
rect 13504 13144 14004 13172
rect 13504 13132 13510 13144
rect 13998 13132 14004 13144
rect 14056 13132 14062 13184
rect 14274 13172 14280 13184
rect 14235 13144 14280 13172
rect 14274 13132 14280 13144
rect 14332 13132 14338 13184
rect 15013 13175 15071 13181
rect 15013 13141 15025 13175
rect 15059 13172 15071 13175
rect 15286 13172 15292 13184
rect 15059 13144 15292 13172
rect 15059 13141 15071 13144
rect 15013 13135 15071 13141
rect 15286 13132 15292 13144
rect 15344 13132 15350 13184
rect 15473 13175 15531 13181
rect 15473 13141 15485 13175
rect 15519 13172 15531 13175
rect 15746 13172 15752 13184
rect 15519 13144 15752 13172
rect 15519 13141 15531 13144
rect 15473 13135 15531 13141
rect 15746 13132 15752 13144
rect 15804 13132 15810 13184
rect 1104 13082 16008 13104
rect 1104 13030 4698 13082
rect 4750 13030 4762 13082
rect 4814 13030 4826 13082
rect 4878 13030 4890 13082
rect 4942 13030 4954 13082
rect 5006 13030 8446 13082
rect 8498 13030 8510 13082
rect 8562 13030 8574 13082
rect 8626 13030 8638 13082
rect 8690 13030 8702 13082
rect 8754 13030 12194 13082
rect 12246 13030 12258 13082
rect 12310 13030 12322 13082
rect 12374 13030 12386 13082
rect 12438 13030 12450 13082
rect 12502 13030 16008 13082
rect 1104 13008 16008 13030
rect 2777 12971 2835 12977
rect 2777 12937 2789 12971
rect 2823 12968 2835 12971
rect 3142 12968 3148 12980
rect 2823 12940 3148 12968
rect 2823 12937 2835 12940
rect 2777 12931 2835 12937
rect 1578 12792 1584 12844
rect 1636 12832 1642 12844
rect 1673 12835 1731 12841
rect 1673 12832 1685 12835
rect 1636 12804 1685 12832
rect 1636 12792 1642 12804
rect 1673 12801 1685 12804
rect 1719 12801 1731 12835
rect 1946 12832 1952 12844
rect 1907 12804 1952 12832
rect 1673 12795 1731 12801
rect 1946 12792 1952 12804
rect 2004 12792 2010 12844
rect 2884 12841 2912 12940
rect 3142 12928 3148 12940
rect 3200 12928 3206 12980
rect 4433 12971 4491 12977
rect 4433 12968 4445 12971
rect 4356 12940 4445 12968
rect 2869 12835 2927 12841
rect 2869 12801 2881 12835
rect 2915 12801 2927 12835
rect 2869 12795 2927 12801
rect 3136 12835 3194 12841
rect 3136 12801 3148 12835
rect 3182 12832 3194 12835
rect 4356 12832 4384 12940
rect 4433 12937 4445 12940
rect 4479 12937 4491 12971
rect 4433 12931 4491 12937
rect 5626 12928 5632 12980
rect 5684 12968 5690 12980
rect 6086 12968 6092 12980
rect 5684 12940 6092 12968
rect 5684 12928 5690 12940
rect 6086 12928 6092 12940
rect 6144 12928 6150 12980
rect 6914 12928 6920 12980
rect 6972 12968 6978 12980
rect 7009 12971 7067 12977
rect 7009 12968 7021 12971
rect 6972 12940 7021 12968
rect 6972 12928 6978 12940
rect 7009 12937 7021 12940
rect 7055 12968 7067 12971
rect 7193 12971 7251 12977
rect 7193 12968 7205 12971
rect 7055 12940 7205 12968
rect 7055 12937 7067 12940
rect 7009 12931 7067 12937
rect 7193 12937 7205 12940
rect 7239 12968 7251 12971
rect 8941 12971 8999 12977
rect 8941 12968 8953 12971
rect 7239 12940 8953 12968
rect 7239 12937 7251 12940
rect 7193 12931 7251 12937
rect 5074 12860 5080 12912
rect 5132 12900 5138 12912
rect 5132 12872 5948 12900
rect 5132 12860 5138 12872
rect 3182 12804 4384 12832
rect 3182 12801 3194 12804
rect 3136 12795 3194 12801
rect 4356 12764 4384 12804
rect 5258 12792 5264 12844
rect 5316 12832 5322 12844
rect 5546 12835 5604 12841
rect 5546 12832 5558 12835
rect 5316 12804 5558 12832
rect 5316 12792 5322 12804
rect 5546 12801 5558 12804
rect 5592 12801 5604 12835
rect 5546 12795 5604 12801
rect 5718 12792 5724 12844
rect 5776 12832 5782 12844
rect 5813 12835 5871 12841
rect 5813 12832 5825 12835
rect 5776 12804 5825 12832
rect 5776 12792 5782 12804
rect 5813 12801 5825 12804
rect 5859 12801 5871 12835
rect 5813 12795 5871 12801
rect 4430 12764 4436 12776
rect 4356 12736 4436 12764
rect 4430 12724 4436 12736
rect 4488 12724 4494 12776
rect 5828 12696 5856 12795
rect 5920 12764 5948 12872
rect 7300 12841 7328 12940
rect 8941 12937 8953 12940
rect 8987 12968 8999 12971
rect 9030 12968 9036 12980
rect 8987 12940 9036 12968
rect 8987 12937 8999 12940
rect 8941 12931 8999 12937
rect 9030 12928 9036 12940
rect 9088 12968 9094 12980
rect 9309 12971 9367 12977
rect 9309 12968 9321 12971
rect 9088 12940 9321 12968
rect 9088 12928 9094 12940
rect 9309 12937 9321 12940
rect 9355 12937 9367 12971
rect 9309 12931 9367 12937
rect 9674 12928 9680 12980
rect 9732 12968 9738 12980
rect 10778 12968 10784 12980
rect 9732 12940 10784 12968
rect 9732 12928 9738 12940
rect 10778 12928 10784 12940
rect 10836 12968 10842 12980
rect 11701 12971 11759 12977
rect 11701 12968 11713 12971
rect 10836 12940 11713 12968
rect 10836 12928 10842 12940
rect 11701 12937 11713 12940
rect 11747 12937 11759 12971
rect 11701 12931 11759 12937
rect 13078 12928 13084 12980
rect 13136 12968 13142 12980
rect 13357 12971 13415 12977
rect 13357 12968 13369 12971
rect 13136 12940 13369 12968
rect 13136 12928 13142 12940
rect 13357 12937 13369 12940
rect 13403 12937 13415 12971
rect 13722 12968 13728 12980
rect 13683 12940 13728 12968
rect 13357 12931 13415 12937
rect 13722 12928 13728 12940
rect 13780 12928 13786 12980
rect 13814 12928 13820 12980
rect 13872 12968 13878 12980
rect 14458 12968 14464 12980
rect 13872 12940 14464 12968
rect 13872 12928 13878 12940
rect 14458 12928 14464 12940
rect 14516 12968 14522 12980
rect 14645 12971 14703 12977
rect 14645 12968 14657 12971
rect 14516 12940 14657 12968
rect 14516 12928 14522 12940
rect 14645 12937 14657 12940
rect 14691 12968 14703 12971
rect 14826 12968 14832 12980
rect 14691 12940 14832 12968
rect 14691 12937 14703 12940
rect 14645 12931 14703 12937
rect 14826 12928 14832 12940
rect 14884 12928 14890 12980
rect 15010 12928 15016 12980
rect 15068 12968 15074 12980
rect 15565 12971 15623 12977
rect 15565 12968 15577 12971
rect 15068 12940 15577 12968
rect 15068 12928 15074 12940
rect 15565 12937 15577 12940
rect 15611 12937 15623 12971
rect 15565 12931 15623 12937
rect 7552 12903 7610 12909
rect 7552 12869 7564 12903
rect 7598 12900 7610 12903
rect 9214 12900 9220 12912
rect 7598 12872 9220 12900
rect 7598 12869 7610 12872
rect 7552 12863 7610 12869
rect 9214 12860 9220 12872
rect 9272 12860 9278 12912
rect 10529 12872 11008 12900
rect 7285 12835 7343 12841
rect 7285 12801 7297 12835
rect 7331 12801 7343 12835
rect 10529 12832 10557 12872
rect 7285 12795 7343 12801
rect 7372 12804 10557 12832
rect 10617 12835 10675 12841
rect 7372 12764 7400 12804
rect 10617 12801 10629 12835
rect 10663 12832 10675 12835
rect 10778 12832 10784 12844
rect 10663 12804 10784 12832
rect 10663 12801 10675 12804
rect 10617 12795 10675 12801
rect 10778 12792 10784 12804
rect 10836 12792 10842 12844
rect 5920 12736 7400 12764
rect 8294 12724 8300 12776
rect 8352 12764 8358 12776
rect 9214 12764 9220 12776
rect 8352 12736 9220 12764
rect 8352 12724 8358 12736
rect 9214 12724 9220 12736
rect 9272 12724 9278 12776
rect 9674 12764 9680 12776
rect 9324 12736 9680 12764
rect 6914 12696 6920 12708
rect 3804 12668 4384 12696
rect 5828 12668 6920 12696
rect 3804 12640 3832 12668
rect 1486 12628 1492 12640
rect 1447 12600 1492 12628
rect 1486 12588 1492 12600
rect 1544 12588 1550 12640
rect 1670 12588 1676 12640
rect 1728 12628 1734 12640
rect 1765 12631 1823 12637
rect 1765 12628 1777 12631
rect 1728 12600 1777 12628
rect 1728 12588 1734 12600
rect 1765 12597 1777 12600
rect 1811 12597 1823 12631
rect 1765 12591 1823 12597
rect 3786 12588 3792 12640
rect 3844 12588 3850 12640
rect 4246 12628 4252 12640
rect 4207 12600 4252 12628
rect 4246 12588 4252 12600
rect 4304 12588 4310 12640
rect 4356 12628 4384 12668
rect 6914 12656 6920 12668
rect 6972 12656 6978 12708
rect 9324 12696 9352 12736
rect 9674 12724 9680 12736
rect 9732 12724 9738 12776
rect 10873 12767 10931 12773
rect 10873 12733 10885 12767
rect 10919 12733 10931 12767
rect 10980 12764 11008 12872
rect 11054 12860 11060 12912
rect 11112 12900 11118 12912
rect 11514 12900 11520 12912
rect 11112 12872 11520 12900
rect 11112 12860 11118 12872
rect 11514 12860 11520 12872
rect 11572 12860 11578 12912
rect 11790 12860 11796 12912
rect 11848 12900 11854 12912
rect 12345 12903 12403 12909
rect 12345 12900 12357 12903
rect 11848 12872 12357 12900
rect 11848 12860 11854 12872
rect 12345 12869 12357 12872
rect 12391 12900 12403 12903
rect 12805 12903 12863 12909
rect 12805 12900 12817 12903
rect 12391 12872 12817 12900
rect 12391 12869 12403 12872
rect 12345 12863 12403 12869
rect 12805 12869 12817 12872
rect 12851 12869 12863 12903
rect 12805 12863 12863 12869
rect 12897 12903 12955 12909
rect 12897 12869 12909 12903
rect 12943 12900 12955 12903
rect 13262 12900 13268 12912
rect 12943 12872 13268 12900
rect 12943 12869 12955 12872
rect 12897 12863 12955 12869
rect 13262 12860 13268 12872
rect 13320 12900 13326 12912
rect 13446 12900 13452 12912
rect 13320 12872 13452 12900
rect 13320 12860 13326 12872
rect 13446 12860 13452 12872
rect 13504 12860 13510 12912
rect 14844 12900 14872 12928
rect 15105 12903 15163 12909
rect 15105 12900 15117 12903
rect 14844 12872 15117 12900
rect 15105 12869 15117 12872
rect 15151 12869 15163 12903
rect 15654 12900 15660 12912
rect 15105 12863 15163 12869
rect 15212 12872 15660 12900
rect 13170 12792 13176 12844
rect 13228 12832 13234 12844
rect 14553 12835 14611 12841
rect 14553 12832 14565 12835
rect 13228 12804 14565 12832
rect 13228 12792 13234 12804
rect 14553 12801 14565 12804
rect 14599 12832 14611 12835
rect 15212 12832 15240 12872
rect 15654 12860 15660 12872
rect 15712 12860 15718 12912
rect 14599 12804 15240 12832
rect 15473 12835 15531 12841
rect 14599 12801 14611 12804
rect 14553 12795 14611 12801
rect 15473 12801 15485 12835
rect 15519 12801 15531 12835
rect 15473 12795 15531 12801
rect 12621 12767 12679 12773
rect 12621 12764 12633 12767
rect 10980 12736 12633 12764
rect 10873 12727 10931 12733
rect 12621 12733 12633 12736
rect 12667 12764 12679 12767
rect 13354 12764 13360 12776
rect 12667 12736 13360 12764
rect 12667 12733 12679 12736
rect 12621 12727 12679 12733
rect 8220 12668 9352 12696
rect 8220 12628 8248 12668
rect 8662 12628 8668 12640
rect 4356 12600 8248 12628
rect 8623 12600 8668 12628
rect 8662 12588 8668 12600
rect 8720 12588 8726 12640
rect 9493 12631 9551 12637
rect 9493 12597 9505 12631
rect 9539 12628 9551 12631
rect 9674 12628 9680 12640
rect 9539 12600 9680 12628
rect 9539 12597 9551 12600
rect 9493 12591 9551 12597
rect 9674 12588 9680 12600
rect 9732 12588 9738 12640
rect 10686 12588 10692 12640
rect 10744 12628 10750 12640
rect 10888 12628 10916 12727
rect 13354 12724 13360 12736
rect 13412 12724 13418 12776
rect 13538 12724 13544 12776
rect 13596 12764 13602 12776
rect 13817 12767 13875 12773
rect 13817 12764 13829 12767
rect 13596 12736 13829 12764
rect 13596 12724 13602 12736
rect 13817 12733 13829 12736
rect 13863 12733 13875 12767
rect 13998 12764 14004 12776
rect 13959 12736 14004 12764
rect 13817 12727 13875 12733
rect 13998 12724 14004 12736
rect 14056 12724 14062 12776
rect 14642 12724 14648 12776
rect 14700 12764 14706 12776
rect 14737 12767 14795 12773
rect 14737 12764 14749 12767
rect 14700 12736 14749 12764
rect 14700 12724 14706 12736
rect 14737 12733 14749 12736
rect 14783 12733 14795 12767
rect 15488 12764 15516 12795
rect 15654 12764 15660 12776
rect 15488 12736 15660 12764
rect 14737 12727 14795 12733
rect 15654 12724 15660 12736
rect 15712 12764 15718 12776
rect 16114 12764 16120 12776
rect 15712 12736 16120 12764
rect 15712 12724 15718 12736
rect 16114 12724 16120 12736
rect 16172 12724 16178 12776
rect 11238 12656 11244 12708
rect 11296 12696 11302 12708
rect 14185 12699 14243 12705
rect 14185 12696 14197 12699
rect 11296 12668 14197 12696
rect 11296 12656 11302 12668
rect 14185 12665 14197 12668
rect 14231 12665 14243 12699
rect 14185 12659 14243 12665
rect 14826 12656 14832 12708
rect 14884 12696 14890 12708
rect 15289 12699 15347 12705
rect 15289 12696 15301 12699
rect 14884 12668 15301 12696
rect 14884 12656 14890 12668
rect 15289 12665 15301 12668
rect 15335 12665 15347 12699
rect 15289 12659 15347 12665
rect 13262 12628 13268 12640
rect 10744 12600 10916 12628
rect 13223 12600 13268 12628
rect 10744 12588 10750 12600
rect 13262 12588 13268 12600
rect 13320 12588 13326 12640
rect 15194 12588 15200 12640
rect 15252 12628 15258 12640
rect 15562 12628 15568 12640
rect 15252 12600 15568 12628
rect 15252 12588 15258 12600
rect 15562 12588 15568 12600
rect 15620 12588 15626 12640
rect 1104 12538 16008 12560
rect 1104 12486 2824 12538
rect 2876 12486 2888 12538
rect 2940 12486 2952 12538
rect 3004 12486 3016 12538
rect 3068 12486 3080 12538
rect 3132 12486 6572 12538
rect 6624 12486 6636 12538
rect 6688 12486 6700 12538
rect 6752 12486 6764 12538
rect 6816 12486 6828 12538
rect 6880 12486 10320 12538
rect 10372 12486 10384 12538
rect 10436 12486 10448 12538
rect 10500 12486 10512 12538
rect 10564 12486 10576 12538
rect 10628 12486 14068 12538
rect 14120 12486 14132 12538
rect 14184 12486 14196 12538
rect 14248 12486 14260 12538
rect 14312 12486 14324 12538
rect 14376 12486 16008 12538
rect 1104 12464 16008 12486
rect 1946 12384 1952 12436
rect 2004 12424 2010 12436
rect 2133 12427 2191 12433
rect 2133 12424 2145 12427
rect 2004 12396 2145 12424
rect 2004 12384 2010 12396
rect 2133 12393 2145 12396
rect 2179 12393 2191 12427
rect 2590 12424 2596 12436
rect 2133 12387 2191 12393
rect 2240 12396 2596 12424
rect 2240 12297 2268 12396
rect 2590 12384 2596 12396
rect 2648 12424 2654 12436
rect 3142 12424 3148 12436
rect 2648 12396 3148 12424
rect 2648 12384 2654 12396
rect 3142 12384 3148 12396
rect 3200 12384 3206 12436
rect 3234 12384 3240 12436
rect 3292 12424 3298 12436
rect 3418 12424 3424 12436
rect 3292 12396 3424 12424
rect 3292 12384 3298 12396
rect 3418 12384 3424 12396
rect 3476 12384 3482 12436
rect 4522 12384 4528 12436
rect 4580 12424 4586 12436
rect 4893 12427 4951 12433
rect 4893 12424 4905 12427
rect 4580 12396 4905 12424
rect 4580 12384 4586 12396
rect 4893 12393 4905 12396
rect 4939 12393 4951 12427
rect 6914 12424 6920 12436
rect 4893 12387 4951 12393
rect 5000 12396 6920 12424
rect 3160 12356 3188 12384
rect 3789 12359 3847 12365
rect 3789 12356 3801 12359
rect 3160 12328 3801 12356
rect 3789 12325 3801 12328
rect 3835 12356 3847 12359
rect 3878 12356 3884 12368
rect 3835 12328 3884 12356
rect 3835 12325 3847 12328
rect 3789 12319 3847 12325
rect 3878 12316 3884 12328
rect 3936 12356 3942 12368
rect 4249 12359 4307 12365
rect 4249 12356 4261 12359
rect 3936 12328 4261 12356
rect 3936 12316 3942 12328
rect 4249 12325 4261 12328
rect 4295 12325 4307 12359
rect 4249 12319 4307 12325
rect 1581 12291 1639 12297
rect 1581 12257 1593 12291
rect 1627 12288 1639 12291
rect 2225 12291 2283 12297
rect 1627 12260 2176 12288
rect 1627 12257 1639 12260
rect 1581 12251 1639 12257
rect 1762 12220 1768 12232
rect 1723 12192 1768 12220
rect 1762 12180 1768 12192
rect 1820 12180 1826 12232
rect 2148 12220 2176 12260
rect 2225 12257 2237 12291
rect 2271 12257 2283 12291
rect 4264 12288 4292 12319
rect 4338 12316 4344 12368
rect 4396 12356 4402 12368
rect 5000 12356 5028 12396
rect 6914 12384 6920 12396
rect 6972 12424 6978 12436
rect 7190 12424 7196 12436
rect 6972 12396 7196 12424
rect 6972 12384 6978 12396
rect 7190 12384 7196 12396
rect 7248 12384 7254 12436
rect 7282 12384 7288 12436
rect 7340 12424 7346 12436
rect 7558 12424 7564 12436
rect 7340 12396 7564 12424
rect 7340 12384 7346 12396
rect 7558 12384 7564 12396
rect 7616 12384 7622 12436
rect 8757 12427 8815 12433
rect 8757 12393 8769 12427
rect 8803 12424 8815 12427
rect 9214 12424 9220 12436
rect 8803 12396 9220 12424
rect 8803 12393 8815 12396
rect 8757 12387 8815 12393
rect 9214 12384 9220 12396
rect 9272 12384 9278 12436
rect 10042 12384 10048 12436
rect 10100 12424 10106 12436
rect 12986 12424 12992 12436
rect 10100 12396 12992 12424
rect 10100 12384 10106 12396
rect 12986 12384 12992 12396
rect 13044 12384 13050 12436
rect 13541 12427 13599 12433
rect 13541 12393 13553 12427
rect 13587 12424 13599 12427
rect 13630 12424 13636 12436
rect 13587 12396 13636 12424
rect 13587 12393 13599 12396
rect 13541 12387 13599 12393
rect 13630 12384 13636 12396
rect 13688 12384 13694 12436
rect 13906 12384 13912 12436
rect 13964 12424 13970 12436
rect 14093 12427 14151 12433
rect 14093 12424 14105 12427
rect 13964 12396 14105 12424
rect 13964 12384 13970 12396
rect 14093 12393 14105 12396
rect 14139 12393 14151 12427
rect 14093 12387 14151 12393
rect 4396 12328 5028 12356
rect 4396 12316 4402 12328
rect 9030 12316 9036 12368
rect 9088 12356 9094 12368
rect 9490 12356 9496 12368
rect 9088 12328 9496 12356
rect 9088 12316 9094 12328
rect 9490 12316 9496 12328
rect 9548 12356 9554 12368
rect 13817 12359 13875 12365
rect 13817 12356 13829 12359
rect 9548 12328 13829 12356
rect 9548 12316 9554 12328
rect 13817 12325 13829 12328
rect 13863 12356 13875 12359
rect 14182 12356 14188 12368
rect 13863 12328 14188 12356
rect 13863 12325 13875 12328
rect 13817 12319 13875 12325
rect 14182 12316 14188 12328
rect 14240 12316 14246 12368
rect 14550 12356 14556 12368
rect 14463 12328 14556 12356
rect 4617 12291 4675 12297
rect 4617 12288 4629 12291
rect 4264 12260 4629 12288
rect 2225 12251 2283 12257
rect 4617 12257 4629 12260
rect 4663 12257 4675 12291
rect 4617 12251 4675 12257
rect 9950 12248 9956 12300
rect 10008 12288 10014 12300
rect 10870 12288 10876 12300
rect 10008 12260 10876 12288
rect 10008 12248 10014 12260
rect 10870 12248 10876 12260
rect 10928 12288 10934 12300
rect 12618 12288 12624 12300
rect 10928 12260 12624 12288
rect 10928 12248 10934 12260
rect 12618 12248 12624 12260
rect 12676 12248 12682 12300
rect 12897 12291 12955 12297
rect 12897 12257 12909 12291
rect 12943 12257 12955 12291
rect 12897 12251 12955 12257
rect 2148 12192 2774 12220
rect 1854 12112 1860 12164
rect 1912 12152 1918 12164
rect 2470 12155 2528 12161
rect 2470 12152 2482 12155
rect 1912 12124 2482 12152
rect 1912 12112 1918 12124
rect 2470 12121 2482 12124
rect 2516 12121 2528 12155
rect 2746 12152 2774 12192
rect 5718 12180 5724 12232
rect 5776 12220 5782 12232
rect 6273 12223 6331 12229
rect 6273 12220 6285 12223
rect 5776 12192 6285 12220
rect 5776 12180 5782 12192
rect 6273 12189 6285 12192
rect 6319 12220 6331 12223
rect 7193 12223 7251 12229
rect 7193 12220 7205 12223
rect 6319 12192 7205 12220
rect 6319 12189 6331 12192
rect 6273 12183 6331 12189
rect 7193 12189 7205 12192
rect 7239 12220 7251 12223
rect 7377 12223 7435 12229
rect 7377 12220 7389 12223
rect 7239 12192 7389 12220
rect 7239 12189 7251 12192
rect 7193 12183 7251 12189
rect 7377 12189 7389 12192
rect 7423 12189 7435 12223
rect 7377 12183 7435 12189
rect 7644 12223 7702 12229
rect 7644 12189 7656 12223
rect 7690 12220 7702 12223
rect 8662 12220 8668 12232
rect 7690 12192 8668 12220
rect 7690 12189 7702 12192
rect 7644 12183 7702 12189
rect 8662 12180 8668 12192
rect 8720 12220 8726 12232
rect 12912 12220 12940 12251
rect 13354 12248 13360 12300
rect 13412 12288 13418 12300
rect 14476 12288 14504 12328
rect 14550 12316 14556 12328
rect 14608 12356 14614 12368
rect 14608 12328 15056 12356
rect 14608 12316 14614 12328
rect 14642 12288 14648 12300
rect 13412 12260 14504 12288
rect 14603 12260 14648 12288
rect 13412 12248 13418 12260
rect 14642 12248 14648 12260
rect 14700 12248 14706 12300
rect 15028 12297 15056 12328
rect 15013 12291 15071 12297
rect 15013 12257 15025 12291
rect 15059 12257 15071 12291
rect 15013 12251 15071 12257
rect 13906 12220 13912 12232
rect 8720 12192 13912 12220
rect 8720 12180 8726 12192
rect 13906 12180 13912 12192
rect 13964 12180 13970 12232
rect 14553 12223 14611 12229
rect 14553 12189 14565 12223
rect 14599 12220 14611 12223
rect 14734 12220 14740 12232
rect 14599 12192 14740 12220
rect 14599 12189 14611 12192
rect 14553 12183 14611 12189
rect 14734 12180 14740 12192
rect 14792 12180 14798 12232
rect 15289 12223 15347 12229
rect 15289 12189 15301 12223
rect 15335 12220 15347 12223
rect 15654 12220 15660 12232
rect 15335 12192 15660 12220
rect 15335 12189 15347 12192
rect 15289 12183 15347 12189
rect 15654 12180 15660 12192
rect 15712 12180 15718 12232
rect 5442 12152 5448 12164
rect 2746 12124 5448 12152
rect 2470 12115 2528 12121
rect 5442 12112 5448 12124
rect 5500 12112 5506 12164
rect 5810 12112 5816 12164
rect 5868 12152 5874 12164
rect 6006 12155 6064 12161
rect 6006 12152 6018 12155
rect 5868 12124 6018 12152
rect 5868 12112 5874 12124
rect 6006 12121 6018 12124
rect 6052 12121 6064 12155
rect 6006 12115 6064 12121
rect 9490 12112 9496 12164
rect 9548 12152 9554 12164
rect 12066 12152 12072 12164
rect 9548 12124 12072 12152
rect 9548 12112 9554 12124
rect 12066 12112 12072 12124
rect 12124 12112 12130 12164
rect 12618 12112 12624 12164
rect 12676 12152 12682 12164
rect 13081 12155 13139 12161
rect 13081 12152 13093 12155
rect 12676 12124 13093 12152
rect 12676 12112 12682 12124
rect 13081 12121 13093 12124
rect 13127 12121 13139 12155
rect 13081 12115 13139 12121
rect 13173 12155 13231 12161
rect 13173 12121 13185 12155
rect 13219 12152 13231 12155
rect 13725 12155 13783 12161
rect 13725 12152 13737 12155
rect 13219 12124 13737 12152
rect 13219 12121 13231 12124
rect 13173 12115 13231 12121
rect 13725 12121 13737 12124
rect 13771 12152 13783 12155
rect 13814 12152 13820 12164
rect 13771 12124 13820 12152
rect 13771 12121 13783 12124
rect 13725 12115 13783 12121
rect 13814 12112 13820 12124
rect 13872 12112 13878 12164
rect 1673 12087 1731 12093
rect 1673 12053 1685 12087
rect 1719 12084 1731 12087
rect 2130 12084 2136 12096
rect 1719 12056 2136 12084
rect 1719 12053 1731 12056
rect 1673 12047 1731 12053
rect 2130 12044 2136 12056
rect 2188 12044 2194 12096
rect 3605 12087 3663 12093
rect 3605 12053 3617 12087
rect 3651 12084 3663 12087
rect 3970 12084 3976 12096
rect 3651 12056 3976 12084
rect 3651 12053 3663 12056
rect 3605 12047 3663 12053
rect 3970 12044 3976 12056
rect 4028 12044 4034 12096
rect 4430 12084 4436 12096
rect 4391 12056 4436 12084
rect 4430 12044 4436 12056
rect 4488 12044 4494 12096
rect 5534 12044 5540 12096
rect 5592 12084 5598 12096
rect 11238 12084 11244 12096
rect 5592 12056 11244 12084
rect 5592 12044 5598 12056
rect 11238 12044 11244 12056
rect 11296 12044 11302 12096
rect 14458 12084 14464 12096
rect 14419 12056 14464 12084
rect 14458 12044 14464 12056
rect 14516 12084 14522 12096
rect 15197 12087 15255 12093
rect 15197 12084 15209 12087
rect 14516 12056 15209 12084
rect 14516 12044 14522 12056
rect 15197 12053 15209 12056
rect 15243 12053 15255 12087
rect 15654 12084 15660 12096
rect 15615 12056 15660 12084
rect 15197 12047 15255 12053
rect 15654 12044 15660 12056
rect 15712 12044 15718 12096
rect 1104 11994 16008 12016
rect 1104 11942 4698 11994
rect 4750 11942 4762 11994
rect 4814 11942 4826 11994
rect 4878 11942 4890 11994
rect 4942 11942 4954 11994
rect 5006 11942 8446 11994
rect 8498 11942 8510 11994
rect 8562 11942 8574 11994
rect 8626 11942 8638 11994
rect 8690 11942 8702 11994
rect 8754 11942 12194 11994
rect 12246 11942 12258 11994
rect 12310 11942 12322 11994
rect 12374 11942 12386 11994
rect 12438 11942 12450 11994
rect 12502 11942 16008 11994
rect 1104 11920 16008 11942
rect 5718 11840 5724 11892
rect 5776 11880 5782 11892
rect 6089 11883 6147 11889
rect 6089 11880 6101 11883
rect 5776 11852 6101 11880
rect 5776 11840 5782 11852
rect 6089 11849 6101 11852
rect 6135 11849 6147 11883
rect 6089 11843 6147 11849
rect 4448 11784 6049 11812
rect 1670 11744 1676 11756
rect 1631 11716 1676 11744
rect 1670 11704 1676 11716
rect 1728 11704 1734 11756
rect 2952 11747 3010 11753
rect 2952 11713 2964 11747
rect 2998 11744 3010 11747
rect 4448 11744 4476 11784
rect 2998 11716 4476 11744
rect 4516 11747 4574 11753
rect 2998 11713 3010 11716
rect 2952 11707 3010 11713
rect 4516 11713 4528 11747
rect 4562 11744 4574 11747
rect 5258 11744 5264 11756
rect 4562 11716 5264 11744
rect 4562 11713 4574 11716
rect 4516 11707 4574 11713
rect 5258 11704 5264 11716
rect 5316 11704 5322 11756
rect 2590 11636 2596 11688
rect 2648 11676 2654 11688
rect 2685 11679 2743 11685
rect 2685 11676 2697 11679
rect 2648 11648 2697 11676
rect 2648 11636 2654 11648
rect 2685 11645 2697 11648
rect 2731 11645 2743 11679
rect 2685 11639 2743 11645
rect 3878 11636 3884 11688
rect 3936 11676 3942 11688
rect 4249 11679 4307 11685
rect 4249 11676 4261 11679
rect 3936 11648 4261 11676
rect 3936 11636 3942 11648
rect 4249 11645 4261 11648
rect 4295 11645 4307 11679
rect 6021 11676 6049 11784
rect 6104 11744 6132 11843
rect 7006 11840 7012 11892
rect 7064 11880 7070 11892
rect 7929 11883 7987 11889
rect 7929 11880 7941 11883
rect 7064 11852 7941 11880
rect 7064 11840 7070 11852
rect 7929 11849 7941 11852
rect 7975 11849 7987 11883
rect 9674 11880 9680 11892
rect 7929 11843 7987 11849
rect 8266 11852 9680 11880
rect 6632 11815 6690 11821
rect 6632 11781 6644 11815
rect 6678 11812 6690 11815
rect 8266 11812 8294 11852
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 10318 11840 10324 11892
rect 10376 11880 10382 11892
rect 11514 11880 11520 11892
rect 10376 11852 10824 11880
rect 11475 11852 11520 11880
rect 10376 11840 10382 11852
rect 6678 11784 8294 11812
rect 6678 11781 6690 11784
rect 6632 11775 6690 11781
rect 9214 11772 9220 11824
rect 9272 11812 9278 11824
rect 9493 11815 9551 11821
rect 9493 11812 9505 11815
rect 9272 11784 9505 11812
rect 9272 11772 9278 11784
rect 9493 11781 9505 11784
rect 9539 11812 9551 11815
rect 9858 11812 9864 11824
rect 9539 11784 9864 11812
rect 9539 11781 9551 11784
rect 9493 11775 9551 11781
rect 9858 11772 9864 11784
rect 9916 11812 9922 11824
rect 10502 11812 10508 11824
rect 9916 11784 10508 11812
rect 9916 11772 9922 11784
rect 10502 11772 10508 11784
rect 10560 11772 10566 11824
rect 10698 11815 10756 11821
rect 10698 11781 10710 11815
rect 10744 11812 10756 11815
rect 10796 11812 10824 11852
rect 11514 11840 11520 11852
rect 11572 11840 11578 11892
rect 11974 11880 11980 11892
rect 11935 11852 11980 11880
rect 11974 11840 11980 11852
rect 12032 11840 12038 11892
rect 14182 11880 14188 11892
rect 14143 11852 14188 11880
rect 14182 11840 14188 11852
rect 14240 11840 14246 11892
rect 15470 11880 15476 11892
rect 15431 11852 15476 11880
rect 15470 11840 15476 11852
rect 15528 11840 15534 11892
rect 15657 11883 15715 11889
rect 15657 11849 15669 11883
rect 15703 11880 15715 11883
rect 16022 11880 16028 11892
rect 15703 11852 16028 11880
rect 15703 11849 15715 11852
rect 15657 11843 15715 11849
rect 16022 11840 16028 11852
rect 16080 11840 16086 11892
rect 10744 11784 10824 11812
rect 10744 11781 10756 11784
rect 10698 11775 10756 11781
rect 10870 11772 10876 11824
rect 10928 11812 10934 11824
rect 10928 11784 11008 11812
rect 10928 11772 10934 11784
rect 6362 11744 6368 11756
rect 6104 11716 6368 11744
rect 6362 11704 6368 11716
rect 6420 11704 6426 11756
rect 6472 11716 7420 11744
rect 6472 11676 6500 11716
rect 6021 11648 6500 11676
rect 7392 11676 7420 11716
rect 7466 11704 7472 11756
rect 7524 11744 7530 11756
rect 10980 11753 11008 11784
rect 11330 11772 11336 11824
rect 11388 11812 11394 11824
rect 12250 11812 12256 11824
rect 11388 11784 12256 11812
rect 11388 11772 11394 11784
rect 12250 11772 12256 11784
rect 12308 11812 12314 11824
rect 12308 11784 12434 11812
rect 12308 11772 12314 11784
rect 10965 11747 11023 11753
rect 7524 11716 10916 11744
rect 7524 11704 7530 11716
rect 9490 11676 9496 11688
rect 7392 11648 9496 11676
rect 4249 11639 4307 11645
rect 9490 11636 9496 11648
rect 9548 11636 9554 11688
rect 10888 11676 10916 11716
rect 10965 11713 10977 11747
rect 11011 11713 11023 11747
rect 10965 11707 11023 11713
rect 11885 11747 11943 11753
rect 11885 11713 11897 11747
rect 11931 11744 11943 11747
rect 11974 11744 11980 11756
rect 11931 11716 11980 11744
rect 11931 11713 11943 11716
rect 11885 11707 11943 11713
rect 11974 11704 11980 11716
rect 12032 11704 12038 11756
rect 12406 11744 12434 11784
rect 13262 11772 13268 11824
rect 13320 11812 13326 11824
rect 14829 11815 14887 11821
rect 14829 11812 14841 11815
rect 13320 11784 14841 11812
rect 13320 11772 13326 11784
rect 14829 11781 14841 11784
rect 14875 11781 14887 11815
rect 14829 11775 14887 11781
rect 12805 11747 12863 11753
rect 12805 11744 12817 11747
rect 12406 11716 12817 11744
rect 12805 11713 12817 11716
rect 12851 11713 12863 11747
rect 12805 11707 12863 11713
rect 12986 11704 12992 11756
rect 13044 11744 13050 11756
rect 14093 11747 14151 11753
rect 14093 11744 14105 11747
rect 13044 11716 14105 11744
rect 13044 11704 13050 11716
rect 14093 11713 14105 11716
rect 14139 11713 14151 11747
rect 14093 11707 14151 11713
rect 14642 11704 14648 11756
rect 14700 11744 14706 11756
rect 14921 11747 14979 11753
rect 14921 11744 14933 11747
rect 14700 11716 14933 11744
rect 14700 11704 14706 11716
rect 14921 11713 14933 11716
rect 14967 11713 14979 11747
rect 14921 11707 14979 11713
rect 12069 11679 12127 11685
rect 12069 11676 12081 11679
rect 10888 11648 12081 11676
rect 12069 11645 12081 11648
rect 12115 11645 12127 11679
rect 12342 11676 12348 11688
rect 12303 11648 12348 11676
rect 12069 11639 12127 11645
rect 12342 11636 12348 11648
rect 12400 11636 12406 11688
rect 13081 11679 13139 11685
rect 13081 11645 13093 11679
rect 13127 11645 13139 11679
rect 14277 11679 14335 11685
rect 14277 11676 14289 11679
rect 13081 11639 13139 11645
rect 13188 11648 14289 11676
rect 7834 11608 7840 11620
rect 5184 11580 6408 11608
rect 1486 11540 1492 11552
rect 1447 11512 1492 11540
rect 1486 11500 1492 11512
rect 1544 11500 1550 11552
rect 4065 11543 4123 11549
rect 4065 11509 4077 11543
rect 4111 11540 4123 11543
rect 4154 11540 4160 11552
rect 4111 11512 4160 11540
rect 4111 11509 4123 11512
rect 4065 11503 4123 11509
rect 4154 11500 4160 11512
rect 4212 11500 4218 11552
rect 4614 11500 4620 11552
rect 4672 11540 4678 11552
rect 5184 11540 5212 11580
rect 5626 11540 5632 11552
rect 4672 11512 5212 11540
rect 5587 11512 5632 11540
rect 4672 11500 4678 11512
rect 5626 11500 5632 11512
rect 5684 11500 5690 11552
rect 6380 11540 6408 11580
rect 7300 11580 7840 11608
rect 7300 11552 7328 11580
rect 7834 11568 7840 11580
rect 7892 11568 7898 11620
rect 11514 11568 11520 11620
rect 11572 11608 11578 11620
rect 13096 11608 13124 11639
rect 11572 11580 13124 11608
rect 11572 11568 11578 11580
rect 7282 11540 7288 11552
rect 6380 11512 7288 11540
rect 7282 11500 7288 11512
rect 7340 11500 7346 11552
rect 7558 11500 7564 11552
rect 7616 11540 7622 11552
rect 7745 11543 7803 11549
rect 7745 11540 7757 11543
rect 7616 11512 7757 11540
rect 7616 11500 7622 11512
rect 7745 11509 7757 11512
rect 7791 11509 7803 11543
rect 7745 11503 7803 11509
rect 9585 11543 9643 11549
rect 9585 11509 9597 11543
rect 9631 11540 9643 11543
rect 10778 11540 10784 11552
rect 9631 11512 10784 11540
rect 9631 11509 9643 11512
rect 9585 11503 9643 11509
rect 10778 11500 10784 11512
rect 10836 11500 10842 11552
rect 12066 11500 12072 11552
rect 12124 11540 12130 11552
rect 13188 11540 13216 11648
rect 14277 11645 14289 11648
rect 14323 11645 14335 11679
rect 14734 11676 14740 11688
rect 14695 11648 14740 11676
rect 14277 11639 14335 11645
rect 14734 11636 14740 11648
rect 14792 11636 14798 11688
rect 12124 11512 13216 11540
rect 12124 11500 12130 11512
rect 13630 11500 13636 11552
rect 13688 11540 13694 11552
rect 13725 11543 13783 11549
rect 13725 11540 13737 11543
rect 13688 11512 13737 11540
rect 13688 11500 13694 11512
rect 13725 11509 13737 11512
rect 13771 11509 13783 11543
rect 15286 11540 15292 11552
rect 15247 11512 15292 11540
rect 13725 11503 13783 11509
rect 15286 11500 15292 11512
rect 15344 11500 15350 11552
rect 1104 11450 16008 11472
rect 1104 11398 2824 11450
rect 2876 11398 2888 11450
rect 2940 11398 2952 11450
rect 3004 11398 3016 11450
rect 3068 11398 3080 11450
rect 3132 11398 6572 11450
rect 6624 11398 6636 11450
rect 6688 11398 6700 11450
rect 6752 11398 6764 11450
rect 6816 11398 6828 11450
rect 6880 11398 10320 11450
rect 10372 11398 10384 11450
rect 10436 11398 10448 11450
rect 10500 11398 10512 11450
rect 10564 11398 10576 11450
rect 10628 11398 14068 11450
rect 14120 11398 14132 11450
rect 14184 11398 14196 11450
rect 14248 11398 14260 11450
rect 14312 11398 14324 11450
rect 14376 11398 16008 11450
rect 1104 11376 16008 11398
rect 1489 11339 1547 11345
rect 1489 11305 1501 11339
rect 1535 11336 1547 11339
rect 1578 11336 1584 11348
rect 1535 11308 1584 11336
rect 1535 11305 1547 11308
rect 1489 11299 1547 11305
rect 1578 11296 1584 11308
rect 1636 11296 1642 11348
rect 2498 11336 2504 11348
rect 2148 11308 2504 11336
rect 2148 11209 2176 11308
rect 2498 11296 2504 11308
rect 2556 11296 2562 11348
rect 3878 11296 3884 11348
rect 3936 11336 3942 11348
rect 4065 11339 4123 11345
rect 4065 11336 4077 11339
rect 3936 11308 4077 11336
rect 3936 11296 3942 11308
rect 4065 11305 4077 11308
rect 4111 11336 4123 11339
rect 4249 11339 4307 11345
rect 4249 11336 4261 11339
rect 4111 11308 4261 11336
rect 4111 11305 4123 11308
rect 4065 11299 4123 11305
rect 4249 11305 4261 11308
rect 4295 11336 4307 11339
rect 4433 11339 4491 11345
rect 4433 11336 4445 11339
rect 4295 11308 4445 11336
rect 4295 11305 4307 11308
rect 4249 11299 4307 11305
rect 4433 11305 4445 11308
rect 4479 11336 4491 11339
rect 5629 11339 5687 11345
rect 5629 11336 5641 11339
rect 4479 11308 5641 11336
rect 4479 11305 4491 11308
rect 4433 11299 4491 11305
rect 5629 11305 5641 11308
rect 5675 11336 5687 11339
rect 7193 11339 7251 11345
rect 5675 11308 5856 11336
rect 5675 11305 5687 11308
rect 5629 11299 5687 11305
rect 3513 11271 3571 11277
rect 3513 11237 3525 11271
rect 3559 11268 3571 11271
rect 5534 11268 5540 11280
rect 3559 11240 5540 11268
rect 3559 11237 3571 11240
rect 3513 11231 3571 11237
rect 5534 11228 5540 11240
rect 5592 11228 5598 11280
rect 5828 11209 5856 11308
rect 7193 11305 7205 11339
rect 7239 11336 7251 11339
rect 10318 11336 10324 11348
rect 7239 11308 10324 11336
rect 7239 11305 7251 11308
rect 7193 11299 7251 11305
rect 10318 11296 10324 11308
rect 10376 11296 10382 11348
rect 11241 11339 11299 11345
rect 11241 11305 11253 11339
rect 11287 11336 11299 11339
rect 11422 11336 11428 11348
rect 11287 11308 11428 11336
rect 11287 11305 11299 11308
rect 11241 11299 11299 11305
rect 11422 11296 11428 11308
rect 11480 11296 11486 11348
rect 11882 11296 11888 11348
rect 11940 11336 11946 11348
rect 13173 11339 13231 11345
rect 13173 11336 13185 11339
rect 11940 11308 13185 11336
rect 11940 11296 11946 11308
rect 13173 11305 13185 11308
rect 13219 11305 13231 11339
rect 13173 11299 13231 11305
rect 13538 11296 13544 11348
rect 13596 11336 13602 11348
rect 14829 11339 14887 11345
rect 14829 11336 14841 11339
rect 13596 11308 14841 11336
rect 13596 11296 13602 11308
rect 14829 11305 14841 11308
rect 14875 11305 14887 11339
rect 14829 11299 14887 11305
rect 9033 11271 9091 11277
rect 9033 11237 9045 11271
rect 9079 11268 9091 11271
rect 9214 11268 9220 11280
rect 9079 11240 9220 11268
rect 9079 11237 9091 11240
rect 9033 11231 9091 11237
rect 2133 11203 2191 11209
rect 2133 11169 2145 11203
rect 2179 11169 2191 11203
rect 2133 11163 2191 11169
rect 5813 11203 5871 11209
rect 5813 11169 5825 11203
rect 5859 11169 5871 11203
rect 5813 11163 5871 11169
rect 1673 11135 1731 11141
rect 1673 11101 1685 11135
rect 1719 11132 1731 11135
rect 3234 11132 3240 11144
rect 1719 11104 3240 11132
rect 1719 11101 1731 11104
rect 1673 11095 1731 11101
rect 3234 11092 3240 11104
rect 3292 11092 3298 11144
rect 3973 11135 4031 11141
rect 3973 11101 3985 11135
rect 4019 11132 4031 11135
rect 4706 11132 4712 11144
rect 4019 11104 4712 11132
rect 4019 11101 4031 11104
rect 3973 11095 4031 11101
rect 2400 11067 2458 11073
rect 2400 11033 2412 11067
rect 2446 11064 2458 11067
rect 3988 11064 4016 11095
rect 4706 11092 4712 11104
rect 4764 11092 4770 11144
rect 6080 11135 6138 11141
rect 6080 11101 6092 11135
rect 6126 11132 6138 11135
rect 7006 11132 7012 11144
rect 6126 11104 7012 11132
rect 6126 11101 6138 11104
rect 6080 11095 6138 11101
rect 7006 11092 7012 11104
rect 7064 11092 7070 11144
rect 7374 11132 7380 11144
rect 7287 11104 7380 11132
rect 7374 11092 7380 11104
rect 7432 11132 7438 11144
rect 9048 11132 9076 11231
rect 9214 11228 9220 11240
rect 9272 11228 9278 11280
rect 12250 11228 12256 11280
rect 12308 11268 12314 11280
rect 13081 11271 13139 11277
rect 12308 11240 12756 11268
rect 12308 11228 12314 11240
rect 10686 11200 10692 11212
rect 10647 11172 10692 11200
rect 10686 11160 10692 11172
rect 10744 11160 10750 11212
rect 11882 11200 11888 11212
rect 11843 11172 11888 11200
rect 11882 11160 11888 11172
rect 11940 11160 11946 11212
rect 12066 11160 12072 11212
rect 12124 11200 12130 11212
rect 12437 11203 12495 11209
rect 12437 11200 12449 11203
rect 12124 11172 12449 11200
rect 12124 11160 12130 11172
rect 12437 11169 12449 11172
rect 12483 11169 12495 11203
rect 12437 11163 12495 11169
rect 7432 11104 9076 11132
rect 11609 11135 11667 11141
rect 7432 11092 7438 11104
rect 11609 11101 11621 11135
rect 11655 11132 11667 11135
rect 12342 11132 12348 11144
rect 11655 11104 12348 11132
rect 11655 11101 11667 11104
rect 11609 11095 11667 11101
rect 12342 11092 12348 11104
rect 12400 11092 12406 11144
rect 12728 11141 12756 11240
rect 13081 11237 13093 11271
rect 13127 11237 13139 11271
rect 13081 11231 13139 11237
rect 12713 11135 12771 11141
rect 12713 11101 12725 11135
rect 12759 11101 12771 11135
rect 13096 11132 13124 11231
rect 13354 11228 13360 11280
rect 13412 11268 13418 11280
rect 13412 11240 13768 11268
rect 13412 11228 13418 11240
rect 13630 11200 13636 11212
rect 13591 11172 13636 11200
rect 13630 11160 13636 11172
rect 13688 11160 13694 11212
rect 13740 11209 13768 11240
rect 13725 11203 13783 11209
rect 13725 11169 13737 11203
rect 13771 11169 13783 11203
rect 13725 11163 13783 11169
rect 13906 11160 13912 11212
rect 13964 11200 13970 11212
rect 15381 11203 15439 11209
rect 15381 11200 15393 11203
rect 13964 11172 15393 11200
rect 13964 11160 13970 11172
rect 15381 11169 15393 11172
rect 15427 11169 15439 11203
rect 15381 11163 15439 11169
rect 15746 11160 15752 11212
rect 15804 11160 15810 11212
rect 13541 11135 13599 11141
rect 13541 11132 13553 11135
rect 13096 11104 13553 11132
rect 12713 11095 12771 11101
rect 13541 11101 13553 11104
rect 13587 11101 13599 11135
rect 14366 11132 14372 11144
rect 14327 11104 14372 11132
rect 13541 11095 13599 11101
rect 14366 11092 14372 11104
rect 14424 11132 14430 11144
rect 14642 11132 14648 11144
rect 14424 11104 14648 11132
rect 14424 11092 14430 11104
rect 14642 11092 14648 11104
rect 14700 11092 14706 11144
rect 15197 11135 15255 11141
rect 15197 11101 15209 11135
rect 15243 11132 15255 11135
rect 15764 11132 15792 11160
rect 15243 11104 15884 11132
rect 15243 11101 15255 11104
rect 15197 11095 15255 11101
rect 7650 11073 7656 11076
rect 7644 11064 7656 11073
rect 2446 11036 4016 11064
rect 7611 11036 7656 11064
rect 2446 11033 2458 11036
rect 2400 11027 2458 11033
rect 7644 11027 7656 11036
rect 7650 11024 7656 11027
rect 7708 11024 7714 11076
rect 7834 11024 7840 11076
rect 7892 11064 7898 11076
rect 10444 11067 10502 11073
rect 7892 11036 9352 11064
rect 7892 11024 7898 11036
rect 1394 10956 1400 11008
rect 1452 10996 1458 11008
rect 2866 10996 2872 11008
rect 1452 10968 2872 10996
rect 1452 10956 1458 10968
rect 2866 10956 2872 10968
rect 2924 10996 2930 11008
rect 5258 10996 5264 11008
rect 2924 10968 5264 10996
rect 2924 10956 2930 10968
rect 5258 10956 5264 10968
rect 5316 10956 5322 11008
rect 8757 10999 8815 11005
rect 8757 10965 8769 10999
rect 8803 10996 8815 10999
rect 9214 10996 9220 11008
rect 8803 10968 9220 10996
rect 8803 10965 8815 10968
rect 8757 10959 8815 10965
rect 9214 10956 9220 10968
rect 9272 10956 9278 11008
rect 9324 11005 9352 11036
rect 10444 11033 10456 11067
rect 10490 11064 10502 11067
rect 10778 11064 10784 11076
rect 10490 11036 10784 11064
rect 10490 11033 10502 11036
rect 10444 11027 10502 11033
rect 10778 11024 10784 11036
rect 10836 11024 10842 11076
rect 11422 11024 11428 11076
rect 11480 11064 11486 11076
rect 12621 11067 12679 11073
rect 12621 11064 12633 11067
rect 11480 11036 12633 11064
rect 11480 11024 11486 11036
rect 12621 11033 12633 11036
rect 12667 11033 12679 11067
rect 12621 11027 12679 11033
rect 15289 11067 15347 11073
rect 15289 11033 15301 11067
rect 15335 11064 15347 11067
rect 15746 11064 15752 11076
rect 15335 11036 15752 11064
rect 15335 11033 15347 11036
rect 15289 11027 15347 11033
rect 15746 11024 15752 11036
rect 15804 11024 15810 11076
rect 15856 11008 15884 11104
rect 9309 10999 9367 11005
rect 9309 10965 9321 10999
rect 9355 10965 9367 10999
rect 9309 10959 9367 10965
rect 10226 10956 10232 11008
rect 10284 10996 10290 11008
rect 11701 10999 11759 11005
rect 11701 10996 11713 10999
rect 10284 10968 11713 10996
rect 10284 10956 10290 10968
rect 11701 10965 11713 10968
rect 11747 10996 11759 10999
rect 12161 10999 12219 11005
rect 12161 10996 12173 10999
rect 11747 10968 12173 10996
rect 11747 10965 11759 10968
rect 11701 10959 11759 10965
rect 12161 10965 12173 10968
rect 12207 10996 12219 10999
rect 14918 10996 14924 11008
rect 12207 10968 14924 10996
rect 12207 10965 12219 10968
rect 12161 10959 12219 10965
rect 14918 10956 14924 10968
rect 14976 10956 14982 11008
rect 15838 10956 15844 11008
rect 15896 10956 15902 11008
rect 1104 10906 16008 10928
rect 1104 10854 4698 10906
rect 4750 10854 4762 10906
rect 4814 10854 4826 10906
rect 4878 10854 4890 10906
rect 4942 10854 4954 10906
rect 5006 10854 8446 10906
rect 8498 10854 8510 10906
rect 8562 10854 8574 10906
rect 8626 10854 8638 10906
rect 8690 10854 8702 10906
rect 8754 10854 12194 10906
rect 12246 10854 12258 10906
rect 12310 10854 12322 10906
rect 12374 10854 12386 10906
rect 12438 10854 12450 10906
rect 12502 10854 16008 10906
rect 1104 10832 16008 10854
rect 1765 10795 1823 10801
rect 1765 10761 1777 10795
rect 1811 10792 1823 10795
rect 2225 10795 2283 10801
rect 2225 10792 2237 10795
rect 1811 10764 2237 10792
rect 1811 10761 1823 10764
rect 1765 10755 1823 10761
rect 2225 10761 2237 10764
rect 2271 10761 2283 10795
rect 3142 10792 3148 10804
rect 3055 10764 3148 10792
rect 2225 10755 2283 10761
rect 3142 10752 3148 10764
rect 3200 10792 3206 10804
rect 3694 10792 3700 10804
rect 3200 10764 3700 10792
rect 3200 10752 3206 10764
rect 3694 10752 3700 10764
rect 3752 10752 3758 10804
rect 3789 10795 3847 10801
rect 3789 10761 3801 10795
rect 3835 10792 3847 10795
rect 3878 10792 3884 10804
rect 3835 10764 3884 10792
rect 3835 10761 3847 10764
rect 3789 10755 3847 10761
rect 3878 10752 3884 10764
rect 3936 10752 3942 10804
rect 6362 10752 6368 10804
rect 6420 10792 6426 10804
rect 7009 10795 7067 10801
rect 7009 10792 7021 10795
rect 6420 10764 7021 10792
rect 6420 10752 6426 10764
rect 7009 10761 7021 10764
rect 7055 10792 7067 10795
rect 7374 10792 7380 10804
rect 7055 10764 7380 10792
rect 7055 10761 7067 10764
rect 7009 10755 7067 10761
rect 5626 10724 5632 10736
rect 1596 10696 5632 10724
rect 1596 10597 1624 10696
rect 5626 10684 5632 10696
rect 5684 10684 5690 10736
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 2038 10656 2044 10668
rect 1719 10628 2044 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 2038 10616 2044 10628
rect 2096 10616 2102 10668
rect 2593 10659 2651 10665
rect 2593 10625 2605 10659
rect 2639 10625 2651 10659
rect 3878 10656 3884 10668
rect 3839 10628 3884 10656
rect 2593 10619 2651 10625
rect 1581 10591 1639 10597
rect 1581 10557 1593 10591
rect 1627 10557 1639 10591
rect 1581 10551 1639 10557
rect 2130 10520 2136 10532
rect 2091 10492 2136 10520
rect 2130 10480 2136 10492
rect 2188 10480 2194 10532
rect 2608 10452 2636 10619
rect 3878 10616 3884 10628
rect 3936 10616 3942 10668
rect 4154 10665 4160 10668
rect 4148 10619 4160 10665
rect 4212 10656 4218 10668
rect 7116 10665 7144 10764
rect 7374 10752 7380 10764
rect 7432 10752 7438 10804
rect 13262 10792 13268 10804
rect 7484 10764 13268 10792
rect 7484 10724 7512 10764
rect 13262 10752 13268 10764
rect 13320 10752 13326 10804
rect 13449 10795 13507 10801
rect 13449 10761 13461 10795
rect 13495 10792 13507 10795
rect 14829 10795 14887 10801
rect 14829 10792 14841 10795
rect 13495 10764 14841 10792
rect 13495 10761 13507 10764
rect 13449 10755 13507 10761
rect 14829 10761 14841 10764
rect 14875 10761 14887 10795
rect 14829 10755 14887 10761
rect 15197 10795 15255 10801
rect 15197 10761 15209 10795
rect 15243 10792 15255 10795
rect 15286 10792 15292 10804
rect 15243 10764 15292 10792
rect 15243 10761 15255 10764
rect 15197 10755 15255 10761
rect 15286 10752 15292 10764
rect 15344 10752 15350 10804
rect 7208 10696 7512 10724
rect 9493 10727 9551 10733
rect 7101 10659 7159 10665
rect 4212 10628 4248 10656
rect 4154 10616 4160 10619
rect 4212 10616 4218 10628
rect 7101 10625 7113 10659
rect 7147 10625 7159 10659
rect 7101 10619 7159 10625
rect 2685 10591 2743 10597
rect 2685 10557 2697 10591
rect 2731 10557 2743 10591
rect 2866 10588 2872 10600
rect 2827 10560 2872 10588
rect 2685 10551 2743 10557
rect 2700 10520 2728 10551
rect 2866 10548 2872 10560
rect 2924 10548 2930 10600
rect 5718 10548 5724 10600
rect 5776 10588 5782 10600
rect 5994 10588 6000 10600
rect 5776 10560 6000 10588
rect 5776 10548 5782 10560
rect 5994 10548 6000 10560
rect 6052 10588 6058 10600
rect 7208 10588 7236 10696
rect 9493 10693 9505 10727
rect 9539 10724 9551 10727
rect 9858 10724 9864 10736
rect 9539 10696 9864 10724
rect 9539 10693 9551 10696
rect 9493 10687 9551 10693
rect 9858 10684 9864 10696
rect 9916 10724 9922 10736
rect 14458 10724 14464 10736
rect 9916 10696 11008 10724
rect 9916 10684 9922 10696
rect 7368 10659 7426 10665
rect 7368 10625 7380 10659
rect 7414 10656 7426 10659
rect 7742 10656 7748 10668
rect 7414 10628 7748 10656
rect 7414 10625 7426 10628
rect 7368 10619 7426 10625
rect 7742 10616 7748 10628
rect 7800 10616 7806 10668
rect 9214 10616 9220 10668
rect 9272 10656 9278 10668
rect 10980 10665 11008 10696
rect 12406 10696 13584 10724
rect 14371 10696 14464 10724
rect 10698 10659 10756 10665
rect 10698 10656 10710 10659
rect 9272 10628 10710 10656
rect 9272 10616 9278 10628
rect 10698 10625 10710 10628
rect 10744 10656 10756 10659
rect 10965 10659 11023 10665
rect 10744 10628 10916 10656
rect 10744 10625 10756 10628
rect 10698 10619 10756 10625
rect 6052 10560 7236 10588
rect 10888 10588 10916 10628
rect 10965 10625 10977 10659
rect 11011 10625 11023 10659
rect 10965 10619 11023 10625
rect 12406 10588 12434 10696
rect 13354 10656 13360 10668
rect 13315 10628 13360 10656
rect 13354 10616 13360 10628
rect 13412 10616 13418 10668
rect 12894 10588 12900 10600
rect 10888 10560 12434 10588
rect 12855 10560 12900 10588
rect 6052 10548 6058 10560
rect 12894 10548 12900 10560
rect 12952 10548 12958 10600
rect 13556 10597 13584 10696
rect 14458 10684 14464 10696
rect 14516 10724 14522 10736
rect 15010 10724 15016 10736
rect 14516 10696 15016 10724
rect 14516 10684 14522 10696
rect 15010 10684 15016 10696
rect 15068 10684 15074 10736
rect 14369 10659 14427 10665
rect 14369 10625 14381 10659
rect 14415 10656 14427 10659
rect 14826 10656 14832 10668
rect 14415 10628 14832 10656
rect 14415 10625 14427 10628
rect 14369 10619 14427 10625
rect 14826 10616 14832 10628
rect 14884 10616 14890 10668
rect 13541 10591 13599 10597
rect 13541 10557 13553 10591
rect 13587 10557 13599 10591
rect 13541 10551 13599 10557
rect 13906 10548 13912 10600
rect 13964 10588 13970 10600
rect 14553 10591 14611 10597
rect 14553 10588 14565 10591
rect 13964 10560 14565 10588
rect 13964 10548 13970 10560
rect 14553 10557 14565 10560
rect 14599 10557 14611 10591
rect 14553 10551 14611 10557
rect 14918 10548 14924 10600
rect 14976 10588 14982 10600
rect 15289 10591 15347 10597
rect 15289 10588 15301 10591
rect 14976 10560 15301 10588
rect 14976 10548 14982 10560
rect 15289 10557 15301 10560
rect 15335 10557 15347 10591
rect 15289 10551 15347 10557
rect 15381 10591 15439 10597
rect 15381 10557 15393 10591
rect 15427 10557 15439 10591
rect 15381 10551 15439 10557
rect 12986 10520 12992 10532
rect 2700 10492 3924 10520
rect 3142 10452 3148 10464
rect 2608 10424 3148 10452
rect 3142 10412 3148 10424
rect 3200 10412 3206 10464
rect 3896 10452 3924 10492
rect 8128 10492 10088 10520
rect 12947 10492 12992 10520
rect 4154 10452 4160 10464
rect 3896 10424 4160 10452
rect 4154 10412 4160 10424
rect 4212 10412 4218 10464
rect 5261 10455 5319 10461
rect 5261 10421 5273 10455
rect 5307 10452 5319 10455
rect 8128 10452 8156 10492
rect 5307 10424 8156 10452
rect 5307 10421 5319 10424
rect 5261 10415 5319 10421
rect 8202 10412 8208 10464
rect 8260 10452 8266 10464
rect 8481 10455 8539 10461
rect 8481 10452 8493 10455
rect 8260 10424 8493 10452
rect 8260 10412 8266 10424
rect 8481 10421 8493 10424
rect 8527 10421 8539 10455
rect 8481 10415 8539 10421
rect 9490 10412 9496 10464
rect 9548 10452 9554 10464
rect 9585 10455 9643 10461
rect 9585 10452 9597 10455
rect 9548 10424 9597 10452
rect 9548 10412 9554 10424
rect 9585 10421 9597 10424
rect 9631 10421 9643 10455
rect 10060 10452 10088 10492
rect 12986 10480 12992 10492
rect 13044 10480 13050 10532
rect 13722 10480 13728 10532
rect 13780 10520 13786 10532
rect 14001 10523 14059 10529
rect 14001 10520 14013 10523
rect 13780 10492 14013 10520
rect 13780 10480 13786 10492
rect 14001 10489 14013 10492
rect 14047 10489 14059 10523
rect 14001 10483 14059 10489
rect 14642 10480 14648 10532
rect 14700 10520 14706 10532
rect 15396 10520 15424 10551
rect 14700 10492 15424 10520
rect 14700 10480 14706 10492
rect 11146 10452 11152 10464
rect 10060 10424 11152 10452
rect 9585 10415 9643 10421
rect 11146 10412 11152 10424
rect 11204 10452 11210 10464
rect 11698 10452 11704 10464
rect 11204 10424 11704 10452
rect 11204 10412 11210 10424
rect 11698 10412 11704 10424
rect 11756 10412 11762 10464
rect 13262 10412 13268 10464
rect 13320 10452 13326 10464
rect 13538 10452 13544 10464
rect 13320 10424 13544 10452
rect 13320 10412 13326 10424
rect 13538 10412 13544 10424
rect 13596 10452 13602 10464
rect 14734 10452 14740 10464
rect 13596 10424 14740 10452
rect 13596 10412 13602 10424
rect 14734 10412 14740 10424
rect 14792 10452 14798 10464
rect 15470 10452 15476 10464
rect 14792 10424 15476 10452
rect 14792 10412 14798 10424
rect 15470 10412 15476 10424
rect 15528 10412 15534 10464
rect 1104 10362 16008 10384
rect 1104 10310 2824 10362
rect 2876 10310 2888 10362
rect 2940 10310 2952 10362
rect 3004 10310 3016 10362
rect 3068 10310 3080 10362
rect 3132 10310 6572 10362
rect 6624 10310 6636 10362
rect 6688 10310 6700 10362
rect 6752 10310 6764 10362
rect 6816 10310 6828 10362
rect 6880 10310 10320 10362
rect 10372 10310 10384 10362
rect 10436 10310 10448 10362
rect 10500 10310 10512 10362
rect 10564 10310 10576 10362
rect 10628 10310 14068 10362
rect 14120 10310 14132 10362
rect 14184 10310 14196 10362
rect 14248 10310 14260 10362
rect 14312 10310 14324 10362
rect 14376 10310 16008 10362
rect 1104 10288 16008 10310
rect 1486 10248 1492 10260
rect 1447 10220 1492 10248
rect 1486 10208 1492 10220
rect 1544 10208 1550 10260
rect 6917 10251 6975 10257
rect 6917 10217 6929 10251
rect 6963 10248 6975 10251
rect 7650 10248 7656 10260
rect 6963 10220 7656 10248
rect 6963 10217 6975 10220
rect 6917 10211 6975 10217
rect 7650 10208 7656 10220
rect 7708 10248 7714 10260
rect 10597 10251 10655 10257
rect 7708 10220 10557 10248
rect 7708 10208 7714 10220
rect 7377 10183 7435 10189
rect 7377 10149 7389 10183
rect 7423 10180 7435 10183
rect 7466 10180 7472 10192
rect 7423 10152 7472 10180
rect 7423 10149 7435 10152
rect 7377 10143 7435 10149
rect 7466 10140 7472 10152
rect 7524 10140 7530 10192
rect 10529 10180 10557 10220
rect 10597 10217 10609 10251
rect 10643 10248 10655 10251
rect 10962 10248 10968 10260
rect 10643 10220 10968 10248
rect 10643 10217 10655 10220
rect 10597 10211 10655 10217
rect 10962 10208 10968 10220
rect 11020 10208 11026 10260
rect 11072 10220 12572 10248
rect 11072 10180 11100 10220
rect 10529 10152 11100 10180
rect 12544 10180 12572 10220
rect 12618 10208 12624 10260
rect 12676 10248 12682 10260
rect 12986 10248 12992 10260
rect 12676 10220 12992 10248
rect 12676 10208 12682 10220
rect 12986 10208 12992 10220
rect 13044 10208 13050 10260
rect 13354 10208 13360 10260
rect 13412 10248 13418 10260
rect 14093 10251 14151 10257
rect 14093 10248 14105 10251
rect 13412 10220 14105 10248
rect 13412 10208 13418 10220
rect 14093 10217 14105 10220
rect 14139 10217 14151 10251
rect 14642 10248 14648 10260
rect 14093 10211 14151 10217
rect 14568 10220 14648 10248
rect 14568 10180 14596 10220
rect 14642 10208 14648 10220
rect 14700 10208 14706 10260
rect 14918 10248 14924 10260
rect 14879 10220 14924 10248
rect 14918 10208 14924 10220
rect 14976 10208 14982 10260
rect 12544 10152 14596 10180
rect 10505 10115 10563 10121
rect 10505 10081 10517 10115
rect 10551 10112 10563 10115
rect 10686 10112 10692 10124
rect 10551 10084 10692 10112
rect 10551 10081 10563 10084
rect 10505 10075 10563 10081
rect 10686 10072 10692 10084
rect 10744 10072 10750 10124
rect 12066 10072 12072 10124
rect 12124 10112 12130 10124
rect 12529 10115 12587 10121
rect 12529 10112 12541 10115
rect 12124 10084 12541 10112
rect 12124 10072 12130 10084
rect 12529 10081 12541 10084
rect 12575 10081 12587 10115
rect 12710 10112 12716 10124
rect 12671 10084 12716 10112
rect 12529 10075 12587 10081
rect 12710 10072 12716 10084
rect 12768 10072 12774 10124
rect 12989 10115 13047 10121
rect 12989 10081 13001 10115
rect 13035 10081 13047 10115
rect 12989 10075 13047 10081
rect 13173 10115 13231 10121
rect 13173 10081 13185 10115
rect 13219 10112 13231 10115
rect 13262 10112 13268 10124
rect 13219 10084 13268 10112
rect 13219 10081 13231 10084
rect 13173 10075 13231 10081
rect 1670 10044 1676 10056
rect 1631 10016 1676 10044
rect 1670 10004 1676 10016
rect 1728 10004 1734 10056
rect 5537 10047 5595 10053
rect 5537 10013 5549 10047
rect 5583 10013 5595 10047
rect 5537 10007 5595 10013
rect 5804 10047 5862 10053
rect 5804 10013 5816 10047
rect 5850 10013 5862 10047
rect 5804 10007 5862 10013
rect 7285 10047 7343 10053
rect 7285 10013 7297 10047
rect 7331 10044 7343 10047
rect 8757 10047 8815 10053
rect 8757 10044 8769 10047
rect 7331 10016 8769 10044
rect 7331 10013 7343 10016
rect 7285 10007 7343 10013
rect 8757 10013 8769 10016
rect 8803 10044 8815 10047
rect 8846 10044 8852 10056
rect 8803 10016 8852 10044
rect 8803 10013 8815 10016
rect 8757 10007 8815 10013
rect 4433 9979 4491 9985
rect 4433 9945 4445 9979
rect 4479 9976 4491 9979
rect 5353 9979 5411 9985
rect 5353 9976 5365 9979
rect 4479 9948 5365 9976
rect 4479 9945 4491 9948
rect 4433 9939 4491 9945
rect 5353 9945 5365 9948
rect 5399 9976 5411 9979
rect 5442 9976 5448 9988
rect 5399 9948 5448 9976
rect 5399 9945 5411 9948
rect 5353 9939 5411 9945
rect 5442 9936 5448 9948
rect 5500 9976 5506 9988
rect 5552 9976 5580 10007
rect 5500 9948 5580 9976
rect 5500 9936 5506 9948
rect 5718 9936 5724 9988
rect 5776 9976 5782 9988
rect 5828 9976 5856 10007
rect 8846 10004 8852 10016
rect 8904 10004 8910 10056
rect 9766 10004 9772 10056
rect 9824 10044 9830 10056
rect 10238 10047 10296 10053
rect 10238 10044 10250 10047
rect 9824 10016 10250 10044
rect 9824 10004 9830 10016
rect 10238 10013 10250 10016
rect 10284 10013 10296 10047
rect 10704 10044 10732 10072
rect 11977 10047 12035 10053
rect 11977 10044 11989 10047
rect 10704 10016 11989 10044
rect 10238 10007 10296 10013
rect 11977 10013 11989 10016
rect 12023 10013 12035 10047
rect 11977 10007 12035 10013
rect 12437 10047 12495 10053
rect 12437 10013 12449 10047
rect 12483 10044 12495 10047
rect 12483 10016 12572 10044
rect 12483 10013 12495 10016
rect 12437 10007 12495 10013
rect 5776 9948 5856 9976
rect 5776 9936 5782 9948
rect 7926 9936 7932 9988
rect 7984 9976 7990 9988
rect 8490 9979 8548 9985
rect 8490 9976 8502 9979
rect 7984 9948 8502 9976
rect 7984 9936 7990 9948
rect 8490 9945 8502 9948
rect 8536 9976 8548 9979
rect 11238 9976 11244 9988
rect 8536 9948 11244 9976
rect 8536 9945 8548 9948
rect 8490 9939 8548 9945
rect 11238 9936 11244 9948
rect 11296 9936 11302 9988
rect 11698 9936 11704 9988
rect 11756 9985 11762 9988
rect 11756 9976 11768 9985
rect 11756 9948 11801 9976
rect 11756 9939 11768 9948
rect 11756 9936 11762 9939
rect 2222 9868 2228 9920
rect 2280 9908 2286 9920
rect 9125 9911 9183 9917
rect 9125 9908 9137 9911
rect 2280 9880 9137 9908
rect 2280 9868 2286 9880
rect 9125 9877 9137 9880
rect 9171 9877 9183 9911
rect 9125 9871 9183 9877
rect 11146 9868 11152 9920
rect 11204 9908 11210 9920
rect 12069 9911 12127 9917
rect 12069 9908 12081 9911
rect 11204 9880 12081 9908
rect 11204 9868 11210 9880
rect 12069 9877 12081 9880
rect 12115 9877 12127 9911
rect 12544 9908 12572 10016
rect 12618 10004 12624 10056
rect 12676 10044 12682 10056
rect 13004 10044 13032 10075
rect 13262 10072 13268 10084
rect 13320 10072 13326 10124
rect 13814 10112 13820 10124
rect 13775 10084 13820 10112
rect 13814 10072 13820 10084
rect 13872 10072 13878 10124
rect 13998 10072 14004 10124
rect 14056 10112 14062 10124
rect 14550 10112 14556 10124
rect 14056 10084 14556 10112
rect 14056 10072 14062 10084
rect 14550 10072 14556 10084
rect 14608 10072 14614 10124
rect 14642 10072 14648 10124
rect 14700 10112 14706 10124
rect 14737 10115 14795 10121
rect 14737 10112 14749 10115
rect 14700 10084 14749 10112
rect 14700 10072 14706 10084
rect 14737 10081 14749 10084
rect 14783 10081 14795 10115
rect 15378 10112 15384 10124
rect 15339 10084 15384 10112
rect 14737 10075 14795 10081
rect 15378 10072 15384 10084
rect 15436 10072 15442 10124
rect 15470 10072 15476 10124
rect 15528 10112 15534 10124
rect 15528 10084 15573 10112
rect 15528 10072 15534 10084
rect 12676 10016 13032 10044
rect 15289 10047 15347 10053
rect 12676 10004 12682 10016
rect 15289 10013 15301 10047
rect 15335 10044 15347 10047
rect 15654 10044 15660 10056
rect 15335 10016 15660 10044
rect 15335 10013 15347 10016
rect 15289 10007 15347 10013
rect 15654 10004 15660 10016
rect 15712 10004 15718 10056
rect 13814 9936 13820 9988
rect 13872 9976 13878 9988
rect 14553 9979 14611 9985
rect 14553 9976 14565 9979
rect 13872 9948 14565 9976
rect 13872 9936 13878 9948
rect 14553 9945 14565 9948
rect 14599 9945 14611 9979
rect 14553 9939 14611 9945
rect 13265 9911 13323 9917
rect 13265 9908 13277 9911
rect 12544 9880 13277 9908
rect 12069 9871 12127 9877
rect 13265 9877 13277 9880
rect 13311 9908 13323 9911
rect 13446 9908 13452 9920
rect 13311 9880 13452 9908
rect 13311 9877 13323 9880
rect 13265 9871 13323 9877
rect 13446 9868 13452 9880
rect 13504 9868 13510 9920
rect 13630 9908 13636 9920
rect 13591 9880 13636 9908
rect 13630 9868 13636 9880
rect 13688 9868 13694 9920
rect 14458 9908 14464 9920
rect 14419 9880 14464 9908
rect 14458 9868 14464 9880
rect 14516 9868 14522 9920
rect 1104 9818 16008 9840
rect 1104 9766 4698 9818
rect 4750 9766 4762 9818
rect 4814 9766 4826 9818
rect 4878 9766 4890 9818
rect 4942 9766 4954 9818
rect 5006 9766 8446 9818
rect 8498 9766 8510 9818
rect 8562 9766 8574 9818
rect 8626 9766 8638 9818
rect 8690 9766 8702 9818
rect 8754 9766 12194 9818
rect 12246 9766 12258 9818
rect 12310 9766 12322 9818
rect 12374 9766 12386 9818
rect 12438 9766 12450 9818
rect 12502 9766 16008 9818
rect 1104 9744 16008 9766
rect 1670 9664 1676 9716
rect 1728 9704 1734 9716
rect 1765 9707 1823 9713
rect 1765 9704 1777 9707
rect 1728 9676 1777 9704
rect 1728 9664 1734 9676
rect 1765 9673 1777 9676
rect 1811 9673 1823 9707
rect 1765 9667 1823 9673
rect 2314 9664 2320 9716
rect 2372 9704 2378 9716
rect 5718 9704 5724 9716
rect 2372 9676 5724 9704
rect 2372 9664 2378 9676
rect 5718 9664 5724 9676
rect 5776 9664 5782 9716
rect 7558 9664 7564 9716
rect 7616 9704 7622 9716
rect 7616 9676 7880 9704
rect 7616 9664 7622 9676
rect 5442 9596 5448 9648
rect 5500 9636 5506 9648
rect 6181 9639 6239 9645
rect 5500 9608 5948 9636
rect 5500 9596 5506 9608
rect 1673 9571 1731 9577
rect 1673 9537 1685 9571
rect 1719 9568 1731 9571
rect 1762 9568 1768 9580
rect 1719 9540 1768 9568
rect 1719 9537 1731 9540
rect 1673 9531 1731 9537
rect 1762 9528 1768 9540
rect 1820 9528 1826 9580
rect 1949 9571 2007 9577
rect 1949 9537 1961 9571
rect 1995 9568 2007 9571
rect 2130 9568 2136 9580
rect 1995 9540 2136 9568
rect 1995 9537 2007 9540
rect 1949 9531 2007 9537
rect 2130 9528 2136 9540
rect 2188 9528 2194 9580
rect 3228 9571 3286 9577
rect 3228 9537 3240 9571
rect 3274 9568 3286 9571
rect 3970 9568 3976 9580
rect 3274 9540 3976 9568
rect 3274 9537 3286 9540
rect 3228 9531 3286 9537
rect 3970 9528 3976 9540
rect 4028 9568 4034 9580
rect 5350 9568 5356 9580
rect 4028 9540 5356 9568
rect 4028 9528 4034 9540
rect 5350 9528 5356 9540
rect 5408 9528 5414 9580
rect 5920 9577 5948 9608
rect 6181 9605 6193 9639
rect 6227 9636 6239 9639
rect 7852 9636 7880 9676
rect 9490 9664 9496 9716
rect 9548 9704 9554 9716
rect 10686 9704 10692 9716
rect 9548 9676 10088 9704
rect 10647 9676 10692 9704
rect 9548 9664 9554 9676
rect 8662 9636 8668 9648
rect 6227 9608 7788 9636
rect 7852 9608 8668 9636
rect 6227 9605 6239 9608
rect 6181 9599 6239 9605
rect 5649 9571 5707 9577
rect 5649 9537 5661 9571
rect 5695 9568 5707 9571
rect 5905 9571 5963 9577
rect 5695 9540 5856 9568
rect 5695 9537 5707 9540
rect 5649 9531 5707 9537
rect 2961 9503 3019 9509
rect 2961 9469 2973 9503
rect 3007 9469 3019 9503
rect 5828 9500 5856 9540
rect 5905 9537 5917 9571
rect 5951 9568 5963 9571
rect 6196 9568 6224 9599
rect 5951 9540 6224 9568
rect 5951 9537 5963 9540
rect 5905 9531 5963 9537
rect 7466 9528 7472 9580
rect 7524 9577 7530 9580
rect 7524 9568 7536 9577
rect 7524 9540 7569 9568
rect 7524 9531 7536 9540
rect 7524 9528 7530 9531
rect 7760 9509 7788 9608
rect 8662 9596 8668 9608
rect 8720 9596 8726 9648
rect 8757 9639 8815 9645
rect 8757 9605 8769 9639
rect 8803 9636 8815 9639
rect 8846 9636 8852 9648
rect 8803 9608 8852 9636
rect 8803 9605 8815 9608
rect 8757 9599 8815 9605
rect 8846 9596 8852 9608
rect 8904 9636 8910 9648
rect 8941 9639 8999 9645
rect 8941 9636 8953 9639
rect 8904 9608 8953 9636
rect 8904 9596 8910 9608
rect 8941 9605 8953 9608
rect 8987 9636 8999 9639
rect 9858 9636 9864 9648
rect 8987 9608 9864 9636
rect 8987 9605 8999 9608
rect 8941 9599 8999 9605
rect 9858 9596 9864 9608
rect 9916 9596 9922 9648
rect 10060 9636 10088 9676
rect 10686 9664 10692 9676
rect 10744 9664 10750 9716
rect 11698 9664 11704 9716
rect 11756 9704 11762 9716
rect 12618 9704 12624 9716
rect 11756 9676 12624 9704
rect 11756 9664 11762 9676
rect 12618 9664 12624 9676
rect 12676 9664 12682 9716
rect 12894 9664 12900 9716
rect 12952 9704 12958 9716
rect 13173 9707 13231 9713
rect 13173 9704 13185 9707
rect 12952 9676 13185 9704
rect 12952 9664 12958 9676
rect 13173 9673 13185 9676
rect 13219 9673 13231 9707
rect 13173 9667 13231 9673
rect 14458 9664 14464 9716
rect 14516 9704 14522 9716
rect 14829 9707 14887 9713
rect 14829 9704 14841 9707
rect 14516 9676 14841 9704
rect 14516 9664 14522 9676
rect 14829 9673 14841 9676
rect 14875 9673 14887 9707
rect 14829 9667 14887 9673
rect 10238 9639 10296 9645
rect 10238 9636 10250 9639
rect 10060 9608 10250 9636
rect 10238 9605 10250 9608
rect 10284 9605 10296 9639
rect 10238 9599 10296 9605
rect 7834 9528 7840 9580
rect 7892 9568 7898 9580
rect 10505 9571 10563 9577
rect 7892 9540 10465 9568
rect 7892 9528 7898 9540
rect 7745 9503 7803 9509
rect 5828 9472 6408 9500
rect 2961 9463 3019 9469
rect 1486 9432 1492 9444
rect 1447 9404 1492 9432
rect 1486 9392 1492 9404
rect 1544 9392 1550 9444
rect 2869 9367 2927 9373
rect 2869 9333 2881 9367
rect 2915 9364 2927 9367
rect 2976 9364 3004 9463
rect 4338 9432 4344 9444
rect 4299 9404 4344 9432
rect 4338 9392 4344 9404
rect 4396 9392 4402 9444
rect 3142 9364 3148 9376
rect 2915 9336 3148 9364
rect 2915 9333 2927 9336
rect 2869 9327 2927 9333
rect 3142 9324 3148 9336
rect 3200 9364 3206 9376
rect 3970 9364 3976 9376
rect 3200 9336 3976 9364
rect 3200 9324 3206 9336
rect 3970 9324 3976 9336
rect 4028 9324 4034 9376
rect 4525 9367 4583 9373
rect 4525 9333 4537 9367
rect 4571 9364 4583 9367
rect 5534 9364 5540 9376
rect 4571 9336 5540 9364
rect 4571 9333 4583 9336
rect 4525 9327 4583 9333
rect 5534 9324 5540 9336
rect 5592 9324 5598 9376
rect 6380 9373 6408 9472
rect 7745 9469 7757 9503
rect 7791 9500 7803 9503
rect 8846 9500 8852 9512
rect 7791 9472 8852 9500
rect 7791 9469 7803 9472
rect 7745 9463 7803 9469
rect 8846 9460 8852 9472
rect 8904 9460 8910 9512
rect 10437 9500 10465 9540
rect 10505 9537 10517 9571
rect 10551 9568 10563 9571
rect 10704 9568 10732 9664
rect 11790 9596 11796 9648
rect 11848 9636 11854 9648
rect 11848 9608 13492 9636
rect 11848 9596 11854 9608
rect 10551 9540 10732 9568
rect 11977 9571 12035 9577
rect 10551 9537 10563 9540
rect 10505 9531 10563 9537
rect 11977 9537 11989 9571
rect 12023 9568 12035 9571
rect 12618 9568 12624 9580
rect 12023 9540 12624 9568
rect 12023 9537 12035 9540
rect 11977 9531 12035 9537
rect 12618 9528 12624 9540
rect 12676 9528 12682 9580
rect 12802 9528 12808 9580
rect 12860 9568 12866 9580
rect 12860 9540 13400 9568
rect 12860 9528 12866 9540
rect 12069 9503 12127 9509
rect 12069 9500 12081 9503
rect 10437 9472 12081 9500
rect 12069 9469 12081 9472
rect 12115 9469 12127 9503
rect 12069 9463 12127 9469
rect 11606 9432 11612 9444
rect 8588 9404 9260 9432
rect 11567 9404 11612 9432
rect 6365 9367 6423 9373
rect 6365 9333 6377 9367
rect 6411 9364 6423 9367
rect 8588 9364 8616 9404
rect 9122 9364 9128 9376
rect 6411 9336 8616 9364
rect 9083 9336 9128 9364
rect 6411 9333 6423 9336
rect 6365 9327 6423 9333
rect 9122 9324 9128 9336
rect 9180 9324 9186 9376
rect 9232 9364 9260 9404
rect 11606 9392 11612 9404
rect 11664 9392 11670 9444
rect 12084 9432 12112 9463
rect 12158 9460 12164 9512
rect 12216 9500 12222 9512
rect 13078 9500 13084 9512
rect 12216 9472 12261 9500
rect 12544 9472 13084 9500
rect 12216 9460 12222 9472
rect 12544 9441 12572 9472
rect 13078 9460 13084 9472
rect 13136 9460 13142 9512
rect 13170 9460 13176 9512
rect 13228 9500 13234 9512
rect 13372 9509 13400 9540
rect 13265 9503 13323 9509
rect 13265 9500 13277 9503
rect 13228 9472 13277 9500
rect 13228 9460 13234 9472
rect 13265 9469 13277 9472
rect 13311 9469 13323 9503
rect 13265 9463 13323 9469
rect 13357 9503 13415 9509
rect 13357 9469 13369 9503
rect 13403 9469 13415 9503
rect 13464 9500 13492 9608
rect 13630 9596 13636 9648
rect 13688 9636 13694 9648
rect 14093 9639 14151 9645
rect 14093 9636 14105 9639
rect 13688 9608 14105 9636
rect 13688 9596 13694 9608
rect 14093 9605 14105 9608
rect 14139 9605 14151 9639
rect 14093 9599 14151 9605
rect 15197 9639 15255 9645
rect 15197 9605 15209 9639
rect 15243 9636 15255 9639
rect 15286 9636 15292 9648
rect 15243 9608 15292 9636
rect 15243 9605 15255 9608
rect 15197 9599 15255 9605
rect 15286 9596 15292 9608
rect 15344 9596 15350 9648
rect 13906 9528 13912 9580
rect 13964 9568 13970 9580
rect 14001 9571 14059 9577
rect 14001 9568 14013 9571
rect 13964 9540 14013 9568
rect 13964 9528 13970 9540
rect 14001 9537 14013 9540
rect 14047 9537 14059 9571
rect 14001 9531 14059 9537
rect 14458 9528 14464 9580
rect 14516 9568 14522 9580
rect 14553 9571 14611 9577
rect 14553 9568 14565 9571
rect 14516 9540 14565 9568
rect 14516 9528 14522 9540
rect 14553 9537 14565 9540
rect 14599 9537 14611 9571
rect 15562 9568 15568 9580
rect 14553 9531 14611 9537
rect 15304 9540 15568 9568
rect 15304 9509 15332 9540
rect 15562 9528 15568 9540
rect 15620 9528 15626 9580
rect 14185 9503 14243 9509
rect 14185 9500 14197 9503
rect 13464 9472 14197 9500
rect 13357 9463 13415 9469
rect 14185 9469 14197 9472
rect 14231 9469 14243 9503
rect 14185 9463 14243 9469
rect 15289 9503 15347 9509
rect 15289 9469 15301 9503
rect 15335 9469 15347 9503
rect 15470 9500 15476 9512
rect 15431 9472 15476 9500
rect 15289 9463 15347 9469
rect 15470 9460 15476 9472
rect 15528 9460 15534 9512
rect 12529 9435 12587 9441
rect 12529 9432 12541 9435
rect 12084 9404 12541 9432
rect 12529 9401 12541 9404
rect 12575 9401 12587 9435
rect 12802 9432 12808 9444
rect 12763 9404 12808 9432
rect 12529 9395 12587 9401
rect 12802 9392 12808 9404
rect 12860 9392 12866 9444
rect 11790 9364 11796 9376
rect 9232 9336 11796 9364
rect 11790 9324 11796 9336
rect 11848 9324 11854 9376
rect 12618 9364 12624 9376
rect 12579 9336 12624 9364
rect 12618 9324 12624 9336
rect 12676 9324 12682 9376
rect 13630 9364 13636 9376
rect 13591 9336 13636 9364
rect 13630 9324 13636 9336
rect 13688 9324 13694 9376
rect 14737 9367 14795 9373
rect 14737 9333 14749 9367
rect 14783 9364 14795 9367
rect 15470 9364 15476 9376
rect 14783 9336 15476 9364
rect 14783 9333 14795 9336
rect 14737 9327 14795 9333
rect 15470 9324 15476 9336
rect 15528 9324 15534 9376
rect 1104 9274 16008 9296
rect 1104 9222 2824 9274
rect 2876 9222 2888 9274
rect 2940 9222 2952 9274
rect 3004 9222 3016 9274
rect 3068 9222 3080 9274
rect 3132 9222 6572 9274
rect 6624 9222 6636 9274
rect 6688 9222 6700 9274
rect 6752 9222 6764 9274
rect 6816 9222 6828 9274
rect 6880 9222 10320 9274
rect 10372 9222 10384 9274
rect 10436 9222 10448 9274
rect 10500 9222 10512 9274
rect 10564 9222 10576 9274
rect 10628 9222 14068 9274
rect 14120 9222 14132 9274
rect 14184 9222 14196 9274
rect 14248 9222 14260 9274
rect 14312 9222 14324 9274
rect 14376 9222 16008 9274
rect 1104 9200 16008 9222
rect 1762 9160 1768 9172
rect 1723 9132 1768 9160
rect 1762 9120 1768 9132
rect 1820 9120 1826 9172
rect 3142 9160 3148 9172
rect 2240 9132 3148 9160
rect 2240 9033 2268 9132
rect 3142 9120 3148 9132
rect 3200 9120 3206 9172
rect 3973 9163 4031 9169
rect 3973 9129 3985 9163
rect 4019 9160 4031 9163
rect 7374 9160 7380 9172
rect 4019 9132 7380 9160
rect 4019 9129 4031 9132
rect 3973 9123 4031 9129
rect 3510 9052 3516 9104
rect 3568 9092 3574 9104
rect 3786 9092 3792 9104
rect 3568 9064 3792 9092
rect 3568 9052 3574 9064
rect 3786 9052 3792 9064
rect 3844 9052 3850 9104
rect 2225 9027 2283 9033
rect 2225 8993 2237 9027
rect 2271 8993 2283 9027
rect 3988 9024 4016 9123
rect 7374 9120 7380 9132
rect 7432 9120 7438 9172
rect 8846 9120 8852 9172
rect 8904 9160 8910 9172
rect 9217 9163 9275 9169
rect 9217 9160 9229 9163
rect 8904 9132 9229 9160
rect 8904 9120 8910 9132
rect 9217 9129 9229 9132
rect 9263 9129 9275 9163
rect 9217 9123 9275 9129
rect 9306 9120 9312 9172
rect 9364 9160 9370 9172
rect 9401 9163 9459 9169
rect 9401 9160 9413 9163
rect 9364 9132 9413 9160
rect 9364 9120 9370 9132
rect 9401 9129 9413 9132
rect 9447 9129 9459 9163
rect 9401 9123 9459 9129
rect 9582 9120 9588 9172
rect 9640 9160 9646 9172
rect 11793 9163 11851 9169
rect 11793 9160 11805 9163
rect 9640 9132 11805 9160
rect 9640 9120 9646 9132
rect 11793 9129 11805 9132
rect 11839 9160 11851 9163
rect 15194 9160 15200 9172
rect 11839 9132 15200 9160
rect 11839 9129 11851 9132
rect 11793 9123 11851 9129
rect 15194 9120 15200 9132
rect 15252 9120 15258 9172
rect 5350 9052 5356 9104
rect 5408 9092 5414 9104
rect 7466 9092 7472 9104
rect 5408 9064 7472 9092
rect 5408 9052 5414 9064
rect 7466 9052 7472 9064
rect 7524 9052 7530 9104
rect 5442 9024 5448 9036
rect 2225 8987 2283 8993
rect 3528 8996 4016 9024
rect 5368 8996 5448 9024
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8956 1731 8959
rect 1762 8956 1768 8968
rect 1719 8928 1768 8956
rect 1719 8925 1731 8928
rect 1673 8919 1731 8925
rect 1762 8916 1768 8928
rect 1820 8916 1826 8968
rect 1946 8956 1952 8968
rect 1907 8928 1952 8956
rect 1946 8916 1952 8928
rect 2004 8916 2010 8968
rect 2038 8848 2044 8900
rect 2096 8888 2102 8900
rect 2222 8888 2228 8900
rect 2096 8860 2228 8888
rect 2096 8848 2102 8860
rect 2222 8848 2228 8860
rect 2280 8888 2286 8900
rect 2470 8891 2528 8897
rect 2470 8888 2482 8891
rect 2280 8860 2482 8888
rect 2280 8848 2286 8860
rect 2470 8857 2482 8860
rect 2516 8857 2528 8891
rect 2470 8851 2528 8857
rect 1486 8820 1492 8832
rect 1447 8792 1492 8820
rect 1486 8780 1492 8792
rect 1544 8780 1550 8832
rect 2314 8780 2320 8832
rect 2372 8820 2378 8832
rect 3528 8820 3556 8996
rect 3881 8959 3939 8965
rect 3881 8925 3893 8959
rect 3927 8956 3939 8959
rect 3970 8956 3976 8968
rect 3927 8928 3976 8956
rect 3927 8925 3939 8928
rect 3881 8919 3939 8925
rect 3970 8916 3976 8928
rect 4028 8956 4034 8968
rect 5368 8965 5396 8996
rect 5442 8984 5448 8996
rect 5500 8984 5506 9036
rect 8757 9027 8815 9033
rect 8757 8993 8769 9027
rect 8803 9024 8815 9027
rect 8864 9024 8892 9120
rect 9030 9052 9036 9104
rect 9088 9092 9094 9104
rect 9490 9092 9496 9104
rect 9088 9064 9496 9092
rect 9088 9052 9094 9064
rect 9490 9052 9496 9064
rect 9548 9052 9554 9104
rect 11606 9052 11612 9104
rect 11664 9092 11670 9104
rect 11882 9092 11888 9104
rect 11664 9064 11888 9092
rect 11664 9052 11670 9064
rect 11882 9052 11888 9064
rect 11940 9092 11946 9104
rect 12158 9092 12164 9104
rect 11940 9064 12164 9092
rect 11940 9052 11946 9064
rect 12158 9052 12164 9064
rect 12216 9052 12222 9104
rect 12526 9092 12532 9104
rect 12487 9064 12532 9092
rect 12526 9052 12532 9064
rect 12584 9092 12590 9104
rect 13078 9092 13084 9104
rect 12584 9064 13084 9092
rect 12584 9052 12590 9064
rect 13078 9052 13084 9064
rect 13136 9052 13142 9104
rect 14918 9092 14924 9104
rect 13188 9064 14924 9092
rect 8803 8996 8892 9024
rect 8803 8993 8815 8996
rect 8757 8987 8815 8993
rect 5353 8959 5411 8965
rect 5353 8956 5365 8959
rect 4028 8928 5365 8956
rect 4028 8916 4034 8928
rect 5353 8925 5365 8928
rect 5399 8925 5411 8959
rect 5353 8919 5411 8925
rect 7285 8959 7343 8965
rect 7285 8925 7297 8959
rect 7331 8956 7343 8959
rect 8864 8956 8892 8996
rect 11974 8984 11980 9036
rect 12032 9024 12038 9036
rect 13188 9024 13216 9064
rect 14918 9052 14924 9064
rect 14976 9052 14982 9104
rect 15102 9052 15108 9104
rect 15160 9092 15166 9104
rect 15565 9095 15623 9101
rect 15565 9092 15577 9095
rect 15160 9064 15577 9092
rect 15160 9052 15166 9064
rect 15565 9061 15577 9064
rect 15611 9061 15623 9095
rect 15565 9055 15623 9061
rect 12032 8996 13216 9024
rect 13541 9027 13599 9033
rect 12032 8984 12038 8996
rect 13541 8993 13553 9027
rect 13587 9024 13599 9027
rect 14734 9024 14740 9036
rect 13587 8996 14740 9024
rect 13587 8993 13599 8996
rect 13541 8987 13599 8993
rect 14734 8984 14740 8996
rect 14792 8984 14798 9036
rect 15286 9024 15292 9036
rect 15247 8996 15292 9024
rect 15286 8984 15292 8996
rect 15344 8984 15350 9036
rect 9030 8956 9036 8968
rect 7331 8928 9036 8956
rect 7331 8925 7343 8928
rect 7285 8919 7343 8925
rect 9030 8916 9036 8928
rect 9088 8916 9094 8968
rect 10686 8916 10692 8968
rect 10744 8956 10750 8968
rect 10781 8959 10839 8965
rect 10781 8956 10793 8959
rect 10744 8928 10793 8956
rect 10744 8916 10750 8928
rect 10781 8925 10793 8928
rect 10827 8925 10839 8959
rect 13262 8956 13268 8968
rect 13223 8928 13268 8956
rect 10781 8919 10839 8925
rect 13262 8916 13268 8928
rect 13320 8916 13326 8968
rect 13817 8959 13875 8965
rect 13817 8925 13829 8959
rect 13863 8956 13875 8959
rect 14550 8956 14556 8968
rect 13863 8928 14556 8956
rect 13863 8925 13875 8928
rect 13817 8919 13875 8925
rect 14550 8916 14556 8928
rect 14608 8916 14614 8968
rect 14645 8959 14703 8965
rect 14645 8925 14657 8959
rect 14691 8956 14703 8959
rect 15102 8956 15108 8968
rect 14691 8928 15108 8956
rect 14691 8925 14703 8928
rect 14645 8919 14703 8925
rect 15102 8916 15108 8928
rect 15160 8916 15166 8968
rect 15381 8959 15439 8965
rect 15381 8925 15393 8959
rect 15427 8956 15439 8959
rect 15470 8956 15476 8968
rect 15427 8928 15476 8956
rect 15427 8925 15439 8928
rect 15381 8919 15439 8925
rect 15470 8916 15476 8928
rect 15528 8916 15534 8968
rect 3694 8848 3700 8900
rect 3752 8888 3758 8900
rect 3752 8860 3924 8888
rect 3752 8848 3758 8860
rect 2372 8792 3556 8820
rect 3605 8823 3663 8829
rect 2372 8780 2378 8792
rect 3605 8789 3617 8823
rect 3651 8820 3663 8823
rect 3786 8820 3792 8832
rect 3651 8792 3792 8820
rect 3651 8789 3663 8792
rect 3605 8783 3663 8789
rect 3786 8780 3792 8792
rect 3844 8780 3850 8832
rect 3896 8820 3924 8860
rect 4338 8848 4344 8900
rect 4396 8888 4402 8900
rect 5086 8891 5144 8897
rect 5086 8888 5098 8891
rect 4396 8860 5098 8888
rect 4396 8848 4402 8860
rect 5086 8857 5098 8860
rect 5132 8857 5144 8891
rect 5086 8851 5144 8857
rect 6086 8848 6092 8900
rect 6144 8888 6150 8900
rect 6454 8888 6460 8900
rect 6144 8860 6460 8888
rect 6144 8848 6150 8860
rect 6454 8848 6460 8860
rect 6512 8848 6518 8900
rect 8294 8848 8300 8900
rect 8352 8888 8358 8900
rect 8490 8891 8548 8897
rect 8490 8888 8502 8891
rect 8352 8860 8502 8888
rect 8352 8848 8358 8860
rect 8490 8857 8502 8860
rect 8536 8888 8548 8891
rect 9214 8888 9220 8900
rect 8536 8860 9220 8888
rect 8536 8857 8548 8860
rect 8490 8851 8548 8857
rect 9214 8848 9220 8860
rect 9272 8848 9278 8900
rect 10318 8848 10324 8900
rect 10376 8888 10382 8900
rect 10514 8891 10572 8897
rect 10514 8888 10526 8891
rect 10376 8860 10526 8888
rect 10376 8848 10382 8860
rect 10514 8857 10526 8860
rect 10560 8857 10572 8891
rect 10514 8851 10572 8857
rect 11330 8848 11336 8900
rect 11388 8888 11394 8900
rect 11977 8891 12035 8897
rect 11977 8888 11989 8891
rect 11388 8860 11989 8888
rect 11388 8848 11394 8860
rect 11977 8857 11989 8860
rect 12023 8888 12035 8891
rect 12805 8891 12863 8897
rect 12023 8860 12480 8888
rect 12023 8857 12035 8860
rect 11977 8851 12035 8857
rect 7377 8823 7435 8829
rect 7377 8820 7389 8823
rect 3896 8792 7389 8820
rect 7377 8789 7389 8792
rect 7423 8820 7435 8823
rect 10686 8820 10692 8832
rect 7423 8792 10692 8820
rect 7423 8789 7435 8792
rect 7377 8783 7435 8789
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 12066 8780 12072 8832
rect 12124 8820 12130 8832
rect 12452 8829 12480 8860
rect 12805 8857 12817 8891
rect 12851 8888 12863 8891
rect 12986 8888 12992 8900
rect 12851 8860 12992 8888
rect 12851 8857 12863 8860
rect 12805 8851 12863 8857
rect 12986 8848 12992 8860
rect 13044 8848 13050 8900
rect 13357 8891 13415 8897
rect 13357 8857 13369 8891
rect 13403 8888 13415 8891
rect 14274 8888 14280 8900
rect 13403 8860 14280 8888
rect 13403 8857 13415 8860
rect 13357 8851 13415 8857
rect 14274 8848 14280 8860
rect 14332 8888 14338 8900
rect 16390 8888 16396 8900
rect 14332 8860 16396 8888
rect 14332 8848 14338 8860
rect 16390 8848 16396 8860
rect 16448 8848 16454 8900
rect 12161 8823 12219 8829
rect 12161 8820 12173 8823
rect 12124 8792 12173 8820
rect 12124 8780 12130 8792
rect 12161 8789 12173 8792
rect 12207 8789 12219 8823
rect 12161 8783 12219 8789
rect 12437 8823 12495 8829
rect 12437 8789 12449 8823
rect 12483 8820 12495 8823
rect 12526 8820 12532 8832
rect 12483 8792 12532 8820
rect 12483 8789 12495 8792
rect 12437 8783 12495 8789
rect 12526 8780 12532 8792
rect 12584 8780 12590 8832
rect 12894 8820 12900 8832
rect 12855 8792 12900 8820
rect 12894 8780 12900 8792
rect 12952 8780 12958 8832
rect 13170 8780 13176 8832
rect 13228 8820 13234 8832
rect 13630 8820 13636 8832
rect 13228 8792 13636 8820
rect 13228 8780 13234 8792
rect 13630 8780 13636 8792
rect 13688 8780 13694 8832
rect 14090 8820 14096 8832
rect 14051 8792 14096 8820
rect 14090 8780 14096 8792
rect 14148 8780 14154 8832
rect 14458 8820 14464 8832
rect 14419 8792 14464 8820
rect 14458 8780 14464 8792
rect 14516 8780 14522 8832
rect 1104 8730 16008 8752
rect 1104 8678 4698 8730
rect 4750 8678 4762 8730
rect 4814 8678 4826 8730
rect 4878 8678 4890 8730
rect 4942 8678 4954 8730
rect 5006 8678 8446 8730
rect 8498 8678 8510 8730
rect 8562 8678 8574 8730
rect 8626 8678 8638 8730
rect 8690 8678 8702 8730
rect 8754 8678 12194 8730
rect 12246 8678 12258 8730
rect 12310 8678 12322 8730
rect 12374 8678 12386 8730
rect 12438 8678 12450 8730
rect 12502 8678 16008 8730
rect 1104 8656 16008 8678
rect 1854 8616 1860 8628
rect 1815 8588 1860 8616
rect 1854 8576 1860 8588
rect 1912 8576 1918 8628
rect 1946 8576 1952 8628
rect 2004 8616 2010 8628
rect 2225 8619 2283 8625
rect 2225 8616 2237 8619
rect 2004 8588 2237 8616
rect 2004 8576 2010 8588
rect 2225 8585 2237 8588
rect 2271 8585 2283 8619
rect 2225 8579 2283 8585
rect 5258 8576 5264 8628
rect 5316 8616 5322 8628
rect 7745 8619 7803 8625
rect 5316 8588 7236 8616
rect 5316 8576 5322 8588
rect 1765 8551 1823 8557
rect 1765 8517 1777 8551
rect 1811 8548 1823 8551
rect 6730 8548 6736 8560
rect 1811 8520 6736 8548
rect 1811 8517 1823 8520
rect 1765 8511 1823 8517
rect 6730 8508 6736 8520
rect 6788 8508 6794 8560
rect 7208 8548 7236 8588
rect 7745 8585 7757 8619
rect 7791 8616 7803 8619
rect 7926 8616 7932 8628
rect 7791 8588 7932 8616
rect 7791 8585 7803 8588
rect 7745 8579 7803 8585
rect 7926 8576 7932 8588
rect 7984 8576 7990 8628
rect 9030 8616 9036 8628
rect 8991 8588 9036 8616
rect 9030 8576 9036 8588
rect 9088 8576 9094 8628
rect 9674 8576 9680 8628
rect 9732 8616 9738 8628
rect 10318 8616 10324 8628
rect 9732 8588 10324 8616
rect 9732 8576 9738 8588
rect 10318 8576 10324 8588
rect 10376 8576 10382 8628
rect 10597 8619 10655 8625
rect 10597 8585 10609 8619
rect 10643 8616 10655 8619
rect 10870 8616 10876 8628
rect 10643 8588 10876 8616
rect 10643 8585 10655 8588
rect 10597 8579 10655 8585
rect 10870 8576 10876 8588
rect 10928 8616 10934 8628
rect 13538 8616 13544 8628
rect 10928 8588 12480 8616
rect 13499 8588 13544 8616
rect 10928 8576 10934 8588
rect 7208 8520 7972 8548
rect 3694 8440 3700 8492
rect 3752 8489 3758 8492
rect 3752 8480 3764 8489
rect 3970 8480 3976 8492
rect 3752 8452 3797 8480
rect 3931 8452 3976 8480
rect 3752 8443 3764 8452
rect 3752 8440 3758 8443
rect 3970 8440 3976 8452
rect 4028 8480 4034 8492
rect 4065 8483 4123 8489
rect 4065 8480 4077 8483
rect 4028 8452 4077 8480
rect 4028 8440 4034 8452
rect 4065 8449 4077 8452
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 4332 8483 4390 8489
rect 4332 8449 4344 8483
rect 4378 8480 4390 8483
rect 4614 8480 4620 8492
rect 4378 8452 4620 8480
rect 4378 8449 4390 8452
rect 4332 8443 4390 8449
rect 4614 8440 4620 8452
rect 4672 8440 4678 8492
rect 6632 8483 6690 8489
rect 6632 8449 6644 8483
rect 6678 8480 6690 8483
rect 6678 8452 7880 8480
rect 6678 8449 6690 8452
rect 6632 8443 6690 8449
rect 1673 8415 1731 8421
rect 1673 8381 1685 8415
rect 1719 8412 1731 8415
rect 6365 8415 6423 8421
rect 1719 8384 3004 8412
rect 1719 8381 1731 8384
rect 1673 8375 1731 8381
rect 2406 8236 2412 8288
rect 2464 8276 2470 8288
rect 2593 8279 2651 8285
rect 2593 8276 2605 8279
rect 2464 8248 2605 8276
rect 2464 8236 2470 8248
rect 2593 8245 2605 8248
rect 2639 8245 2651 8279
rect 2976 8276 3004 8384
rect 6365 8381 6377 8415
rect 6411 8381 6423 8415
rect 6365 8375 6423 8381
rect 5534 8344 5540 8356
rect 5000 8316 5540 8344
rect 5000 8276 5028 8316
rect 5534 8304 5540 8316
rect 5592 8304 5598 8356
rect 2976 8248 5028 8276
rect 2593 8239 2651 8245
rect 5350 8236 5356 8288
rect 5408 8276 5414 8288
rect 5445 8279 5503 8285
rect 5445 8276 5457 8279
rect 5408 8248 5457 8276
rect 5408 8236 5414 8248
rect 5445 8245 5457 8248
rect 5491 8245 5503 8279
rect 5445 8239 5503 8245
rect 6181 8279 6239 8285
rect 6181 8245 6193 8279
rect 6227 8276 6239 8279
rect 6380 8276 6408 8375
rect 7650 8276 7656 8288
rect 6227 8248 7656 8276
rect 6227 8245 6239 8248
rect 6181 8239 6239 8245
rect 7650 8236 7656 8248
rect 7708 8236 7714 8288
rect 7852 8276 7880 8452
rect 7944 8424 7972 8520
rect 9048 8480 9076 8576
rect 9122 8508 9128 8560
rect 9180 8548 9186 8560
rect 9462 8551 9520 8557
rect 9462 8548 9474 8551
rect 9180 8520 9474 8548
rect 9180 8508 9186 8520
rect 9462 8517 9474 8520
rect 9508 8517 9520 8551
rect 11606 8548 11612 8560
rect 9462 8511 9520 8517
rect 9600 8520 11612 8548
rect 9217 8483 9275 8489
rect 9217 8480 9229 8483
rect 9048 8452 9229 8480
rect 9217 8449 9229 8452
rect 9263 8449 9275 8483
rect 9600 8480 9628 8520
rect 11606 8508 11612 8520
rect 11664 8508 11670 8560
rect 11698 8508 11704 8560
rect 11756 8548 11762 8560
rect 11756 8520 12112 8548
rect 11756 8508 11762 8520
rect 9217 8443 9275 8449
rect 9324 8452 9628 8480
rect 7926 8372 7932 8424
rect 7984 8412 7990 8424
rect 9324 8412 9352 8452
rect 11054 8440 11060 8492
rect 11112 8480 11118 8492
rect 11882 8480 11888 8492
rect 11112 8452 11888 8480
rect 11112 8440 11118 8452
rect 11882 8440 11888 8452
rect 11940 8440 11946 8492
rect 7984 8384 9352 8412
rect 11333 8415 11391 8421
rect 7984 8372 7990 8384
rect 11333 8381 11345 8415
rect 11379 8412 11391 8415
rect 11698 8412 11704 8424
rect 11379 8384 11704 8412
rect 11379 8381 11391 8384
rect 11333 8375 11391 8381
rect 11698 8372 11704 8384
rect 11756 8372 11762 8424
rect 11974 8412 11980 8424
rect 11935 8384 11980 8412
rect 11974 8372 11980 8384
rect 12032 8372 12038 8424
rect 12084 8421 12112 8520
rect 12452 8480 12480 8588
rect 13538 8576 13544 8588
rect 13596 8576 13602 8628
rect 13906 8576 13912 8628
rect 13964 8616 13970 8628
rect 14185 8619 14243 8625
rect 14185 8616 14197 8619
rect 13964 8588 14197 8616
rect 13964 8576 13970 8588
rect 14185 8585 14197 8588
rect 14231 8585 14243 8619
rect 14185 8579 14243 8585
rect 14553 8619 14611 8625
rect 14553 8585 14565 8619
rect 14599 8616 14611 8619
rect 14599 8588 14780 8616
rect 14599 8585 14611 8588
rect 14553 8579 14611 8585
rect 12713 8551 12771 8557
rect 12713 8517 12725 8551
rect 12759 8548 12771 8551
rect 12802 8548 12808 8560
rect 12759 8520 12808 8548
rect 12759 8517 12771 8520
rect 12713 8511 12771 8517
rect 12802 8508 12808 8520
rect 12860 8508 12866 8560
rect 13446 8508 13452 8560
rect 13504 8508 13510 8560
rect 14274 8548 14280 8560
rect 14016 8520 14280 8548
rect 13464 8480 13492 8508
rect 14016 8480 14044 8520
rect 14274 8508 14280 8520
rect 14332 8508 14338 8560
rect 14642 8508 14648 8560
rect 14700 8508 14706 8560
rect 14752 8548 14780 8588
rect 14918 8576 14924 8628
rect 14976 8616 14982 8628
rect 15565 8619 15623 8625
rect 15565 8616 15577 8619
rect 14976 8588 15577 8616
rect 14976 8576 14982 8588
rect 15565 8585 15577 8588
rect 15611 8585 15623 8619
rect 15565 8579 15623 8585
rect 15102 8548 15108 8560
rect 14752 8520 15108 8548
rect 15102 8508 15108 8520
rect 15160 8508 15166 8560
rect 12452 8452 12940 8480
rect 12069 8415 12127 8421
rect 12069 8381 12081 8415
rect 12115 8412 12127 8415
rect 12802 8412 12808 8424
rect 12115 8384 12664 8412
rect 12763 8384 12808 8412
rect 12115 8381 12127 8384
rect 12069 8375 12127 8381
rect 10594 8304 10600 8356
rect 10652 8344 10658 8356
rect 11882 8344 11888 8356
rect 10652 8316 11888 8344
rect 10652 8304 10658 8316
rect 11882 8304 11888 8316
rect 11940 8344 11946 8356
rect 12084 8344 12112 8375
rect 12342 8344 12348 8356
rect 11940 8316 12112 8344
rect 12303 8316 12348 8344
rect 11940 8304 11946 8316
rect 12342 8304 12348 8316
rect 12400 8304 12406 8356
rect 12636 8344 12664 8384
rect 12802 8372 12808 8384
rect 12860 8372 12866 8424
rect 12912 8421 12940 8452
rect 13372 8452 13492 8480
rect 13556 8452 14044 8480
rect 14093 8483 14151 8489
rect 13372 8421 13400 8452
rect 12897 8415 12955 8421
rect 12897 8381 12909 8415
rect 12943 8381 12955 8415
rect 12897 8375 12955 8381
rect 13357 8415 13415 8421
rect 13357 8381 13369 8415
rect 13403 8381 13415 8415
rect 13357 8375 13415 8381
rect 13449 8415 13507 8421
rect 13449 8381 13461 8415
rect 13495 8412 13507 8415
rect 13556 8412 13584 8452
rect 14093 8449 14105 8483
rect 14139 8480 14151 8483
rect 14182 8480 14188 8492
rect 14139 8452 14188 8480
rect 14139 8449 14151 8452
rect 14093 8443 14151 8449
rect 14182 8440 14188 8452
rect 14240 8480 14246 8492
rect 14458 8480 14464 8492
rect 14240 8452 14464 8480
rect 14240 8440 14246 8452
rect 14458 8440 14464 8452
rect 14516 8440 14522 8492
rect 14660 8480 14688 8508
rect 14918 8480 14924 8492
rect 14660 8452 14924 8480
rect 14918 8440 14924 8452
rect 14976 8440 14982 8492
rect 13495 8384 13584 8412
rect 13495 8381 13507 8384
rect 13449 8375 13507 8381
rect 13630 8372 13636 8424
rect 13688 8412 13694 8424
rect 14645 8415 14703 8421
rect 14645 8412 14657 8415
rect 13688 8384 14657 8412
rect 13688 8372 13694 8384
rect 14645 8381 14657 8384
rect 14691 8381 14703 8415
rect 14645 8375 14703 8381
rect 14737 8415 14795 8421
rect 14737 8381 14749 8415
rect 14783 8381 14795 8415
rect 15102 8412 15108 8424
rect 15063 8384 15108 8412
rect 14737 8375 14795 8381
rect 14752 8344 14780 8375
rect 15102 8372 15108 8384
rect 15160 8372 15166 8424
rect 12636 8316 14780 8344
rect 15473 8347 15531 8353
rect 15473 8313 15485 8347
rect 15519 8344 15531 8347
rect 15654 8344 15660 8356
rect 15519 8316 15660 8344
rect 15519 8313 15531 8316
rect 15473 8307 15531 8313
rect 15654 8304 15660 8316
rect 15712 8304 15718 8356
rect 9398 8276 9404 8288
rect 7852 8248 9404 8276
rect 9398 8236 9404 8248
rect 9456 8236 9462 8288
rect 11330 8236 11336 8288
rect 11388 8276 11394 8288
rect 11517 8279 11575 8285
rect 11517 8276 11529 8279
rect 11388 8248 11529 8276
rect 11388 8236 11394 8248
rect 11517 8245 11529 8248
rect 11563 8245 11575 8279
rect 11517 8239 11575 8245
rect 13814 8236 13820 8288
rect 13872 8276 13878 8288
rect 13909 8279 13967 8285
rect 13909 8276 13921 8279
rect 13872 8248 13921 8276
rect 13872 8236 13878 8248
rect 13909 8245 13921 8248
rect 13955 8245 13967 8279
rect 13909 8239 13967 8245
rect 14366 8236 14372 8288
rect 14424 8276 14430 8288
rect 14642 8276 14648 8288
rect 14424 8248 14648 8276
rect 14424 8236 14430 8248
rect 14642 8236 14648 8248
rect 14700 8236 14706 8288
rect 1104 8186 16008 8208
rect 1104 8134 2824 8186
rect 2876 8134 2888 8186
rect 2940 8134 2952 8186
rect 3004 8134 3016 8186
rect 3068 8134 3080 8186
rect 3132 8134 6572 8186
rect 6624 8134 6636 8186
rect 6688 8134 6700 8186
rect 6752 8134 6764 8186
rect 6816 8134 6828 8186
rect 6880 8134 10320 8186
rect 10372 8134 10384 8186
rect 10436 8134 10448 8186
rect 10500 8134 10512 8186
rect 10564 8134 10576 8186
rect 10628 8134 14068 8186
rect 14120 8134 14132 8186
rect 14184 8134 14196 8186
rect 14248 8134 14260 8186
rect 14312 8134 14324 8186
rect 14376 8134 16008 8186
rect 1104 8112 16008 8134
rect 2130 8072 2136 8084
rect 2091 8044 2136 8072
rect 2130 8032 2136 8044
rect 2188 8032 2194 8084
rect 2240 8044 4016 8072
rect 2240 7945 2268 8044
rect 3605 8007 3663 8013
rect 3605 7973 3617 8007
rect 3651 8004 3663 8007
rect 3878 8004 3884 8016
rect 3651 7976 3884 8004
rect 3651 7973 3663 7976
rect 3605 7967 3663 7973
rect 3878 7964 3884 7976
rect 3936 7964 3942 8016
rect 1581 7939 1639 7945
rect 1581 7905 1593 7939
rect 1627 7905 1639 7939
rect 1581 7899 1639 7905
rect 2225 7939 2283 7945
rect 2225 7905 2237 7939
rect 2271 7905 2283 7939
rect 2225 7899 2283 7905
rect 1596 7868 1624 7899
rect 2489 7868 2495 7880
rect 1596 7840 2360 7868
rect 2450 7840 2495 7868
rect 1765 7803 1823 7809
rect 1765 7769 1777 7803
rect 1811 7800 1823 7803
rect 2332 7800 2360 7840
rect 2489 7828 2495 7840
rect 2547 7828 2553 7880
rect 3988 7877 4016 8044
rect 4816 8044 7696 8072
rect 4816 7936 4844 8044
rect 6288 8013 6316 8044
rect 6273 8007 6331 8013
rect 6273 7973 6285 8007
rect 6319 7973 6331 8007
rect 7668 8004 7696 8044
rect 9030 8032 9036 8084
rect 9088 8072 9094 8084
rect 9214 8072 9220 8084
rect 9088 8044 9220 8072
rect 9088 8032 9094 8044
rect 9214 8032 9220 8044
rect 9272 8072 9278 8084
rect 12529 8075 12587 8081
rect 9272 8044 10824 8072
rect 9272 8032 9278 8044
rect 9674 8004 9680 8016
rect 7668 7976 9680 8004
rect 6273 7967 6331 7973
rect 9674 7964 9680 7976
rect 9732 7964 9738 8016
rect 4816 7908 4936 7936
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7868 4031 7871
rect 4157 7871 4215 7877
rect 4157 7868 4169 7871
rect 4019 7840 4169 7868
rect 4019 7837 4031 7840
rect 3973 7831 4031 7837
rect 4157 7837 4169 7840
rect 4203 7868 4215 7871
rect 4341 7871 4399 7877
rect 4341 7868 4353 7871
rect 4203 7840 4353 7868
rect 4203 7837 4215 7840
rect 4157 7831 4215 7837
rect 4341 7837 4353 7840
rect 4387 7868 4399 7871
rect 4614 7868 4620 7880
rect 4387 7840 4620 7868
rect 4387 7837 4399 7840
rect 4341 7831 4399 7837
rect 4614 7828 4620 7840
rect 4672 7868 4678 7880
rect 4801 7871 4859 7877
rect 4801 7868 4813 7871
rect 4672 7840 4813 7868
rect 4672 7828 4678 7840
rect 4801 7837 4813 7840
rect 4847 7837 4859 7871
rect 4801 7831 4859 7837
rect 4908 7800 4936 7908
rect 7650 7896 7656 7948
rect 7708 7936 7714 7948
rect 9030 7936 9036 7948
rect 7708 7908 9036 7936
rect 7708 7896 7714 7908
rect 9030 7896 9036 7908
rect 9088 7896 9094 7948
rect 10796 7945 10824 8044
rect 12529 8041 12541 8075
rect 12575 8072 12587 8075
rect 12710 8072 12716 8084
rect 12575 8044 12716 8072
rect 12575 8041 12587 8044
rect 12529 8035 12587 8041
rect 12710 8032 12716 8044
rect 12768 8032 12774 8084
rect 13909 8075 13967 8081
rect 13909 8041 13921 8075
rect 13955 8072 13967 8075
rect 14458 8072 14464 8084
rect 13955 8044 14464 8072
rect 13955 8041 13967 8044
rect 13909 8035 13967 8041
rect 14458 8032 14464 8044
rect 14516 8072 14522 8084
rect 14734 8072 14740 8084
rect 14516 8044 14740 8072
rect 14516 8032 14522 8044
rect 14734 8032 14740 8044
rect 14792 8072 14798 8084
rect 15565 8075 15623 8081
rect 15565 8072 15577 8075
rect 14792 8044 15577 8072
rect 14792 8032 14798 8044
rect 15565 8041 15577 8044
rect 15611 8041 15623 8075
rect 15565 8035 15623 8041
rect 11330 7964 11336 8016
rect 11388 7964 11394 8016
rect 12066 8004 12072 8016
rect 12027 7976 12072 8004
rect 12066 7964 12072 7976
rect 12124 7964 12130 8016
rect 13814 7964 13820 8016
rect 13872 8004 13878 8016
rect 14277 8007 14335 8013
rect 14277 8004 14289 8007
rect 13872 7976 14289 8004
rect 13872 7964 13878 7976
rect 14277 7973 14289 7976
rect 14323 7973 14335 8007
rect 14277 7967 14335 7973
rect 10781 7939 10839 7945
rect 10781 7905 10793 7939
rect 10827 7905 10839 7939
rect 10781 7899 10839 7905
rect 7742 7828 7748 7880
rect 7800 7868 7806 7880
rect 7800 7840 9444 7868
rect 7800 7828 7806 7840
rect 1811 7772 2268 7800
rect 2332 7772 4936 7800
rect 5068 7803 5126 7809
rect 1811 7769 1823 7772
rect 1765 7763 1823 7769
rect 1670 7732 1676 7744
rect 1631 7704 1676 7732
rect 1670 7692 1676 7704
rect 1728 7692 1734 7744
rect 2240 7732 2268 7772
rect 5068 7769 5080 7803
rect 5114 7800 5126 7803
rect 5350 7800 5356 7812
rect 5114 7772 5356 7800
rect 5114 7769 5126 7772
rect 5068 7763 5126 7769
rect 5350 7760 5356 7772
rect 5408 7760 5414 7812
rect 5506 7772 7328 7800
rect 5506 7732 5534 7772
rect 2240 7704 5534 7732
rect 6181 7735 6239 7741
rect 6181 7701 6193 7735
rect 6227 7732 6239 7735
rect 6270 7732 6276 7744
rect 6227 7704 6276 7732
rect 6227 7701 6239 7704
rect 6181 7695 6239 7701
rect 6270 7692 6276 7704
rect 6328 7692 6334 7744
rect 7300 7732 7328 7772
rect 7374 7760 7380 7812
rect 7432 7809 7438 7812
rect 7432 7800 7444 7809
rect 7432 7772 7477 7800
rect 7432 7763 7444 7772
rect 7432 7760 7438 7763
rect 8294 7732 8300 7744
rect 7300 7704 8300 7732
rect 8294 7692 8300 7704
rect 8352 7692 8358 7744
rect 8573 7735 8631 7741
rect 8573 7701 8585 7735
rect 8619 7732 8631 7735
rect 8846 7732 8852 7744
rect 8619 7704 8852 7732
rect 8619 7701 8631 7704
rect 8573 7695 8631 7701
rect 8846 7692 8852 7704
rect 8904 7692 8910 7744
rect 9416 7741 9444 7840
rect 10134 7828 10140 7880
rect 10192 7868 10198 7880
rect 10525 7871 10583 7877
rect 10192 7840 10456 7868
rect 10192 7828 10198 7840
rect 10428 7812 10456 7840
rect 10525 7837 10537 7871
rect 10571 7868 10583 7871
rect 10962 7868 10968 7880
rect 10571 7840 10968 7868
rect 10571 7837 10583 7840
rect 10525 7831 10583 7837
rect 10962 7828 10968 7840
rect 11020 7828 11026 7880
rect 11348 7877 11376 7964
rect 11609 7939 11667 7945
rect 11609 7905 11621 7939
rect 11655 7936 11667 7939
rect 11790 7936 11796 7948
rect 11655 7908 11796 7936
rect 11655 7905 11667 7908
rect 11609 7899 11667 7905
rect 11790 7896 11796 7908
rect 11848 7896 11854 7948
rect 12158 7936 12164 7948
rect 12119 7908 12164 7936
rect 12158 7896 12164 7908
rect 12216 7896 12222 7948
rect 12894 7896 12900 7948
rect 12952 7936 12958 7948
rect 12989 7939 13047 7945
rect 12989 7936 13001 7939
rect 12952 7908 13001 7936
rect 12952 7896 12958 7908
rect 12989 7905 13001 7908
rect 13035 7905 13047 7939
rect 13170 7936 13176 7948
rect 13131 7908 13176 7936
rect 12989 7899 13047 7905
rect 13170 7896 13176 7908
rect 13228 7896 13234 7948
rect 13538 7896 13544 7948
rect 13596 7936 13602 7948
rect 13725 7939 13783 7945
rect 13725 7936 13737 7939
rect 13596 7908 13737 7936
rect 13596 7896 13602 7908
rect 13725 7905 13737 7908
rect 13771 7936 13783 7939
rect 13906 7936 13912 7948
rect 13771 7908 13912 7936
rect 13771 7905 13783 7908
rect 13725 7899 13783 7905
rect 13906 7896 13912 7908
rect 13964 7896 13970 7948
rect 14550 7936 14556 7948
rect 14108 7908 14556 7936
rect 14108 7880 14136 7908
rect 14550 7896 14556 7908
rect 14608 7936 14614 7948
rect 15289 7939 15347 7945
rect 15289 7936 15301 7939
rect 14608 7908 15301 7936
rect 14608 7896 14614 7908
rect 15289 7905 15301 7908
rect 15335 7905 15347 7939
rect 15289 7899 15347 7905
rect 11333 7871 11391 7877
rect 11333 7837 11345 7871
rect 11379 7837 11391 7871
rect 11333 7831 11391 7837
rect 11514 7828 11520 7880
rect 11572 7868 11578 7880
rect 14090 7868 14096 7880
rect 11572 7840 14096 7868
rect 11572 7828 11578 7840
rect 14090 7828 14096 7840
rect 14148 7828 14154 7880
rect 14366 7828 14372 7880
rect 14424 7868 14430 7880
rect 15102 7868 15108 7880
rect 14424 7840 14872 7868
rect 15063 7840 15108 7868
rect 14424 7828 14430 7840
rect 10410 7760 10416 7812
rect 10468 7760 10474 7812
rect 10686 7760 10692 7812
rect 10744 7800 10750 7812
rect 10870 7800 10876 7812
rect 10744 7772 10876 7800
rect 10744 7760 10750 7772
rect 10870 7760 10876 7772
rect 10928 7760 10934 7812
rect 12897 7803 12955 7809
rect 12897 7769 12909 7803
rect 12943 7800 12955 7803
rect 14844 7800 14872 7840
rect 15102 7828 15108 7840
rect 15160 7828 15166 7880
rect 15197 7803 15255 7809
rect 15197 7800 15209 7803
rect 12943 7772 14780 7800
rect 14844 7772 15209 7800
rect 12943 7769 12955 7772
rect 12897 7763 12955 7769
rect 9401 7735 9459 7741
rect 9401 7701 9413 7735
rect 9447 7701 9459 7735
rect 9401 7695 9459 7701
rect 9582 7692 9588 7744
rect 9640 7732 9646 7744
rect 10965 7735 11023 7741
rect 10965 7732 10977 7735
rect 9640 7704 10977 7732
rect 9640 7692 9646 7704
rect 10965 7701 10977 7704
rect 11011 7701 11023 7735
rect 11422 7732 11428 7744
rect 11383 7704 11428 7732
rect 10965 7695 11023 7701
rect 11422 7692 11428 7704
rect 11480 7692 11486 7744
rect 11606 7692 11612 7744
rect 11664 7732 11670 7744
rect 11793 7735 11851 7741
rect 11793 7732 11805 7735
rect 11664 7704 11805 7732
rect 11664 7692 11670 7704
rect 11793 7701 11805 7704
rect 11839 7701 11851 7735
rect 11793 7695 11851 7701
rect 12437 7735 12495 7741
rect 12437 7701 12449 7735
rect 12483 7732 12495 7735
rect 12526 7732 12532 7744
rect 12483 7704 12532 7732
rect 12483 7701 12495 7704
rect 12437 7695 12495 7701
rect 12526 7692 12532 7704
rect 12584 7692 12590 7744
rect 13446 7732 13452 7744
rect 13407 7704 13452 7732
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 13906 7692 13912 7744
rect 13964 7732 13970 7744
rect 14093 7735 14151 7741
rect 14093 7732 14105 7735
rect 13964 7704 14105 7732
rect 13964 7692 13970 7704
rect 14093 7701 14105 7704
rect 14139 7701 14151 7735
rect 14093 7695 14151 7701
rect 14366 7692 14372 7744
rect 14424 7732 14430 7744
rect 14752 7741 14780 7772
rect 15197 7769 15209 7772
rect 15243 7769 15255 7803
rect 15197 7763 15255 7769
rect 14553 7735 14611 7741
rect 14553 7732 14565 7735
rect 14424 7704 14565 7732
rect 14424 7692 14430 7704
rect 14553 7701 14565 7704
rect 14599 7701 14611 7735
rect 14553 7695 14611 7701
rect 14737 7735 14795 7741
rect 14737 7701 14749 7735
rect 14783 7701 14795 7735
rect 14737 7695 14795 7701
rect 1104 7642 16008 7664
rect 1104 7590 4698 7642
rect 4750 7590 4762 7642
rect 4814 7590 4826 7642
rect 4878 7590 4890 7642
rect 4942 7590 4954 7642
rect 5006 7590 8446 7642
rect 8498 7590 8510 7642
rect 8562 7590 8574 7642
rect 8626 7590 8638 7642
rect 8690 7590 8702 7642
rect 8754 7590 12194 7642
rect 12246 7590 12258 7642
rect 12310 7590 12322 7642
rect 12374 7590 12386 7642
rect 12438 7590 12450 7642
rect 12502 7590 16008 7642
rect 1104 7568 16008 7590
rect 1486 7528 1492 7540
rect 1447 7500 1492 7528
rect 1486 7488 1492 7500
rect 1544 7488 1550 7540
rect 1762 7528 1768 7540
rect 1723 7500 1768 7528
rect 1762 7488 1768 7500
rect 1820 7488 1826 7540
rect 6181 7531 6239 7537
rect 6181 7497 6193 7531
rect 6227 7528 6239 7531
rect 7469 7531 7527 7537
rect 7469 7528 7481 7531
rect 6227 7500 7481 7528
rect 6227 7497 6239 7500
rect 6181 7491 6239 7497
rect 7469 7497 7481 7500
rect 7515 7528 7527 7531
rect 7650 7528 7656 7540
rect 7515 7500 7656 7528
rect 7515 7497 7527 7500
rect 7469 7491 7527 7497
rect 3053 7463 3111 7469
rect 3053 7429 3065 7463
rect 3099 7460 3111 7463
rect 3099 7432 4568 7460
rect 3099 7429 3111 7432
rect 3053 7423 3111 7429
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7392 1731 7395
rect 1762 7392 1768 7404
rect 1719 7364 1768 7392
rect 1719 7361 1731 7364
rect 1673 7355 1731 7361
rect 1762 7352 1768 7364
rect 1820 7352 1826 7404
rect 1946 7392 1952 7404
rect 1907 7364 1952 7392
rect 1946 7352 1952 7364
rect 2004 7352 2010 7404
rect 3970 7352 3976 7404
rect 4028 7392 4034 7404
rect 4540 7401 4568 7432
rect 5534 7420 5540 7472
rect 5592 7460 5598 7472
rect 5730 7463 5788 7469
rect 5730 7460 5742 7463
rect 5592 7432 5742 7460
rect 5592 7420 5598 7432
rect 5730 7429 5742 7432
rect 5776 7429 5788 7463
rect 5730 7423 5788 7429
rect 4258 7395 4316 7401
rect 4258 7392 4270 7395
rect 4028 7364 4270 7392
rect 4028 7352 4034 7364
rect 4258 7361 4270 7364
rect 4304 7392 4316 7395
rect 4525 7395 4583 7401
rect 4304 7364 4476 7392
rect 4304 7361 4316 7364
rect 4258 7355 4316 7361
rect 4448 7324 4476 7364
rect 4525 7361 4537 7395
rect 4571 7392 4583 7395
rect 4614 7392 4620 7404
rect 4571 7364 4620 7392
rect 4571 7361 4583 7364
rect 4525 7355 4583 7361
rect 4614 7352 4620 7364
rect 4672 7392 4678 7404
rect 5997 7395 6055 7401
rect 5997 7392 6009 7395
rect 4672 7364 6009 7392
rect 4672 7352 4678 7364
rect 5997 7361 6009 7364
rect 6043 7392 6055 7395
rect 6196 7392 6224 7491
rect 7650 7488 7656 7500
rect 7708 7488 7714 7540
rect 9214 7528 9220 7540
rect 9175 7500 9220 7528
rect 9214 7488 9220 7500
rect 9272 7488 9278 7540
rect 9309 7531 9367 7537
rect 9309 7497 9321 7531
rect 9355 7528 9367 7531
rect 9398 7528 9404 7540
rect 9355 7500 9404 7528
rect 9355 7497 9367 7500
rect 9309 7491 9367 7497
rect 9398 7488 9404 7500
rect 9456 7488 9462 7540
rect 9950 7488 9956 7540
rect 10008 7528 10014 7540
rect 10962 7528 10968 7540
rect 10008 7500 10968 7528
rect 10008 7488 10014 7500
rect 10962 7488 10968 7500
rect 11020 7488 11026 7540
rect 11054 7488 11060 7540
rect 11112 7528 11118 7540
rect 11149 7531 11207 7537
rect 11149 7528 11161 7531
rect 11112 7500 11161 7528
rect 11112 7488 11118 7500
rect 11149 7497 11161 7500
rect 11195 7528 11207 7531
rect 11790 7528 11796 7540
rect 11195 7500 11796 7528
rect 11195 7497 11207 7500
rect 11149 7491 11207 7497
rect 11790 7488 11796 7500
rect 11848 7488 11854 7540
rect 11885 7531 11943 7537
rect 11885 7497 11897 7531
rect 11931 7528 11943 7531
rect 12158 7528 12164 7540
rect 11931 7500 12164 7528
rect 11931 7497 11943 7500
rect 11885 7491 11943 7497
rect 12158 7488 12164 7500
rect 12216 7488 12222 7540
rect 12342 7488 12348 7540
rect 12400 7528 12406 7540
rect 15473 7531 15531 7537
rect 15473 7528 15485 7531
rect 12400 7500 15485 7528
rect 12400 7488 12406 7500
rect 15473 7497 15485 7500
rect 15519 7497 15531 7531
rect 15473 7491 15531 7497
rect 6043 7364 6224 7392
rect 6043 7361 6055 7364
rect 5997 7355 6055 7361
rect 7190 7352 7196 7404
rect 7248 7392 7254 7404
rect 8478 7392 8484 7404
rect 7248 7364 8484 7392
rect 7248 7352 7254 7364
rect 8478 7352 8484 7364
rect 8536 7352 8542 7404
rect 8777 7395 8835 7401
rect 8777 7361 8789 7395
rect 8823 7392 8835 7395
rect 9033 7395 9091 7401
rect 8823 7364 8984 7392
rect 8823 7361 8835 7364
rect 8777 7355 8835 7361
rect 4448 7296 4660 7324
rect 4632 7265 4660 7296
rect 6454 7284 6460 7336
rect 6512 7324 6518 7336
rect 7834 7324 7840 7336
rect 6512 7296 7840 7324
rect 6512 7284 6518 7296
rect 7834 7284 7840 7296
rect 7892 7284 7898 7336
rect 8956 7324 8984 7364
rect 9033 7361 9045 7395
rect 9079 7392 9091 7395
rect 9232 7392 9260 7488
rect 10410 7420 10416 7472
rect 10468 7469 10474 7472
rect 10468 7460 10480 7469
rect 10980 7460 11008 7488
rect 12894 7460 12900 7472
rect 10468 7432 10513 7460
rect 10980 7432 12112 7460
rect 12855 7432 12900 7460
rect 10468 7423 10480 7432
rect 10468 7420 10474 7423
rect 10689 7395 10747 7401
rect 10689 7392 10701 7395
rect 9079 7364 10701 7392
rect 9079 7361 9091 7364
rect 9033 7355 9091 7361
rect 10689 7361 10701 7364
rect 10735 7361 10747 7395
rect 11238 7392 11244 7404
rect 10689 7355 10747 7361
rect 10888 7364 11244 7392
rect 9306 7324 9312 7336
rect 8956 7296 9312 7324
rect 9306 7284 9312 7296
rect 9364 7284 9370 7336
rect 4617 7259 4675 7265
rect 4617 7225 4629 7259
rect 4663 7225 4675 7259
rect 4617 7219 4675 7225
rect 7653 7259 7711 7265
rect 7653 7225 7665 7259
rect 7699 7256 7711 7259
rect 7926 7256 7932 7268
rect 7699 7228 7932 7256
rect 7699 7225 7711 7228
rect 7653 7219 7711 7225
rect 7926 7216 7932 7228
rect 7984 7216 7990 7268
rect 10686 7216 10692 7268
rect 10744 7256 10750 7268
rect 10888 7256 10916 7364
rect 11238 7352 11244 7364
rect 11296 7392 11302 7404
rect 11977 7395 12035 7401
rect 11977 7392 11989 7395
rect 11296 7364 11989 7392
rect 11296 7352 11302 7364
rect 11977 7361 11989 7364
rect 12023 7361 12035 7395
rect 11977 7355 12035 7361
rect 10965 7327 11023 7333
rect 10965 7293 10977 7327
rect 11011 7324 11023 7327
rect 11054 7324 11060 7336
rect 11011 7296 11060 7324
rect 11011 7293 11023 7296
rect 10965 7287 11023 7293
rect 11054 7284 11060 7296
rect 11112 7284 11118 7336
rect 11514 7284 11520 7336
rect 11572 7284 11578 7336
rect 12084 7333 12112 7432
rect 12894 7420 12900 7432
rect 12952 7460 12958 7472
rect 13078 7460 13084 7472
rect 12952 7432 13084 7460
rect 12952 7420 12958 7432
rect 13078 7420 13084 7432
rect 13136 7460 13142 7472
rect 14366 7460 14372 7472
rect 13136 7432 14372 7460
rect 13136 7420 13142 7432
rect 14366 7420 14372 7432
rect 14424 7420 14430 7472
rect 16758 7460 16764 7472
rect 14660 7432 16764 7460
rect 14553 7404 14611 7405
rect 12529 7395 12587 7401
rect 12529 7361 12541 7395
rect 12575 7392 12587 7395
rect 12710 7392 12716 7404
rect 12575 7364 12716 7392
rect 12575 7361 12587 7364
rect 12529 7355 12587 7361
rect 12710 7352 12716 7364
rect 12768 7392 12774 7404
rect 12986 7392 12992 7404
rect 12768 7364 12992 7392
rect 12768 7352 12774 7364
rect 12986 7352 12992 7364
rect 13044 7352 13050 7404
rect 13449 7395 13507 7401
rect 13449 7361 13461 7395
rect 13495 7392 13507 7395
rect 13538 7392 13544 7404
rect 13495 7364 13544 7392
rect 13495 7361 13507 7364
rect 13449 7355 13507 7361
rect 13538 7352 13544 7364
rect 13596 7352 13602 7404
rect 13909 7395 13967 7401
rect 13909 7361 13921 7395
rect 13955 7361 13967 7395
rect 13909 7355 13967 7361
rect 14001 7395 14059 7401
rect 14001 7361 14013 7395
rect 14047 7392 14059 7395
rect 14458 7392 14464 7404
rect 14047 7364 14464 7392
rect 14047 7361 14059 7364
rect 14001 7355 14059 7361
rect 12069 7327 12127 7333
rect 12069 7293 12081 7327
rect 12115 7293 12127 7327
rect 12069 7287 12127 7293
rect 11532 7256 11560 7284
rect 10744 7228 10916 7256
rect 10980 7228 11560 7256
rect 10744 7216 10750 7228
rect 3142 7188 3148 7200
rect 3103 7160 3148 7188
rect 3142 7148 3148 7160
rect 3200 7148 3206 7200
rect 6362 7148 6368 7200
rect 6420 7188 6426 7200
rect 10980 7188 11008 7228
rect 12618 7216 12624 7268
rect 12676 7256 12682 7268
rect 12713 7259 12771 7265
rect 12713 7256 12725 7259
rect 12676 7228 12725 7256
rect 12676 7216 12682 7228
rect 12713 7225 12725 7228
rect 12759 7256 12771 7259
rect 12894 7256 12900 7268
rect 12759 7228 12900 7256
rect 12759 7225 12771 7228
rect 12713 7219 12771 7225
rect 12894 7216 12900 7228
rect 12952 7216 12958 7268
rect 13265 7259 13323 7265
rect 13265 7225 13277 7259
rect 13311 7256 13323 7259
rect 13446 7256 13452 7268
rect 13311 7228 13452 7256
rect 13311 7225 13323 7228
rect 13265 7219 13323 7225
rect 13446 7216 13452 7228
rect 13504 7216 13510 7268
rect 13924 7256 13952 7355
rect 14458 7352 14464 7364
rect 14516 7352 14522 7404
rect 14550 7352 14556 7404
rect 14608 7392 14614 7404
rect 14660 7392 14688 7432
rect 16758 7420 16764 7432
rect 16816 7420 16822 7472
rect 15013 7395 15071 7401
rect 14608 7364 14701 7392
rect 14608 7352 14614 7364
rect 15013 7361 15025 7395
rect 15059 7361 15071 7395
rect 15013 7355 15071 7361
rect 15105 7395 15163 7401
rect 15105 7361 15117 7395
rect 15151 7392 15163 7395
rect 15286 7392 15292 7404
rect 15151 7364 15292 7392
rect 15151 7361 15163 7364
rect 15105 7355 15163 7361
rect 14090 7324 14096 7336
rect 14051 7296 14096 7324
rect 14090 7284 14096 7296
rect 14148 7324 14154 7336
rect 15028 7324 15056 7355
rect 15286 7352 15292 7364
rect 15344 7352 15350 7404
rect 15562 7352 15568 7404
rect 15620 7392 15626 7404
rect 15657 7395 15715 7401
rect 15657 7392 15669 7395
rect 15620 7364 15669 7392
rect 15620 7352 15626 7364
rect 15657 7361 15669 7364
rect 15703 7361 15715 7395
rect 15657 7355 15715 7361
rect 15197 7327 15255 7333
rect 14148 7296 14964 7324
rect 15028 7296 15148 7324
rect 14148 7284 14154 7296
rect 14550 7256 14556 7268
rect 13924 7228 14556 7256
rect 14550 7216 14556 7228
rect 14608 7216 14614 7268
rect 11330 7188 11336 7200
rect 6420 7160 11008 7188
rect 11291 7160 11336 7188
rect 6420 7148 6426 7160
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 11514 7188 11520 7200
rect 11475 7160 11520 7188
rect 11514 7148 11520 7160
rect 11572 7148 11578 7200
rect 13078 7188 13084 7200
rect 13039 7160 13084 7188
rect 13078 7148 13084 7160
rect 13136 7148 13142 7200
rect 13538 7188 13544 7200
rect 13499 7160 13544 7188
rect 13538 7148 13544 7160
rect 13596 7148 13602 7200
rect 14366 7188 14372 7200
rect 14327 7160 14372 7188
rect 14366 7148 14372 7160
rect 14424 7148 14430 7200
rect 14642 7188 14648 7200
rect 14603 7160 14648 7188
rect 14642 7148 14648 7160
rect 14700 7148 14706 7200
rect 14936 7188 14964 7296
rect 15120 7268 15148 7296
rect 15197 7293 15209 7327
rect 15243 7293 15255 7327
rect 15197 7287 15255 7293
rect 15102 7216 15108 7268
rect 15160 7216 15166 7268
rect 15212 7188 15240 7287
rect 14936 7160 15240 7188
rect 1104 7098 16008 7120
rect 1104 7046 2824 7098
rect 2876 7046 2888 7098
rect 2940 7046 2952 7098
rect 3004 7046 3016 7098
rect 3068 7046 3080 7098
rect 3132 7046 6572 7098
rect 6624 7046 6636 7098
rect 6688 7046 6700 7098
rect 6752 7046 6764 7098
rect 6816 7046 6828 7098
rect 6880 7046 10320 7098
rect 10372 7046 10384 7098
rect 10436 7046 10448 7098
rect 10500 7046 10512 7098
rect 10564 7046 10576 7098
rect 10628 7046 14068 7098
rect 14120 7046 14132 7098
rect 14184 7046 14196 7098
rect 14248 7046 14260 7098
rect 14312 7046 14324 7098
rect 14376 7046 16008 7098
rect 1104 7024 16008 7046
rect 4525 6987 4583 6993
rect 4525 6953 4537 6987
rect 4571 6984 4583 6987
rect 4614 6984 4620 6996
rect 4571 6956 4620 6984
rect 4571 6953 4583 6956
rect 4525 6947 4583 6953
rect 4614 6944 4620 6956
rect 4672 6944 4678 6996
rect 6457 6987 6515 6993
rect 6457 6953 6469 6987
rect 6503 6984 6515 6987
rect 7558 6984 7564 6996
rect 6503 6956 7564 6984
rect 6503 6953 6515 6956
rect 6457 6947 6515 6953
rect 2590 6876 2596 6928
rect 2648 6916 2654 6928
rect 3418 6916 3424 6928
rect 2648 6888 3424 6916
rect 2648 6876 2654 6888
rect 3418 6876 3424 6888
rect 3476 6876 3482 6928
rect 1946 6848 1952 6860
rect 1907 6820 1952 6848
rect 1946 6808 1952 6820
rect 2004 6808 2010 6860
rect 6564 6857 6592 6956
rect 7558 6944 7564 6956
rect 7616 6944 7622 6996
rect 8021 6987 8079 6993
rect 8021 6984 8033 6987
rect 7944 6956 8033 6984
rect 7650 6876 7656 6928
rect 7708 6916 7714 6928
rect 7944 6916 7972 6956
rect 8021 6953 8033 6956
rect 8067 6953 8079 6987
rect 8386 6984 8392 6996
rect 8299 6956 8392 6984
rect 8021 6947 8079 6953
rect 8386 6944 8392 6956
rect 8444 6984 8450 6996
rect 9214 6984 9220 6996
rect 8444 6956 9220 6984
rect 8444 6944 8450 6956
rect 9214 6944 9220 6956
rect 9272 6944 9278 6996
rect 10962 6944 10968 6996
rect 11020 6944 11026 6996
rect 11149 6987 11207 6993
rect 11149 6953 11161 6987
rect 11195 6984 11207 6987
rect 11422 6984 11428 6996
rect 11195 6956 11428 6984
rect 11195 6953 11207 6956
rect 11149 6947 11207 6953
rect 11422 6944 11428 6956
rect 11480 6944 11486 6996
rect 11790 6944 11796 6996
rect 11848 6984 11854 6996
rect 13814 6984 13820 6996
rect 11848 6956 13820 6984
rect 11848 6944 11854 6956
rect 13814 6944 13820 6956
rect 13872 6984 13878 6996
rect 14182 6984 14188 6996
rect 13872 6956 14188 6984
rect 13872 6944 13878 6956
rect 14182 6944 14188 6956
rect 14240 6944 14246 6996
rect 15102 6984 15108 6996
rect 14292 6956 15108 6984
rect 8481 6919 8539 6925
rect 8481 6916 8493 6919
rect 7708 6888 7972 6916
rect 8036 6888 8493 6916
rect 7708 6876 7714 6888
rect 6549 6851 6607 6857
rect 6549 6817 6561 6851
rect 6595 6817 6607 6851
rect 6549 6811 6607 6817
rect 7558 6808 7564 6860
rect 7616 6848 7622 6860
rect 7926 6848 7932 6860
rect 7616 6820 7932 6848
rect 7616 6808 7622 6820
rect 7926 6808 7932 6820
rect 7984 6808 7990 6860
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 3418 6780 3424 6792
rect 1719 6752 3424 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 3418 6740 3424 6752
rect 3476 6740 3482 6792
rect 6638 6740 6644 6792
rect 6696 6780 6702 6792
rect 6805 6783 6863 6789
rect 6805 6780 6817 6783
rect 6696 6752 6817 6780
rect 6696 6740 6702 6752
rect 6805 6749 6817 6752
rect 6851 6749 6863 6783
rect 8036 6780 8064 6888
rect 8481 6885 8493 6888
rect 8527 6885 8539 6919
rect 8481 6879 8539 6885
rect 8757 6919 8815 6925
rect 8757 6885 8769 6919
rect 8803 6916 8815 6919
rect 9674 6916 9680 6928
rect 8803 6888 9680 6916
rect 8803 6885 8815 6888
rect 8757 6879 8815 6885
rect 9674 6876 9680 6888
rect 9732 6916 9738 6928
rect 10226 6916 10232 6928
rect 9732 6888 10232 6916
rect 9732 6876 9738 6888
rect 10226 6876 10232 6888
rect 10284 6916 10290 6928
rect 10873 6919 10931 6925
rect 10873 6916 10885 6919
rect 10284 6888 10885 6916
rect 10284 6876 10290 6888
rect 10873 6885 10885 6888
rect 10919 6885 10931 6919
rect 10873 6879 10931 6885
rect 9122 6848 9128 6860
rect 6805 6743 6863 6749
rect 7024 6752 8064 6780
rect 8128 6820 9128 6848
rect 2222 6712 2228 6724
rect 2183 6684 2228 6712
rect 2222 6672 2228 6684
rect 2280 6672 2286 6724
rect 5442 6672 5448 6724
rect 5500 6712 5506 6724
rect 7024 6712 7052 6752
rect 8128 6712 8156 6820
rect 9122 6808 9128 6820
rect 9180 6808 9186 6860
rect 9490 6808 9496 6860
rect 9548 6848 9554 6860
rect 9858 6848 9864 6860
rect 9548 6820 9593 6848
rect 9819 6820 9864 6848
rect 9548 6808 9554 6820
rect 9858 6808 9864 6820
rect 9916 6808 9922 6860
rect 10980 6848 11008 6944
rect 11882 6916 11888 6928
rect 11716 6888 11888 6916
rect 11330 6848 11336 6860
rect 10704 6820 11336 6848
rect 8205 6759 8263 6765
rect 8205 6725 8217 6759
rect 8251 6725 8263 6759
rect 8478 6740 8484 6792
rect 8536 6780 8542 6792
rect 8536 6752 8984 6780
rect 8536 6740 8542 6752
rect 8205 6719 8263 6725
rect 5500 6684 7052 6712
rect 7944 6684 8156 6712
rect 5500 6672 5506 6684
rect 1486 6644 1492 6656
rect 1447 6616 1492 6644
rect 1486 6604 1492 6616
rect 1544 6604 1550 6656
rect 2133 6647 2191 6653
rect 2133 6613 2145 6647
rect 2179 6644 2191 6647
rect 2498 6644 2504 6656
rect 2179 6616 2504 6644
rect 2179 6613 2191 6616
rect 2133 6607 2191 6613
rect 2498 6604 2504 6616
rect 2556 6604 2562 6656
rect 2593 6647 2651 6653
rect 2593 6613 2605 6647
rect 2639 6644 2651 6647
rect 2682 6644 2688 6656
rect 2639 6616 2688 6644
rect 2639 6613 2651 6616
rect 2593 6607 2651 6613
rect 2682 6604 2688 6616
rect 2740 6604 2746 6656
rect 3602 6604 3608 6656
rect 3660 6644 3666 6656
rect 5626 6644 5632 6656
rect 3660 6616 5632 6644
rect 3660 6604 3666 6616
rect 5626 6604 5632 6616
rect 5684 6604 5690 6656
rect 6914 6604 6920 6656
rect 6972 6644 6978 6656
rect 7190 6644 7196 6656
rect 6972 6616 7196 6644
rect 6972 6604 6978 6616
rect 7190 6604 7196 6616
rect 7248 6604 7254 6656
rect 7944 6653 7972 6684
rect 7929 6647 7987 6653
rect 7929 6613 7941 6647
rect 7975 6613 7987 6647
rect 8220 6644 8248 6719
rect 8754 6644 8760 6656
rect 8220 6616 8760 6644
rect 7929 6607 7987 6613
rect 8754 6604 8760 6616
rect 8812 6604 8818 6656
rect 8956 6653 8984 6752
rect 9140 6712 9168 6808
rect 10704 6792 10732 6820
rect 11330 6808 11336 6820
rect 11388 6808 11394 6860
rect 11716 6857 11744 6888
rect 11882 6876 11888 6888
rect 11940 6876 11946 6928
rect 11701 6851 11759 6857
rect 11701 6817 11713 6851
rect 11747 6817 11759 6851
rect 11701 6811 11759 6817
rect 11790 6808 11796 6860
rect 11848 6848 11854 6860
rect 12529 6851 12587 6857
rect 12529 6848 12541 6851
rect 11848 6820 12541 6848
rect 11848 6808 11854 6820
rect 12529 6817 12541 6820
rect 12575 6817 12587 6851
rect 13170 6848 13176 6860
rect 13083 6820 13176 6848
rect 12529 6811 12587 6817
rect 13170 6808 13176 6820
rect 13228 6848 13234 6860
rect 13357 6851 13415 6857
rect 13357 6848 13369 6851
rect 13228 6820 13369 6848
rect 13228 6808 13234 6820
rect 13357 6817 13369 6820
rect 13403 6817 13415 6851
rect 13357 6811 13415 6817
rect 13998 6808 14004 6860
rect 14056 6848 14062 6860
rect 14292 6848 14320 6956
rect 15102 6944 15108 6956
rect 15160 6944 15166 6996
rect 14366 6876 14372 6928
rect 14424 6916 14430 6928
rect 14734 6916 14740 6928
rect 14424 6888 14740 6916
rect 14424 6876 14430 6888
rect 14734 6876 14740 6888
rect 14792 6876 14798 6928
rect 14461 6851 14519 6857
rect 14461 6848 14473 6851
rect 14056 6820 14473 6848
rect 14056 6808 14062 6820
rect 14461 6817 14473 6820
rect 14507 6817 14519 6851
rect 14461 6811 14519 6817
rect 14829 6851 14887 6857
rect 14829 6817 14841 6851
rect 14875 6848 14887 6851
rect 15838 6848 15844 6860
rect 14875 6820 15844 6848
rect 14875 6817 14887 6820
rect 14829 6811 14887 6817
rect 15838 6808 15844 6820
rect 15896 6808 15902 6860
rect 9214 6740 9220 6792
rect 9272 6780 9278 6792
rect 9401 6783 9459 6789
rect 9401 6780 9413 6783
rect 9272 6752 9413 6780
rect 9272 6740 9278 6752
rect 9401 6749 9413 6752
rect 9447 6749 9459 6783
rect 9401 6743 9459 6749
rect 10686 6740 10692 6792
rect 10744 6740 10750 6792
rect 10781 6783 10839 6789
rect 10781 6749 10793 6783
rect 10827 6780 10839 6783
rect 10870 6780 10876 6792
rect 10827 6752 10876 6780
rect 10827 6749 10839 6752
rect 10781 6743 10839 6749
rect 10870 6740 10876 6752
rect 10928 6740 10934 6792
rect 11514 6780 11520 6792
rect 11475 6752 11520 6780
rect 11514 6740 11520 6752
rect 11572 6740 11578 6792
rect 13188 6780 13216 6808
rect 12268 6752 13216 6780
rect 13265 6783 13323 6789
rect 12268 6712 12296 6752
rect 13265 6749 13277 6783
rect 13311 6780 13323 6783
rect 13538 6780 13544 6792
rect 13311 6752 13544 6780
rect 13311 6749 13323 6752
rect 13265 6743 13323 6749
rect 13538 6740 13544 6752
rect 13596 6740 13602 6792
rect 13814 6740 13820 6792
rect 13872 6740 13878 6792
rect 13909 6783 13967 6789
rect 13909 6749 13921 6783
rect 13955 6749 13967 6783
rect 13909 6743 13967 6749
rect 9140 6684 12296 6712
rect 12345 6715 12403 6721
rect 12345 6681 12357 6715
rect 12391 6712 12403 6715
rect 12986 6712 12992 6724
rect 12391 6684 12992 6712
rect 12391 6681 12403 6684
rect 12345 6675 12403 6681
rect 12986 6672 12992 6684
rect 13044 6672 13050 6724
rect 13173 6715 13231 6721
rect 13173 6681 13185 6715
rect 13219 6712 13231 6715
rect 13832 6712 13860 6740
rect 13219 6684 13860 6712
rect 13924 6712 13952 6743
rect 14090 6740 14096 6792
rect 14148 6740 14154 6792
rect 14274 6740 14280 6792
rect 14332 6780 14338 6792
rect 14553 6783 14611 6789
rect 14332 6752 14504 6780
rect 14332 6740 14338 6752
rect 14108 6712 14136 6740
rect 13924 6684 14136 6712
rect 13219 6681 13231 6684
rect 13173 6675 13231 6681
rect 8941 6647 8999 6653
rect 8941 6613 8953 6647
rect 8987 6613 8999 6647
rect 8941 6607 8999 6613
rect 9122 6604 9128 6656
rect 9180 6644 9186 6656
rect 9309 6647 9367 6653
rect 9309 6644 9321 6647
rect 9180 6616 9321 6644
rect 9180 6604 9186 6616
rect 9309 6613 9321 6616
rect 9355 6613 9367 6647
rect 9309 6607 9367 6613
rect 9398 6604 9404 6656
rect 9456 6644 9462 6656
rect 9582 6644 9588 6656
rect 9456 6616 9588 6644
rect 9456 6604 9462 6616
rect 9582 6604 9588 6616
rect 9640 6644 9646 6656
rect 10134 6644 10140 6656
rect 9640 6616 10140 6644
rect 9640 6604 9646 6616
rect 10134 6604 10140 6616
rect 10192 6604 10198 6656
rect 10226 6604 10232 6656
rect 10284 6644 10290 6656
rect 10321 6647 10379 6653
rect 10321 6644 10333 6647
rect 10284 6616 10333 6644
rect 10284 6604 10290 6616
rect 10321 6613 10333 6616
rect 10367 6613 10379 6647
rect 10321 6607 10379 6613
rect 10597 6647 10655 6653
rect 10597 6613 10609 6647
rect 10643 6644 10655 6647
rect 10686 6644 10692 6656
rect 10643 6616 10692 6644
rect 10643 6613 10655 6616
rect 10597 6607 10655 6613
rect 10686 6604 10692 6616
rect 10744 6604 10750 6656
rect 11609 6647 11667 6653
rect 11609 6613 11621 6647
rect 11655 6644 11667 6647
rect 11790 6644 11796 6656
rect 11655 6616 11796 6644
rect 11655 6613 11667 6616
rect 11609 6607 11667 6613
rect 11790 6604 11796 6616
rect 11848 6604 11854 6656
rect 11882 6604 11888 6656
rect 11940 6644 11946 6656
rect 11977 6647 12035 6653
rect 11977 6644 11989 6647
rect 11940 6616 11989 6644
rect 11940 6604 11946 6616
rect 11977 6613 11989 6616
rect 12023 6613 12035 6647
rect 11977 6607 12035 6613
rect 12437 6647 12495 6653
rect 12437 6613 12449 6647
rect 12483 6644 12495 6647
rect 12618 6644 12624 6656
rect 12483 6616 12624 6644
rect 12483 6613 12495 6616
rect 12437 6607 12495 6613
rect 12618 6604 12624 6616
rect 12676 6604 12682 6656
rect 12802 6644 12808 6656
rect 12763 6616 12808 6644
rect 12802 6604 12808 6616
rect 12860 6604 12866 6656
rect 13630 6604 13636 6656
rect 13688 6644 13694 6656
rect 13725 6647 13783 6653
rect 13725 6644 13737 6647
rect 13688 6616 13737 6644
rect 13688 6604 13694 6616
rect 13725 6613 13737 6616
rect 13771 6613 13783 6647
rect 13725 6607 13783 6613
rect 13814 6604 13820 6656
rect 13872 6644 13878 6656
rect 14093 6647 14151 6653
rect 14093 6644 14105 6647
rect 13872 6616 14105 6644
rect 13872 6604 13878 6616
rect 14093 6613 14105 6616
rect 14139 6613 14151 6647
rect 14476 6644 14504 6752
rect 14553 6749 14565 6783
rect 14599 6780 14611 6783
rect 14734 6780 14740 6792
rect 14599 6752 14740 6780
rect 14599 6749 14611 6752
rect 14553 6743 14611 6749
rect 14734 6740 14740 6752
rect 14792 6740 14798 6792
rect 15102 6780 15108 6792
rect 15063 6752 15108 6780
rect 15102 6740 15108 6752
rect 15160 6740 15166 6792
rect 14737 6647 14795 6653
rect 14737 6644 14749 6647
rect 14476 6616 14749 6644
rect 14093 6607 14151 6613
rect 14737 6613 14749 6616
rect 14783 6644 14795 6647
rect 15746 6644 15752 6656
rect 14783 6616 15752 6644
rect 14783 6613 14795 6616
rect 14737 6607 14795 6613
rect 15746 6604 15752 6616
rect 15804 6604 15810 6656
rect 1104 6554 16008 6576
rect 1104 6502 4698 6554
rect 4750 6502 4762 6554
rect 4814 6502 4826 6554
rect 4878 6502 4890 6554
rect 4942 6502 4954 6554
rect 5006 6502 8446 6554
rect 8498 6502 8510 6554
rect 8562 6502 8574 6554
rect 8626 6502 8638 6554
rect 8690 6502 8702 6554
rect 8754 6502 12194 6554
rect 12246 6502 12258 6554
rect 12310 6502 12322 6554
rect 12374 6502 12386 6554
rect 12438 6502 12450 6554
rect 12502 6502 16008 6554
rect 1104 6480 16008 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 1670 6440 1676 6452
rect 1627 6412 1676 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 1670 6400 1676 6412
rect 1728 6400 1734 6452
rect 1949 6443 2007 6449
rect 1949 6409 1961 6443
rect 1995 6440 2007 6443
rect 2961 6443 3019 6449
rect 2961 6440 2973 6443
rect 1995 6412 2973 6440
rect 1995 6409 2007 6412
rect 1949 6403 2007 6409
rect 2961 6409 2973 6412
rect 3007 6409 3019 6443
rect 2961 6403 3019 6409
rect 3329 6443 3387 6449
rect 3329 6409 3341 6443
rect 3375 6440 3387 6443
rect 3881 6443 3939 6449
rect 3881 6440 3893 6443
rect 3375 6412 3893 6440
rect 3375 6409 3387 6412
rect 3329 6403 3387 6409
rect 3881 6409 3893 6412
rect 3927 6440 3939 6443
rect 4246 6440 4252 6452
rect 3927 6412 4252 6440
rect 3927 6409 3939 6412
rect 3881 6403 3939 6409
rect 4246 6400 4252 6412
rect 4304 6440 4310 6452
rect 4614 6440 4620 6452
rect 4304 6412 4620 6440
rect 4304 6400 4310 6412
rect 4614 6400 4620 6412
rect 4672 6400 4678 6452
rect 4706 6400 4712 6452
rect 4764 6440 4770 6452
rect 5166 6440 5172 6452
rect 4764 6412 5172 6440
rect 4764 6400 4770 6412
rect 5166 6400 5172 6412
rect 5224 6400 5230 6452
rect 5626 6400 5632 6452
rect 5684 6440 5690 6452
rect 5684 6412 5729 6440
rect 5684 6400 5690 6412
rect 5902 6400 5908 6452
rect 5960 6440 5966 6452
rect 6181 6443 6239 6449
rect 6181 6440 6193 6443
rect 5960 6412 6193 6440
rect 5960 6400 5966 6412
rect 6181 6409 6193 6412
rect 6227 6440 6239 6443
rect 6454 6440 6460 6452
rect 6227 6412 6460 6440
rect 6227 6409 6239 6412
rect 6181 6403 6239 6409
rect 6454 6400 6460 6412
rect 6512 6400 6518 6452
rect 7009 6443 7067 6449
rect 7009 6409 7021 6443
rect 7055 6440 7067 6443
rect 7742 6440 7748 6452
rect 7055 6412 7748 6440
rect 7055 6409 7067 6412
rect 7009 6403 7067 6409
rect 7742 6400 7748 6412
rect 7800 6400 7806 6452
rect 9030 6400 9036 6452
rect 9088 6440 9094 6452
rect 10042 6440 10048 6452
rect 9088 6412 10048 6440
rect 9088 6400 9094 6412
rect 10042 6400 10048 6412
rect 10100 6440 10106 6452
rect 10597 6443 10655 6449
rect 10597 6440 10609 6443
rect 10100 6412 10609 6440
rect 10100 6400 10106 6412
rect 10597 6409 10609 6412
rect 10643 6409 10655 6443
rect 10597 6403 10655 6409
rect 10965 6443 11023 6449
rect 10965 6409 10977 6443
rect 11011 6409 11023 6443
rect 10965 6403 11023 6409
rect 11149 6443 11207 6449
rect 11149 6409 11161 6443
rect 11195 6440 11207 6443
rect 11238 6440 11244 6452
rect 11195 6412 11244 6440
rect 11195 6409 11207 6412
rect 11149 6403 11207 6409
rect 3510 6332 3516 6384
rect 3568 6372 3574 6384
rect 4982 6372 4988 6384
rect 3568 6344 4988 6372
rect 3568 6332 3574 6344
rect 4982 6332 4988 6344
rect 5040 6372 5046 6384
rect 5442 6372 5448 6384
rect 5040 6344 5448 6372
rect 5040 6332 5046 6344
rect 5442 6332 5448 6344
rect 5500 6332 5506 6384
rect 6914 6332 6920 6384
rect 6972 6372 6978 6384
rect 7653 6375 7711 6381
rect 7653 6372 7665 6375
rect 6972 6344 7665 6372
rect 6972 6332 6978 6344
rect 7653 6341 7665 6344
rect 7699 6341 7711 6375
rect 7834 6372 7840 6384
rect 7795 6344 7840 6372
rect 7653 6335 7711 6341
rect 7834 6332 7840 6344
rect 7892 6332 7898 6384
rect 8202 6381 8208 6384
rect 8196 6335 8208 6381
rect 8260 6372 8266 6384
rect 8260 6344 8296 6372
rect 8202 6332 8208 6335
rect 8260 6332 8266 6344
rect 8846 6332 8852 6384
rect 8904 6372 8910 6384
rect 9766 6372 9772 6384
rect 8904 6344 9772 6372
rect 8904 6332 8910 6344
rect 9766 6332 9772 6344
rect 9824 6332 9830 6384
rect 9861 6375 9919 6381
rect 9861 6341 9873 6375
rect 9907 6372 9919 6375
rect 10318 6372 10324 6384
rect 9907 6344 10324 6372
rect 9907 6341 9919 6344
rect 9861 6335 9919 6341
rect 10318 6332 10324 6344
rect 10376 6332 10382 6384
rect 10980 6372 11008 6403
rect 11238 6400 11244 6412
rect 11296 6400 11302 6452
rect 12066 6400 12072 6452
rect 12124 6440 12130 6452
rect 12253 6443 12311 6449
rect 12253 6440 12265 6443
rect 12124 6412 12265 6440
rect 12124 6400 12130 6412
rect 12253 6409 12265 6412
rect 12299 6409 12311 6443
rect 12618 6440 12624 6452
rect 12579 6412 12624 6440
rect 12253 6403 12311 6409
rect 12618 6400 12624 6412
rect 12676 6400 12682 6452
rect 12986 6400 12992 6452
rect 13044 6440 13050 6452
rect 13449 6443 13507 6449
rect 13449 6440 13461 6443
rect 13044 6412 13461 6440
rect 13044 6400 13050 6412
rect 13449 6409 13461 6412
rect 13495 6409 13507 6443
rect 13814 6440 13820 6452
rect 13775 6412 13820 6440
rect 13449 6403 13507 6409
rect 13814 6400 13820 6412
rect 13872 6400 13878 6452
rect 13909 6443 13967 6449
rect 13909 6409 13921 6443
rect 13955 6440 13967 6443
rect 14090 6440 14096 6452
rect 13955 6412 14096 6440
rect 13955 6409 13967 6412
rect 13909 6403 13967 6409
rect 14090 6400 14096 6412
rect 14148 6400 14154 6452
rect 14461 6443 14519 6449
rect 14461 6409 14473 6443
rect 14507 6440 14519 6443
rect 14642 6440 14648 6452
rect 14507 6412 14648 6440
rect 14507 6409 14519 6412
rect 14461 6403 14519 6409
rect 14642 6400 14648 6412
rect 14700 6400 14706 6452
rect 14918 6440 14924 6452
rect 14879 6412 14924 6440
rect 14918 6400 14924 6412
rect 14976 6400 14982 6452
rect 15286 6440 15292 6452
rect 15247 6412 15292 6440
rect 15286 6400 15292 6412
rect 15344 6400 15350 6452
rect 10980 6344 11284 6372
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6304 3479 6307
rect 3878 6304 3884 6316
rect 3467 6276 3884 6304
rect 3467 6273 3479 6276
rect 3421 6267 3479 6273
rect 3878 6264 3884 6276
rect 3936 6264 3942 6316
rect 4062 6264 4068 6316
rect 4120 6304 4126 6316
rect 5534 6304 5540 6316
rect 4120 6276 5540 6304
rect 4120 6264 4126 6276
rect 5534 6264 5540 6276
rect 5592 6264 5598 6316
rect 6457 6307 6515 6313
rect 6457 6273 6469 6307
rect 6503 6304 6515 6307
rect 7006 6304 7012 6316
rect 6503 6276 7012 6304
rect 6503 6273 6515 6276
rect 6457 6267 6515 6273
rect 7006 6264 7012 6276
rect 7064 6264 7070 6316
rect 7098 6264 7104 6316
rect 7156 6304 7162 6316
rect 7156 6276 7201 6304
rect 7156 6264 7162 6276
rect 7374 6264 7380 6316
rect 7432 6304 7438 6316
rect 7929 6307 7987 6313
rect 7929 6304 7941 6307
rect 7432 6276 7941 6304
rect 7432 6264 7438 6276
rect 7929 6273 7941 6276
rect 7975 6273 7987 6307
rect 8312 6304 8432 6308
rect 7929 6267 7987 6273
rect 8036 6280 8984 6304
rect 8036 6276 8340 6280
rect 8404 6276 8984 6280
rect 2038 6236 2044 6248
rect 1999 6208 2044 6236
rect 2038 6196 2044 6208
rect 2096 6196 2102 6248
rect 2225 6239 2283 6245
rect 2225 6205 2237 6239
rect 2271 6236 2283 6239
rect 2314 6236 2320 6248
rect 2271 6208 2320 6236
rect 2271 6205 2283 6208
rect 2225 6199 2283 6205
rect 2314 6196 2320 6208
rect 2372 6196 2378 6248
rect 3605 6239 3663 6245
rect 3605 6205 3617 6239
rect 3651 6205 3663 6239
rect 3605 6199 3663 6205
rect 3142 6128 3148 6180
rect 3200 6168 3206 6180
rect 3620 6168 3648 6199
rect 4522 6196 4528 6248
rect 4580 6236 4586 6248
rect 5442 6236 5448 6248
rect 4580 6208 5448 6236
rect 4580 6196 4586 6208
rect 5442 6196 5448 6208
rect 5500 6196 5506 6248
rect 5810 6236 5816 6248
rect 5771 6208 5816 6236
rect 5810 6196 5816 6208
rect 5868 6196 5874 6248
rect 6822 6236 6828 6248
rect 6783 6208 6828 6236
rect 6822 6196 6828 6208
rect 6880 6196 6886 6248
rect 8036 6236 8064 6276
rect 7116 6208 8064 6236
rect 4338 6168 4344 6180
rect 3200 6140 4344 6168
rect 3200 6128 3206 6140
rect 4338 6128 4344 6140
rect 4396 6168 4402 6180
rect 7116 6168 7144 6208
rect 7558 6168 7564 6180
rect 4396 6140 7144 6168
rect 7208 6140 7564 6168
rect 4396 6128 4402 6140
rect 1394 6100 1400 6112
rect 1355 6072 1400 6100
rect 1394 6060 1400 6072
rect 1452 6060 1458 6112
rect 3694 6060 3700 6112
rect 3752 6100 3758 6112
rect 3973 6103 4031 6109
rect 3973 6100 3985 6103
rect 3752 6072 3985 6100
rect 3752 6060 3758 6072
rect 3973 6069 3985 6072
rect 4019 6069 4031 6103
rect 4614 6100 4620 6112
rect 4575 6072 4620 6100
rect 3973 6063 4031 6069
rect 4614 6060 4620 6072
rect 4672 6060 4678 6112
rect 5166 6100 5172 6112
rect 5127 6072 5172 6100
rect 5166 6060 5172 6072
rect 5224 6060 5230 6112
rect 6454 6060 6460 6112
rect 6512 6100 6518 6112
rect 6641 6103 6699 6109
rect 6641 6100 6653 6103
rect 6512 6072 6653 6100
rect 6512 6060 6518 6072
rect 6641 6069 6653 6072
rect 6687 6100 6699 6103
rect 7098 6100 7104 6112
rect 6687 6072 7104 6100
rect 6687 6069 6699 6072
rect 6641 6063 6699 6069
rect 7098 6060 7104 6072
rect 7156 6100 7162 6112
rect 7208 6100 7236 6140
rect 7558 6128 7564 6140
rect 7616 6128 7622 6180
rect 7466 6100 7472 6112
rect 7156 6072 7236 6100
rect 7427 6072 7472 6100
rect 7156 6060 7162 6072
rect 7466 6060 7472 6072
rect 7524 6060 7530 6112
rect 7834 6060 7840 6112
rect 7892 6100 7898 6112
rect 8662 6100 8668 6112
rect 7892 6072 8668 6100
rect 7892 6060 7898 6072
rect 8662 6060 8668 6072
rect 8720 6060 8726 6112
rect 8956 6100 8984 6276
rect 9030 6264 9036 6316
rect 9088 6304 9094 6316
rect 9324 6304 9505 6308
rect 9088 6280 9527 6304
rect 9088 6276 9352 6280
rect 9477 6276 9527 6280
rect 9088 6264 9094 6276
rect 9306 6168 9312 6180
rect 9267 6140 9312 6168
rect 9306 6128 9312 6140
rect 9364 6128 9370 6180
rect 9401 6171 9459 6177
rect 9401 6137 9413 6171
rect 9447 6168 9459 6171
rect 9499 6168 9527 6276
rect 10134 6264 10140 6316
rect 10192 6304 10198 6316
rect 10505 6307 10563 6313
rect 10505 6304 10517 6307
rect 10192 6276 10517 6304
rect 10192 6264 10198 6276
rect 10505 6273 10517 6276
rect 10551 6273 10563 6307
rect 11256 6304 11284 6344
rect 11422 6332 11428 6384
rect 11480 6372 11486 6384
rect 15102 6372 15108 6384
rect 11480 6344 15108 6372
rect 11480 6332 11486 6344
rect 15102 6332 15108 6344
rect 15160 6332 15166 6384
rect 11790 6304 11796 6316
rect 11256 6276 11796 6304
rect 10505 6267 10563 6273
rect 11790 6264 11796 6276
rect 11848 6264 11854 6316
rect 12158 6264 12164 6316
rect 12216 6304 12222 6316
rect 12216 6276 12261 6304
rect 12216 6264 12222 6276
rect 12710 6264 12716 6316
rect 12768 6304 12774 6316
rect 12989 6307 13047 6313
rect 12989 6304 13001 6307
rect 12768 6276 13001 6304
rect 12768 6264 12774 6276
rect 12989 6273 13001 6276
rect 13035 6273 13047 6307
rect 13722 6304 13728 6316
rect 12989 6267 13047 6273
rect 13096 6276 13728 6304
rect 9582 6196 9588 6248
rect 9640 6236 9646 6248
rect 9953 6239 10011 6245
rect 9953 6236 9965 6239
rect 9640 6208 9965 6236
rect 9640 6196 9646 6208
rect 9953 6205 9965 6208
rect 9999 6205 10011 6239
rect 9953 6199 10011 6205
rect 10413 6239 10471 6245
rect 10413 6205 10425 6239
rect 10459 6236 10471 6239
rect 10594 6236 10600 6248
rect 10459 6208 10600 6236
rect 10459 6205 10471 6208
rect 10413 6199 10471 6205
rect 10594 6196 10600 6208
rect 10652 6196 10658 6248
rect 11701 6239 11759 6245
rect 11701 6205 11713 6239
rect 11747 6236 11759 6239
rect 12437 6239 12495 6245
rect 12437 6236 12449 6239
rect 11747 6208 12449 6236
rect 11747 6205 11759 6208
rect 11701 6199 11759 6205
rect 12437 6205 12449 6208
rect 12483 6236 12495 6239
rect 12618 6236 12624 6248
rect 12483 6208 12624 6236
rect 12483 6205 12495 6208
rect 12437 6199 12495 6205
rect 12618 6196 12624 6208
rect 12676 6196 12682 6248
rect 12894 6196 12900 6248
rect 12952 6236 12958 6248
rect 13096 6245 13124 6276
rect 13722 6264 13728 6276
rect 13780 6264 13786 6316
rect 13906 6264 13912 6316
rect 13964 6304 13970 6316
rect 14277 6307 14335 6313
rect 14277 6304 14289 6307
rect 13964 6276 14289 6304
rect 13964 6264 13970 6276
rect 14277 6273 14289 6276
rect 14323 6273 14335 6307
rect 15562 6304 15568 6316
rect 14277 6267 14335 6273
rect 14660 6276 15148 6304
rect 15475 6276 15568 6304
rect 13081 6239 13139 6245
rect 13081 6236 13093 6239
rect 12952 6208 13093 6236
rect 12952 6196 12958 6208
rect 13081 6205 13093 6208
rect 13127 6205 13139 6239
rect 13081 6199 13139 6205
rect 13173 6239 13231 6245
rect 13173 6205 13185 6239
rect 13219 6236 13231 6239
rect 14001 6239 14059 6245
rect 14001 6236 14013 6239
rect 13219 6208 14013 6236
rect 13219 6205 13231 6208
rect 13173 6199 13231 6205
rect 14001 6205 14013 6208
rect 14047 6205 14059 6239
rect 14001 6199 14059 6205
rect 13188 6168 13216 6199
rect 14366 6196 14372 6248
rect 14424 6236 14430 6248
rect 14660 6245 14688 6276
rect 15120 6248 15148 6276
rect 15562 6264 15568 6276
rect 15620 6304 15626 6316
rect 16574 6304 16580 6316
rect 15620 6276 16580 6304
rect 15620 6264 15626 6276
rect 16574 6264 16580 6276
rect 16632 6264 16638 6316
rect 14645 6239 14703 6245
rect 14645 6236 14657 6239
rect 14424 6208 14657 6236
rect 14424 6196 14430 6208
rect 14645 6205 14657 6208
rect 14691 6205 14703 6239
rect 14645 6199 14703 6205
rect 14829 6239 14887 6245
rect 14829 6205 14841 6239
rect 14875 6205 14887 6239
rect 14829 6199 14887 6205
rect 9447 6140 9527 6168
rect 10060 6140 13216 6168
rect 9447 6137 9459 6140
rect 9401 6131 9459 6137
rect 10060 6100 10088 6140
rect 8956 6072 10088 6100
rect 10134 6060 10140 6112
rect 10192 6100 10198 6112
rect 10962 6100 10968 6112
rect 10192 6072 10968 6100
rect 10192 6060 10198 6072
rect 10962 6060 10968 6072
rect 11020 6060 11026 6112
rect 11238 6100 11244 6112
rect 11199 6072 11244 6100
rect 11238 6060 11244 6072
rect 11296 6060 11302 6112
rect 11330 6060 11336 6112
rect 11388 6100 11394 6112
rect 11793 6103 11851 6109
rect 11793 6100 11805 6103
rect 11388 6072 11805 6100
rect 11388 6060 11394 6072
rect 11793 6069 11805 6072
rect 11839 6069 11851 6103
rect 11793 6063 11851 6069
rect 11974 6060 11980 6112
rect 12032 6100 12038 6112
rect 12342 6100 12348 6112
rect 12032 6072 12348 6100
rect 12032 6060 12038 6072
rect 12342 6060 12348 6072
rect 12400 6060 12406 6112
rect 13814 6060 13820 6112
rect 13872 6100 13878 6112
rect 13998 6100 14004 6112
rect 13872 6072 14004 6100
rect 13872 6060 13878 6072
rect 13998 6060 14004 6072
rect 14056 6060 14062 6112
rect 14182 6060 14188 6112
rect 14240 6100 14246 6112
rect 14642 6100 14648 6112
rect 14240 6072 14648 6100
rect 14240 6060 14246 6072
rect 14642 6060 14648 6072
rect 14700 6100 14706 6112
rect 14844 6100 14872 6199
rect 15102 6196 15108 6248
rect 15160 6196 15166 6248
rect 15378 6100 15384 6112
rect 14700 6072 14872 6100
rect 15339 6072 15384 6100
rect 14700 6060 14706 6072
rect 15378 6060 15384 6072
rect 15436 6060 15442 6112
rect 1104 6010 16008 6032
rect 1104 5958 2824 6010
rect 2876 5958 2888 6010
rect 2940 5958 2952 6010
rect 3004 5958 3016 6010
rect 3068 5958 3080 6010
rect 3132 5958 6572 6010
rect 6624 5958 6636 6010
rect 6688 5958 6700 6010
rect 6752 5958 6764 6010
rect 6816 5958 6828 6010
rect 6880 5958 10320 6010
rect 10372 5958 10384 6010
rect 10436 5958 10448 6010
rect 10500 5958 10512 6010
rect 10564 5958 10576 6010
rect 10628 5958 14068 6010
rect 14120 5958 14132 6010
rect 14184 5958 14196 6010
rect 14248 5958 14260 6010
rect 14312 5958 14324 6010
rect 14376 5958 16008 6010
rect 1104 5936 16008 5958
rect 1762 5896 1768 5908
rect 1723 5868 1768 5896
rect 1762 5856 1768 5868
rect 1820 5856 1826 5908
rect 2038 5856 2044 5908
rect 2096 5896 2102 5908
rect 2317 5899 2375 5905
rect 2317 5896 2329 5899
rect 2096 5868 2329 5896
rect 2096 5856 2102 5868
rect 2317 5865 2329 5868
rect 2363 5865 2375 5899
rect 4617 5899 4675 5905
rect 4617 5896 4629 5899
rect 2317 5859 2375 5865
rect 2746 5868 4629 5896
rect 2746 5828 2774 5868
rect 4617 5865 4629 5868
rect 4663 5865 4675 5899
rect 4617 5859 4675 5865
rect 5258 5856 5264 5908
rect 5316 5896 5322 5908
rect 5810 5896 5816 5908
rect 5316 5868 5816 5896
rect 5316 5856 5322 5868
rect 5810 5856 5816 5868
rect 5868 5856 5874 5908
rect 6270 5856 6276 5908
rect 6328 5896 6334 5908
rect 6730 5896 6736 5908
rect 6328 5868 6736 5896
rect 6328 5856 6334 5868
rect 6730 5856 6736 5868
rect 6788 5896 6794 5908
rect 6788 5868 11008 5896
rect 6788 5856 6794 5868
rect 10980 5840 11008 5868
rect 12618 5856 12624 5908
rect 12676 5896 12682 5908
rect 13998 5896 14004 5908
rect 12676 5868 14004 5896
rect 12676 5856 12682 5868
rect 13998 5856 14004 5868
rect 14056 5856 14062 5908
rect 14277 5899 14335 5905
rect 14277 5865 14289 5899
rect 14323 5896 14335 5899
rect 15562 5896 15568 5908
rect 14323 5868 15568 5896
rect 14323 5865 14335 5868
rect 14277 5859 14335 5865
rect 15562 5856 15568 5868
rect 15620 5856 15626 5908
rect 3142 5828 3148 5840
rect 1688 5800 2774 5828
rect 2884 5800 3148 5828
rect 1688 5701 1716 5800
rect 2130 5720 2136 5772
rect 2188 5760 2194 5772
rect 2884 5769 2912 5800
rect 3142 5788 3148 5800
rect 3200 5788 3206 5840
rect 3418 5828 3424 5840
rect 3379 5800 3424 5828
rect 3418 5788 3424 5800
rect 3476 5788 3482 5840
rect 3789 5831 3847 5837
rect 3789 5797 3801 5831
rect 3835 5797 3847 5831
rect 5074 5828 5080 5840
rect 3789 5791 3847 5797
rect 4448 5800 5080 5828
rect 2869 5763 2927 5769
rect 2188 5732 2774 5760
rect 2188 5720 2194 5732
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5661 1731 5695
rect 1673 5655 1731 5661
rect 1949 5695 2007 5701
rect 1949 5661 1961 5695
rect 1995 5692 2007 5695
rect 2314 5692 2320 5704
rect 1995 5664 2320 5692
rect 1995 5661 2007 5664
rect 1949 5655 2007 5661
rect 2314 5652 2320 5664
rect 2372 5652 2378 5704
rect 2746 5692 2774 5732
rect 2869 5729 2881 5763
rect 2915 5729 2927 5763
rect 3804 5760 3832 5791
rect 4338 5760 4344 5772
rect 2869 5723 2927 5729
rect 2976 5732 3832 5760
rect 4080 5732 4344 5760
rect 2976 5692 3004 5732
rect 2746 5664 3004 5692
rect 3605 5695 3663 5701
rect 3605 5661 3617 5695
rect 3651 5692 3663 5695
rect 4080 5692 4108 5732
rect 4338 5720 4344 5732
rect 4396 5720 4402 5772
rect 4448 5769 4476 5800
rect 5074 5788 5080 5800
rect 5132 5788 5138 5840
rect 5534 5788 5540 5840
rect 5592 5828 5598 5840
rect 7834 5828 7840 5840
rect 5592 5800 7840 5828
rect 5592 5788 5598 5800
rect 7834 5788 7840 5800
rect 7892 5788 7898 5840
rect 7926 5788 7932 5840
rect 7984 5828 7990 5840
rect 9030 5828 9036 5840
rect 7984 5800 8029 5828
rect 8266 5800 9036 5828
rect 7984 5788 7990 5800
rect 4433 5763 4491 5769
rect 4433 5729 4445 5763
rect 4479 5729 4491 5763
rect 4433 5723 4491 5729
rect 5258 5720 5264 5772
rect 5316 5760 5322 5772
rect 5316 5732 5361 5760
rect 5316 5720 5322 5732
rect 5442 5720 5448 5772
rect 5500 5760 5506 5772
rect 5994 5760 6000 5772
rect 5500 5732 6000 5760
rect 5500 5720 5506 5732
rect 5994 5720 6000 5732
rect 6052 5760 6058 5772
rect 6454 5760 6460 5772
rect 6052 5732 6460 5760
rect 6052 5720 6058 5732
rect 6454 5720 6460 5732
rect 6512 5720 6518 5772
rect 6730 5760 6736 5772
rect 6691 5732 6736 5760
rect 6730 5720 6736 5732
rect 6788 5720 6794 5772
rect 7098 5760 7104 5772
rect 7059 5732 7104 5760
rect 7098 5720 7104 5732
rect 7156 5720 7162 5772
rect 7190 5720 7196 5772
rect 7248 5760 7254 5772
rect 7285 5763 7343 5769
rect 7285 5760 7297 5763
rect 7248 5732 7297 5760
rect 7248 5720 7254 5732
rect 7285 5729 7297 5732
rect 7331 5729 7343 5763
rect 8266 5760 8294 5800
rect 9030 5788 9036 5800
rect 9088 5788 9094 5840
rect 9217 5831 9275 5837
rect 9217 5797 9229 5831
rect 9263 5828 9275 5831
rect 9306 5828 9312 5840
rect 9263 5800 9312 5828
rect 9263 5797 9275 5800
rect 9217 5791 9275 5797
rect 9306 5788 9312 5800
rect 9364 5788 9370 5840
rect 9401 5831 9459 5837
rect 9401 5797 9413 5831
rect 9447 5828 9459 5831
rect 9490 5828 9496 5840
rect 9447 5800 9496 5828
rect 9447 5797 9459 5800
rect 9401 5791 9459 5797
rect 9490 5788 9496 5800
rect 9548 5788 9554 5840
rect 9766 5788 9772 5840
rect 9824 5828 9830 5840
rect 10410 5828 10416 5840
rect 9824 5800 10416 5828
rect 9824 5788 9830 5800
rect 10410 5788 10416 5800
rect 10468 5828 10474 5840
rect 10505 5831 10563 5837
rect 10505 5828 10517 5831
rect 10468 5800 10517 5828
rect 10468 5788 10474 5800
rect 10505 5797 10517 5800
rect 10551 5797 10563 5831
rect 10505 5791 10563 5797
rect 10962 5788 10968 5840
rect 11020 5828 11026 5840
rect 11020 5800 11376 5828
rect 11020 5788 11026 5800
rect 7285 5723 7343 5729
rect 8211 5732 8294 5760
rect 3651 5664 4108 5692
rect 4157 5695 4215 5701
rect 3651 5661 3663 5664
rect 3605 5655 3663 5661
rect 4157 5661 4169 5695
rect 4203 5692 4215 5695
rect 4706 5692 4712 5704
rect 4203 5664 4712 5692
rect 4203 5661 4215 5664
rect 4157 5655 4215 5661
rect 4706 5652 4712 5664
rect 4764 5652 4770 5704
rect 4801 5695 4859 5701
rect 4801 5661 4813 5695
rect 4847 5692 4859 5695
rect 5074 5692 5080 5704
rect 4847 5664 5080 5692
rect 4847 5661 4859 5664
rect 4801 5655 4859 5661
rect 5074 5652 5080 5664
rect 5132 5652 5138 5704
rect 5169 5695 5227 5701
rect 5169 5661 5181 5695
rect 5215 5692 5227 5695
rect 5460 5692 5488 5720
rect 5215 5664 5488 5692
rect 5537 5695 5595 5701
rect 5215 5661 5227 5664
rect 5169 5655 5227 5661
rect 5537 5661 5549 5695
rect 5583 5661 5595 5695
rect 5537 5655 5595 5661
rect 2222 5624 2228 5636
rect 2183 5596 2228 5624
rect 2222 5584 2228 5596
rect 2280 5584 2286 5636
rect 2590 5584 2596 5636
rect 2648 5624 2654 5636
rect 2685 5627 2743 5633
rect 2685 5624 2697 5627
rect 2648 5596 2697 5624
rect 2648 5584 2654 5596
rect 2685 5593 2697 5596
rect 2731 5593 2743 5627
rect 2685 5587 2743 5593
rect 2777 5627 2835 5633
rect 2777 5593 2789 5627
rect 2823 5624 2835 5627
rect 5552 5624 5580 5655
rect 6270 5652 6276 5704
rect 6328 5692 6334 5704
rect 6549 5695 6607 5701
rect 6549 5692 6561 5695
rect 6328 5664 6561 5692
rect 6328 5652 6334 5664
rect 6549 5661 6561 5664
rect 6595 5661 6607 5695
rect 7300 5692 7328 5723
rect 8211 5708 8239 5732
rect 8386 5720 8392 5772
rect 8444 5760 8450 5772
rect 8573 5763 8631 5769
rect 8573 5760 8585 5763
rect 8444 5732 8585 5760
rect 8444 5720 8450 5732
rect 8573 5729 8585 5732
rect 8619 5760 8631 5763
rect 9122 5760 9128 5772
rect 8619 5732 9128 5760
rect 8619 5729 8631 5732
rect 8573 5723 8631 5729
rect 9122 5720 9128 5732
rect 9180 5760 9186 5772
rect 9582 5760 9588 5772
rect 9180 5732 9588 5760
rect 9180 5720 9186 5732
rect 9582 5720 9588 5732
rect 9640 5720 9646 5772
rect 9677 5763 9735 5769
rect 9677 5729 9689 5763
rect 9723 5760 9735 5763
rect 10134 5760 10140 5772
rect 9723 5732 10140 5760
rect 9723 5729 9735 5732
rect 9677 5723 9735 5729
rect 10134 5720 10140 5732
rect 10192 5720 10198 5772
rect 11348 5769 11376 5800
rect 11790 5788 11796 5840
rect 11848 5828 11854 5840
rect 14734 5828 14740 5840
rect 11848 5800 14740 5828
rect 11848 5788 11854 5800
rect 14734 5788 14740 5800
rect 14792 5788 14798 5840
rect 11333 5763 11391 5769
rect 11333 5729 11345 5763
rect 11379 5729 11391 5763
rect 12345 5763 12403 5769
rect 12345 5760 12357 5763
rect 11333 5723 11391 5729
rect 11440 5732 12357 5760
rect 7561 5695 7619 5701
rect 7300 5664 7521 5692
rect 6549 5655 6607 5661
rect 2823 5596 3556 5624
rect 2823 5593 2835 5596
rect 2777 5587 2835 5593
rect 1486 5556 1492 5568
rect 1447 5528 1492 5556
rect 1486 5516 1492 5528
rect 1544 5516 1550 5568
rect 2700 5556 2728 5587
rect 3528 5568 3556 5596
rect 4172 5596 5580 5624
rect 6641 5627 6699 5633
rect 4172 5568 4200 5596
rect 6641 5593 6653 5627
rect 6687 5624 6699 5627
rect 7374 5624 7380 5636
rect 6687 5596 7380 5624
rect 6687 5593 6699 5596
rect 6641 5587 6699 5593
rect 7374 5584 7380 5596
rect 7432 5584 7438 5636
rect 7493 5624 7521 5664
rect 7561 5661 7573 5695
rect 7607 5692 7619 5695
rect 8128 5692 8239 5708
rect 7607 5680 8239 5692
rect 7607 5664 8156 5680
rect 7607 5661 7619 5664
rect 7561 5655 7619 5661
rect 8294 5652 8300 5704
rect 8352 5692 8358 5704
rect 8846 5692 8852 5704
rect 8352 5664 8852 5692
rect 8352 5652 8358 5664
rect 8846 5652 8852 5664
rect 8904 5652 8910 5704
rect 9030 5692 9036 5704
rect 8991 5664 9036 5692
rect 9030 5652 9036 5664
rect 9088 5652 9094 5704
rect 9499 5668 9904 5692
rect 9232 5664 9904 5668
rect 9232 5640 9527 5664
rect 7834 5624 7840 5636
rect 7493 5596 7840 5624
rect 7834 5584 7840 5596
rect 7892 5584 7898 5636
rect 8389 5627 8447 5633
rect 8389 5593 8401 5627
rect 8435 5624 8447 5627
rect 8570 5624 8576 5636
rect 8435 5596 8576 5624
rect 8435 5593 8447 5596
rect 8389 5587 8447 5593
rect 8570 5584 8576 5596
rect 8628 5584 8634 5636
rect 8662 5584 8668 5636
rect 8720 5624 8726 5636
rect 9232 5624 9260 5640
rect 8720 5596 9260 5624
rect 8720 5584 8726 5596
rect 9582 5584 9588 5636
rect 9640 5624 9646 5636
rect 9876 5633 9904 5664
rect 10042 5652 10048 5704
rect 10100 5692 10106 5704
rect 10321 5695 10379 5701
rect 10321 5692 10333 5695
rect 10100 5664 10333 5692
rect 10100 5652 10106 5664
rect 10321 5661 10333 5664
rect 10367 5692 10379 5695
rect 10962 5692 10968 5704
rect 10367 5664 10968 5692
rect 10367 5661 10379 5664
rect 10321 5655 10379 5661
rect 10962 5652 10968 5664
rect 11020 5652 11026 5704
rect 11146 5692 11152 5704
rect 11107 5664 11152 5692
rect 11146 5652 11152 5664
rect 11204 5652 11210 5704
rect 11238 5652 11244 5704
rect 11296 5692 11302 5704
rect 11440 5692 11468 5732
rect 12345 5729 12357 5732
rect 12391 5729 12403 5763
rect 12345 5723 12403 5729
rect 12434 5720 12440 5772
rect 12492 5760 12498 5772
rect 13354 5760 13360 5772
rect 12492 5732 12537 5760
rect 13315 5732 13360 5760
rect 12492 5720 12498 5732
rect 13354 5720 13360 5732
rect 13412 5720 13418 5772
rect 14274 5720 14280 5772
rect 14332 5760 14338 5772
rect 15105 5763 15163 5769
rect 15105 5760 15117 5763
rect 14332 5732 15117 5760
rect 14332 5720 14338 5732
rect 15105 5729 15117 5732
rect 15151 5729 15163 5763
rect 15105 5723 15163 5729
rect 11296 5664 11468 5692
rect 11609 5695 11667 5701
rect 11296 5652 11302 5664
rect 11609 5661 11621 5695
rect 11655 5692 11667 5695
rect 11974 5692 11980 5704
rect 11655 5664 11980 5692
rect 11655 5661 11667 5664
rect 11609 5655 11667 5661
rect 11974 5652 11980 5664
rect 12032 5652 12038 5704
rect 12253 5695 12311 5701
rect 12253 5661 12265 5695
rect 12299 5692 12311 5695
rect 14090 5692 14096 5704
rect 12299 5664 13952 5692
rect 14051 5664 14096 5692
rect 12299 5661 12311 5664
rect 12253 5655 12311 5661
rect 13924 5633 13952 5664
rect 14090 5652 14096 5664
rect 14148 5652 14154 5704
rect 14553 5695 14611 5701
rect 14553 5661 14565 5695
rect 14599 5692 14611 5695
rect 14642 5692 14648 5704
rect 14599 5664 14648 5692
rect 14599 5661 14611 5664
rect 14553 5655 14611 5661
rect 14642 5652 14648 5664
rect 14700 5652 14706 5704
rect 14826 5692 14832 5704
rect 14787 5664 14832 5692
rect 14826 5652 14832 5664
rect 14884 5652 14890 5704
rect 9861 5627 9919 5633
rect 9640 5584 9674 5624
rect 9861 5593 9873 5627
rect 9907 5624 9919 5627
rect 11057 5627 11115 5633
rect 9907 5596 11008 5624
rect 9907 5593 9919 5596
rect 9861 5587 9919 5593
rect 3145 5559 3203 5565
rect 3145 5556 3157 5559
rect 2700 5528 3157 5556
rect 3145 5525 3157 5528
rect 3191 5525 3203 5559
rect 3145 5519 3203 5525
rect 3510 5516 3516 5568
rect 3568 5516 3574 5568
rect 4154 5516 4160 5568
rect 4212 5516 4218 5568
rect 4246 5516 4252 5568
rect 4304 5556 4310 5568
rect 4985 5559 5043 5565
rect 4304 5528 4349 5556
rect 4304 5516 4310 5528
rect 4985 5525 4997 5559
rect 5031 5556 5043 5559
rect 5258 5556 5264 5568
rect 5031 5528 5264 5556
rect 5031 5525 5043 5528
rect 4985 5519 5043 5525
rect 5258 5516 5264 5528
rect 5316 5516 5322 5568
rect 5442 5516 5448 5568
rect 5500 5556 5506 5568
rect 6181 5559 6239 5565
rect 6181 5556 6193 5559
rect 5500 5528 6193 5556
rect 5500 5516 5506 5528
rect 6181 5525 6193 5528
rect 6227 5525 6239 5559
rect 6181 5519 6239 5525
rect 7469 5559 7527 5565
rect 7469 5525 7481 5559
rect 7515 5556 7527 5559
rect 8021 5559 8079 5565
rect 8021 5556 8033 5559
rect 7515 5528 8033 5556
rect 7515 5525 7527 5528
rect 7469 5519 7527 5525
rect 8021 5525 8033 5528
rect 8067 5525 8079 5559
rect 8021 5519 8079 5525
rect 8202 5516 8208 5568
rect 8260 5556 8266 5568
rect 8481 5559 8539 5565
rect 8481 5556 8493 5559
rect 8260 5528 8493 5556
rect 8260 5516 8266 5528
rect 8481 5525 8493 5528
rect 8527 5556 8539 5559
rect 9030 5556 9036 5568
rect 8527 5528 9036 5556
rect 8527 5525 8539 5528
rect 8481 5519 8539 5525
rect 9030 5516 9036 5528
rect 9088 5516 9094 5568
rect 9646 5556 9674 5584
rect 9766 5556 9772 5568
rect 9646 5528 9772 5556
rect 9766 5516 9772 5528
rect 9824 5516 9830 5568
rect 10226 5556 10232 5568
rect 10187 5528 10232 5556
rect 10226 5516 10232 5528
rect 10284 5516 10290 5568
rect 10686 5556 10692 5568
rect 10647 5528 10692 5556
rect 10686 5516 10692 5528
rect 10744 5516 10750 5568
rect 10980 5556 11008 5596
rect 11057 5593 11069 5627
rect 11103 5624 11115 5627
rect 13081 5627 13139 5633
rect 11103 5596 12756 5624
rect 11103 5593 11115 5596
rect 11057 5587 11115 5593
rect 11422 5556 11428 5568
rect 10980 5528 11428 5556
rect 11422 5516 11428 5528
rect 11480 5516 11486 5568
rect 11790 5556 11796 5568
rect 11751 5528 11796 5556
rect 11790 5516 11796 5528
rect 11848 5516 11854 5568
rect 11885 5559 11943 5565
rect 11885 5525 11897 5559
rect 11931 5556 11943 5559
rect 12342 5556 12348 5568
rect 11931 5528 12348 5556
rect 11931 5525 11943 5528
rect 11885 5519 11943 5525
rect 12342 5516 12348 5528
rect 12400 5516 12406 5568
rect 12728 5565 12756 5596
rect 13081 5593 13093 5627
rect 13127 5624 13139 5627
rect 13541 5627 13599 5633
rect 13541 5624 13553 5627
rect 13127 5596 13553 5624
rect 13127 5593 13139 5596
rect 13081 5587 13139 5593
rect 13541 5593 13553 5596
rect 13587 5593 13599 5627
rect 13541 5587 13599 5593
rect 13909 5627 13967 5633
rect 13909 5593 13921 5627
rect 13955 5624 13967 5627
rect 14182 5624 14188 5636
rect 13955 5596 14188 5624
rect 13955 5593 13967 5596
rect 13909 5587 13967 5593
rect 14182 5584 14188 5596
rect 14240 5584 14246 5636
rect 12713 5559 12771 5565
rect 12713 5525 12725 5559
rect 12759 5525 12771 5559
rect 12713 5519 12771 5525
rect 13173 5559 13231 5565
rect 13173 5525 13185 5559
rect 13219 5556 13231 5559
rect 13722 5556 13728 5568
rect 13219 5528 13728 5556
rect 13219 5525 13231 5528
rect 13173 5519 13231 5525
rect 13722 5516 13728 5528
rect 13780 5516 13786 5568
rect 14366 5556 14372 5568
rect 14327 5528 14372 5556
rect 14366 5516 14372 5528
rect 14424 5516 14430 5568
rect 14737 5559 14795 5565
rect 14737 5525 14749 5559
rect 14783 5556 14795 5559
rect 15010 5556 15016 5568
rect 14783 5528 15016 5556
rect 14783 5525 14795 5528
rect 14737 5519 14795 5525
rect 15010 5516 15016 5528
rect 15068 5516 15074 5568
rect 1104 5466 16008 5488
rect 1104 5414 4698 5466
rect 4750 5414 4762 5466
rect 4814 5414 4826 5466
rect 4878 5414 4890 5466
rect 4942 5414 4954 5466
rect 5006 5414 8446 5466
rect 8498 5414 8510 5466
rect 8562 5414 8574 5466
rect 8626 5414 8638 5466
rect 8690 5414 8702 5466
rect 8754 5414 12194 5466
rect 12246 5414 12258 5466
rect 12310 5414 12322 5466
rect 12374 5414 12386 5466
rect 12438 5414 12450 5466
rect 12502 5414 16008 5466
rect 1104 5392 16008 5414
rect 2593 5355 2651 5361
rect 2593 5321 2605 5355
rect 2639 5352 2651 5355
rect 3053 5355 3111 5361
rect 3053 5352 3065 5355
rect 2639 5324 3065 5352
rect 2639 5321 2651 5324
rect 2593 5315 2651 5321
rect 3053 5321 3065 5324
rect 3099 5321 3111 5355
rect 3053 5315 3111 5321
rect 3510 5312 3516 5364
rect 3568 5352 3574 5364
rect 3605 5355 3663 5361
rect 3605 5352 3617 5355
rect 3568 5324 3617 5352
rect 3568 5312 3574 5324
rect 3605 5321 3617 5324
rect 3651 5321 3663 5355
rect 3605 5315 3663 5321
rect 3970 5312 3976 5364
rect 4028 5352 4034 5364
rect 4028 5324 4292 5352
rect 4028 5312 4034 5324
rect 2133 5287 2191 5293
rect 2133 5253 2145 5287
rect 2179 5284 2191 5287
rect 2179 5256 2636 5284
rect 2179 5253 2191 5256
rect 2133 5247 2191 5253
rect 1670 5216 1676 5228
rect 1631 5188 1676 5216
rect 1670 5176 1676 5188
rect 1728 5176 1734 5228
rect 2225 5219 2283 5225
rect 2225 5185 2237 5219
rect 2271 5216 2283 5219
rect 2498 5216 2504 5228
rect 2271 5188 2504 5216
rect 2271 5185 2283 5188
rect 2225 5179 2283 5185
rect 2498 5176 2504 5188
rect 2556 5176 2562 5228
rect 2608 5216 2636 5256
rect 2682 5244 2688 5296
rect 2740 5284 2746 5296
rect 3145 5287 3203 5293
rect 3145 5284 3157 5287
rect 2740 5256 3157 5284
rect 2740 5244 2746 5256
rect 3145 5253 3157 5256
rect 3191 5253 3203 5287
rect 4154 5284 4160 5296
rect 3145 5247 3203 5253
rect 3344 5256 4160 5284
rect 3344 5216 3372 5256
rect 4154 5244 4160 5256
rect 4212 5244 4218 5296
rect 3786 5216 3792 5228
rect 2608 5188 3372 5216
rect 3436 5188 3792 5216
rect 3436 5160 3464 5188
rect 3786 5176 3792 5188
rect 3844 5176 3850 5228
rect 3970 5216 3976 5228
rect 3931 5188 3976 5216
rect 3970 5176 3976 5188
rect 4028 5176 4034 5228
rect 1946 5148 1952 5160
rect 1907 5120 1952 5148
rect 1946 5108 1952 5120
rect 2004 5108 2010 5160
rect 3329 5151 3387 5157
rect 3329 5117 3341 5151
rect 3375 5148 3387 5151
rect 3418 5148 3424 5160
rect 3375 5120 3424 5148
rect 3375 5117 3387 5120
rect 3329 5111 3387 5117
rect 3418 5108 3424 5120
rect 3476 5108 3482 5160
rect 3602 5108 3608 5160
rect 3660 5148 3666 5160
rect 4264 5157 4292 5324
rect 4982 5312 4988 5364
rect 5040 5352 5046 5364
rect 5350 5352 5356 5364
rect 5040 5324 5356 5352
rect 5040 5312 5046 5324
rect 5350 5312 5356 5324
rect 5408 5312 5414 5364
rect 5442 5312 5448 5364
rect 5500 5352 5506 5364
rect 5537 5355 5595 5361
rect 5537 5352 5549 5355
rect 5500 5324 5549 5352
rect 5500 5312 5506 5324
rect 5537 5321 5549 5324
rect 5583 5321 5595 5355
rect 7285 5355 7343 5361
rect 7285 5352 7297 5355
rect 5537 5315 5595 5321
rect 5644 5324 7297 5352
rect 5258 5244 5264 5296
rect 5316 5284 5322 5296
rect 5644 5284 5672 5324
rect 7285 5321 7297 5324
rect 7331 5352 7343 5355
rect 7650 5352 7656 5364
rect 7331 5324 7656 5352
rect 7331 5321 7343 5324
rect 7285 5315 7343 5321
rect 7650 5312 7656 5324
rect 7708 5312 7714 5364
rect 7742 5312 7748 5364
rect 7800 5352 7806 5364
rect 8573 5355 8631 5361
rect 8573 5352 8585 5355
rect 7800 5324 8585 5352
rect 7800 5312 7806 5324
rect 8573 5321 8585 5324
rect 8619 5321 8631 5355
rect 8573 5315 8631 5321
rect 8941 5355 8999 5361
rect 8941 5321 8953 5355
rect 8987 5352 8999 5355
rect 9766 5352 9772 5364
rect 8987 5324 9772 5352
rect 8987 5321 8999 5324
rect 8941 5315 8999 5321
rect 9766 5312 9772 5324
rect 9824 5312 9830 5364
rect 10045 5355 10103 5361
rect 10045 5321 10057 5355
rect 10091 5352 10103 5355
rect 10226 5352 10232 5364
rect 10091 5324 10232 5352
rect 10091 5321 10103 5324
rect 10045 5315 10103 5321
rect 10226 5312 10232 5324
rect 10284 5312 10290 5364
rect 10505 5355 10563 5361
rect 10505 5321 10517 5355
rect 10551 5352 10563 5355
rect 10873 5355 10931 5361
rect 10873 5352 10885 5355
rect 10551 5324 10885 5352
rect 10551 5321 10563 5324
rect 10505 5315 10563 5321
rect 10873 5321 10885 5324
rect 10919 5321 10931 5355
rect 10873 5315 10931 5321
rect 10962 5312 10968 5364
rect 11020 5352 11026 5364
rect 11793 5355 11851 5361
rect 11020 5324 11065 5352
rect 11020 5312 11026 5324
rect 11793 5321 11805 5355
rect 11839 5352 11851 5355
rect 11882 5352 11888 5364
rect 11839 5324 11888 5352
rect 11839 5321 11851 5324
rect 11793 5315 11851 5321
rect 11882 5312 11888 5324
rect 11940 5312 11946 5364
rect 12250 5352 12256 5364
rect 12211 5324 12256 5352
rect 12250 5312 12256 5324
rect 12308 5312 12314 5364
rect 12342 5312 12348 5364
rect 12400 5352 12406 5364
rect 13357 5355 13415 5361
rect 13357 5352 13369 5355
rect 12400 5324 13369 5352
rect 12400 5312 12406 5324
rect 13357 5321 13369 5324
rect 13403 5352 13415 5355
rect 13814 5352 13820 5364
rect 13403 5324 13820 5352
rect 13403 5321 13415 5324
rect 13357 5315 13415 5321
rect 13814 5312 13820 5324
rect 13872 5312 13878 5364
rect 14090 5352 14096 5364
rect 14051 5324 14096 5352
rect 14090 5312 14096 5324
rect 14148 5312 14154 5364
rect 14458 5312 14464 5364
rect 14516 5352 14522 5364
rect 14645 5355 14703 5361
rect 14645 5352 14657 5355
rect 14516 5324 14657 5352
rect 14516 5312 14522 5324
rect 14645 5321 14657 5324
rect 14691 5321 14703 5355
rect 14645 5315 14703 5321
rect 14734 5312 14740 5364
rect 14792 5352 14798 5364
rect 15105 5355 15163 5361
rect 15105 5352 15117 5355
rect 14792 5324 15117 5352
rect 14792 5312 14798 5324
rect 15105 5321 15117 5324
rect 15151 5321 15163 5355
rect 15470 5352 15476 5364
rect 15431 5324 15476 5352
rect 15105 5315 15163 5321
rect 15470 5312 15476 5324
rect 15528 5312 15534 5364
rect 5902 5284 5908 5296
rect 5316 5256 5672 5284
rect 5863 5256 5908 5284
rect 5316 5244 5322 5256
rect 5902 5244 5908 5256
rect 5960 5244 5966 5296
rect 6178 5244 6184 5296
rect 6236 5284 6242 5296
rect 6454 5284 6460 5296
rect 6236 5256 6460 5284
rect 6236 5244 6242 5256
rect 6454 5244 6460 5256
rect 6512 5244 6518 5296
rect 6641 5287 6699 5293
rect 6641 5253 6653 5287
rect 6687 5284 6699 5287
rect 6730 5284 6736 5296
rect 6687 5256 6736 5284
rect 6687 5253 6699 5256
rect 6641 5247 6699 5253
rect 6730 5244 6736 5256
rect 6788 5244 6794 5296
rect 6825 5287 6883 5293
rect 6825 5253 6837 5287
rect 6871 5284 6883 5287
rect 6914 5284 6920 5296
rect 6871 5256 6920 5284
rect 6871 5253 6883 5256
rect 6825 5247 6883 5253
rect 6914 5244 6920 5256
rect 6972 5284 6978 5296
rect 8113 5287 8171 5293
rect 6972 5256 8064 5284
rect 6972 5244 6978 5256
rect 5445 5219 5503 5225
rect 5445 5185 5457 5219
rect 5491 5216 5503 5219
rect 5534 5216 5540 5228
rect 5491 5188 5540 5216
rect 5491 5185 5503 5188
rect 5445 5179 5503 5185
rect 5534 5176 5540 5188
rect 5592 5176 5598 5228
rect 5810 5176 5816 5228
rect 5868 5216 5874 5228
rect 7190 5216 7196 5228
rect 5868 5188 7196 5216
rect 5868 5176 5874 5188
rect 7190 5176 7196 5188
rect 7248 5176 7254 5228
rect 7282 5176 7288 5228
rect 7340 5216 7346 5228
rect 8036 5216 8064 5256
rect 8113 5253 8125 5287
rect 8159 5284 8171 5287
rect 9401 5287 9459 5293
rect 9401 5284 9413 5287
rect 8159 5256 9413 5284
rect 8159 5253 8171 5256
rect 8113 5247 8171 5253
rect 9401 5253 9413 5256
rect 9447 5253 9459 5287
rect 11330 5284 11336 5296
rect 9401 5247 9459 5253
rect 10060 5256 11336 5284
rect 10060 5228 10088 5256
rect 11330 5244 11336 5256
rect 11388 5244 11394 5296
rect 12434 5284 12440 5296
rect 11900 5256 12440 5284
rect 9030 5216 9036 5228
rect 7340 5188 7604 5216
rect 8036 5188 8800 5216
rect 8991 5188 9036 5216
rect 7340 5176 7346 5188
rect 4065 5151 4123 5157
rect 4065 5148 4077 5151
rect 3660 5120 4077 5148
rect 3660 5108 3666 5120
rect 4065 5117 4077 5120
rect 4111 5117 4123 5151
rect 4065 5111 4123 5117
rect 4249 5151 4307 5157
rect 4249 5117 4261 5151
rect 4295 5117 4307 5151
rect 4249 5111 4307 5117
rect 4525 5151 4583 5157
rect 4525 5117 4537 5151
rect 4571 5148 4583 5151
rect 5629 5151 5687 5157
rect 5629 5148 5641 5151
rect 4571 5120 5396 5148
rect 4571 5117 4583 5120
rect 4525 5111 4583 5117
rect 2314 5040 2320 5092
rect 2372 5080 2378 5092
rect 5077 5083 5135 5089
rect 5077 5080 5089 5083
rect 2372 5052 5089 5080
rect 2372 5040 2378 5052
rect 5077 5049 5089 5052
rect 5123 5049 5135 5083
rect 5077 5043 5135 5049
rect 1486 5012 1492 5024
rect 1447 4984 1492 5012
rect 1486 4972 1492 4984
rect 1544 4972 1550 5024
rect 1854 4972 1860 5024
rect 1912 5012 1918 5024
rect 2685 5015 2743 5021
rect 2685 5012 2697 5015
rect 1912 4984 2697 5012
rect 1912 4972 1918 4984
rect 2685 4981 2697 4984
rect 2731 4981 2743 5015
rect 2685 4975 2743 4981
rect 3142 4972 3148 5024
rect 3200 5012 3206 5024
rect 3694 5012 3700 5024
rect 3200 4984 3700 5012
rect 3200 4972 3206 4984
rect 3694 4972 3700 4984
rect 3752 4972 3758 5024
rect 4062 4972 4068 5024
rect 4120 5012 4126 5024
rect 4709 5015 4767 5021
rect 4709 5012 4721 5015
rect 4120 4984 4721 5012
rect 4120 4972 4126 4984
rect 4709 4981 4721 4984
rect 4755 4981 4767 5015
rect 4890 5012 4896 5024
rect 4851 4984 4896 5012
rect 4709 4975 4767 4981
rect 4890 4972 4896 4984
rect 4948 4972 4954 5024
rect 5368 5012 5396 5120
rect 5460 5120 5641 5148
rect 5460 5092 5488 5120
rect 5629 5117 5641 5120
rect 5675 5117 5687 5151
rect 5629 5111 5687 5117
rect 7098 5108 7104 5160
rect 7156 5148 7162 5160
rect 7576 5157 7604 5188
rect 7377 5151 7435 5157
rect 7377 5148 7389 5151
rect 7156 5120 7389 5148
rect 7156 5108 7162 5120
rect 7377 5117 7389 5120
rect 7423 5117 7435 5151
rect 7377 5111 7435 5117
rect 7561 5151 7619 5157
rect 7561 5117 7573 5151
rect 7607 5117 7619 5151
rect 7834 5148 7840 5160
rect 7795 5120 7840 5148
rect 7561 5111 7619 5117
rect 7834 5108 7840 5120
rect 7892 5108 7898 5160
rect 8021 5151 8079 5157
rect 8021 5117 8033 5151
rect 8067 5148 8079 5151
rect 8478 5148 8484 5160
rect 8067 5120 8484 5148
rect 8067 5117 8079 5120
rect 8021 5111 8079 5117
rect 5442 5040 5448 5092
rect 5500 5040 5506 5092
rect 6181 5083 6239 5089
rect 6181 5049 6193 5083
rect 6227 5080 6239 5083
rect 6227 5052 7420 5080
rect 6227 5049 6239 5052
rect 6181 5043 6239 5049
rect 7392 5024 7420 5052
rect 5994 5012 6000 5024
rect 5368 4984 6000 5012
rect 5994 4972 6000 4984
rect 6052 4972 6058 5024
rect 6362 5012 6368 5024
rect 6323 4984 6368 5012
rect 6362 4972 6368 4984
rect 6420 4972 6426 5024
rect 6917 5015 6975 5021
rect 6917 4981 6929 5015
rect 6963 5012 6975 5015
rect 7098 5012 7104 5024
rect 6963 4984 7104 5012
rect 6963 4981 6975 4984
rect 6917 4975 6975 4981
rect 7098 4972 7104 4984
rect 7156 4972 7162 5024
rect 7374 4972 7380 5024
rect 7432 5012 7438 5024
rect 8036 5012 8064 5111
rect 8478 5108 8484 5120
rect 8536 5108 8542 5160
rect 8772 5148 8800 5188
rect 9030 5176 9036 5188
rect 9088 5176 9094 5228
rect 10042 5176 10048 5228
rect 10100 5176 10106 5228
rect 10137 5219 10195 5225
rect 10137 5185 10149 5219
rect 10183 5216 10195 5219
rect 10226 5216 10232 5228
rect 10183 5188 10232 5216
rect 10183 5185 10195 5188
rect 10137 5179 10195 5185
rect 10226 5176 10232 5188
rect 10284 5176 10290 5228
rect 10594 5176 10600 5228
rect 10652 5216 10658 5228
rect 11900 5225 11928 5256
rect 12434 5244 12440 5256
rect 12492 5244 12498 5296
rect 13538 5284 13544 5296
rect 12544 5256 13308 5284
rect 13499 5256 13544 5284
rect 10980 5216 11100 5220
rect 11885 5219 11943 5225
rect 10652 5192 11744 5216
rect 10652 5188 11008 5192
rect 11072 5188 11744 5192
rect 10652 5176 10658 5188
rect 9122 5148 9128 5160
rect 8772 5120 8892 5148
rect 9083 5120 9128 5148
rect 8202 5040 8208 5092
rect 8260 5080 8266 5092
rect 8386 5080 8392 5092
rect 8260 5052 8392 5080
rect 8260 5040 8266 5052
rect 8386 5040 8392 5052
rect 8444 5040 8450 5092
rect 7432 4984 8064 5012
rect 8481 5015 8539 5021
rect 7432 4972 7438 4984
rect 8481 4981 8493 5015
rect 8527 5012 8539 5015
rect 8754 5012 8760 5024
rect 8527 4984 8760 5012
rect 8527 4981 8539 4984
rect 8481 4975 8539 4981
rect 8754 4972 8760 4984
rect 8812 4972 8818 5024
rect 8864 5012 8892 5120
rect 9122 5108 9128 5120
rect 9180 5108 9186 5160
rect 9858 5148 9864 5160
rect 9819 5120 9864 5148
rect 9858 5108 9864 5120
rect 9916 5108 9922 5160
rect 9950 5108 9956 5160
rect 10008 5148 10014 5160
rect 10502 5148 10508 5160
rect 10008 5120 10508 5148
rect 10008 5108 10014 5120
rect 10502 5108 10508 5120
rect 10560 5108 10566 5160
rect 10686 5148 10692 5160
rect 10647 5120 10692 5148
rect 10686 5108 10692 5120
rect 10744 5108 10750 5160
rect 11422 5108 11428 5160
rect 11480 5148 11486 5160
rect 11609 5151 11667 5157
rect 11609 5148 11621 5151
rect 11480 5120 11621 5148
rect 11480 5108 11486 5120
rect 11609 5117 11621 5120
rect 11655 5117 11667 5151
rect 11716 5148 11744 5188
rect 11885 5185 11897 5219
rect 11931 5185 11943 5219
rect 11885 5179 11943 5185
rect 12544 5148 12572 5256
rect 12710 5216 12716 5228
rect 12671 5188 12716 5216
rect 12710 5176 12716 5188
rect 12768 5176 12774 5228
rect 12894 5176 12900 5228
rect 12952 5176 12958 5228
rect 13078 5176 13084 5228
rect 13136 5216 13142 5228
rect 13173 5219 13231 5225
rect 13173 5216 13185 5219
rect 13136 5188 13185 5216
rect 13136 5176 13142 5188
rect 13173 5185 13185 5188
rect 13219 5185 13231 5219
rect 13280 5216 13308 5256
rect 13538 5244 13544 5256
rect 13596 5244 13602 5296
rect 14274 5284 14280 5296
rect 13648 5256 14280 5284
rect 13648 5216 13676 5256
rect 14274 5244 14280 5256
rect 14332 5244 14338 5296
rect 15013 5287 15071 5293
rect 15013 5253 15025 5287
rect 15059 5284 15071 5287
rect 15838 5284 15844 5296
rect 15059 5256 15844 5284
rect 15059 5253 15071 5256
rect 15013 5247 15071 5253
rect 13280 5188 13676 5216
rect 14001 5219 14059 5225
rect 13173 5179 13231 5185
rect 14001 5185 14013 5219
rect 14047 5216 14059 5219
rect 15286 5216 15292 5228
rect 14047 5188 14780 5216
rect 14047 5185 14059 5188
rect 14001 5179 14059 5185
rect 12802 5148 12808 5160
rect 11716 5120 12572 5148
rect 12763 5120 12808 5148
rect 11609 5111 11667 5117
rect 12802 5108 12808 5120
rect 12860 5108 12866 5160
rect 12912 5148 12940 5176
rect 12989 5151 13047 5157
rect 12989 5148 13001 5151
rect 12912 5120 13001 5148
rect 12989 5117 13001 5120
rect 13035 5117 13047 5151
rect 13188 5148 13216 5179
rect 13538 5148 13544 5160
rect 13188 5120 13544 5148
rect 12989 5111 13047 5117
rect 13538 5108 13544 5120
rect 13596 5108 13602 5160
rect 14090 5108 14096 5160
rect 14148 5148 14154 5160
rect 14277 5151 14335 5157
rect 14277 5148 14289 5151
rect 14148 5120 14289 5148
rect 14148 5108 14154 5120
rect 14277 5117 14289 5120
rect 14323 5148 14335 5151
rect 14642 5148 14648 5160
rect 14323 5120 14648 5148
rect 14323 5117 14335 5120
rect 14277 5111 14335 5117
rect 14642 5108 14648 5120
rect 14700 5108 14706 5160
rect 14752 5148 14780 5188
rect 15120 5188 15292 5216
rect 15120 5148 15148 5188
rect 15286 5176 15292 5188
rect 15344 5176 15350 5228
rect 14752 5120 15148 5148
rect 15197 5151 15255 5157
rect 15197 5117 15209 5151
rect 15243 5117 15255 5151
rect 15197 5111 15255 5117
rect 9490 5040 9496 5092
rect 9548 5080 9554 5092
rect 13633 5083 13691 5089
rect 13633 5080 13645 5083
rect 9548 5052 13645 5080
rect 9548 5040 9554 5052
rect 13633 5049 13645 5052
rect 13679 5049 13691 5083
rect 13633 5043 13691 5049
rect 13740 5052 14596 5080
rect 10318 5012 10324 5024
rect 8864 4984 10324 5012
rect 10318 4972 10324 4984
rect 10376 4972 10382 5024
rect 11330 5012 11336 5024
rect 11291 4984 11336 5012
rect 11330 4972 11336 4984
rect 11388 4972 11394 5024
rect 12342 5012 12348 5024
rect 12303 4984 12348 5012
rect 12342 4972 12348 4984
rect 12400 4972 12406 5024
rect 12434 4972 12440 5024
rect 12492 5012 12498 5024
rect 13740 5012 13768 5052
rect 14458 5012 14464 5024
rect 12492 4984 13768 5012
rect 14419 4984 14464 5012
rect 12492 4972 12498 4984
rect 14458 4972 14464 4984
rect 14516 4972 14522 5024
rect 14568 5012 14596 5052
rect 15102 5040 15108 5092
rect 15160 5080 15166 5092
rect 15212 5080 15240 5111
rect 15160 5052 15240 5080
rect 15160 5040 15166 5052
rect 15396 5012 15424 5256
rect 15838 5244 15844 5256
rect 15896 5244 15902 5296
rect 15654 5216 15660 5228
rect 15615 5188 15660 5216
rect 15654 5176 15660 5188
rect 15712 5176 15718 5228
rect 14568 4984 15424 5012
rect 1104 4922 16008 4944
rect 1104 4870 2824 4922
rect 2876 4870 2888 4922
rect 2940 4870 2952 4922
rect 3004 4870 3016 4922
rect 3068 4870 3080 4922
rect 3132 4870 6572 4922
rect 6624 4870 6636 4922
rect 6688 4870 6700 4922
rect 6752 4870 6764 4922
rect 6816 4870 6828 4922
rect 6880 4870 10320 4922
rect 10372 4870 10384 4922
rect 10436 4870 10448 4922
rect 10500 4870 10512 4922
rect 10564 4870 10576 4922
rect 10628 4870 14068 4922
rect 14120 4870 14132 4922
rect 14184 4870 14196 4922
rect 14248 4870 14260 4922
rect 14312 4870 14324 4922
rect 14376 4870 16008 4922
rect 1104 4848 16008 4870
rect 1670 4808 1676 4820
rect 1631 4780 1676 4808
rect 1670 4768 1676 4780
rect 1728 4768 1734 4820
rect 2406 4808 2412 4820
rect 2367 4780 2412 4808
rect 2406 4768 2412 4780
rect 2464 4768 2470 4820
rect 2590 4768 2596 4820
rect 2648 4808 2654 4820
rect 3789 4811 3847 4817
rect 3789 4808 3801 4811
rect 2648 4780 3801 4808
rect 2648 4768 2654 4780
rect 3789 4777 3801 4780
rect 3835 4777 3847 4811
rect 3789 4771 3847 4777
rect 4522 4768 4528 4820
rect 4580 4808 4586 4820
rect 5442 4808 5448 4820
rect 4580 4780 5448 4808
rect 4580 4768 4586 4780
rect 5442 4768 5448 4780
rect 5500 4768 5506 4820
rect 5537 4811 5595 4817
rect 5537 4777 5549 4811
rect 5583 4808 5595 4811
rect 6270 4808 6276 4820
rect 5583 4780 6276 4808
rect 5583 4777 5595 4780
rect 5537 4771 5595 4777
rect 6270 4768 6276 4780
rect 6328 4768 6334 4820
rect 6362 4768 6368 4820
rect 6420 4808 6426 4820
rect 6546 4808 6552 4820
rect 6420 4780 6552 4808
rect 6420 4768 6426 4780
rect 6546 4768 6552 4780
rect 6604 4768 6610 4820
rect 6641 4811 6699 4817
rect 6641 4777 6653 4811
rect 6687 4808 6699 4811
rect 7282 4808 7288 4820
rect 6687 4780 7288 4808
rect 6687 4777 6699 4780
rect 6641 4771 6699 4777
rect 7282 4768 7288 4780
rect 7340 4768 7346 4820
rect 8297 4811 8355 4817
rect 8297 4777 8309 4811
rect 8343 4808 8355 4811
rect 8343 4780 8984 4808
rect 8343 4777 8355 4780
rect 8297 4771 8355 4777
rect 8956 4752 8984 4780
rect 9030 4768 9036 4820
rect 9088 4808 9094 4820
rect 9401 4811 9459 4817
rect 9401 4808 9413 4811
rect 9088 4780 9413 4808
rect 9088 4768 9094 4780
rect 9401 4777 9413 4780
rect 9447 4777 9459 4811
rect 9401 4771 9459 4777
rect 9677 4811 9735 4817
rect 9677 4777 9689 4811
rect 9723 4808 9735 4811
rect 9766 4808 9772 4820
rect 9723 4780 9772 4808
rect 9723 4777 9735 4780
rect 9677 4771 9735 4777
rect 9766 4768 9772 4780
rect 9824 4768 9830 4820
rect 10505 4811 10563 4817
rect 10505 4777 10517 4811
rect 10551 4808 10563 4811
rect 10962 4808 10968 4820
rect 10551 4780 10968 4808
rect 10551 4777 10563 4780
rect 10505 4771 10563 4777
rect 10962 4768 10968 4780
rect 11020 4768 11026 4820
rect 11054 4768 11060 4820
rect 11112 4808 11118 4820
rect 11330 4808 11336 4820
rect 11112 4780 11336 4808
rect 11112 4768 11118 4780
rect 11330 4768 11336 4780
rect 11388 4768 11394 4820
rect 12342 4808 12348 4820
rect 11716 4780 12348 4808
rect 1578 4740 1584 4752
rect 1539 4712 1584 4740
rect 1578 4700 1584 4712
rect 1636 4700 1642 4752
rect 3326 4700 3332 4752
rect 3384 4740 3390 4752
rect 3421 4743 3479 4749
rect 3421 4740 3433 4743
rect 3384 4712 3433 4740
rect 3384 4700 3390 4712
rect 3421 4709 3433 4712
rect 3467 4740 3479 4743
rect 3602 4740 3608 4752
rect 3467 4712 3608 4740
rect 3467 4709 3479 4712
rect 3421 4703 3479 4709
rect 3602 4700 3608 4712
rect 3660 4700 3666 4752
rect 6822 4740 6828 4752
rect 4273 4712 6828 4740
rect 2590 4672 2596 4684
rect 2148 4644 2596 4672
rect 1394 4604 1400 4616
rect 1355 4576 1400 4604
rect 1394 4564 1400 4576
rect 1452 4564 1458 4616
rect 2148 4613 2176 4644
rect 2590 4632 2596 4644
rect 2648 4632 2654 4684
rect 3237 4675 3295 4681
rect 3237 4641 3249 4675
rect 3283 4672 3295 4675
rect 4273 4672 4301 4712
rect 6822 4700 6828 4712
rect 6880 4700 6886 4752
rect 8754 4700 8760 4752
rect 8812 4740 8818 4752
rect 8812 4712 8892 4740
rect 8812 4700 8818 4712
rect 4430 4672 4436 4684
rect 3283 4644 4301 4672
rect 4391 4644 4436 4672
rect 3283 4641 3295 4644
rect 3237 4635 3295 4641
rect 4430 4632 4436 4644
rect 4488 4632 4494 4684
rect 4982 4672 4988 4684
rect 4943 4644 4988 4672
rect 4982 4632 4988 4644
rect 5040 4632 5046 4684
rect 5077 4675 5135 4681
rect 5077 4641 5089 4675
rect 5123 4672 5135 4675
rect 5810 4672 5816 4684
rect 5123 4644 5816 4672
rect 5123 4641 5135 4644
rect 5077 4635 5135 4641
rect 5810 4632 5816 4644
rect 5868 4632 5874 4684
rect 6270 4672 6276 4684
rect 6231 4644 6276 4672
rect 6270 4632 6276 4644
rect 6328 4632 6334 4684
rect 6454 4672 6460 4684
rect 6415 4644 6460 4672
rect 6454 4632 6460 4644
rect 6512 4632 6518 4684
rect 7098 4672 7104 4684
rect 7059 4644 7104 4672
rect 7098 4632 7104 4644
rect 7156 4632 7162 4684
rect 7282 4672 7288 4684
rect 7243 4644 7288 4672
rect 7282 4632 7288 4644
rect 7340 4632 7346 4684
rect 7926 4672 7932 4684
rect 7887 4644 7932 4672
rect 7926 4632 7932 4644
rect 7984 4632 7990 4684
rect 8018 4632 8024 4684
rect 8076 4672 8082 4684
rect 8864 4672 8892 4712
rect 8938 4700 8944 4752
rect 8996 4700 9002 4752
rect 9490 4700 9496 4752
rect 9548 4740 9554 4752
rect 11425 4743 11483 4749
rect 11425 4740 11437 4743
rect 9548 4712 11437 4740
rect 9548 4700 9554 4712
rect 11425 4709 11437 4712
rect 11471 4709 11483 4743
rect 11425 4703 11483 4709
rect 9858 4672 9864 4684
rect 8076 4644 8121 4672
rect 8864 4644 9864 4672
rect 8076 4632 8082 4644
rect 9858 4632 9864 4644
rect 9916 4632 9922 4684
rect 10045 4675 10103 4681
rect 10045 4641 10057 4675
rect 10091 4672 10103 4675
rect 10686 4672 10692 4684
rect 10091 4644 10692 4672
rect 10091 4641 10103 4644
rect 10045 4635 10103 4641
rect 10686 4632 10692 4644
rect 10744 4632 10750 4684
rect 10778 4632 10784 4684
rect 10836 4672 10842 4684
rect 11149 4675 11207 4681
rect 11149 4672 11161 4675
rect 10836 4644 11161 4672
rect 10836 4632 10842 4644
rect 11149 4641 11161 4644
rect 11195 4641 11207 4675
rect 11149 4635 11207 4641
rect 1857 4607 1915 4613
rect 1857 4573 1869 4607
rect 1903 4573 1915 4607
rect 1857 4567 1915 4573
rect 2133 4607 2191 4613
rect 2133 4573 2145 4607
rect 2179 4573 2191 4607
rect 2133 4567 2191 4573
rect 1872 4536 1900 4567
rect 2222 4564 2228 4616
rect 2280 4604 2286 4616
rect 4249 4607 4307 4613
rect 2280 4576 2325 4604
rect 2280 4564 2286 4576
rect 4249 4573 4261 4607
rect 4295 4604 4307 4607
rect 5718 4604 5724 4616
rect 4295 4576 5724 4604
rect 4295 4573 4307 4576
rect 4249 4567 4307 4573
rect 5718 4564 5724 4576
rect 5776 4564 5782 4616
rect 5902 4564 5908 4616
rect 5960 4604 5966 4616
rect 6181 4607 6239 4613
rect 6181 4604 6193 4607
rect 5960 4576 6193 4604
rect 5960 4564 5966 4576
rect 6181 4573 6193 4576
rect 6227 4573 6239 4607
rect 6181 4567 6239 4573
rect 6914 4564 6920 4616
rect 6972 4604 6978 4616
rect 7009 4607 7067 4613
rect 7009 4604 7021 4607
rect 6972 4576 7021 4604
rect 6972 4564 6978 4576
rect 7009 4573 7021 4576
rect 7055 4573 7067 4607
rect 7009 4567 7067 4573
rect 7466 4564 7472 4616
rect 7524 4604 7530 4616
rect 7837 4607 7895 4613
rect 7837 4604 7849 4607
rect 7524 4576 7849 4604
rect 7524 4564 7530 4576
rect 7837 4573 7849 4576
rect 7883 4573 7895 4607
rect 8457 4607 8515 4613
rect 8457 4604 8469 4607
rect 7944 4592 8469 4604
rect 7837 4567 7895 4573
rect 2406 4536 2412 4548
rect 1872 4508 2412 4536
rect 2406 4496 2412 4508
rect 2464 4496 2470 4548
rect 2593 4539 2651 4545
rect 2593 4505 2605 4539
rect 2639 4536 2651 4539
rect 2682 4536 2688 4548
rect 2639 4508 2688 4536
rect 2639 4505 2651 4508
rect 2593 4499 2651 4505
rect 2682 4496 2688 4508
rect 2740 4496 2746 4548
rect 2777 4539 2835 4545
rect 2777 4505 2789 4539
rect 2823 4536 2835 4539
rect 3234 4536 3240 4548
rect 2823 4508 3240 4536
rect 2823 4505 2835 4508
rect 2777 4499 2835 4505
rect 1949 4471 2007 4477
rect 1949 4437 1961 4471
rect 1995 4468 2007 4471
rect 2038 4468 2044 4480
rect 1995 4440 2044 4468
rect 1995 4437 2007 4440
rect 1949 4431 2007 4437
rect 2038 4428 2044 4440
rect 2096 4428 2102 4480
rect 2498 4428 2504 4480
rect 2556 4468 2562 4480
rect 2792 4468 2820 4499
rect 3234 4496 3240 4508
rect 3292 4536 3298 4548
rect 3510 4536 3516 4548
rect 3292 4508 3516 4536
rect 3292 4496 3298 4508
rect 3510 4496 3516 4508
rect 3568 4496 3574 4548
rect 4709 4539 4767 4545
rect 4709 4505 4721 4539
rect 4755 4536 4767 4539
rect 5534 4536 5540 4548
rect 4755 4508 5540 4536
rect 4755 4505 4767 4508
rect 4709 4499 4767 4505
rect 5534 4496 5540 4508
rect 5592 4496 5598 4548
rect 5629 4539 5687 4545
rect 7926 4540 7932 4592
rect 7984 4576 8469 4592
rect 7984 4540 7990 4576
rect 8457 4573 8469 4576
rect 8503 4573 8515 4607
rect 8457 4567 8515 4573
rect 5629 4505 5641 4539
rect 5675 4536 5687 4539
rect 5675 4508 6132 4536
rect 5675 4505 5687 4508
rect 5629 4499 5687 4505
rect 3050 4468 3056 4480
rect 2556 4440 2820 4468
rect 3011 4440 3056 4468
rect 2556 4428 2562 4440
rect 3050 4428 3056 4440
rect 3108 4428 3114 4480
rect 3605 4471 3663 4477
rect 3605 4437 3617 4471
rect 3651 4468 3663 4471
rect 3786 4468 3792 4480
rect 3651 4440 3792 4468
rect 3651 4437 3663 4440
rect 3605 4431 3663 4437
rect 3786 4428 3792 4440
rect 3844 4428 3850 4480
rect 4154 4468 4160 4480
rect 4115 4440 4160 4468
rect 4154 4428 4160 4440
rect 4212 4428 4218 4480
rect 5169 4471 5227 4477
rect 5169 4437 5181 4471
rect 5215 4468 5227 4471
rect 5442 4468 5448 4480
rect 5215 4440 5448 4468
rect 5215 4437 5227 4440
rect 5169 4431 5227 4437
rect 5442 4428 5448 4440
rect 5500 4428 5506 4480
rect 5813 4471 5871 4477
rect 5813 4437 5825 4471
rect 5859 4468 5871 4471
rect 5902 4468 5908 4480
rect 5859 4440 5908 4468
rect 5859 4437 5871 4440
rect 5813 4431 5871 4437
rect 5902 4428 5908 4440
rect 5960 4428 5966 4480
rect 6104 4468 6132 4508
rect 8294 4496 8300 4548
rect 8352 4536 8358 4548
rect 8570 4540 8576 4592
rect 8628 4580 8634 4592
rect 8628 4552 8673 4580
rect 8754 4564 8760 4616
rect 8812 4600 8818 4616
rect 9309 4607 9367 4613
rect 8864 4600 9076 4604
rect 8812 4576 9076 4600
rect 8812 4572 8892 4576
rect 8812 4564 8818 4572
rect 8628 4540 8634 4552
rect 8352 4508 8524 4536
rect 8352 4496 8358 4508
rect 7098 4468 7104 4480
rect 6104 4440 7104 4468
rect 7098 4428 7104 4440
rect 7156 4428 7162 4480
rect 7282 4428 7288 4480
rect 7340 4468 7346 4480
rect 7469 4471 7527 4477
rect 7469 4468 7481 4471
rect 7340 4440 7481 4468
rect 7340 4428 7346 4440
rect 7469 4437 7481 4440
rect 7515 4437 7527 4471
rect 7469 4431 7527 4437
rect 7742 4428 7748 4480
rect 7800 4468 7806 4480
rect 8386 4468 8392 4480
rect 7800 4440 8392 4468
rect 7800 4428 7806 4440
rect 8386 4428 8392 4440
rect 8444 4428 8450 4480
rect 8496 4468 8524 4508
rect 9048 4477 9076 4576
rect 9309 4573 9321 4607
rect 9355 4604 9367 4607
rect 9582 4604 9588 4616
rect 9355 4576 9588 4604
rect 9355 4573 9367 4576
rect 9309 4567 9367 4573
rect 9582 4564 9588 4576
rect 9640 4604 9646 4616
rect 10965 4607 11023 4613
rect 9640 4576 9904 4604
rect 9640 4564 9646 4576
rect 9876 4548 9904 4576
rect 10965 4573 10977 4607
rect 11011 4604 11023 4607
rect 11716 4604 11744 4780
rect 12342 4768 12348 4780
rect 12400 4768 12406 4820
rect 12710 4808 12716 4820
rect 12671 4780 12716 4808
rect 12710 4768 12716 4780
rect 12768 4768 12774 4820
rect 13906 4808 13912 4820
rect 13867 4780 13912 4808
rect 13906 4768 13912 4780
rect 13964 4768 13970 4820
rect 14550 4808 14556 4820
rect 14511 4780 14556 4808
rect 14550 4768 14556 4780
rect 14608 4768 14614 4820
rect 14642 4768 14648 4820
rect 14700 4808 14706 4820
rect 15470 4808 15476 4820
rect 14700 4780 15476 4808
rect 14700 4768 14706 4780
rect 15470 4768 15476 4780
rect 15528 4768 15534 4820
rect 12066 4700 12072 4752
rect 12124 4740 12130 4752
rect 12124 4712 14320 4740
rect 12124 4700 12130 4712
rect 11977 4675 12035 4681
rect 11977 4641 11989 4675
rect 12023 4672 12035 4675
rect 12529 4675 12587 4681
rect 12529 4672 12541 4675
rect 12023 4644 12541 4672
rect 12023 4641 12035 4644
rect 11977 4635 12035 4641
rect 12529 4641 12541 4644
rect 12575 4672 12587 4675
rect 12894 4672 12900 4684
rect 12575 4644 12900 4672
rect 12575 4641 12587 4644
rect 12529 4635 12587 4641
rect 12894 4632 12900 4644
rect 12952 4632 12958 4684
rect 13170 4632 13176 4684
rect 13228 4632 13234 4684
rect 13354 4672 13360 4684
rect 13315 4644 13360 4672
rect 13354 4632 13360 4644
rect 13412 4632 13418 4684
rect 13446 4632 13452 4684
rect 13504 4672 13510 4684
rect 13722 4672 13728 4684
rect 13504 4644 13728 4672
rect 13504 4632 13510 4644
rect 13722 4632 13728 4644
rect 13780 4632 13786 4684
rect 14292 4681 14320 4712
rect 14277 4675 14335 4681
rect 14277 4641 14289 4675
rect 14323 4641 14335 4675
rect 15010 4672 15016 4684
rect 14971 4644 15016 4672
rect 14277 4635 14335 4641
rect 15010 4632 15016 4644
rect 15068 4632 15074 4684
rect 15102 4632 15108 4684
rect 15160 4672 15166 4684
rect 15160 4644 15205 4672
rect 15160 4632 15166 4644
rect 11011 4576 11744 4604
rect 11793 4607 11851 4613
rect 11011 4573 11023 4576
rect 10965 4567 11023 4573
rect 11793 4573 11805 4607
rect 11839 4604 11851 4607
rect 12066 4604 12072 4616
rect 11839 4576 12072 4604
rect 11839 4573 11851 4576
rect 11793 4567 11851 4573
rect 12066 4564 12072 4576
rect 12124 4564 12130 4616
rect 12250 4564 12256 4616
rect 12308 4564 12314 4616
rect 12437 4607 12495 4613
rect 12437 4573 12449 4607
rect 12483 4604 12495 4607
rect 13188 4604 13216 4632
rect 12483 4576 13216 4604
rect 12483 4573 12495 4576
rect 12437 4567 12495 4573
rect 14090 4564 14096 4616
rect 14148 4604 14154 4616
rect 15381 4607 15439 4613
rect 15381 4604 15393 4607
rect 14148 4576 15393 4604
rect 14148 4564 14154 4576
rect 15381 4573 15393 4576
rect 15427 4573 15439 4607
rect 15381 4567 15439 4573
rect 9858 4496 9864 4548
rect 9916 4536 9922 4548
rect 10137 4539 10195 4545
rect 10137 4536 10149 4539
rect 9916 4508 10149 4536
rect 9916 4496 9922 4508
rect 10137 4505 10149 4508
rect 10183 4505 10195 4539
rect 11054 4536 11060 4548
rect 10137 4499 10195 4505
rect 10437 4508 10732 4536
rect 11015 4508 11060 4536
rect 8757 4471 8815 4477
rect 8757 4468 8769 4471
rect 8496 4440 8769 4468
rect 8757 4437 8769 4440
rect 8803 4437 8815 4471
rect 8757 4431 8815 4437
rect 9033 4471 9091 4477
rect 9033 4437 9045 4471
rect 9079 4468 9091 4471
rect 10437 4468 10465 4508
rect 10594 4468 10600 4480
rect 9079 4440 10465 4468
rect 10555 4440 10600 4468
rect 9079 4437 9091 4440
rect 9033 4431 9091 4437
rect 10594 4428 10600 4440
rect 10652 4428 10658 4480
rect 10704 4468 10732 4508
rect 11054 4496 11060 4508
rect 11112 4496 11118 4548
rect 12158 4536 12164 4548
rect 11164 4508 12164 4536
rect 11164 4468 11192 4508
rect 12158 4496 12164 4508
rect 12216 4496 12222 4548
rect 12268 4536 12296 4564
rect 12710 4536 12716 4548
rect 12268 4508 12716 4536
rect 12710 4496 12716 4508
rect 12768 4496 12774 4548
rect 13081 4539 13139 4545
rect 13081 4505 13093 4539
rect 13127 4536 13139 4539
rect 13541 4539 13599 4545
rect 13541 4536 13553 4539
rect 13127 4508 13553 4536
rect 13127 4505 13139 4508
rect 13081 4499 13139 4505
rect 13541 4505 13553 4508
rect 13587 4505 13599 4539
rect 13541 4499 13599 4505
rect 13722 4496 13728 4548
rect 13780 4536 13786 4548
rect 14185 4539 14243 4545
rect 14185 4536 14197 4539
rect 13780 4508 14197 4536
rect 13780 4496 13786 4508
rect 14185 4505 14197 4508
rect 14231 4505 14243 4539
rect 14185 4499 14243 4505
rect 14826 4496 14832 4548
rect 14884 4536 14890 4548
rect 14921 4539 14979 4545
rect 14921 4536 14933 4539
rect 14884 4508 14933 4536
rect 14884 4496 14890 4508
rect 14921 4505 14933 4508
rect 14967 4505 14979 4539
rect 14921 4499 14979 4505
rect 10704 4440 11192 4468
rect 11330 4428 11336 4480
rect 11388 4468 11394 4480
rect 11885 4471 11943 4477
rect 11885 4468 11897 4471
rect 11388 4440 11897 4468
rect 11388 4428 11394 4440
rect 11885 4437 11897 4440
rect 11931 4437 11943 4471
rect 11885 4431 11943 4437
rect 11974 4428 11980 4480
rect 12032 4468 12038 4480
rect 12253 4471 12311 4477
rect 12253 4468 12265 4471
rect 12032 4440 12265 4468
rect 12032 4428 12038 4440
rect 12253 4437 12265 4440
rect 12299 4437 12311 4471
rect 12253 4431 12311 4437
rect 12986 4428 12992 4480
rect 13044 4468 13050 4480
rect 13173 4471 13231 4477
rect 13173 4468 13185 4471
rect 13044 4440 13185 4468
rect 13044 4428 13050 4440
rect 13173 4437 13185 4440
rect 13219 4437 13231 4471
rect 13173 4431 13231 4437
rect 15102 4428 15108 4480
rect 15160 4468 15166 4480
rect 15565 4471 15623 4477
rect 15565 4468 15577 4471
rect 15160 4440 15577 4468
rect 15160 4428 15166 4440
rect 15565 4437 15577 4440
rect 15611 4437 15623 4471
rect 15565 4431 15623 4437
rect 1104 4378 16008 4400
rect 1104 4326 4698 4378
rect 4750 4326 4762 4378
rect 4814 4326 4826 4378
rect 4878 4326 4890 4378
rect 4942 4326 4954 4378
rect 5006 4326 8446 4378
rect 8498 4326 8510 4378
rect 8562 4326 8574 4378
rect 8626 4326 8638 4378
rect 8690 4326 8702 4378
rect 8754 4326 12194 4378
rect 12246 4326 12258 4378
rect 12310 4326 12322 4378
rect 12374 4326 12386 4378
rect 12438 4326 12450 4378
rect 12502 4326 16008 4378
rect 1104 4304 16008 4326
rect 1854 4264 1860 4276
rect 1815 4236 1860 4264
rect 1854 4224 1860 4236
rect 1912 4224 1918 4276
rect 1946 4224 1952 4276
rect 2004 4264 2010 4276
rect 2314 4264 2320 4276
rect 2004 4236 2320 4264
rect 2004 4224 2010 4236
rect 2314 4224 2320 4236
rect 2372 4224 2378 4276
rect 3050 4224 3056 4276
rect 3108 4264 3114 4276
rect 3694 4264 3700 4276
rect 3108 4236 3700 4264
rect 3108 4224 3114 4236
rect 3694 4224 3700 4236
rect 3752 4224 3758 4276
rect 4338 4224 4344 4276
rect 4396 4264 4402 4276
rect 4522 4264 4528 4276
rect 4396 4236 4528 4264
rect 4396 4224 4402 4236
rect 4522 4224 4528 4236
rect 4580 4224 4586 4276
rect 5534 4224 5540 4276
rect 5592 4264 5598 4276
rect 8846 4264 8852 4276
rect 5592 4236 6316 4264
rect 5592 4224 5598 4236
rect 1489 4199 1547 4205
rect 1489 4165 1501 4199
rect 1535 4196 1547 4199
rect 3068 4196 3096 4224
rect 3970 4196 3976 4208
rect 1535 4168 3096 4196
rect 3436 4168 3976 4196
rect 1535 4165 1547 4168
rect 1489 4159 1547 4165
rect 1946 4128 1952 4140
rect 1907 4100 1952 4128
rect 1946 4088 1952 4100
rect 2004 4088 2010 4140
rect 2593 4131 2651 4137
rect 2593 4128 2605 4131
rect 2332 4100 2605 4128
rect 1762 4060 1768 4072
rect 1723 4032 1768 4060
rect 1762 4020 1768 4032
rect 1820 4020 1826 4072
rect 2332 4001 2360 4100
rect 2593 4097 2605 4100
rect 2639 4097 2651 4131
rect 2866 4128 2872 4140
rect 2827 4100 2872 4128
rect 2593 4091 2651 4097
rect 2866 4088 2872 4100
rect 2924 4088 2930 4140
rect 3145 4131 3203 4137
rect 3145 4097 3157 4131
rect 3191 4128 3203 4131
rect 3234 4128 3240 4140
rect 3191 4100 3240 4128
rect 3191 4097 3203 4100
rect 3145 4091 3203 4097
rect 3234 4088 3240 4100
rect 3292 4088 3298 4140
rect 3326 4088 3332 4140
rect 3384 4088 3390 4140
rect 3436 4137 3464 4168
rect 3970 4156 3976 4168
rect 4028 4156 4034 4208
rect 4154 4156 4160 4208
rect 4212 4196 4218 4208
rect 5629 4199 5687 4205
rect 4212 4168 5304 4196
rect 4212 4156 4218 4168
rect 5276 4140 5304 4168
rect 5629 4165 5641 4199
rect 5675 4196 5687 4199
rect 5718 4196 5724 4208
rect 5675 4168 5724 4196
rect 5675 4165 5687 4168
rect 5629 4159 5687 4165
rect 5718 4156 5724 4168
rect 5776 4156 5782 4208
rect 6288 4196 6316 4236
rect 6656 4236 8852 4264
rect 6656 4196 6684 4236
rect 8846 4224 8852 4236
rect 8904 4224 8910 4276
rect 10042 4224 10048 4276
rect 10100 4264 10106 4276
rect 10137 4267 10195 4273
rect 10137 4264 10149 4267
rect 10100 4236 10149 4264
rect 10100 4224 10106 4236
rect 10137 4233 10149 4236
rect 10183 4233 10195 4267
rect 10137 4227 10195 4233
rect 10505 4267 10563 4273
rect 10505 4233 10517 4267
rect 10551 4264 10563 4267
rect 11885 4267 11943 4273
rect 11885 4264 11897 4267
rect 10551 4236 11897 4264
rect 10551 4233 10563 4236
rect 10505 4227 10563 4233
rect 11885 4233 11897 4236
rect 11931 4233 11943 4267
rect 11885 4227 11943 4233
rect 12894 4224 12900 4276
rect 12952 4264 12958 4276
rect 13173 4267 13231 4273
rect 13173 4264 13185 4267
rect 12952 4236 13185 4264
rect 12952 4224 12958 4236
rect 13173 4233 13185 4236
rect 13219 4233 13231 4267
rect 13173 4227 13231 4233
rect 13446 4224 13452 4276
rect 13504 4264 13510 4276
rect 13906 4264 13912 4276
rect 13504 4236 13912 4264
rect 13504 4224 13510 4236
rect 13906 4224 13912 4236
rect 13964 4224 13970 4276
rect 14826 4224 14832 4276
rect 14884 4264 14890 4276
rect 14921 4267 14979 4273
rect 14921 4264 14933 4267
rect 14884 4236 14933 4264
rect 14884 4224 14890 4236
rect 14921 4233 14933 4236
rect 14967 4233 14979 4267
rect 14921 4227 14979 4233
rect 6288 4168 6684 4196
rect 6733 4199 6791 4205
rect 6733 4165 6745 4199
rect 6779 4196 6791 4199
rect 7558 4196 7564 4208
rect 6779 4168 7564 4196
rect 6779 4165 6791 4168
rect 6733 4159 6791 4165
rect 7558 4156 7564 4168
rect 7616 4156 7622 4208
rect 8941 4199 8999 4205
rect 8941 4165 8953 4199
rect 8987 4196 8999 4199
rect 10594 4196 10600 4208
rect 8987 4168 10600 4196
rect 8987 4165 8999 4168
rect 3421 4131 3479 4137
rect 3421 4097 3433 4131
rect 3467 4097 3479 4131
rect 3421 4091 3479 4097
rect 3881 4131 3939 4137
rect 3881 4097 3893 4131
rect 3927 4097 3939 4131
rect 3881 4091 3939 4097
rect 3344 4060 3372 4088
rect 3605 4063 3663 4069
rect 3605 4060 3617 4063
rect 3344 4032 3617 4060
rect 3605 4029 3617 4032
rect 3651 4029 3663 4063
rect 3786 4060 3792 4072
rect 3747 4032 3792 4060
rect 3605 4023 3663 4029
rect 3786 4020 3792 4032
rect 3844 4020 3850 4072
rect 2317 3995 2375 4001
rect 2317 3961 2329 3995
rect 2363 3961 2375 3995
rect 2317 3955 2375 3961
rect 2961 3995 3019 4001
rect 2961 3961 2973 3995
rect 3007 3992 3019 3995
rect 3326 3992 3332 4004
rect 3007 3964 3332 3992
rect 3007 3961 3019 3964
rect 2961 3955 3019 3961
rect 3326 3952 3332 3964
rect 3384 3952 3390 4004
rect 3896 3936 3924 4091
rect 4062 4088 4068 4140
rect 4120 4128 4126 4140
rect 4709 4131 4767 4137
rect 4709 4128 4721 4131
rect 4120 4100 4721 4128
rect 4120 4088 4126 4100
rect 4709 4097 4721 4100
rect 4755 4097 4767 4131
rect 4709 4091 4767 4097
rect 4801 4131 4859 4137
rect 4801 4097 4813 4131
rect 4847 4128 4859 4131
rect 4847 4100 5212 4128
rect 4847 4097 4859 4100
rect 4801 4091 4859 4097
rect 4985 4063 5043 4069
rect 4985 4029 4997 4063
rect 5031 4029 5043 4063
rect 5184 4060 5212 4100
rect 5258 4088 5264 4140
rect 5316 4128 5322 4140
rect 5537 4131 5595 4137
rect 5537 4128 5549 4131
rect 5316 4100 5549 4128
rect 5316 4088 5322 4100
rect 5537 4097 5549 4100
rect 5583 4097 5595 4131
rect 6173 4131 6231 4137
rect 5537 4091 5595 4097
rect 5745 4100 6049 4128
rect 5745 4060 5773 4100
rect 5184 4032 5773 4060
rect 5813 4063 5871 4069
rect 4985 4023 5043 4029
rect 5813 4029 5825 4063
rect 5859 4029 5871 4063
rect 6021 4060 6049 4100
rect 6173 4097 6185 4131
rect 6219 4128 6231 4131
rect 6362 4128 6368 4140
rect 6219 4100 6368 4128
rect 6219 4097 6231 4100
rect 6173 4091 6231 4097
rect 6362 4088 6368 4100
rect 6420 4088 6426 4140
rect 7374 4128 7380 4140
rect 7335 4100 7380 4128
rect 7374 4088 7380 4100
rect 7432 4088 7438 4140
rect 7466 4088 7472 4140
rect 7524 4128 7530 4140
rect 7653 4131 7711 4137
rect 7653 4128 7665 4131
rect 7524 4100 7665 4128
rect 7524 4088 7530 4100
rect 7653 4097 7665 4100
rect 7699 4097 7711 4131
rect 8110 4128 8116 4140
rect 8071 4100 8116 4128
rect 7653 4091 7711 4097
rect 8110 4088 8116 4100
rect 8168 4088 8174 4140
rect 8202 4112 8208 4164
rect 8260 4128 8266 4164
rect 8941 4159 8999 4165
rect 10594 4156 10600 4168
rect 10652 4156 10658 4208
rect 12805 4199 12863 4205
rect 10796 4168 12388 4196
rect 8260 4112 9168 4128
rect 8220 4100 9168 4112
rect 6825 4063 6883 4069
rect 6021 4032 6132 4060
rect 5813 4023 5871 4029
rect 4246 3992 4252 4004
rect 4207 3964 4252 3992
rect 4246 3952 4252 3964
rect 4304 3952 4310 4004
rect 5000 3992 5028 4023
rect 5350 3992 5356 4004
rect 5000 3964 5356 3992
rect 5350 3952 5356 3964
rect 5408 3992 5414 4004
rect 5828 3992 5856 4023
rect 6104 4004 6132 4032
rect 6825 4029 6837 4063
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 6917 4063 6975 4069
rect 6917 4029 6929 4063
rect 6963 4029 6975 4063
rect 6917 4023 6975 4029
rect 5408 3964 5856 3992
rect 5408 3952 5414 3964
rect 6086 3952 6092 4004
rect 6144 3952 6150 4004
rect 6840 3992 6868 4023
rect 6472 3964 6868 3992
rect 6472 3936 6500 3964
rect 1670 3884 1676 3936
rect 1728 3924 1734 3936
rect 2409 3927 2467 3933
rect 2409 3924 2421 3927
rect 1728 3896 2421 3924
rect 1728 3884 1734 3896
rect 2409 3893 2421 3896
rect 2455 3893 2467 3927
rect 2409 3887 2467 3893
rect 2590 3884 2596 3936
rect 2648 3924 2654 3936
rect 2685 3927 2743 3933
rect 2685 3924 2697 3927
rect 2648 3896 2697 3924
rect 2648 3884 2654 3896
rect 2685 3893 2697 3896
rect 2731 3893 2743 3927
rect 3234 3924 3240 3936
rect 3195 3896 3240 3924
rect 2685 3887 2743 3893
rect 3234 3884 3240 3896
rect 3292 3884 3298 3936
rect 3878 3884 3884 3936
rect 3936 3884 3942 3936
rect 4341 3927 4399 3933
rect 4341 3893 4353 3927
rect 4387 3924 4399 3927
rect 4430 3924 4436 3936
rect 4387 3896 4436 3924
rect 4387 3893 4399 3896
rect 4341 3887 4399 3893
rect 4430 3884 4436 3896
rect 4488 3884 4494 3936
rect 4522 3884 4528 3936
rect 4580 3924 4586 3936
rect 5169 3927 5227 3933
rect 5169 3924 5181 3927
rect 4580 3896 5181 3924
rect 4580 3884 4586 3896
rect 5169 3893 5181 3896
rect 5215 3893 5227 3927
rect 5169 3887 5227 3893
rect 5258 3884 5264 3936
rect 5316 3924 5322 3936
rect 5997 3927 6055 3933
rect 5997 3924 6009 3927
rect 5316 3896 6009 3924
rect 5316 3884 5322 3896
rect 5997 3893 6009 3896
rect 6043 3893 6055 3927
rect 5997 3887 6055 3893
rect 6270 3884 6276 3936
rect 6328 3924 6334 3936
rect 6365 3927 6423 3933
rect 6365 3924 6377 3927
rect 6328 3896 6377 3924
rect 6328 3884 6334 3896
rect 6365 3893 6377 3896
rect 6411 3893 6423 3927
rect 6365 3887 6423 3893
rect 6454 3884 6460 3936
rect 6512 3884 6518 3936
rect 6638 3884 6644 3936
rect 6696 3924 6702 3936
rect 6932 3924 6960 4023
rect 7190 4020 7196 4072
rect 7248 4060 7254 4072
rect 7834 4060 7840 4072
rect 7248 4032 7840 4060
rect 7248 4020 7254 4032
rect 7834 4020 7840 4032
rect 7892 4020 7898 4072
rect 8021 4063 8079 4069
rect 8021 4029 8033 4063
rect 8067 4060 8079 4063
rect 8202 4060 8208 4072
rect 8067 4032 8208 4060
rect 8067 4029 8079 4032
rect 8021 4023 8079 4029
rect 8202 4020 8208 4032
rect 8260 4020 8266 4072
rect 8662 4060 8668 4072
rect 8404 4032 8668 4060
rect 7098 3952 7104 4004
rect 7156 3992 7162 4004
rect 8404 3992 8432 4032
rect 8662 4020 8668 4032
rect 8720 4020 8726 4072
rect 9030 4060 9036 4072
rect 8991 4032 9036 4060
rect 9030 4020 9036 4032
rect 9088 4020 9094 4072
rect 9140 4069 9168 4100
rect 9398 4088 9404 4140
rect 9456 4128 9462 4140
rect 9493 4131 9551 4137
rect 9493 4128 9505 4131
rect 9456 4100 9505 4128
rect 9456 4088 9462 4100
rect 9493 4097 9505 4100
rect 9539 4097 9551 4131
rect 9493 4091 9551 4097
rect 9766 4088 9772 4140
rect 9824 4128 9830 4140
rect 10045 4131 10103 4137
rect 10045 4128 10057 4131
rect 9824 4100 10057 4128
rect 9824 4088 9830 4100
rect 10045 4097 10057 4100
rect 10091 4097 10103 4131
rect 10796 4128 10824 4168
rect 10962 4128 10968 4140
rect 10045 4091 10103 4097
rect 10336 4100 10824 4128
rect 10923 4100 10968 4128
rect 10336 4072 10364 4100
rect 10962 4088 10968 4100
rect 11020 4088 11026 4140
rect 11330 4088 11336 4140
rect 11388 4128 11394 4140
rect 12250 4128 12256 4140
rect 11388 4100 12256 4128
rect 11388 4088 11394 4100
rect 12250 4088 12256 4100
rect 12308 4088 12314 4140
rect 9125 4063 9183 4069
rect 9125 4029 9137 4063
rect 9171 4029 9183 4063
rect 9953 4063 10011 4069
rect 9953 4060 9965 4063
rect 9125 4023 9183 4029
rect 9600 4032 9965 4060
rect 7156 3964 8432 3992
rect 8481 3995 8539 4001
rect 7156 3952 7162 3964
rect 8481 3961 8493 3995
rect 8527 3992 8539 3995
rect 9214 3992 9220 4004
rect 8527 3964 9220 3992
rect 8527 3961 8539 3964
rect 8481 3955 8539 3961
rect 9214 3952 9220 3964
rect 9272 3952 9278 4004
rect 7190 3924 7196 3936
rect 6696 3896 6960 3924
rect 7151 3896 7196 3924
rect 6696 3884 6702 3896
rect 7190 3884 7196 3896
rect 7248 3884 7254 3936
rect 7374 3884 7380 3936
rect 7432 3924 7438 3936
rect 7469 3927 7527 3933
rect 7469 3924 7481 3927
rect 7432 3896 7481 3924
rect 7432 3884 7438 3896
rect 7469 3893 7481 3896
rect 7515 3893 7527 3927
rect 7469 3887 7527 3893
rect 7834 3884 7840 3936
rect 7892 3924 7898 3936
rect 8573 3927 8631 3933
rect 8573 3924 8585 3927
rect 7892 3896 8585 3924
rect 7892 3884 7898 3896
rect 8573 3893 8585 3896
rect 8619 3893 8631 3927
rect 8573 3887 8631 3893
rect 8938 3884 8944 3936
rect 8996 3924 9002 3936
rect 9600 3924 9628 4032
rect 9953 4029 9965 4032
rect 9999 4060 10011 4063
rect 10318 4060 10324 4072
rect 9999 4032 10324 4060
rect 9999 4029 10011 4032
rect 9953 4023 10011 4029
rect 10318 4020 10324 4032
rect 10376 4020 10382 4072
rect 10778 4020 10784 4072
rect 10836 4060 10842 4072
rect 11057 4063 11115 4069
rect 11057 4060 11069 4063
rect 10836 4032 11069 4060
rect 10836 4020 10842 4032
rect 11057 4029 11069 4032
rect 11103 4029 11115 4063
rect 11057 4023 11115 4029
rect 11241 4063 11299 4069
rect 11241 4029 11253 4063
rect 11287 4060 11299 4063
rect 11422 4060 11428 4072
rect 11287 4032 11428 4060
rect 11287 4029 11299 4032
rect 11241 4023 11299 4029
rect 11422 4020 11428 4032
rect 11480 4020 11486 4072
rect 11977 4063 12035 4069
rect 11977 4029 11989 4063
rect 12023 4029 12035 4063
rect 12158 4060 12164 4072
rect 12119 4032 12164 4060
rect 11977 4023 12035 4029
rect 9677 3995 9735 4001
rect 9677 3961 9689 3995
rect 9723 3992 9735 3995
rect 11992 3992 12020 4023
rect 12158 4020 12164 4032
rect 12216 4020 12222 4072
rect 12360 4060 12388 4168
rect 12805 4165 12817 4199
rect 12851 4196 12863 4199
rect 13078 4196 13084 4208
rect 12851 4168 13084 4196
rect 12851 4165 12863 4168
rect 12805 4159 12863 4165
rect 13078 4156 13084 4168
rect 13136 4156 13142 4208
rect 15286 4196 15292 4208
rect 14108 4168 15292 4196
rect 12713 4131 12771 4137
rect 12713 4097 12725 4131
rect 12759 4128 12771 4131
rect 12986 4128 12992 4140
rect 12759 4100 12992 4128
rect 12759 4097 12771 4100
rect 12713 4091 12771 4097
rect 12986 4088 12992 4100
rect 13044 4088 13050 4140
rect 13170 4088 13176 4140
rect 13228 4128 13234 4140
rect 13372 4128 13492 4132
rect 13541 4131 13599 4137
rect 13541 4128 13553 4131
rect 13228 4104 13553 4128
rect 13228 4100 13400 4104
rect 13464 4100 13553 4104
rect 13228 4088 13234 4100
rect 13541 4097 13553 4100
rect 13587 4097 13599 4131
rect 13541 4091 13599 4097
rect 13814 4088 13820 4140
rect 13872 4128 13878 4140
rect 14001 4131 14059 4137
rect 14001 4128 14013 4131
rect 13872 4100 14013 4128
rect 13872 4088 13878 4100
rect 14001 4097 14013 4100
rect 14047 4097 14059 4131
rect 14001 4091 14059 4097
rect 12897 4063 12955 4069
rect 12360 4032 12664 4060
rect 12345 3995 12403 4001
rect 12345 3992 12357 3995
rect 9723 3964 11652 3992
rect 11992 3964 12357 3992
rect 9723 3961 9735 3964
rect 9677 3955 9735 3961
rect 10594 3924 10600 3936
rect 8996 3896 9628 3924
rect 10555 3896 10600 3924
rect 8996 3884 9002 3896
rect 10594 3884 10600 3896
rect 10652 3884 10658 3936
rect 11514 3924 11520 3936
rect 11475 3896 11520 3924
rect 11514 3884 11520 3896
rect 11572 3884 11578 3936
rect 11624 3924 11652 3964
rect 12345 3961 12357 3964
rect 12391 3961 12403 3995
rect 12636 3992 12664 4032
rect 12897 4029 12909 4063
rect 12943 4029 12955 4063
rect 13633 4063 13691 4069
rect 13633 4060 13645 4063
rect 12897 4023 12955 4029
rect 13280 4032 13645 4060
rect 12912 3992 12940 4023
rect 13280 4004 13308 4032
rect 13633 4029 13645 4032
rect 13679 4029 13691 4063
rect 13633 4023 13691 4029
rect 13725 4063 13783 4069
rect 13725 4029 13737 4063
rect 13771 4029 13783 4063
rect 13725 4023 13783 4029
rect 12636 3964 12940 3992
rect 12345 3955 12403 3961
rect 13262 3952 13268 4004
rect 13320 3952 13326 4004
rect 13354 3952 13360 4004
rect 13412 3992 13418 4004
rect 13740 3992 13768 4023
rect 13412 3964 13768 3992
rect 13412 3952 13418 3964
rect 13814 3952 13820 4004
rect 13872 3992 13878 4004
rect 14108 3992 14136 4168
rect 15286 4156 15292 4168
rect 15344 4156 15350 4208
rect 14461 4131 14519 4137
rect 14461 4097 14473 4131
rect 14507 4128 14519 4131
rect 15381 4131 15439 4137
rect 14507 4100 14964 4128
rect 14507 4097 14519 4100
rect 14461 4091 14519 4097
rect 14642 4060 14648 4072
rect 14603 4032 14648 4060
rect 14642 4020 14648 4032
rect 14700 4020 14706 4072
rect 14826 4060 14832 4072
rect 14787 4032 14832 4060
rect 14826 4020 14832 4032
rect 14884 4020 14890 4072
rect 14936 4060 14964 4100
rect 15381 4097 15393 4131
rect 15427 4128 15439 4131
rect 16114 4128 16120 4140
rect 15427 4100 16120 4128
rect 15427 4097 15439 4100
rect 15381 4091 15439 4097
rect 16114 4088 16120 4100
rect 16172 4088 16178 4140
rect 16390 4060 16396 4072
rect 14936 4032 16396 4060
rect 16390 4020 16396 4032
rect 16448 4020 16454 4072
rect 13872 3964 14136 3992
rect 14185 3995 14243 4001
rect 13872 3952 13878 3964
rect 14185 3961 14197 3995
rect 14231 3992 14243 3995
rect 15010 3992 15016 4004
rect 14231 3964 15016 3992
rect 14231 3961 14243 3964
rect 14185 3955 14243 3961
rect 15010 3952 15016 3964
rect 15068 3952 15074 4004
rect 14090 3924 14096 3936
rect 11624 3896 14096 3924
rect 14090 3884 14096 3896
rect 14148 3884 14154 3936
rect 14277 3927 14335 3933
rect 14277 3893 14289 3927
rect 14323 3924 14335 3927
rect 14642 3924 14648 3936
rect 14323 3896 14648 3924
rect 14323 3893 14335 3896
rect 14277 3887 14335 3893
rect 14642 3884 14648 3896
rect 14700 3884 14706 3936
rect 15286 3924 15292 3936
rect 15247 3896 15292 3924
rect 15286 3884 15292 3896
rect 15344 3884 15350 3936
rect 15562 3924 15568 3936
rect 15523 3896 15568 3924
rect 15562 3884 15568 3896
rect 15620 3884 15626 3936
rect 1104 3834 16008 3856
rect 1104 3782 2824 3834
rect 2876 3782 2888 3834
rect 2940 3782 2952 3834
rect 3004 3782 3016 3834
rect 3068 3782 3080 3834
rect 3132 3782 6572 3834
rect 6624 3782 6636 3834
rect 6688 3782 6700 3834
rect 6752 3782 6764 3834
rect 6816 3782 6828 3834
rect 6880 3782 10320 3834
rect 10372 3782 10384 3834
rect 10436 3782 10448 3834
rect 10500 3782 10512 3834
rect 10564 3782 10576 3834
rect 10628 3782 14068 3834
rect 14120 3782 14132 3834
rect 14184 3782 14196 3834
rect 14248 3782 14260 3834
rect 14312 3782 14324 3834
rect 14376 3782 16008 3834
rect 1104 3760 16008 3782
rect 1486 3720 1492 3732
rect 1447 3692 1492 3720
rect 1486 3680 1492 3692
rect 1544 3680 1550 3732
rect 2498 3680 2504 3732
rect 2556 3720 2562 3732
rect 3970 3720 3976 3732
rect 2556 3692 3976 3720
rect 2556 3680 2562 3692
rect 3970 3680 3976 3692
rect 4028 3680 4034 3732
rect 4062 3680 4068 3732
rect 4120 3720 4126 3732
rect 6273 3723 6331 3729
rect 6273 3720 6285 3723
rect 4120 3692 6285 3720
rect 4120 3680 4126 3692
rect 6273 3689 6285 3692
rect 6319 3689 6331 3723
rect 6273 3683 6331 3689
rect 6362 3680 6368 3732
rect 6420 3720 6426 3732
rect 6825 3723 6883 3729
rect 6825 3720 6837 3723
rect 6420 3692 6837 3720
rect 6420 3680 6426 3692
rect 6825 3689 6837 3692
rect 6871 3689 6883 3723
rect 6825 3683 6883 3689
rect 7098 3680 7104 3732
rect 7156 3720 7162 3732
rect 7837 3723 7895 3729
rect 7837 3720 7849 3723
rect 7156 3692 7849 3720
rect 7156 3680 7162 3692
rect 7837 3689 7849 3692
rect 7883 3689 7895 3723
rect 7837 3683 7895 3689
rect 8018 3680 8024 3732
rect 8076 3720 8082 3732
rect 8570 3720 8576 3732
rect 8076 3692 8576 3720
rect 8076 3680 8082 3692
rect 8570 3680 8576 3692
rect 8628 3680 8634 3732
rect 8938 3720 8944 3732
rect 8899 3692 8944 3720
rect 8938 3680 8944 3692
rect 8996 3680 9002 3732
rect 9030 3680 9036 3732
rect 9088 3720 9094 3732
rect 9953 3723 10011 3729
rect 9953 3720 9965 3723
rect 9088 3692 9965 3720
rect 9088 3680 9094 3692
rect 9953 3689 9965 3692
rect 9999 3689 10011 3723
rect 11054 3720 11060 3732
rect 11015 3692 11060 3720
rect 9953 3683 10011 3689
rect 11054 3680 11060 3692
rect 11112 3680 11118 3732
rect 11146 3680 11152 3732
rect 11204 3720 11210 3732
rect 12710 3720 12716 3732
rect 11204 3692 12716 3720
rect 11204 3680 11210 3692
rect 12710 3680 12716 3692
rect 12768 3680 12774 3732
rect 13538 3680 13544 3732
rect 13596 3720 13602 3732
rect 14458 3720 14464 3732
rect 13596 3692 14464 3720
rect 13596 3680 13602 3692
rect 14458 3680 14464 3692
rect 14516 3680 14522 3732
rect 14921 3723 14979 3729
rect 14921 3689 14933 3723
rect 14967 3689 14979 3723
rect 14921 3683 14979 3689
rect 3050 3612 3056 3664
rect 3108 3652 3114 3664
rect 3329 3655 3387 3661
rect 3329 3652 3341 3655
rect 3108 3624 3341 3652
rect 3108 3612 3114 3624
rect 3329 3621 3341 3624
rect 3375 3621 3387 3655
rect 3789 3655 3847 3661
rect 3789 3652 3801 3655
rect 3329 3615 3387 3621
rect 3528 3624 3801 3652
rect 2682 3544 2688 3596
rect 2740 3584 2746 3596
rect 2740 3556 3271 3584
rect 2740 3544 2746 3556
rect 1670 3516 1676 3528
rect 1631 3488 1676 3516
rect 1670 3476 1676 3488
rect 1728 3476 1734 3528
rect 2038 3516 2044 3528
rect 1999 3488 2044 3516
rect 2038 3476 2044 3488
rect 2096 3476 2102 3528
rect 2130 3476 2136 3528
rect 2188 3516 2194 3528
rect 2317 3519 2375 3525
rect 2317 3516 2329 3519
rect 2188 3488 2329 3516
rect 2188 3476 2194 3488
rect 2317 3485 2329 3488
rect 2363 3485 2375 3519
rect 2317 3479 2375 3485
rect 2593 3519 2651 3525
rect 2593 3485 2605 3519
rect 2639 3485 2651 3519
rect 2866 3516 2872 3528
rect 2827 3488 2872 3516
rect 2593 3479 2651 3485
rect 2608 3448 2636 3479
rect 2866 3476 2872 3488
rect 2924 3476 2930 3528
rect 3142 3516 3148 3528
rect 3103 3488 3148 3516
rect 3142 3476 3148 3488
rect 3200 3476 3206 3528
rect 3243 3448 3271 3556
rect 3528 3525 3556 3624
rect 3789 3621 3801 3624
rect 3835 3621 3847 3655
rect 3789 3615 3847 3621
rect 4264 3624 4660 3652
rect 3694 3544 3700 3596
rect 3752 3584 3758 3596
rect 4264 3593 4292 3624
rect 4249 3587 4307 3593
rect 4249 3584 4261 3587
rect 3752 3556 4261 3584
rect 3752 3544 3758 3556
rect 4249 3553 4261 3556
rect 4295 3553 4307 3587
rect 4249 3547 4307 3553
rect 4341 3587 4399 3593
rect 4341 3553 4353 3587
rect 4387 3584 4399 3587
rect 4522 3584 4528 3596
rect 4387 3556 4528 3584
rect 4387 3553 4399 3556
rect 4341 3547 4399 3553
rect 4522 3544 4528 3556
rect 4580 3544 4586 3596
rect 4632 3584 4660 3624
rect 5074 3612 5080 3664
rect 5132 3652 5138 3664
rect 5445 3655 5503 3661
rect 5445 3652 5457 3655
rect 5132 3624 5457 3652
rect 5132 3612 5138 3624
rect 5445 3621 5457 3624
rect 5491 3621 5503 3655
rect 9125 3655 9183 3661
rect 9125 3652 9137 3655
rect 5445 3615 5503 3621
rect 5828 3624 9137 3652
rect 5718 3584 5724 3596
rect 4632 3556 5724 3584
rect 5718 3544 5724 3556
rect 5776 3544 5782 3596
rect 3513 3519 3571 3525
rect 3513 3485 3525 3519
rect 3559 3485 3571 3519
rect 3513 3479 3571 3485
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3485 4031 3519
rect 4430 3516 4436 3528
rect 4391 3488 4436 3516
rect 3973 3479 4031 3485
rect 3988 3448 4016 3479
rect 4430 3476 4436 3488
rect 4488 3476 4494 3528
rect 5169 3519 5227 3525
rect 5169 3485 5181 3519
rect 5215 3516 5227 3519
rect 5350 3516 5356 3528
rect 5215 3488 5356 3516
rect 5215 3485 5227 3488
rect 5169 3479 5227 3485
rect 5350 3476 5356 3488
rect 5408 3476 5414 3528
rect 5828 3525 5856 3624
rect 9125 3621 9137 3624
rect 9171 3621 9183 3655
rect 10410 3652 10416 3664
rect 9125 3615 9183 3621
rect 9232 3624 10416 3652
rect 5997 3587 6055 3593
rect 5997 3553 6009 3587
rect 6043 3584 6055 3587
rect 6822 3584 6828 3596
rect 6043 3556 6828 3584
rect 6043 3553 6055 3556
rect 5997 3547 6055 3553
rect 6822 3544 6828 3556
rect 6880 3544 6886 3596
rect 7282 3584 7288 3596
rect 7243 3556 7288 3584
rect 7282 3544 7288 3556
rect 7340 3544 7346 3596
rect 7469 3587 7527 3593
rect 7469 3553 7481 3587
rect 7515 3553 7527 3587
rect 7469 3547 7527 3553
rect 5813 3519 5871 3525
rect 5813 3485 5825 3519
rect 5859 3485 5871 3519
rect 5813 3479 5871 3485
rect 6270 3476 6276 3528
rect 6328 3516 6334 3528
rect 6457 3519 6515 3525
rect 6328 3512 6408 3516
rect 6457 3512 6469 3519
rect 6328 3488 6469 3512
rect 6328 3476 6334 3488
rect 6380 3485 6469 3488
rect 6503 3485 6515 3519
rect 6380 3484 6515 3485
rect 6457 3479 6515 3484
rect 6549 3495 6607 3501
rect 6549 3461 6561 3495
rect 6595 3492 6607 3495
rect 6638 3492 6644 3528
rect 6595 3476 6644 3492
rect 6696 3476 6702 3528
rect 7193 3519 7251 3525
rect 7193 3485 7205 3519
rect 7239 3485 7251 3519
rect 7193 3479 7251 3485
rect 6595 3464 6675 3476
rect 6595 3461 6607 3464
rect 5442 3448 5448 3460
rect 2608 3420 3096 3448
rect 3243 3420 5448 3448
rect 1854 3380 1860 3392
rect 1815 3352 1860 3380
rect 1854 3340 1860 3352
rect 1912 3340 1918 3392
rect 1946 3340 1952 3392
rect 2004 3380 2010 3392
rect 2133 3383 2191 3389
rect 2133 3380 2145 3383
rect 2004 3352 2145 3380
rect 2004 3340 2010 3352
rect 2133 3349 2145 3352
rect 2179 3349 2191 3383
rect 2133 3343 2191 3349
rect 2222 3340 2228 3392
rect 2280 3380 2286 3392
rect 2409 3383 2467 3389
rect 2409 3380 2421 3383
rect 2280 3352 2421 3380
rect 2280 3340 2286 3352
rect 2409 3349 2421 3352
rect 2455 3349 2467 3383
rect 2409 3343 2467 3349
rect 2498 3340 2504 3392
rect 2556 3380 2562 3392
rect 2685 3383 2743 3389
rect 2685 3380 2697 3383
rect 2556 3352 2697 3380
rect 2556 3340 2562 3352
rect 2685 3349 2697 3352
rect 2731 3349 2743 3383
rect 2958 3380 2964 3392
rect 2919 3352 2964 3380
rect 2685 3343 2743 3349
rect 2958 3340 2964 3352
rect 3016 3340 3022 3392
rect 3068 3380 3096 3420
rect 5442 3408 5448 3420
rect 5500 3408 5506 3460
rect 5534 3408 5540 3460
rect 5592 3448 5598 3460
rect 5905 3451 5963 3457
rect 6549 3455 6607 3461
rect 5905 3448 5917 3451
rect 5592 3420 5917 3448
rect 5592 3408 5598 3420
rect 5905 3417 5917 3420
rect 5951 3417 5963 3451
rect 7208 3448 7236 3479
rect 7484 3460 7512 3547
rect 8018 3544 8024 3596
rect 8076 3584 8082 3596
rect 8076 3556 8340 3584
rect 8076 3544 8082 3556
rect 7929 3519 7987 3525
rect 7929 3485 7941 3519
rect 7975 3516 7987 3519
rect 8202 3516 8208 3528
rect 7975 3488 8208 3516
rect 7975 3485 7987 3488
rect 7929 3479 7987 3485
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 8312 3525 8340 3556
rect 8386 3544 8392 3596
rect 8444 3584 8450 3596
rect 8573 3587 8631 3593
rect 8573 3584 8585 3587
rect 8444 3556 8585 3584
rect 8444 3544 8450 3556
rect 8573 3553 8585 3556
rect 8619 3553 8631 3587
rect 9232 3584 9260 3624
rect 10410 3612 10416 3624
rect 10468 3612 10474 3664
rect 11330 3652 11336 3664
rect 10520 3624 11336 3652
rect 8573 3547 8631 3553
rect 8680 3556 9260 3584
rect 8297 3519 8355 3525
rect 8297 3485 8309 3519
rect 8343 3485 8355 3519
rect 8680 3516 8708 3556
rect 9490 3544 9496 3596
rect 9548 3584 9554 3596
rect 9585 3587 9643 3593
rect 9585 3584 9597 3587
rect 9548 3556 9597 3584
rect 9548 3544 9554 3556
rect 9585 3553 9597 3556
rect 9631 3553 9643 3587
rect 9585 3547 9643 3553
rect 9677 3587 9735 3593
rect 9677 3553 9689 3587
rect 9723 3553 9735 3587
rect 9677 3547 9735 3553
rect 8297 3479 8355 3485
rect 8404 3488 8708 3516
rect 7282 3448 7288 3460
rect 7208 3420 7288 3448
rect 5905 3411 5963 3417
rect 7282 3408 7288 3420
rect 7340 3408 7346 3460
rect 7466 3408 7472 3460
rect 7524 3408 7530 3460
rect 7742 3408 7748 3460
rect 7800 3448 7806 3460
rect 8113 3451 8171 3457
rect 8113 3448 8125 3451
rect 7800 3420 8125 3448
rect 7800 3408 7806 3420
rect 8113 3417 8125 3420
rect 8159 3417 8171 3451
rect 8113 3411 8171 3417
rect 4154 3380 4160 3392
rect 3068 3352 4160 3380
rect 4154 3340 4160 3352
rect 4212 3340 4218 3392
rect 4614 3340 4620 3392
rect 4672 3380 4678 3392
rect 4801 3383 4859 3389
rect 4801 3380 4813 3383
rect 4672 3352 4813 3380
rect 4672 3340 4678 3352
rect 4801 3349 4813 3352
rect 4847 3349 4859 3383
rect 4801 3343 4859 3349
rect 4985 3383 5043 3389
rect 4985 3349 4997 3383
rect 5031 3380 5043 3383
rect 5074 3380 5080 3392
rect 5031 3352 5080 3380
rect 5031 3349 5043 3352
rect 4985 3343 5043 3349
rect 5074 3340 5080 3352
rect 5132 3340 5138 3392
rect 5353 3383 5411 3389
rect 5353 3349 5365 3383
rect 5399 3380 5411 3383
rect 5810 3380 5816 3392
rect 5399 3352 5816 3380
rect 5399 3349 5411 3352
rect 5353 3343 5411 3349
rect 5810 3340 5816 3352
rect 5868 3340 5874 3392
rect 6362 3340 6368 3392
rect 6420 3380 6426 3392
rect 6733 3383 6791 3389
rect 6733 3380 6745 3383
rect 6420 3352 6745 3380
rect 6420 3340 6426 3352
rect 6733 3349 6745 3352
rect 6779 3349 6791 3383
rect 6733 3343 6791 3349
rect 6822 3340 6828 3392
rect 6880 3380 6886 3392
rect 8404 3380 8432 3488
rect 9214 3476 9220 3528
rect 9272 3516 9278 3528
rect 9692 3516 9720 3547
rect 10042 3544 10048 3596
rect 10100 3584 10106 3596
rect 10520 3593 10548 3624
rect 11330 3612 11336 3624
rect 11388 3612 11394 3664
rect 11422 3612 11428 3664
rect 11480 3652 11486 3664
rect 14936 3652 14964 3683
rect 11480 3624 12388 3652
rect 11480 3612 11486 3624
rect 10505 3587 10563 3593
rect 10505 3584 10517 3587
rect 10100 3556 10517 3584
rect 10100 3544 10106 3556
rect 10505 3553 10517 3556
rect 10551 3553 10563 3587
rect 10505 3547 10563 3553
rect 10594 3544 10600 3596
rect 10652 3584 10658 3596
rect 10652 3556 10916 3584
rect 10652 3544 10658 3556
rect 9272 3488 9720 3516
rect 10321 3519 10379 3525
rect 9272 3476 9278 3488
rect 10321 3485 10333 3519
rect 10367 3516 10379 3519
rect 10778 3516 10784 3528
rect 10367 3488 10784 3516
rect 10367 3485 10379 3488
rect 10321 3479 10379 3485
rect 10778 3476 10784 3488
rect 10836 3476 10842 3528
rect 10888 3516 10916 3556
rect 10962 3544 10968 3596
rect 11020 3584 11026 3596
rect 11241 3587 11299 3593
rect 11241 3584 11253 3587
rect 11020 3556 11253 3584
rect 11020 3544 11026 3556
rect 11241 3553 11253 3556
rect 11287 3553 11299 3587
rect 11241 3547 11299 3553
rect 11974 3544 11980 3596
rect 12032 3584 12038 3596
rect 12360 3593 12388 3624
rect 13464 3624 14964 3652
rect 12069 3587 12127 3593
rect 12069 3584 12081 3587
rect 12032 3556 12081 3584
rect 12032 3544 12038 3556
rect 12069 3553 12081 3556
rect 12115 3553 12127 3587
rect 12069 3547 12127 3553
rect 12345 3587 12403 3593
rect 12345 3553 12357 3587
rect 12391 3553 12403 3587
rect 12345 3547 12403 3553
rect 12437 3587 12495 3593
rect 12437 3553 12449 3587
rect 12483 3584 12495 3587
rect 12618 3584 12624 3596
rect 12483 3556 12624 3584
rect 12483 3553 12495 3556
rect 12437 3547 12495 3553
rect 12618 3544 12624 3556
rect 12676 3544 12682 3596
rect 12713 3587 12771 3593
rect 12713 3553 12725 3587
rect 12759 3553 12771 3587
rect 12713 3547 12771 3553
rect 11882 3516 11888 3528
rect 10888 3488 11888 3516
rect 11882 3476 11888 3488
rect 11940 3476 11946 3528
rect 10226 3448 10232 3460
rect 8496 3420 10232 3448
rect 8496 3389 8524 3420
rect 10226 3408 10232 3420
rect 10284 3448 10290 3460
rect 10284 3420 11928 3448
rect 10284 3408 10290 3420
rect 11900 3392 11928 3420
rect 11974 3408 11980 3460
rect 12032 3448 12038 3460
rect 12636 3448 12664 3544
rect 12728 3516 12756 3547
rect 13078 3544 13084 3596
rect 13136 3584 13142 3596
rect 13464 3584 13492 3624
rect 13906 3584 13912 3596
rect 13136 3556 13492 3584
rect 13556 3556 13912 3584
rect 13136 3544 13142 3556
rect 13170 3516 13176 3528
rect 12728 3488 13176 3516
rect 13170 3476 13176 3488
rect 13228 3476 13234 3528
rect 13556 3525 13584 3556
rect 13906 3544 13912 3556
rect 13964 3544 13970 3596
rect 14277 3587 14335 3593
rect 14277 3553 14289 3587
rect 14323 3584 14335 3587
rect 14550 3584 14556 3596
rect 14323 3556 14556 3584
rect 14323 3553 14335 3556
rect 14277 3547 14335 3553
rect 14550 3544 14556 3556
rect 14608 3544 14614 3596
rect 14918 3544 14924 3596
rect 14976 3584 14982 3596
rect 15381 3587 15439 3593
rect 15381 3584 15393 3587
rect 14976 3556 15393 3584
rect 14976 3544 14982 3556
rect 15381 3553 15393 3556
rect 15427 3553 15439 3587
rect 15381 3547 15439 3553
rect 15470 3544 15476 3596
rect 15528 3584 15534 3596
rect 15528 3556 15573 3584
rect 15528 3544 15534 3556
rect 13541 3519 13599 3525
rect 13541 3485 13553 3519
rect 13587 3485 13599 3519
rect 13633 3519 13691 3525
rect 13633 3504 13645 3519
rect 13679 3504 13691 3519
rect 13541 3479 13599 3485
rect 12032 3420 12664 3448
rect 12032 3408 12038 3420
rect 13078 3408 13084 3460
rect 13136 3448 13142 3460
rect 13446 3448 13452 3460
rect 13136 3420 13452 3448
rect 13136 3408 13142 3420
rect 13446 3408 13452 3420
rect 13504 3408 13510 3460
rect 13630 3452 13636 3504
rect 13688 3452 13694 3504
rect 13998 3476 14004 3528
rect 14056 3516 14062 3528
rect 14826 3516 14832 3528
rect 14056 3488 14832 3516
rect 14056 3476 14062 3488
rect 14826 3476 14832 3488
rect 14884 3476 14890 3528
rect 15286 3516 15292 3528
rect 15247 3488 15292 3516
rect 15286 3476 15292 3488
rect 15344 3476 15350 3528
rect 13832 3420 15332 3448
rect 6880 3352 8432 3380
rect 8481 3383 8539 3389
rect 6880 3340 6886 3352
rect 8481 3349 8493 3383
rect 8527 3349 8539 3383
rect 8481 3343 8539 3349
rect 8662 3340 8668 3392
rect 8720 3380 8726 3392
rect 9122 3380 9128 3392
rect 8720 3352 9128 3380
rect 8720 3340 8726 3352
rect 9122 3340 9128 3352
rect 9180 3340 9186 3392
rect 9490 3380 9496 3392
rect 9451 3352 9496 3380
rect 9490 3340 9496 3352
rect 9548 3340 9554 3392
rect 10410 3340 10416 3392
rect 10468 3380 10474 3392
rect 10778 3380 10784 3392
rect 10468 3352 10513 3380
rect 10739 3352 10784 3380
rect 10468 3340 10474 3352
rect 10778 3340 10784 3352
rect 10836 3340 10842 3392
rect 11882 3340 11888 3392
rect 11940 3340 11946 3392
rect 12618 3340 12624 3392
rect 12676 3380 12682 3392
rect 13832 3389 13860 3420
rect 15304 3392 15332 3420
rect 13357 3383 13415 3389
rect 13357 3380 13369 3383
rect 12676 3352 13369 3380
rect 12676 3340 12682 3352
rect 13357 3349 13369 3352
rect 13403 3349 13415 3383
rect 13357 3343 13415 3349
rect 13817 3383 13875 3389
rect 13817 3349 13829 3383
rect 13863 3349 13875 3383
rect 14366 3380 14372 3392
rect 14327 3352 14372 3380
rect 13817 3343 13875 3349
rect 14366 3340 14372 3352
rect 14424 3340 14430 3392
rect 14458 3340 14464 3392
rect 14516 3380 14522 3392
rect 14826 3380 14832 3392
rect 14516 3352 14561 3380
rect 14787 3352 14832 3380
rect 14516 3340 14522 3352
rect 14826 3340 14832 3352
rect 14884 3340 14890 3392
rect 15286 3340 15292 3392
rect 15344 3340 15350 3392
rect 1104 3290 16008 3312
rect 1104 3238 4698 3290
rect 4750 3238 4762 3290
rect 4814 3238 4826 3290
rect 4878 3238 4890 3290
rect 4942 3238 4954 3290
rect 5006 3238 8446 3290
rect 8498 3238 8510 3290
rect 8562 3238 8574 3290
rect 8626 3238 8638 3290
rect 8690 3238 8702 3290
rect 8754 3238 12194 3290
rect 12246 3238 12258 3290
rect 12310 3238 12322 3290
rect 12374 3238 12386 3290
rect 12438 3238 12450 3290
rect 12502 3238 16008 3290
rect 1104 3216 16008 3238
rect 3789 3179 3847 3185
rect 3789 3145 3801 3179
rect 3835 3176 3847 3179
rect 3878 3176 3884 3188
rect 3835 3148 3884 3176
rect 3835 3145 3847 3148
rect 3789 3139 3847 3145
rect 3878 3136 3884 3148
rect 3936 3136 3942 3188
rect 3970 3136 3976 3188
rect 4028 3176 4034 3188
rect 4028 3148 4375 3176
rect 4028 3136 4034 3148
rect 2593 3111 2651 3117
rect 2593 3077 2605 3111
rect 2639 3108 2651 3111
rect 4157 3111 4215 3117
rect 2639 3080 4108 3108
rect 2639 3077 2651 3080
rect 2593 3071 2651 3077
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3040 1731 3043
rect 1946 3040 1952 3052
rect 1719 3012 1952 3040
rect 1719 3009 1731 3012
rect 1673 3003 1731 3009
rect 1946 3000 1952 3012
rect 2004 3000 2010 3052
rect 2041 3043 2099 3049
rect 2041 3009 2053 3043
rect 2087 3009 2099 3043
rect 2041 3003 2099 3009
rect 2409 3043 2467 3049
rect 2409 3009 2421 3043
rect 2455 3040 2467 3043
rect 2958 3040 2964 3052
rect 2455 3012 2774 3040
rect 2919 3012 2964 3040
rect 2455 3009 2467 3012
rect 2409 3003 2467 3009
rect 2056 2972 2084 3003
rect 2590 2972 2596 2984
rect 2056 2944 2596 2972
rect 2590 2932 2596 2944
rect 2648 2932 2654 2984
rect 2746 2972 2774 3012
rect 2958 3000 2964 3012
rect 3016 3000 3022 3052
rect 3329 3043 3387 3049
rect 3329 3009 3341 3043
rect 3375 3009 3387 3043
rect 3329 3003 3387 3009
rect 3690 3043 3748 3049
rect 3690 3009 3702 3043
rect 3736 3040 3748 3043
rect 3970 3040 3976 3052
rect 3736 3012 3976 3040
rect 3736 3009 3748 3012
rect 3690 3003 3748 3009
rect 3234 2972 3240 2984
rect 2746 2944 3240 2972
rect 3234 2932 3240 2944
rect 3292 2932 3298 2984
rect 3344 2972 3372 3003
rect 3970 3000 3976 3012
rect 4028 3000 4034 3052
rect 4080 3040 4108 3080
rect 4157 3077 4169 3111
rect 4203 3108 4215 3111
rect 4246 3108 4252 3120
rect 4203 3080 4252 3108
rect 4203 3077 4215 3080
rect 4157 3071 4215 3077
rect 4246 3068 4252 3080
rect 4304 3068 4310 3120
rect 4347 3108 4375 3148
rect 4614 3136 4620 3188
rect 4672 3176 4678 3188
rect 4893 3179 4951 3185
rect 4893 3176 4905 3179
rect 4672 3148 4905 3176
rect 4672 3136 4678 3148
rect 4893 3145 4905 3148
rect 4939 3145 4951 3179
rect 4893 3139 4951 3145
rect 4985 3179 5043 3185
rect 4985 3145 4997 3179
rect 5031 3176 5043 3179
rect 5445 3179 5503 3185
rect 5445 3176 5457 3179
rect 5031 3148 5457 3176
rect 5031 3145 5043 3148
rect 4985 3139 5043 3145
rect 5445 3145 5457 3148
rect 5491 3145 5503 3179
rect 5902 3176 5908 3188
rect 5863 3148 5908 3176
rect 5445 3139 5503 3145
rect 5902 3136 5908 3148
rect 5960 3136 5966 3188
rect 6454 3136 6460 3188
rect 6512 3176 6518 3188
rect 6512 3148 7512 3176
rect 6512 3136 6518 3148
rect 5258 3108 5264 3120
rect 4347 3080 5264 3108
rect 5258 3068 5264 3080
rect 5316 3068 5322 3120
rect 5813 3111 5871 3117
rect 5813 3077 5825 3111
rect 5859 3108 5871 3111
rect 6086 3108 6092 3120
rect 5859 3080 6092 3108
rect 5859 3077 5871 3080
rect 5813 3071 5871 3077
rect 6086 3068 6092 3080
rect 6144 3068 6150 3120
rect 6546 3068 6552 3120
rect 6604 3068 6610 3120
rect 7484 3108 7512 3148
rect 7558 3136 7564 3188
rect 7616 3176 7622 3188
rect 7653 3179 7711 3185
rect 7653 3176 7665 3179
rect 7616 3148 7665 3176
rect 7616 3136 7622 3148
rect 7653 3145 7665 3148
rect 7699 3145 7711 3179
rect 7653 3139 7711 3145
rect 7760 3148 9168 3176
rect 7760 3108 7788 3148
rect 6932 3080 7429 3108
rect 7484 3080 7788 3108
rect 8021 3111 8079 3117
rect 6454 3040 6460 3052
rect 4080 3012 5773 3040
rect 3344 2944 4108 2972
rect 3145 2907 3203 2913
rect 3145 2873 3157 2907
rect 3191 2904 3203 2907
rect 3694 2904 3700 2916
rect 3191 2876 3700 2904
rect 3191 2873 3203 2876
rect 3145 2867 3203 2873
rect 3694 2864 3700 2876
rect 3752 2864 3758 2916
rect 4080 2904 4108 2944
rect 4154 2932 4160 2984
rect 4212 2972 4218 2984
rect 4249 2975 4307 2981
rect 4249 2972 4261 2975
rect 4212 2944 4261 2972
rect 4212 2932 4218 2944
rect 4249 2941 4261 2944
rect 4295 2941 4307 2975
rect 4249 2935 4307 2941
rect 4433 2975 4491 2981
rect 4433 2941 4445 2975
rect 4479 2972 4491 2975
rect 4522 2972 4528 2984
rect 4479 2944 4528 2972
rect 4479 2941 4491 2944
rect 4433 2935 4491 2941
rect 4522 2932 4528 2944
rect 4580 2932 4586 2984
rect 4801 2975 4859 2981
rect 4801 2941 4813 2975
rect 4847 2972 4859 2975
rect 5442 2972 5448 2984
rect 4847 2944 5448 2972
rect 4847 2941 4859 2944
rect 4801 2935 4859 2941
rect 5442 2932 5448 2944
rect 5500 2932 5506 2984
rect 5258 2904 5264 2916
rect 4080 2876 5264 2904
rect 5258 2864 5264 2876
rect 5316 2864 5322 2916
rect 5353 2907 5411 2913
rect 5353 2873 5365 2907
rect 5399 2904 5411 2907
rect 5534 2904 5540 2916
rect 5399 2876 5540 2904
rect 5399 2873 5411 2876
rect 5353 2867 5411 2873
rect 5534 2864 5540 2876
rect 5592 2864 5598 2916
rect 5745 2904 5773 3012
rect 6104 3012 6460 3040
rect 5810 2932 5816 2984
rect 5868 2972 5874 2984
rect 6104 2981 6132 3012
rect 6454 3000 6460 3012
rect 6512 3000 6518 3052
rect 6089 2975 6147 2981
rect 6089 2972 6101 2975
rect 5868 2944 6101 2972
rect 5868 2932 5874 2944
rect 6089 2941 6101 2944
rect 6135 2941 6147 2975
rect 6564 2972 6592 3068
rect 6634 3043 6692 3049
rect 6634 3009 6646 3043
rect 6680 3040 6692 3043
rect 6932 3040 6960 3080
rect 6680 3012 6960 3040
rect 6680 3009 6692 3012
rect 6634 3003 6692 3009
rect 7006 3000 7012 3052
rect 7064 3040 7070 3052
rect 7101 3043 7159 3049
rect 7101 3040 7113 3043
rect 7064 3012 7113 3040
rect 7064 3000 7070 3012
rect 7101 3009 7113 3012
rect 7147 3009 7159 3043
rect 7101 3003 7159 3009
rect 7193 3043 7251 3049
rect 7193 3009 7205 3043
rect 7239 3040 7251 3043
rect 7282 3040 7288 3052
rect 7239 3012 7288 3040
rect 7239 3009 7251 3012
rect 7193 3003 7251 3009
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 7401 3040 7429 3080
rect 8021 3077 8033 3111
rect 8067 3108 8079 3111
rect 8202 3108 8208 3120
rect 8067 3080 8208 3108
rect 8067 3077 8079 3080
rect 8021 3071 8079 3077
rect 8202 3068 8208 3080
rect 8260 3068 8266 3120
rect 7834 3040 7840 3052
rect 7401 3012 7840 3040
rect 7834 3000 7840 3012
rect 7892 3000 7898 3052
rect 7926 3000 7932 3052
rect 7984 3040 7990 3052
rect 8110 3040 8116 3052
rect 7984 3012 8116 3040
rect 7984 3000 7990 3012
rect 8110 3000 8116 3012
rect 8168 3000 8174 3052
rect 8386 3000 8392 3052
rect 8444 3040 8450 3052
rect 8481 3043 8539 3049
rect 8481 3040 8493 3043
rect 8444 3012 8493 3040
rect 8444 3000 8450 3012
rect 8481 3009 8493 3012
rect 8527 3040 8539 3043
rect 8846 3040 8852 3052
rect 8527 3012 8852 3040
rect 8527 3009 8539 3012
rect 8481 3003 8539 3009
rect 8846 3000 8852 3012
rect 8904 3000 8910 3052
rect 7377 2975 7435 2981
rect 6564 2944 6776 2972
rect 6089 2935 6147 2941
rect 6748 2913 6776 2944
rect 7377 2941 7389 2975
rect 7423 2941 7435 2975
rect 8205 2975 8263 2981
rect 8205 2972 8217 2975
rect 7377 2935 7435 2941
rect 7760 2944 8217 2972
rect 6733 2907 6791 2913
rect 5745 2876 6684 2904
rect 1486 2836 1492 2848
rect 1447 2808 1492 2836
rect 1486 2796 1492 2808
rect 1544 2796 1550 2848
rect 1762 2796 1768 2848
rect 1820 2836 1826 2848
rect 1857 2839 1915 2845
rect 1857 2836 1869 2839
rect 1820 2808 1869 2836
rect 1820 2796 1826 2808
rect 1857 2805 1869 2808
rect 1903 2805 1915 2839
rect 1857 2799 1915 2805
rect 2038 2796 2044 2848
rect 2096 2836 2102 2848
rect 2225 2839 2283 2845
rect 2225 2836 2237 2839
rect 2096 2808 2237 2836
rect 2096 2796 2102 2808
rect 2225 2805 2237 2808
rect 2271 2805 2283 2839
rect 2225 2799 2283 2805
rect 2682 2796 2688 2848
rect 2740 2836 2746 2848
rect 2777 2839 2835 2845
rect 2777 2836 2789 2839
rect 2740 2808 2789 2836
rect 2740 2796 2746 2808
rect 2777 2805 2789 2808
rect 2823 2805 2835 2839
rect 2777 2799 2835 2805
rect 3513 2839 3571 2845
rect 3513 2805 3525 2839
rect 3559 2836 3571 2839
rect 4246 2836 4252 2848
rect 3559 2808 4252 2836
rect 3559 2805 3571 2808
rect 3513 2799 3571 2805
rect 4246 2796 4252 2808
rect 4304 2796 4310 2848
rect 6178 2796 6184 2848
rect 6236 2836 6242 2848
rect 6457 2839 6515 2845
rect 6457 2836 6469 2839
rect 6236 2808 6469 2836
rect 6236 2796 6242 2808
rect 6457 2805 6469 2808
rect 6503 2805 6515 2839
rect 6656 2836 6684 2876
rect 6733 2873 6745 2907
rect 6779 2873 6791 2907
rect 6733 2867 6791 2873
rect 6822 2864 6828 2916
rect 6880 2904 6886 2916
rect 7392 2904 7420 2935
rect 7760 2904 7788 2944
rect 8205 2941 8217 2944
rect 8251 2941 8263 2975
rect 8754 2972 8760 2984
rect 8715 2944 8760 2972
rect 8205 2935 8263 2941
rect 8754 2932 8760 2944
rect 8812 2932 8818 2984
rect 9140 2972 9168 3148
rect 9490 3136 9496 3188
rect 9548 3176 9554 3188
rect 10045 3179 10103 3185
rect 10045 3176 10057 3179
rect 9548 3148 10057 3176
rect 9548 3136 9554 3148
rect 10045 3145 10057 3148
rect 10091 3145 10103 3179
rect 10045 3139 10103 3145
rect 10413 3179 10471 3185
rect 10413 3145 10425 3179
rect 10459 3176 10471 3179
rect 10778 3176 10784 3188
rect 10459 3148 10784 3176
rect 10459 3145 10471 3148
rect 10413 3139 10471 3145
rect 10778 3136 10784 3148
rect 10836 3136 10842 3188
rect 10962 3176 10968 3188
rect 10923 3148 10968 3176
rect 10962 3136 10968 3148
rect 11020 3136 11026 3188
rect 11790 3136 11796 3188
rect 11848 3176 11854 3188
rect 14734 3176 14740 3188
rect 11848 3148 14740 3176
rect 11848 3136 11854 3148
rect 14734 3136 14740 3148
rect 14792 3136 14798 3188
rect 10686 3108 10692 3120
rect 9968 3080 10692 3108
rect 9214 3000 9220 3052
rect 9272 3040 9278 3052
rect 9968 3049 9996 3080
rect 10686 3068 10692 3080
rect 10744 3068 10750 3120
rect 10870 3068 10876 3120
rect 10928 3108 10934 3120
rect 10928 3080 11560 3108
rect 10928 3068 10934 3080
rect 9493 3043 9551 3049
rect 9493 3040 9505 3043
rect 9272 3012 9505 3040
rect 9272 3000 9278 3012
rect 9493 3009 9505 3012
rect 9539 3009 9551 3043
rect 9493 3003 9551 3009
rect 9953 3043 10011 3049
rect 9953 3009 9965 3043
rect 9999 3009 10011 3043
rect 9953 3003 10011 3009
rect 10042 3000 10048 3052
rect 10100 3040 10106 3052
rect 11532 3049 11560 3080
rect 12526 3068 12532 3120
rect 12584 3108 12590 3120
rect 15381 3111 15439 3117
rect 15381 3108 15393 3111
rect 12584 3080 15393 3108
rect 12584 3068 12590 3080
rect 15381 3077 15393 3080
rect 15427 3077 15439 3111
rect 15381 3071 15439 3077
rect 11057 3043 11115 3049
rect 11057 3040 11069 3043
rect 10100 3012 11069 3040
rect 10100 3000 10106 3012
rect 11057 3009 11069 3012
rect 11103 3009 11115 3043
rect 11057 3003 11115 3009
rect 11517 3043 11575 3049
rect 11517 3009 11529 3043
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 10502 2972 10508 2984
rect 9140 2944 10364 2972
rect 10463 2944 10508 2972
rect 6880 2876 7788 2904
rect 6880 2864 6886 2876
rect 9674 2864 9680 2916
rect 9732 2904 9738 2916
rect 10336 2904 10364 2944
rect 10502 2932 10508 2944
rect 10560 2932 10566 2984
rect 10597 2975 10655 2981
rect 10597 2941 10609 2975
rect 10643 2941 10655 2975
rect 10597 2935 10655 2941
rect 10612 2904 10640 2935
rect 9732 2876 9777 2904
rect 10336 2876 10640 2904
rect 11072 2904 11100 3003
rect 11698 3000 11704 3052
rect 11756 3040 11762 3052
rect 11756 3012 12204 3040
rect 11756 3000 11762 3012
rect 11146 2932 11152 2984
rect 11204 2972 11210 2984
rect 11793 2975 11851 2981
rect 11793 2972 11805 2975
rect 11204 2944 11805 2972
rect 11204 2932 11210 2944
rect 11793 2941 11805 2944
rect 11839 2941 11851 2975
rect 12176 2972 12204 3012
rect 12250 3000 12256 3052
rect 12308 3040 12314 3052
rect 12437 3043 12495 3049
rect 12437 3040 12449 3043
rect 12308 3012 12449 3040
rect 12308 3000 12314 3012
rect 12437 3009 12449 3012
rect 12483 3009 12495 3043
rect 12437 3003 12495 3009
rect 12713 3043 12771 3049
rect 12713 3009 12725 3043
rect 12759 3040 12771 3043
rect 12894 3040 12900 3052
rect 12759 3012 12900 3040
rect 12759 3009 12771 3012
rect 12713 3003 12771 3009
rect 12894 3000 12900 3012
rect 12952 3000 12958 3052
rect 12986 3000 12992 3052
rect 13044 3040 13050 3052
rect 13633 3043 13691 3049
rect 13044 3012 13576 3040
rect 13044 3000 13050 3012
rect 13170 2972 13176 2984
rect 12176 2944 13176 2972
rect 11793 2935 11851 2941
rect 13170 2932 13176 2944
rect 13228 2932 13234 2984
rect 13357 2975 13415 2981
rect 13357 2941 13369 2975
rect 13403 2941 13415 2975
rect 13548 2972 13576 3012
rect 13633 3009 13645 3043
rect 13679 3040 13691 3043
rect 13814 3040 13820 3052
rect 13679 3012 13820 3040
rect 13679 3009 13691 3012
rect 13633 3003 13691 3009
rect 13814 3000 13820 3012
rect 13872 3000 13878 3052
rect 14090 3000 14096 3052
rect 14148 3040 14154 3052
rect 14645 3043 14703 3049
rect 14645 3040 14657 3043
rect 14148 3012 14657 3040
rect 14148 3000 14154 3012
rect 14645 3009 14657 3012
rect 14691 3009 14703 3043
rect 14645 3003 14703 3009
rect 14737 3043 14795 3049
rect 14737 3009 14749 3043
rect 14783 3040 14795 3043
rect 14918 3040 14924 3052
rect 14783 3012 14924 3040
rect 14783 3009 14795 3012
rect 14737 3003 14795 3009
rect 14918 3000 14924 3012
rect 14976 3000 14982 3052
rect 15105 3043 15163 3049
rect 15105 3009 15117 3043
rect 15151 3040 15163 3043
rect 15194 3040 15200 3052
rect 15151 3012 15200 3040
rect 15151 3009 15163 3012
rect 15105 3003 15163 3009
rect 15194 3000 15200 3012
rect 15252 3000 15258 3052
rect 14829 2975 14887 2981
rect 13548 2944 14320 2972
rect 13357 2935 13415 2941
rect 11072 2876 12434 2904
rect 9732 2864 9738 2876
rect 8202 2836 8208 2848
rect 6656 2808 8208 2836
rect 6457 2799 6515 2805
rect 8202 2796 8208 2808
rect 8260 2796 8266 2848
rect 8294 2796 8300 2848
rect 8352 2836 8358 2848
rect 9769 2839 9827 2845
rect 9769 2836 9781 2839
rect 8352 2808 9781 2836
rect 8352 2796 8358 2808
rect 9769 2805 9781 2808
rect 9815 2805 9827 2839
rect 10612 2836 10640 2876
rect 11241 2839 11299 2845
rect 11241 2836 11253 2839
rect 10612 2808 11253 2836
rect 9769 2799 9827 2805
rect 11241 2805 11253 2808
rect 11287 2836 11299 2839
rect 11330 2836 11336 2848
rect 11287 2808 11336 2836
rect 11287 2805 11299 2808
rect 11241 2799 11299 2805
rect 11330 2796 11336 2808
rect 11388 2796 11394 2848
rect 11698 2796 11704 2848
rect 11756 2836 11762 2848
rect 12250 2836 12256 2848
rect 11756 2808 12256 2836
rect 11756 2796 11762 2808
rect 12250 2796 12256 2808
rect 12308 2796 12314 2848
rect 12406 2836 12434 2876
rect 12526 2864 12532 2916
rect 12584 2904 12590 2916
rect 12802 2904 12808 2916
rect 12584 2876 12808 2904
rect 12584 2864 12590 2876
rect 12802 2864 12808 2876
rect 12860 2904 12866 2916
rect 13372 2904 13400 2935
rect 12860 2876 13400 2904
rect 12860 2864 12866 2876
rect 13446 2864 13452 2916
rect 13504 2904 13510 2916
rect 14292 2913 14320 2944
rect 14829 2941 14841 2975
rect 14875 2972 14887 2975
rect 15470 2972 15476 2984
rect 14875 2944 15476 2972
rect 14875 2941 14887 2944
rect 14829 2935 14887 2941
rect 15470 2932 15476 2944
rect 15528 2932 15534 2984
rect 14277 2907 14335 2913
rect 13504 2876 13860 2904
rect 13504 2864 13510 2876
rect 13722 2836 13728 2848
rect 12406 2808 13728 2836
rect 13722 2796 13728 2808
rect 13780 2796 13786 2848
rect 13832 2836 13860 2876
rect 14277 2873 14289 2907
rect 14323 2873 14335 2907
rect 14277 2867 14335 2873
rect 15654 2836 15660 2848
rect 13832 2808 15660 2836
rect 15654 2796 15660 2808
rect 15712 2796 15718 2848
rect 1104 2746 16008 2768
rect 1104 2694 2824 2746
rect 2876 2694 2888 2746
rect 2940 2694 2952 2746
rect 3004 2694 3016 2746
rect 3068 2694 3080 2746
rect 3132 2694 6572 2746
rect 6624 2694 6636 2746
rect 6688 2694 6700 2746
rect 6752 2694 6764 2746
rect 6816 2694 6828 2746
rect 6880 2694 10320 2746
rect 10372 2694 10384 2746
rect 10436 2694 10448 2746
rect 10500 2694 10512 2746
rect 10564 2694 10576 2746
rect 10628 2694 14068 2746
rect 14120 2694 14132 2746
rect 14184 2694 14196 2746
rect 14248 2694 14260 2746
rect 14312 2694 14324 2746
rect 14376 2694 16008 2746
rect 1104 2672 16008 2694
rect 2317 2635 2375 2641
rect 2317 2601 2329 2635
rect 2363 2632 2375 2635
rect 3418 2632 3424 2644
rect 2363 2604 3424 2632
rect 2363 2601 2375 2604
rect 2317 2595 2375 2601
rect 3418 2592 3424 2604
rect 3476 2592 3482 2644
rect 3786 2592 3792 2644
rect 3844 2632 3850 2644
rect 4525 2635 4583 2641
rect 4525 2632 4537 2635
rect 3844 2604 4537 2632
rect 3844 2592 3850 2604
rect 4525 2601 4537 2604
rect 4571 2601 4583 2635
rect 4525 2595 4583 2601
rect 5994 2592 6000 2644
rect 6052 2632 6058 2644
rect 6549 2635 6607 2641
rect 6549 2632 6561 2635
rect 6052 2604 6561 2632
rect 6052 2592 6058 2604
rect 6549 2601 6561 2604
rect 6595 2632 6607 2635
rect 7190 2632 7196 2644
rect 6595 2604 7196 2632
rect 6595 2601 6607 2604
rect 6549 2595 6607 2601
rect 7190 2592 7196 2604
rect 7248 2592 7254 2644
rect 7834 2592 7840 2644
rect 7892 2632 7898 2644
rect 8294 2632 8300 2644
rect 7892 2604 8300 2632
rect 7892 2592 7898 2604
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 9309 2635 9367 2641
rect 9309 2601 9321 2635
rect 9355 2632 9367 2635
rect 9766 2632 9772 2644
rect 9355 2604 9772 2632
rect 9355 2601 9367 2604
rect 9309 2595 9367 2601
rect 9766 2592 9772 2604
rect 9824 2592 9830 2644
rect 12618 2632 12624 2644
rect 9876 2604 12624 2632
rect 1949 2567 2007 2573
rect 1949 2533 1961 2567
rect 1995 2564 2007 2567
rect 2590 2564 2596 2576
rect 1995 2536 2596 2564
rect 1995 2533 2007 2536
rect 1949 2527 2007 2533
rect 2590 2524 2596 2536
rect 2648 2524 2654 2576
rect 2685 2567 2743 2573
rect 2685 2533 2697 2567
rect 2731 2564 2743 2567
rect 3970 2564 3976 2576
rect 2731 2536 3976 2564
rect 2731 2533 2743 2536
rect 2685 2527 2743 2533
rect 3970 2524 3976 2536
rect 4028 2524 4034 2576
rect 4062 2524 4068 2576
rect 4120 2524 4126 2576
rect 4154 2524 4160 2576
rect 4212 2564 4218 2576
rect 4249 2567 4307 2573
rect 4249 2564 4261 2567
rect 4212 2536 4261 2564
rect 4212 2524 4218 2536
rect 4249 2533 4261 2536
rect 4295 2533 4307 2567
rect 4249 2527 4307 2533
rect 4706 2524 4712 2576
rect 4764 2524 4770 2576
rect 5626 2524 5632 2576
rect 5684 2564 5690 2576
rect 6454 2564 6460 2576
rect 5684 2536 6460 2564
rect 5684 2524 5690 2536
rect 6454 2524 6460 2536
rect 6512 2564 6518 2576
rect 7377 2567 7435 2573
rect 7377 2564 7389 2567
rect 6512 2536 7389 2564
rect 6512 2524 6518 2536
rect 7377 2533 7389 2536
rect 7423 2533 7435 2567
rect 7377 2527 7435 2533
rect 7466 2524 7472 2576
rect 7524 2564 7530 2576
rect 8113 2567 8171 2573
rect 8113 2564 8125 2567
rect 7524 2536 8125 2564
rect 7524 2524 7530 2536
rect 8113 2533 8125 2536
rect 8159 2533 8171 2567
rect 8113 2527 8171 2533
rect 8202 2524 8208 2576
rect 8260 2564 8266 2576
rect 8662 2564 8668 2576
rect 8260 2536 8668 2564
rect 8260 2524 8266 2536
rect 8662 2524 8668 2536
rect 8720 2524 8726 2576
rect 3326 2496 3332 2508
rect 1780 2468 3332 2496
rect 1780 2437 1808 2468
rect 3326 2456 3332 2468
rect 3384 2456 3390 2508
rect 4080 2496 4108 2524
rect 3528 2468 4108 2496
rect 4724 2496 4752 2524
rect 5077 2499 5135 2505
rect 5077 2496 5089 2499
rect 4724 2468 5089 2496
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 2133 2431 2191 2437
rect 2133 2397 2145 2431
rect 2179 2428 2191 2431
rect 2222 2428 2228 2440
rect 2179 2400 2228 2428
rect 2179 2397 2191 2400
rect 2133 2391 2191 2397
rect 2222 2388 2228 2400
rect 2280 2388 2286 2440
rect 2498 2428 2504 2440
rect 2459 2400 2504 2428
rect 2498 2388 2504 2400
rect 2556 2388 2562 2440
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2428 2927 2431
rect 2958 2428 2964 2440
rect 2915 2400 2964 2428
rect 2915 2397 2927 2400
rect 2869 2391 2927 2397
rect 2958 2388 2964 2400
rect 3016 2388 3022 2440
rect 3237 2431 3295 2437
rect 3237 2397 3249 2431
rect 3283 2428 3295 2431
rect 3528 2428 3556 2468
rect 5077 2465 5089 2468
rect 5123 2465 5135 2499
rect 5077 2459 5135 2465
rect 5258 2456 5264 2508
rect 5316 2496 5322 2508
rect 9876 2496 9904 2604
rect 12618 2592 12624 2604
rect 12676 2592 12682 2644
rect 13722 2632 13728 2644
rect 13096 2604 13728 2632
rect 9950 2524 9956 2576
rect 10008 2564 10014 2576
rect 10594 2564 10600 2576
rect 10008 2536 10600 2564
rect 10008 2524 10014 2536
rect 10594 2524 10600 2536
rect 10652 2564 10658 2576
rect 10652 2536 10916 2564
rect 10652 2524 10658 2536
rect 10778 2496 10784 2508
rect 5316 2468 6132 2496
rect 5316 2456 5322 2468
rect 3283 2400 3556 2428
rect 3605 2431 3663 2437
rect 3283 2397 3295 2400
rect 3237 2391 3295 2397
rect 3605 2397 3617 2431
rect 3651 2428 3663 2431
rect 3878 2428 3884 2440
rect 3651 2400 3884 2428
rect 3651 2397 3663 2400
rect 3605 2391 3663 2397
rect 3878 2388 3884 2400
rect 3936 2388 3942 2440
rect 4062 2428 4068 2440
rect 4023 2400 4068 2428
rect 4062 2388 4068 2400
rect 4120 2388 4126 2440
rect 4430 2428 4436 2440
rect 4391 2400 4436 2428
rect 4430 2388 4436 2400
rect 4488 2388 4494 2440
rect 4890 2428 4896 2440
rect 4851 2400 4896 2428
rect 4890 2388 4896 2400
rect 4948 2388 4954 2440
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2428 5043 2431
rect 5166 2428 5172 2440
rect 5031 2400 5172 2428
rect 5031 2397 5043 2400
rect 4985 2391 5043 2397
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 5810 2428 5816 2440
rect 5771 2400 5816 2428
rect 5810 2388 5816 2400
rect 5868 2388 5874 2440
rect 4338 2360 4344 2372
rect 3068 2332 4344 2360
rect 1581 2295 1639 2301
rect 1581 2261 1593 2295
rect 1627 2292 1639 2295
rect 2222 2292 2228 2304
rect 1627 2264 2228 2292
rect 1627 2261 1639 2264
rect 1581 2255 1639 2261
rect 2222 2252 2228 2264
rect 2280 2252 2286 2304
rect 3068 2301 3096 2332
rect 4338 2320 4344 2332
rect 4396 2320 4402 2372
rect 5258 2360 5264 2372
rect 4816 2332 5264 2360
rect 3053 2295 3111 2301
rect 3053 2261 3065 2295
rect 3099 2261 3111 2295
rect 3053 2255 3111 2261
rect 3421 2295 3479 2301
rect 3421 2261 3433 2295
rect 3467 2292 3479 2295
rect 3786 2292 3792 2304
rect 3467 2264 3792 2292
rect 3467 2261 3479 2264
rect 3421 2255 3479 2261
rect 3786 2252 3792 2264
rect 3844 2252 3850 2304
rect 3881 2295 3939 2301
rect 3881 2261 3893 2295
rect 3927 2292 3939 2295
rect 4816 2292 4844 2332
rect 5258 2320 5264 2332
rect 5316 2320 5322 2372
rect 6104 2360 6132 2468
rect 6932 2468 9904 2496
rect 10437 2468 10660 2496
rect 10739 2468 10784 2496
rect 6181 2431 6239 2437
rect 6181 2397 6193 2431
rect 6227 2428 6239 2431
rect 6270 2428 6276 2440
rect 6227 2400 6276 2428
rect 6227 2397 6239 2400
rect 6181 2391 6239 2397
rect 6270 2388 6276 2400
rect 6328 2388 6334 2440
rect 6365 2431 6423 2437
rect 6365 2397 6377 2431
rect 6411 2428 6423 2431
rect 6822 2428 6828 2440
rect 6411 2400 6828 2428
rect 6411 2397 6423 2400
rect 6365 2391 6423 2397
rect 6822 2388 6828 2400
rect 6880 2388 6886 2440
rect 6932 2437 6960 2468
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2397 6975 2431
rect 7282 2428 7288 2440
rect 7243 2400 7288 2428
rect 6917 2391 6975 2397
rect 7282 2388 7288 2400
rect 7340 2388 7346 2440
rect 8294 2428 8300 2440
rect 7392 2400 8156 2428
rect 8255 2400 8300 2428
rect 7392 2360 7420 2400
rect 6104 2332 7420 2360
rect 7466 2320 7472 2372
rect 7524 2360 7530 2372
rect 7561 2363 7619 2369
rect 7561 2360 7573 2363
rect 7524 2332 7573 2360
rect 7524 2320 7530 2332
rect 7561 2329 7573 2332
rect 7607 2360 7619 2363
rect 7650 2360 7656 2372
rect 7607 2332 7656 2360
rect 7607 2329 7619 2332
rect 7561 2323 7619 2329
rect 7650 2320 7656 2332
rect 7708 2320 7714 2372
rect 7742 2320 7748 2372
rect 7800 2360 7806 2372
rect 7837 2363 7895 2369
rect 7837 2360 7849 2363
rect 7800 2332 7849 2360
rect 7800 2320 7806 2332
rect 7837 2329 7849 2332
rect 7883 2329 7895 2363
rect 7837 2323 7895 2329
rect 5442 2292 5448 2304
rect 3927 2264 4844 2292
rect 5403 2264 5448 2292
rect 3927 2261 3939 2264
rect 3881 2255 3939 2261
rect 5442 2252 5448 2264
rect 5500 2252 5506 2304
rect 5629 2295 5687 2301
rect 5629 2261 5641 2295
rect 5675 2292 5687 2295
rect 5902 2292 5908 2304
rect 5675 2264 5908 2292
rect 5675 2261 5687 2264
rect 5629 2255 5687 2261
rect 5902 2252 5908 2264
rect 5960 2252 5966 2304
rect 5997 2295 6055 2301
rect 5997 2261 6009 2295
rect 6043 2292 6055 2295
rect 6454 2292 6460 2304
rect 6043 2264 6460 2292
rect 6043 2261 6055 2264
rect 5997 2255 6055 2261
rect 6454 2252 6460 2264
rect 6512 2252 6518 2304
rect 6730 2292 6736 2304
rect 6691 2264 6736 2292
rect 6730 2252 6736 2264
rect 6788 2252 6794 2304
rect 7006 2252 7012 2304
rect 7064 2292 7070 2304
rect 7101 2295 7159 2301
rect 7101 2292 7113 2295
rect 7064 2264 7113 2292
rect 7064 2252 7070 2264
rect 7101 2261 7113 2264
rect 7147 2261 7159 2295
rect 7926 2292 7932 2304
rect 7887 2264 7932 2292
rect 7101 2255 7159 2261
rect 7926 2252 7932 2264
rect 7984 2252 7990 2304
rect 8128 2292 8156 2400
rect 8294 2388 8300 2400
rect 8352 2388 8358 2440
rect 8938 2388 8944 2440
rect 8996 2388 9002 2440
rect 9122 2428 9128 2440
rect 9083 2400 9128 2428
rect 9122 2388 9128 2400
rect 9180 2388 9186 2440
rect 9398 2428 9404 2440
rect 9359 2400 9404 2428
rect 9398 2388 9404 2400
rect 9456 2388 9462 2440
rect 9582 2428 9588 2440
rect 9543 2400 9588 2428
rect 9582 2388 9588 2400
rect 9640 2388 9646 2440
rect 9858 2428 9864 2440
rect 9819 2400 9864 2428
rect 9858 2388 9864 2400
rect 9916 2428 9922 2440
rect 10437 2428 10465 2468
rect 9916 2400 10465 2428
rect 10505 2431 10563 2437
rect 9916 2388 9922 2400
rect 10505 2397 10517 2431
rect 10551 2397 10563 2431
rect 10632 2428 10660 2468
rect 10778 2456 10784 2468
rect 10836 2456 10842 2508
rect 10888 2496 10916 2536
rect 11517 2499 11575 2505
rect 11517 2496 11529 2499
rect 10888 2468 11529 2496
rect 11517 2465 11529 2468
rect 11563 2465 11575 2499
rect 11790 2496 11796 2508
rect 11751 2468 11796 2496
rect 11517 2459 11575 2465
rect 11790 2456 11796 2468
rect 11848 2456 11854 2508
rect 11882 2456 11888 2508
rect 11940 2496 11946 2508
rect 13096 2496 13124 2604
rect 13722 2592 13728 2604
rect 13780 2592 13786 2644
rect 13633 2567 13691 2573
rect 13633 2533 13645 2567
rect 13679 2564 13691 2567
rect 13814 2564 13820 2576
rect 13679 2536 13820 2564
rect 13679 2533 13691 2536
rect 13633 2527 13691 2533
rect 13814 2524 13820 2536
rect 13872 2524 13878 2576
rect 14458 2524 14464 2576
rect 14516 2564 14522 2576
rect 15565 2567 15623 2573
rect 15565 2564 15577 2567
rect 14516 2536 15577 2564
rect 14516 2524 14522 2536
rect 15565 2533 15577 2536
rect 15611 2533 15623 2567
rect 15565 2527 15623 2533
rect 11940 2468 13124 2496
rect 11940 2456 11946 2468
rect 13170 2456 13176 2508
rect 13228 2496 13234 2508
rect 14093 2499 14151 2505
rect 14093 2496 14105 2499
rect 13228 2468 14105 2496
rect 13228 2456 13234 2468
rect 14093 2465 14105 2468
rect 14139 2465 14151 2499
rect 14366 2496 14372 2508
rect 14327 2468 14372 2496
rect 14093 2459 14151 2465
rect 14366 2456 14372 2468
rect 14424 2456 14430 2508
rect 11238 2428 11244 2440
rect 10632 2400 11244 2428
rect 10505 2391 10563 2397
rect 8202 2320 8208 2372
rect 8260 2360 8266 2372
rect 8481 2363 8539 2369
rect 8481 2360 8493 2363
rect 8260 2332 8493 2360
rect 8260 2320 8266 2332
rect 8481 2329 8493 2332
rect 8527 2329 8539 2363
rect 8662 2360 8668 2372
rect 8623 2332 8668 2360
rect 8481 2323 8539 2329
rect 8662 2320 8668 2332
rect 8720 2360 8726 2372
rect 8956 2360 8984 2388
rect 8720 2332 8984 2360
rect 8720 2320 8726 2332
rect 10134 2320 10140 2372
rect 10192 2360 10198 2372
rect 10318 2360 10324 2372
rect 10192 2332 10324 2360
rect 10192 2320 10198 2332
rect 10318 2320 10324 2332
rect 10376 2360 10382 2372
rect 10520 2360 10548 2391
rect 11238 2388 11244 2400
rect 11296 2388 11302 2440
rect 11606 2388 11612 2440
rect 11664 2428 11670 2440
rect 12437 2431 12495 2437
rect 12437 2428 12449 2431
rect 11664 2400 12449 2428
rect 11664 2388 11670 2400
rect 12437 2397 12449 2400
rect 12483 2397 12495 2431
rect 12437 2391 12495 2397
rect 12713 2431 12771 2437
rect 12713 2397 12725 2431
rect 12759 2397 12771 2431
rect 12713 2391 12771 2397
rect 10376 2332 10548 2360
rect 10376 2320 10382 2332
rect 10778 2320 10784 2372
rect 10836 2360 10842 2372
rect 12066 2360 12072 2372
rect 10836 2332 12072 2360
rect 10836 2320 10842 2332
rect 12066 2320 12072 2332
rect 12124 2360 12130 2372
rect 12728 2360 12756 2391
rect 12802 2388 12808 2440
rect 12860 2428 12866 2440
rect 13449 2431 13507 2437
rect 13449 2428 13461 2431
rect 12860 2400 13461 2428
rect 12860 2388 12866 2400
rect 13449 2397 13461 2400
rect 13495 2397 13507 2431
rect 13449 2391 13507 2397
rect 13630 2388 13636 2440
rect 13688 2428 13694 2440
rect 13909 2431 13967 2437
rect 13909 2428 13921 2431
rect 13688 2400 13921 2428
rect 13688 2388 13694 2400
rect 13909 2397 13921 2400
rect 13955 2397 13967 2431
rect 15010 2428 15016 2440
rect 14971 2400 15016 2428
rect 13909 2391 13967 2397
rect 15010 2388 15016 2400
rect 15068 2388 15074 2440
rect 15378 2428 15384 2440
rect 15339 2400 15384 2428
rect 15378 2388 15384 2400
rect 15436 2388 15442 2440
rect 14550 2360 14556 2372
rect 12124 2332 12756 2360
rect 13556 2332 14556 2360
rect 12124 2320 12130 2332
rect 8941 2295 8999 2301
rect 8941 2292 8953 2295
rect 8128 2264 8953 2292
rect 8941 2261 8953 2264
rect 8987 2261 8999 2295
rect 8941 2255 8999 2261
rect 9674 2252 9680 2304
rect 9732 2292 9738 2304
rect 13556 2292 13584 2332
rect 14550 2320 14556 2332
rect 14608 2320 14614 2372
rect 13722 2292 13728 2304
rect 9732 2264 13584 2292
rect 13683 2264 13728 2292
rect 9732 2252 9738 2264
rect 13722 2252 13728 2264
rect 13780 2252 13786 2304
rect 14182 2252 14188 2304
rect 14240 2292 14246 2304
rect 15197 2295 15255 2301
rect 15197 2292 15209 2295
rect 14240 2264 15209 2292
rect 14240 2252 14246 2264
rect 15197 2261 15209 2264
rect 15243 2261 15255 2295
rect 15197 2255 15255 2261
rect 1104 2202 16008 2224
rect 1104 2150 4698 2202
rect 4750 2150 4762 2202
rect 4814 2150 4826 2202
rect 4878 2150 4890 2202
rect 4942 2150 4954 2202
rect 5006 2150 8446 2202
rect 8498 2150 8510 2202
rect 8562 2150 8574 2202
rect 8626 2150 8638 2202
rect 8690 2150 8702 2202
rect 8754 2150 12194 2202
rect 12246 2150 12258 2202
rect 12310 2150 12322 2202
rect 12374 2150 12386 2202
rect 12438 2150 12450 2202
rect 12502 2150 16008 2202
rect 1104 2128 16008 2150
rect 3786 2048 3792 2100
rect 3844 2088 3850 2100
rect 5166 2088 5172 2100
rect 3844 2060 5172 2088
rect 3844 2048 3850 2060
rect 5166 2048 5172 2060
rect 5224 2048 5230 2100
rect 6270 2048 6276 2100
rect 6328 2088 6334 2100
rect 6328 2060 12434 2088
rect 6328 2048 6334 2060
rect 4062 1980 4068 2032
rect 4120 2020 4126 2032
rect 7098 2020 7104 2032
rect 4120 1992 7104 2020
rect 4120 1980 4126 1992
rect 7098 1980 7104 1992
rect 7156 1980 7162 2032
rect 9398 2020 9404 2032
rect 7208 1992 9404 2020
rect 4154 1912 4160 1964
rect 4212 1952 4218 1964
rect 5626 1952 5632 1964
rect 4212 1924 5632 1952
rect 4212 1912 4218 1924
rect 5626 1912 5632 1924
rect 5684 1912 5690 1964
rect 5994 1912 6000 1964
rect 6052 1952 6058 1964
rect 7208 1952 7236 1992
rect 9398 1980 9404 1992
rect 9456 2020 9462 2032
rect 9582 2020 9588 2032
rect 9456 1992 9588 2020
rect 9456 1980 9462 1992
rect 9582 1980 9588 1992
rect 9640 1980 9646 2032
rect 12406 2020 12434 2060
rect 13722 2020 13728 2032
rect 12406 1992 13728 2020
rect 13722 1980 13728 1992
rect 13780 1980 13786 2032
rect 6052 1924 7236 1952
rect 6052 1912 6058 1924
rect 7282 1912 7288 1964
rect 7340 1952 7346 1964
rect 16022 1952 16028 1964
rect 7340 1924 16028 1952
rect 7340 1912 7346 1924
rect 16022 1912 16028 1924
rect 16080 1912 16086 1964
rect 4430 1844 4436 1896
rect 4488 1884 4494 1896
rect 9306 1884 9312 1896
rect 4488 1856 9312 1884
rect 4488 1844 4494 1856
rect 9306 1844 9312 1856
rect 9364 1844 9370 1896
rect 12250 1844 12256 1896
rect 12308 1884 12314 1896
rect 13170 1884 13176 1896
rect 12308 1856 13176 1884
rect 12308 1844 12314 1856
rect 13170 1844 13176 1856
rect 13228 1844 13234 1896
rect 2958 1776 2964 1828
rect 3016 1816 3022 1828
rect 7374 1816 7380 1828
rect 3016 1788 7380 1816
rect 3016 1776 3022 1788
rect 7374 1776 7380 1788
rect 7432 1776 7438 1828
rect 5534 1708 5540 1760
rect 5592 1748 5598 1760
rect 7926 1748 7932 1760
rect 5592 1720 7932 1748
rect 5592 1708 5598 1720
rect 7926 1708 7932 1720
rect 7984 1708 7990 1760
rect 11146 1708 11152 1760
rect 11204 1748 11210 1760
rect 11606 1748 11612 1760
rect 11204 1720 11612 1748
rect 11204 1708 11210 1720
rect 11606 1708 11612 1720
rect 11664 1708 11670 1760
rect 3510 1640 3516 1692
rect 3568 1680 3574 1692
rect 8202 1680 8208 1692
rect 3568 1652 8208 1680
rect 3568 1640 3574 1652
rect 8202 1640 8208 1652
rect 8260 1640 8266 1692
rect 5442 1572 5448 1624
rect 5500 1612 5506 1624
rect 9214 1612 9220 1624
rect 5500 1584 9220 1612
rect 5500 1572 5506 1584
rect 9214 1572 9220 1584
rect 9272 1572 9278 1624
rect 6914 1300 6920 1352
rect 6972 1340 6978 1352
rect 7834 1340 7840 1352
rect 6972 1312 7840 1340
rect 6972 1300 6978 1312
rect 7834 1300 7840 1312
rect 7892 1300 7898 1352
<< via1 >>
rect 11704 17892 11756 17944
rect 13084 17892 13136 17944
rect 9680 17824 9732 17876
rect 10232 17824 10284 17876
rect 13728 17824 13780 17876
rect 12440 17756 12492 17808
rect 13360 17756 13412 17808
rect 9220 17688 9272 17740
rect 13452 17688 13504 17740
rect 12624 17620 12676 17672
rect 15660 17620 15712 17672
rect 16120 17620 16172 17672
rect 11336 17552 11388 17604
rect 16488 17552 16540 17604
rect 12808 17484 12860 17536
rect 13636 17484 13688 17536
rect 4698 17382 4750 17434
rect 4762 17382 4814 17434
rect 4826 17382 4878 17434
rect 4890 17382 4942 17434
rect 4954 17382 5006 17434
rect 8446 17382 8498 17434
rect 8510 17382 8562 17434
rect 8574 17382 8626 17434
rect 8638 17382 8690 17434
rect 8702 17382 8754 17434
rect 12194 17382 12246 17434
rect 12258 17382 12310 17434
rect 12322 17382 12374 17434
rect 12386 17382 12438 17434
rect 12450 17382 12502 17434
rect 1400 17280 1452 17332
rect 6920 17280 6972 17332
rect 7288 17280 7340 17332
rect 7656 17280 7708 17332
rect 8024 17280 8076 17332
rect 8300 17280 8352 17332
rect 8852 17280 8904 17332
rect 9128 17280 9180 17332
rect 9496 17280 9548 17332
rect 2320 17212 2372 17264
rect 2044 17144 2096 17196
rect 2504 17187 2556 17196
rect 2504 17153 2513 17187
rect 2513 17153 2547 17187
rect 2547 17153 2556 17187
rect 2504 17144 2556 17153
rect 3332 17187 3384 17196
rect 2596 17076 2648 17128
rect 3332 17153 3341 17187
rect 3341 17153 3375 17187
rect 3375 17153 3384 17187
rect 3332 17144 3384 17153
rect 3792 17187 3844 17196
rect 3792 17153 3801 17187
rect 3801 17153 3835 17187
rect 3835 17153 3844 17187
rect 3792 17144 3844 17153
rect 3884 17144 3936 17196
rect 4344 17144 4396 17196
rect 3424 17076 3476 17128
rect 1676 17008 1728 17060
rect 3240 17008 3292 17060
rect 3608 17008 3660 17060
rect 3976 17051 4028 17060
rect 3976 17017 3985 17051
rect 3985 17017 4019 17051
rect 4019 17017 4028 17051
rect 3976 17008 4028 17017
rect 4620 17008 4672 17060
rect 5448 17212 5500 17264
rect 6276 17212 6328 17264
rect 9312 17212 9364 17264
rect 11152 17280 11204 17332
rect 11520 17280 11572 17332
rect 5172 17187 5224 17196
rect 5172 17153 5181 17187
rect 5181 17153 5215 17187
rect 5215 17153 5224 17187
rect 5172 17144 5224 17153
rect 5632 17187 5684 17196
rect 5632 17153 5641 17187
rect 5641 17153 5675 17187
rect 5675 17153 5684 17187
rect 5632 17144 5684 17153
rect 6000 17144 6052 17196
rect 7288 17187 7340 17196
rect 2136 16940 2188 16992
rect 2412 16940 2464 16992
rect 2872 16940 2924 16992
rect 7288 17153 7297 17187
rect 7297 17153 7331 17187
rect 7331 17153 7340 17187
rect 7288 17144 7340 17153
rect 7656 17187 7708 17196
rect 7656 17153 7665 17187
rect 7665 17153 7699 17187
rect 7699 17153 7708 17187
rect 7656 17144 7708 17153
rect 8392 17187 8444 17196
rect 6184 17008 6236 17060
rect 5264 16983 5316 16992
rect 5264 16949 5273 16983
rect 5273 16949 5307 16983
rect 5307 16949 5316 16983
rect 5264 16940 5316 16949
rect 5540 16940 5592 16992
rect 7564 17076 7616 17128
rect 8392 17153 8401 17187
rect 8401 17153 8435 17187
rect 8435 17153 8444 17187
rect 8392 17144 8444 17153
rect 9220 17187 9272 17196
rect 8300 17076 8352 17128
rect 9220 17153 9229 17187
rect 9229 17153 9263 17187
rect 9263 17153 9272 17187
rect 9220 17144 9272 17153
rect 11336 17187 11388 17196
rect 9772 17119 9824 17128
rect 9772 17085 9781 17119
rect 9781 17085 9815 17119
rect 9815 17085 9824 17119
rect 9772 17076 9824 17085
rect 9956 17119 10008 17128
rect 9956 17085 9965 17119
rect 9965 17085 9999 17119
rect 9999 17085 10008 17119
rect 9956 17076 10008 17085
rect 10784 17076 10836 17128
rect 11336 17153 11345 17187
rect 11345 17153 11379 17187
rect 11379 17153 11388 17187
rect 11336 17144 11388 17153
rect 11520 17119 11572 17128
rect 11520 17085 11529 17119
rect 11529 17085 11563 17119
rect 11563 17085 11572 17119
rect 11796 17119 11848 17128
rect 11520 17076 11572 17085
rect 11796 17085 11805 17119
rect 11805 17085 11839 17119
rect 11839 17085 11848 17119
rect 11796 17076 11848 17085
rect 12072 17144 12124 17196
rect 13268 17187 13320 17196
rect 13268 17153 13277 17187
rect 13277 17153 13311 17187
rect 13311 17153 13320 17187
rect 13268 17144 13320 17153
rect 13728 17187 13780 17196
rect 12900 17076 12952 17128
rect 12992 17119 13044 17128
rect 12992 17085 13001 17119
rect 13001 17085 13035 17119
rect 13035 17085 13044 17119
rect 12992 17076 13044 17085
rect 9220 16940 9272 16992
rect 10140 16940 10192 16992
rect 12716 17008 12768 17060
rect 13084 17008 13136 17060
rect 13728 17153 13737 17187
rect 13737 17153 13771 17187
rect 13771 17153 13780 17187
rect 13728 17144 13780 17153
rect 13912 17144 13964 17196
rect 16028 17144 16080 17196
rect 13636 17076 13688 17128
rect 16580 17076 16632 17128
rect 12256 16940 12308 16992
rect 13728 16940 13780 16992
rect 15200 16940 15252 16992
rect 16396 16940 16448 16992
rect 2824 16838 2876 16890
rect 2888 16838 2940 16890
rect 2952 16838 3004 16890
rect 3016 16838 3068 16890
rect 3080 16838 3132 16890
rect 6572 16838 6624 16890
rect 6636 16838 6688 16890
rect 6700 16838 6752 16890
rect 6764 16838 6816 16890
rect 6828 16838 6880 16890
rect 10320 16838 10372 16890
rect 10384 16838 10436 16890
rect 10448 16838 10500 16890
rect 10512 16838 10564 16890
rect 10576 16838 10628 16890
rect 14068 16838 14120 16890
rect 14132 16838 14184 16890
rect 14196 16838 14248 16890
rect 14260 16838 14312 16890
rect 14324 16838 14376 16890
rect 1768 16668 1820 16720
rect 6000 16736 6052 16788
rect 6276 16736 6328 16788
rect 7288 16736 7340 16788
rect 8392 16736 8444 16788
rect 3792 16668 3844 16720
rect 4344 16711 4396 16720
rect 4344 16677 4353 16711
rect 4353 16677 4387 16711
rect 4387 16677 4396 16711
rect 4344 16668 4396 16677
rect 7932 16668 7984 16720
rect 9864 16736 9916 16788
rect 10232 16779 10284 16788
rect 10232 16745 10241 16779
rect 10241 16745 10275 16779
rect 10275 16745 10284 16779
rect 10232 16736 10284 16745
rect 10324 16736 10376 16788
rect 7472 16643 7524 16652
rect 296 16532 348 16584
rect 1492 16575 1544 16584
rect 1492 16541 1501 16575
rect 1501 16541 1535 16575
rect 1535 16541 1544 16575
rect 1768 16575 1820 16584
rect 1492 16532 1544 16541
rect 1768 16541 1777 16575
rect 1777 16541 1811 16575
rect 1811 16541 1820 16575
rect 1768 16532 1820 16541
rect 2044 16464 2096 16516
rect 1584 16396 1636 16448
rect 2412 16575 2464 16584
rect 2412 16541 2421 16575
rect 2421 16541 2455 16575
rect 2455 16541 2464 16575
rect 3056 16575 3108 16584
rect 2412 16532 2464 16541
rect 3056 16541 3065 16575
rect 3065 16541 3099 16575
rect 3099 16541 3108 16575
rect 3056 16532 3108 16541
rect 3148 16575 3200 16584
rect 3148 16541 3157 16575
rect 3157 16541 3191 16575
rect 3191 16541 3200 16575
rect 3148 16532 3200 16541
rect 3792 16532 3844 16584
rect 4068 16532 4120 16584
rect 2688 16464 2740 16516
rect 2872 16439 2924 16448
rect 2872 16405 2881 16439
rect 2881 16405 2915 16439
rect 2915 16405 2924 16439
rect 2872 16396 2924 16405
rect 3884 16396 3936 16448
rect 4252 16532 4304 16584
rect 7472 16609 7481 16643
rect 7481 16609 7515 16643
rect 7515 16609 7524 16643
rect 7472 16600 7524 16609
rect 5632 16575 5684 16584
rect 5632 16541 5666 16575
rect 5666 16541 5684 16575
rect 5632 16532 5684 16541
rect 7840 16575 7892 16584
rect 7840 16541 7849 16575
rect 7849 16541 7883 16575
rect 7883 16541 7892 16575
rect 7840 16532 7892 16541
rect 10508 16668 10560 16720
rect 11796 16668 11848 16720
rect 4344 16396 4396 16448
rect 4436 16396 4488 16448
rect 4712 16396 4764 16448
rect 9864 16600 9916 16652
rect 10048 16532 10100 16584
rect 5080 16396 5132 16448
rect 7012 16396 7064 16448
rect 8392 16396 8444 16448
rect 9312 16396 9364 16448
rect 9496 16464 9548 16516
rect 11152 16600 11204 16652
rect 12440 16736 12492 16788
rect 12900 16736 12952 16788
rect 16488 16736 16540 16788
rect 12256 16668 12308 16720
rect 11244 16532 11296 16584
rect 13360 16643 13412 16652
rect 13360 16609 13369 16643
rect 13369 16609 13403 16643
rect 13403 16609 13412 16643
rect 14096 16643 14148 16652
rect 13360 16600 13412 16609
rect 14096 16609 14105 16643
rect 14105 16609 14139 16643
rect 14139 16609 14148 16643
rect 14096 16600 14148 16609
rect 14832 16600 14884 16652
rect 10416 16464 10468 16516
rect 12624 16532 12676 16584
rect 12716 16532 12768 16584
rect 12992 16532 13044 16584
rect 13084 16575 13136 16584
rect 13084 16541 13093 16575
rect 13093 16541 13127 16575
rect 13127 16541 13136 16575
rect 13084 16532 13136 16541
rect 13636 16532 13688 16584
rect 12900 16464 12952 16516
rect 13268 16464 13320 16516
rect 13820 16464 13872 16516
rect 9588 16396 9640 16448
rect 11152 16396 11204 16448
rect 12072 16396 12124 16448
rect 12624 16396 12676 16448
rect 15016 16439 15068 16448
rect 15016 16405 15025 16439
rect 15025 16405 15059 16439
rect 15059 16405 15068 16439
rect 15016 16396 15068 16405
rect 15844 16532 15896 16584
rect 16580 16464 16632 16516
rect 15568 16396 15620 16448
rect 4698 16294 4750 16346
rect 4762 16294 4814 16346
rect 4826 16294 4878 16346
rect 4890 16294 4942 16346
rect 4954 16294 5006 16346
rect 8446 16294 8498 16346
rect 8510 16294 8562 16346
rect 8574 16294 8626 16346
rect 8638 16294 8690 16346
rect 8702 16294 8754 16346
rect 12194 16294 12246 16346
rect 12258 16294 12310 16346
rect 12322 16294 12374 16346
rect 12386 16294 12438 16346
rect 12450 16294 12502 16346
rect 1492 16235 1544 16244
rect 1492 16201 1501 16235
rect 1501 16201 1535 16235
rect 1535 16201 1544 16235
rect 1492 16192 1544 16201
rect 1860 16235 1912 16244
rect 1860 16201 1869 16235
rect 1869 16201 1903 16235
rect 1903 16201 1912 16235
rect 1860 16192 1912 16201
rect 2320 16235 2372 16244
rect 2320 16201 2329 16235
rect 2329 16201 2363 16235
rect 2363 16201 2372 16235
rect 2320 16192 2372 16201
rect 3332 16192 3384 16244
rect 4252 16192 4304 16244
rect 5172 16192 5224 16244
rect 5816 16192 5868 16244
rect 6460 16192 6512 16244
rect 7564 16235 7616 16244
rect 1768 16056 1820 16108
rect 2136 16099 2188 16108
rect 2136 16065 2145 16099
rect 2145 16065 2179 16099
rect 2179 16065 2188 16099
rect 4068 16124 4120 16176
rect 4620 16124 4672 16176
rect 2136 16056 2188 16065
rect 3240 16056 3292 16108
rect 664 15988 716 16040
rect 2872 15988 2924 16040
rect 3608 16099 3660 16108
rect 3608 16065 3617 16099
rect 3617 16065 3651 16099
rect 3651 16065 3660 16099
rect 3608 16056 3660 16065
rect 4528 16056 4580 16108
rect 5632 16099 5684 16108
rect 5632 16065 5641 16099
rect 5641 16065 5675 16099
rect 5675 16065 5684 16099
rect 5632 16056 5684 16065
rect 7104 16124 7156 16176
rect 3700 15988 3752 16040
rect 3424 15920 3476 15972
rect 7564 16201 7573 16235
rect 7573 16201 7607 16235
rect 7607 16201 7616 16235
rect 7564 16192 7616 16201
rect 7656 16192 7708 16244
rect 8300 16192 8352 16244
rect 8576 16192 8628 16244
rect 9588 16192 9640 16244
rect 9772 16192 9824 16244
rect 12072 16192 12124 16244
rect 13176 16192 13228 16244
rect 14096 16192 14148 16244
rect 9128 16124 9180 16176
rect 10048 16124 10100 16176
rect 10324 16124 10376 16176
rect 10692 16124 10744 16176
rect 7656 16056 7708 16108
rect 7564 15988 7616 16040
rect 8208 16099 8260 16108
rect 8208 16065 8217 16099
rect 8217 16065 8251 16099
rect 8251 16065 8260 16099
rect 8208 16056 8260 16065
rect 9588 16056 9640 16108
rect 10232 16099 10284 16108
rect 10232 16065 10241 16099
rect 10241 16065 10275 16099
rect 10275 16065 10284 16099
rect 10232 16056 10284 16065
rect 10968 16099 11020 16108
rect 10968 16065 10977 16099
rect 10977 16065 11011 16099
rect 11011 16065 11020 16099
rect 10968 16056 11020 16065
rect 11888 16099 11940 16108
rect 11888 16065 11897 16099
rect 11897 16065 11931 16099
rect 11931 16065 11940 16099
rect 11888 16056 11940 16065
rect 12164 16056 12216 16108
rect 13544 16124 13596 16176
rect 12532 16099 12584 16108
rect 12532 16065 12541 16099
rect 12541 16065 12575 16099
rect 12575 16065 12584 16099
rect 12532 16056 12584 16065
rect 12900 16056 12952 16108
rect 8116 15988 8168 16040
rect 7656 15920 7708 15972
rect 8944 15920 8996 15972
rect 2320 15852 2372 15904
rect 3608 15852 3660 15904
rect 3884 15895 3936 15904
rect 3884 15861 3893 15895
rect 3893 15861 3927 15895
rect 3927 15861 3936 15895
rect 3884 15852 3936 15861
rect 7104 15852 7156 15904
rect 8208 15852 8260 15904
rect 8300 15852 8352 15904
rect 10692 15988 10744 16040
rect 10876 15988 10928 16040
rect 11980 16031 12032 16040
rect 10232 15920 10284 15972
rect 10784 15920 10836 15972
rect 11980 15997 11989 16031
rect 11989 15997 12023 16031
rect 12023 15997 12032 16031
rect 11980 15988 12032 15997
rect 12072 16031 12124 16040
rect 12072 15997 12081 16031
rect 12081 15997 12115 16031
rect 12115 15997 12124 16031
rect 12072 15988 12124 15997
rect 12716 15988 12768 16040
rect 11336 15920 11388 15972
rect 12900 15920 12952 15972
rect 14740 16124 14792 16176
rect 15752 16124 15804 16176
rect 14464 16056 14516 16108
rect 15384 16056 15436 16108
rect 14004 15988 14056 16040
rect 13636 15920 13688 15972
rect 10416 15895 10468 15904
rect 10416 15861 10425 15895
rect 10425 15861 10459 15895
rect 10459 15861 10468 15895
rect 10416 15852 10468 15861
rect 11428 15852 11480 15904
rect 13268 15852 13320 15904
rect 15292 15852 15344 15904
rect 2824 15750 2876 15802
rect 2888 15750 2940 15802
rect 2952 15750 3004 15802
rect 3016 15750 3068 15802
rect 3080 15750 3132 15802
rect 6572 15750 6624 15802
rect 6636 15750 6688 15802
rect 6700 15750 6752 15802
rect 6764 15750 6816 15802
rect 6828 15750 6880 15802
rect 10320 15750 10372 15802
rect 10384 15750 10436 15802
rect 10448 15750 10500 15802
rect 10512 15750 10564 15802
rect 10576 15750 10628 15802
rect 14068 15750 14120 15802
rect 14132 15750 14184 15802
rect 14196 15750 14248 15802
rect 14260 15750 14312 15802
rect 14324 15750 14376 15802
rect 5264 15648 5316 15700
rect 7380 15691 7432 15700
rect 7380 15657 7389 15691
rect 7389 15657 7423 15691
rect 7423 15657 7432 15691
rect 10968 15691 11020 15700
rect 7380 15648 7432 15657
rect 7656 15580 7708 15632
rect 8760 15580 8812 15632
rect 9036 15580 9088 15632
rect 9220 15580 9272 15632
rect 10968 15657 10977 15691
rect 10977 15657 11011 15691
rect 11011 15657 11020 15691
rect 10968 15648 11020 15657
rect 12532 15648 12584 15700
rect 13912 15648 13964 15700
rect 11336 15580 11388 15632
rect 11612 15580 11664 15632
rect 13084 15580 13136 15632
rect 13452 15623 13504 15632
rect 13452 15589 13461 15623
rect 13461 15589 13495 15623
rect 13495 15589 13504 15623
rect 13452 15580 13504 15589
rect 14464 15623 14516 15632
rect 14464 15589 14473 15623
rect 14473 15589 14507 15623
rect 14507 15589 14516 15623
rect 14464 15580 14516 15589
rect 14648 15580 14700 15632
rect 3976 15512 4028 15564
rect 11428 15555 11480 15564
rect 2320 15376 2372 15428
rect 2780 15376 2832 15428
rect 3148 15376 3200 15428
rect 3516 15376 3568 15428
rect 1492 15351 1544 15360
rect 1492 15317 1501 15351
rect 1501 15317 1535 15351
rect 1535 15317 1544 15351
rect 1492 15308 1544 15317
rect 2228 15351 2280 15360
rect 2228 15317 2237 15351
rect 2237 15317 2271 15351
rect 2271 15317 2280 15351
rect 2228 15308 2280 15317
rect 4620 15444 4672 15496
rect 7472 15444 7524 15496
rect 8944 15444 8996 15496
rect 11428 15521 11437 15555
rect 11437 15521 11471 15555
rect 11471 15521 11480 15555
rect 11428 15512 11480 15521
rect 11520 15555 11572 15564
rect 11520 15521 11529 15555
rect 11529 15521 11563 15555
rect 11563 15521 11572 15555
rect 11520 15512 11572 15521
rect 12072 15512 12124 15564
rect 12900 15512 12952 15564
rect 13912 15512 13964 15564
rect 10600 15444 10652 15496
rect 12164 15444 12216 15496
rect 3884 15351 3936 15360
rect 3884 15317 3893 15351
rect 3893 15317 3927 15351
rect 3927 15317 3936 15351
rect 3884 15308 3936 15317
rect 5172 15376 5224 15428
rect 6920 15376 6972 15428
rect 8116 15376 8168 15428
rect 8668 15376 8720 15428
rect 9956 15376 10008 15428
rect 10968 15376 11020 15428
rect 12808 15376 12860 15428
rect 13268 15444 13320 15496
rect 14648 15487 14700 15496
rect 5908 15308 5960 15360
rect 6828 15351 6880 15360
rect 6828 15317 6837 15351
rect 6837 15317 6871 15351
rect 6871 15317 6880 15351
rect 6828 15308 6880 15317
rect 7840 15308 7892 15360
rect 8852 15308 8904 15360
rect 9772 15308 9824 15360
rect 11336 15351 11388 15360
rect 11336 15317 11345 15351
rect 11345 15317 11379 15351
rect 11379 15317 11388 15351
rect 11336 15308 11388 15317
rect 11796 15351 11848 15360
rect 11796 15317 11805 15351
rect 11805 15317 11839 15351
rect 11839 15317 11848 15351
rect 11796 15308 11848 15317
rect 11980 15308 12032 15360
rect 12992 15351 13044 15360
rect 12992 15317 13001 15351
rect 13001 15317 13035 15351
rect 13035 15317 13044 15351
rect 12992 15308 13044 15317
rect 13084 15351 13136 15360
rect 13084 15317 13093 15351
rect 13093 15317 13127 15351
rect 13127 15317 13136 15351
rect 13084 15308 13136 15317
rect 13452 15308 13504 15360
rect 13636 15308 13688 15360
rect 13820 15376 13872 15428
rect 14004 15376 14056 15428
rect 14648 15453 14657 15487
rect 14657 15453 14691 15487
rect 14691 15453 14700 15487
rect 14648 15444 14700 15453
rect 16212 15444 16264 15496
rect 15936 15376 15988 15428
rect 16672 15308 16724 15360
rect 4698 15206 4750 15258
rect 4762 15206 4814 15258
rect 4826 15206 4878 15258
rect 4890 15206 4942 15258
rect 4954 15206 5006 15258
rect 8446 15206 8498 15258
rect 8510 15206 8562 15258
rect 8574 15206 8626 15258
rect 8638 15206 8690 15258
rect 8702 15206 8754 15258
rect 12194 15206 12246 15258
rect 12258 15206 12310 15258
rect 12322 15206 12374 15258
rect 12386 15206 12438 15258
rect 12450 15206 12502 15258
rect 2136 15104 2188 15156
rect 2504 15147 2556 15156
rect 2504 15113 2513 15147
rect 2513 15113 2547 15147
rect 2547 15113 2556 15147
rect 2504 15104 2556 15113
rect 4160 15036 4212 15088
rect 4804 15036 4856 15088
rect 2412 15011 2464 15020
rect 2412 14977 2421 15011
rect 2421 14977 2455 15011
rect 2455 14977 2464 15011
rect 2412 14968 2464 14977
rect 2504 14968 2556 15020
rect 2780 15011 2832 15020
rect 2780 14977 2789 15011
rect 2789 14977 2823 15011
rect 2823 14977 2832 15011
rect 2780 14968 2832 14977
rect 4252 14968 4304 15020
rect 6092 14968 6144 15020
rect 6920 14968 6972 15020
rect 1400 14900 1452 14952
rect 1676 14943 1728 14952
rect 1676 14909 1685 14943
rect 1685 14909 1719 14943
rect 1719 14909 1728 14943
rect 1676 14900 1728 14909
rect 4620 14900 4672 14952
rect 7656 15104 7708 15156
rect 8944 15147 8996 15156
rect 8944 15113 8953 15147
rect 8953 15113 8987 15147
rect 8987 15113 8996 15147
rect 8944 15104 8996 15113
rect 7380 15079 7432 15088
rect 7380 15045 7414 15079
rect 7414 15045 7432 15079
rect 7380 15036 7432 15045
rect 7564 15036 7616 15088
rect 10140 15036 10192 15088
rect 10876 15104 10928 15156
rect 11888 15104 11940 15156
rect 12164 15104 12216 15156
rect 9864 14968 9916 15020
rect 11060 15036 11112 15088
rect 13360 15147 13412 15156
rect 13360 15113 13369 15147
rect 13369 15113 13403 15147
rect 13403 15113 13412 15147
rect 13360 15104 13412 15113
rect 1860 14832 1912 14884
rect 6000 14832 6052 14884
rect 2044 14764 2096 14816
rect 3424 14764 3476 14816
rect 4344 14764 4396 14816
rect 4804 14807 4856 14816
rect 4804 14773 4813 14807
rect 4813 14773 4847 14807
rect 4847 14773 4856 14807
rect 4804 14764 4856 14773
rect 5356 14764 5408 14816
rect 5632 14764 5684 14816
rect 6460 14764 6512 14816
rect 8116 14900 8168 14952
rect 9128 14900 9180 14952
rect 10600 14900 10652 14952
rect 9496 14832 9548 14884
rect 11244 14900 11296 14952
rect 9128 14807 9180 14816
rect 9128 14773 9137 14807
rect 9137 14773 9171 14807
rect 9171 14773 9180 14807
rect 9128 14764 9180 14773
rect 10140 14764 10192 14816
rect 13820 15036 13872 15088
rect 15200 15104 15252 15156
rect 11888 14832 11940 14884
rect 11152 14764 11204 14816
rect 11520 14764 11572 14816
rect 12072 14764 12124 14816
rect 14004 14968 14056 15020
rect 12716 14900 12768 14952
rect 12256 14832 12308 14884
rect 13360 14900 13412 14952
rect 14924 15036 14976 15088
rect 15660 14968 15712 15020
rect 15844 14832 15896 14884
rect 12532 14807 12584 14816
rect 12532 14773 12541 14807
rect 12541 14773 12575 14807
rect 12575 14773 12584 14807
rect 12532 14764 12584 14773
rect 12992 14764 13044 14816
rect 13544 14764 13596 14816
rect 14740 14807 14792 14816
rect 14740 14773 14749 14807
rect 14749 14773 14783 14807
rect 14783 14773 14792 14807
rect 14740 14764 14792 14773
rect 14924 14764 14976 14816
rect 2824 14662 2876 14714
rect 2888 14662 2940 14714
rect 2952 14662 3004 14714
rect 3016 14662 3068 14714
rect 3080 14662 3132 14714
rect 6572 14662 6624 14714
rect 6636 14662 6688 14714
rect 6700 14662 6752 14714
rect 6764 14662 6816 14714
rect 6828 14662 6880 14714
rect 10320 14662 10372 14714
rect 10384 14662 10436 14714
rect 10448 14662 10500 14714
rect 10512 14662 10564 14714
rect 10576 14662 10628 14714
rect 14068 14662 14120 14714
rect 14132 14662 14184 14714
rect 14196 14662 14248 14714
rect 14260 14662 14312 14714
rect 14324 14662 14376 14714
rect 1768 14603 1820 14612
rect 1768 14569 1777 14603
rect 1777 14569 1811 14603
rect 1811 14569 1820 14603
rect 1768 14560 1820 14569
rect 1768 14356 1820 14408
rect 1952 14399 2004 14408
rect 1952 14365 1961 14399
rect 1961 14365 1995 14399
rect 1995 14365 2004 14399
rect 1952 14356 2004 14365
rect 2228 14399 2280 14408
rect 2228 14365 2237 14399
rect 2237 14365 2271 14399
rect 2271 14365 2280 14399
rect 9588 14560 9640 14612
rect 10968 14560 11020 14612
rect 11336 14560 11388 14612
rect 3792 14492 3844 14544
rect 11520 14492 11572 14544
rect 12164 14492 12216 14544
rect 2872 14467 2924 14476
rect 2872 14433 2881 14467
rect 2881 14433 2915 14467
rect 2915 14433 2924 14467
rect 3148 14467 3200 14476
rect 2872 14424 2924 14433
rect 3148 14433 3157 14467
rect 3157 14433 3191 14467
rect 3191 14433 3200 14467
rect 3148 14424 3200 14433
rect 4160 14424 4212 14476
rect 4620 14424 4672 14476
rect 5448 14424 5500 14476
rect 12624 14492 12676 14544
rect 13544 14560 13596 14612
rect 13636 14560 13688 14612
rect 14648 14560 14700 14612
rect 12808 14467 12860 14476
rect 6460 14399 6512 14408
rect 2228 14356 2280 14365
rect 6460 14365 6469 14399
rect 6469 14365 6503 14399
rect 6503 14365 6512 14399
rect 6460 14356 6512 14365
rect 8208 14356 8260 14408
rect 9956 14356 10008 14408
rect 10968 14399 11020 14408
rect 10968 14365 10977 14399
rect 10977 14365 11011 14399
rect 11011 14365 11020 14399
rect 10968 14356 11020 14365
rect 2780 14288 2832 14340
rect 6092 14288 6144 14340
rect 6368 14288 6420 14340
rect 6644 14288 6696 14340
rect 7656 14331 7708 14340
rect 7656 14297 7674 14331
rect 7674 14297 7708 14331
rect 7656 14288 7708 14297
rect 8300 14288 8352 14340
rect 9036 14288 9088 14340
rect 12808 14433 12817 14467
rect 12817 14433 12851 14467
rect 12851 14433 12860 14467
rect 12808 14424 12860 14433
rect 12992 14424 13044 14476
rect 13176 14424 13228 14476
rect 14004 14424 14056 14476
rect 15660 14467 15712 14476
rect 15660 14433 15669 14467
rect 15669 14433 15703 14467
rect 15703 14433 15712 14467
rect 15660 14424 15712 14433
rect 16856 14424 16908 14476
rect 11704 14356 11756 14408
rect 15384 14399 15436 14408
rect 15384 14365 15393 14399
rect 15393 14365 15427 14399
rect 15427 14365 15436 14399
rect 15384 14356 15436 14365
rect 16764 14356 16816 14408
rect 13176 14288 13228 14340
rect 13544 14331 13596 14340
rect 13544 14297 13553 14331
rect 13553 14297 13587 14331
rect 13587 14297 13596 14331
rect 13544 14288 13596 14297
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 3240 14220 3292 14272
rect 4068 14220 4120 14272
rect 5172 14220 5224 14272
rect 5816 14220 5868 14272
rect 7196 14220 7248 14272
rect 10692 14220 10744 14272
rect 11428 14263 11480 14272
rect 11428 14229 11437 14263
rect 11437 14229 11471 14263
rect 11471 14229 11480 14263
rect 11428 14220 11480 14229
rect 11520 14220 11572 14272
rect 11704 14220 11756 14272
rect 12256 14263 12308 14272
rect 12256 14229 12265 14263
rect 12265 14229 12299 14263
rect 12299 14229 12308 14263
rect 12256 14220 12308 14229
rect 12440 14220 12492 14272
rect 12624 14220 12676 14272
rect 14096 14220 14148 14272
rect 4698 14118 4750 14170
rect 4762 14118 4814 14170
rect 4826 14118 4878 14170
rect 4890 14118 4942 14170
rect 4954 14118 5006 14170
rect 8446 14118 8498 14170
rect 8510 14118 8562 14170
rect 8574 14118 8626 14170
rect 8638 14118 8690 14170
rect 8702 14118 8754 14170
rect 12194 14118 12246 14170
rect 12258 14118 12310 14170
rect 12322 14118 12374 14170
rect 12386 14118 12438 14170
rect 12450 14118 12502 14170
rect 1676 14016 1728 14068
rect 1768 14016 1820 14068
rect 2596 14016 2648 14068
rect 2872 14059 2924 14068
rect 2872 14025 2881 14059
rect 2881 14025 2915 14059
rect 2915 14025 2924 14059
rect 2872 14016 2924 14025
rect 3148 14059 3200 14068
rect 3148 14025 3157 14059
rect 3157 14025 3191 14059
rect 3191 14025 3200 14059
rect 3148 14016 3200 14025
rect 4620 14059 4672 14068
rect 4620 14025 4629 14059
rect 4629 14025 4663 14059
rect 4663 14025 4672 14059
rect 4620 14016 4672 14025
rect 5448 14016 5500 14068
rect 5724 14016 5776 14068
rect 6460 14016 6512 14068
rect 6920 14059 6972 14068
rect 6920 14025 6929 14059
rect 6929 14025 6963 14059
rect 6963 14025 6972 14059
rect 6920 14016 6972 14025
rect 7288 14016 7340 14068
rect 8024 14016 8076 14068
rect 2320 13948 2372 14000
rect 2412 13923 2464 13932
rect 2412 13889 2421 13923
rect 2421 13889 2455 13923
rect 2455 13889 2464 13923
rect 2412 13880 2464 13889
rect 2872 13880 2924 13932
rect 2780 13812 2832 13864
rect 3884 13948 3936 14000
rect 6092 13948 6144 14000
rect 9680 14016 9732 14068
rect 11612 14016 11664 14068
rect 12624 14016 12676 14068
rect 13176 14059 13228 14068
rect 13176 14025 13185 14059
rect 13185 14025 13219 14059
rect 13219 14025 13228 14059
rect 13176 14016 13228 14025
rect 13452 14059 13504 14068
rect 13452 14025 13461 14059
rect 13461 14025 13495 14059
rect 13495 14025 13504 14059
rect 13452 14016 13504 14025
rect 13820 14059 13872 14068
rect 13820 14025 13829 14059
rect 13829 14025 13863 14059
rect 13863 14025 13872 14059
rect 13820 14016 13872 14025
rect 15200 14016 15252 14068
rect 15384 14016 15436 14068
rect 15660 14059 15712 14068
rect 15660 14025 15669 14059
rect 15669 14025 15703 14059
rect 15703 14025 15712 14059
rect 15660 14016 15712 14025
rect 3976 13880 4028 13932
rect 5908 13880 5960 13932
rect 10600 13948 10652 14000
rect 12440 13948 12492 14000
rect 6920 13880 6972 13932
rect 7196 13880 7248 13932
rect 8300 13880 8352 13932
rect 9036 13880 9088 13932
rect 10232 13880 10284 13932
rect 11060 13880 11112 13932
rect 11520 13880 11572 13932
rect 14648 13880 14700 13932
rect 6460 13812 6512 13864
rect 11796 13855 11848 13864
rect 2320 13676 2372 13728
rect 4712 13744 4764 13796
rect 6184 13676 6236 13728
rect 8116 13744 8168 13796
rect 11796 13821 11805 13855
rect 11805 13821 11839 13855
rect 11839 13821 11848 13855
rect 11796 13812 11848 13821
rect 12900 13855 12952 13864
rect 12900 13821 12909 13855
rect 12909 13821 12943 13855
rect 12943 13821 12952 13855
rect 12900 13812 12952 13821
rect 13820 13812 13872 13864
rect 13912 13812 13964 13864
rect 11704 13744 11756 13796
rect 12072 13744 12124 13796
rect 13452 13744 13504 13796
rect 14004 13744 14056 13796
rect 15844 13812 15896 13864
rect 15108 13744 15160 13796
rect 11612 13676 11664 13728
rect 11980 13676 12032 13728
rect 13636 13676 13688 13728
rect 14096 13676 14148 13728
rect 14464 13676 14516 13728
rect 2824 13574 2876 13626
rect 2888 13574 2940 13626
rect 2952 13574 3004 13626
rect 3016 13574 3068 13626
rect 3080 13574 3132 13626
rect 6572 13574 6624 13626
rect 6636 13574 6688 13626
rect 6700 13574 6752 13626
rect 6764 13574 6816 13626
rect 6828 13574 6880 13626
rect 10320 13574 10372 13626
rect 10384 13574 10436 13626
rect 10448 13574 10500 13626
rect 10512 13574 10564 13626
rect 10576 13574 10628 13626
rect 14068 13574 14120 13626
rect 14132 13574 14184 13626
rect 14196 13574 14248 13626
rect 14260 13574 14312 13626
rect 14324 13574 14376 13626
rect 2228 13472 2280 13524
rect 4160 13515 4212 13524
rect 4160 13481 4169 13515
rect 4169 13481 4203 13515
rect 4203 13481 4212 13515
rect 4160 13472 4212 13481
rect 6184 13472 6236 13524
rect 9312 13472 9364 13524
rect 10140 13472 10192 13524
rect 10876 13472 10928 13524
rect 11612 13472 11664 13524
rect 3608 13336 3660 13388
rect 4160 13336 4212 13388
rect 4712 13336 4764 13388
rect 5724 13379 5776 13388
rect 5724 13345 5733 13379
rect 5733 13345 5767 13379
rect 5767 13345 5776 13379
rect 5724 13336 5776 13345
rect 1860 13268 1912 13320
rect 5448 13243 5500 13252
rect 5448 13209 5488 13243
rect 5488 13209 5500 13243
rect 9036 13311 9088 13320
rect 9036 13277 9045 13311
rect 9045 13277 9079 13311
rect 9079 13277 9088 13311
rect 9036 13268 9088 13277
rect 11796 13472 11848 13524
rect 12256 13472 12308 13524
rect 13544 13515 13596 13524
rect 13544 13481 13553 13515
rect 13553 13481 13587 13515
rect 13587 13481 13596 13515
rect 13544 13472 13596 13481
rect 13728 13515 13780 13524
rect 13728 13481 13737 13515
rect 13737 13481 13771 13515
rect 13771 13481 13780 13515
rect 13728 13472 13780 13481
rect 13820 13472 13872 13524
rect 14556 13515 14608 13524
rect 14556 13481 14565 13515
rect 14565 13481 14599 13515
rect 14599 13481 14608 13515
rect 14556 13472 14608 13481
rect 14648 13515 14700 13524
rect 14648 13481 14657 13515
rect 14657 13481 14691 13515
rect 14691 13481 14700 13515
rect 14648 13472 14700 13481
rect 15200 13472 15252 13524
rect 11980 13404 12032 13456
rect 12992 13404 13044 13456
rect 13176 13404 13228 13456
rect 15108 13404 15160 13456
rect 15568 13404 15620 13456
rect 11796 13336 11848 13388
rect 12072 13336 12124 13388
rect 12808 13336 12860 13388
rect 14556 13336 14608 13388
rect 5448 13200 5500 13209
rect 6092 13243 6144 13252
rect 6092 13209 6126 13243
rect 6126 13209 6144 13243
rect 6092 13200 6144 13209
rect 6368 13200 6420 13252
rect 1492 13175 1544 13184
rect 1492 13141 1501 13175
rect 1501 13141 1535 13175
rect 1535 13141 1544 13175
rect 1492 13132 1544 13141
rect 4252 13132 4304 13184
rect 5080 13132 5132 13184
rect 5908 13132 5960 13184
rect 6184 13132 6236 13184
rect 7288 13132 7340 13184
rect 8944 13132 8996 13184
rect 9680 13200 9732 13252
rect 10784 13200 10836 13252
rect 12256 13243 12308 13252
rect 12256 13209 12265 13243
rect 12265 13209 12299 13243
rect 12299 13209 12308 13243
rect 12256 13200 12308 13209
rect 13268 13200 13320 13252
rect 11060 13175 11112 13184
rect 11060 13141 11069 13175
rect 11069 13141 11103 13175
rect 11103 13141 11112 13175
rect 11060 13132 11112 13141
rect 11428 13175 11480 13184
rect 11428 13141 11437 13175
rect 11437 13141 11471 13175
rect 11471 13141 11480 13175
rect 11428 13132 11480 13141
rect 11612 13132 11664 13184
rect 13820 13200 13872 13252
rect 15200 13200 15252 13252
rect 13452 13132 13504 13184
rect 14004 13132 14056 13184
rect 14280 13175 14332 13184
rect 14280 13141 14289 13175
rect 14289 13141 14323 13175
rect 14323 13141 14332 13175
rect 14280 13132 14332 13141
rect 15292 13132 15344 13184
rect 15752 13132 15804 13184
rect 4698 13030 4750 13082
rect 4762 13030 4814 13082
rect 4826 13030 4878 13082
rect 4890 13030 4942 13082
rect 4954 13030 5006 13082
rect 8446 13030 8498 13082
rect 8510 13030 8562 13082
rect 8574 13030 8626 13082
rect 8638 13030 8690 13082
rect 8702 13030 8754 13082
rect 12194 13030 12246 13082
rect 12258 13030 12310 13082
rect 12322 13030 12374 13082
rect 12386 13030 12438 13082
rect 12450 13030 12502 13082
rect 1584 12792 1636 12844
rect 1952 12835 2004 12844
rect 1952 12801 1961 12835
rect 1961 12801 1995 12835
rect 1995 12801 2004 12835
rect 1952 12792 2004 12801
rect 3148 12928 3200 12980
rect 5632 12928 5684 12980
rect 6092 12928 6144 12980
rect 6920 12928 6972 12980
rect 5080 12860 5132 12912
rect 5264 12792 5316 12844
rect 5724 12792 5776 12844
rect 4436 12724 4488 12776
rect 9036 12928 9088 12980
rect 9680 12928 9732 12980
rect 10784 12928 10836 12980
rect 13084 12928 13136 12980
rect 13728 12971 13780 12980
rect 13728 12937 13737 12971
rect 13737 12937 13771 12971
rect 13771 12937 13780 12971
rect 13728 12928 13780 12937
rect 13820 12928 13872 12980
rect 14464 12928 14516 12980
rect 14832 12928 14884 12980
rect 15016 12928 15068 12980
rect 9220 12860 9272 12912
rect 10784 12792 10836 12844
rect 8300 12724 8352 12776
rect 9220 12724 9272 12776
rect 1492 12631 1544 12640
rect 1492 12597 1501 12631
rect 1501 12597 1535 12631
rect 1535 12597 1544 12631
rect 1492 12588 1544 12597
rect 1676 12588 1728 12640
rect 3792 12588 3844 12640
rect 4252 12631 4304 12640
rect 4252 12597 4261 12631
rect 4261 12597 4295 12631
rect 4295 12597 4304 12631
rect 4252 12588 4304 12597
rect 6920 12656 6972 12708
rect 9680 12724 9732 12776
rect 11060 12860 11112 12912
rect 11520 12860 11572 12912
rect 11796 12860 11848 12912
rect 13268 12860 13320 12912
rect 13452 12860 13504 12912
rect 13176 12792 13228 12844
rect 15660 12860 15712 12912
rect 8668 12631 8720 12640
rect 8668 12597 8677 12631
rect 8677 12597 8711 12631
rect 8711 12597 8720 12631
rect 8668 12588 8720 12597
rect 9680 12588 9732 12640
rect 10692 12588 10744 12640
rect 13360 12724 13412 12776
rect 13544 12724 13596 12776
rect 14004 12767 14056 12776
rect 14004 12733 14013 12767
rect 14013 12733 14047 12767
rect 14047 12733 14056 12767
rect 14004 12724 14056 12733
rect 14648 12724 14700 12776
rect 15660 12724 15712 12776
rect 16120 12724 16172 12776
rect 11244 12656 11296 12708
rect 14832 12656 14884 12708
rect 13268 12631 13320 12640
rect 13268 12597 13277 12631
rect 13277 12597 13311 12631
rect 13311 12597 13320 12631
rect 13268 12588 13320 12597
rect 15200 12588 15252 12640
rect 15568 12588 15620 12640
rect 2824 12486 2876 12538
rect 2888 12486 2940 12538
rect 2952 12486 3004 12538
rect 3016 12486 3068 12538
rect 3080 12486 3132 12538
rect 6572 12486 6624 12538
rect 6636 12486 6688 12538
rect 6700 12486 6752 12538
rect 6764 12486 6816 12538
rect 6828 12486 6880 12538
rect 10320 12486 10372 12538
rect 10384 12486 10436 12538
rect 10448 12486 10500 12538
rect 10512 12486 10564 12538
rect 10576 12486 10628 12538
rect 14068 12486 14120 12538
rect 14132 12486 14184 12538
rect 14196 12486 14248 12538
rect 14260 12486 14312 12538
rect 14324 12486 14376 12538
rect 1952 12384 2004 12436
rect 2596 12384 2648 12436
rect 3148 12384 3200 12436
rect 3240 12384 3292 12436
rect 3424 12384 3476 12436
rect 4528 12384 4580 12436
rect 3884 12316 3936 12368
rect 1768 12223 1820 12232
rect 1768 12189 1777 12223
rect 1777 12189 1811 12223
rect 1811 12189 1820 12223
rect 1768 12180 1820 12189
rect 4344 12316 4396 12368
rect 6920 12384 6972 12436
rect 7196 12384 7248 12436
rect 7288 12384 7340 12436
rect 7564 12384 7616 12436
rect 9220 12384 9272 12436
rect 10048 12384 10100 12436
rect 12992 12384 13044 12436
rect 13636 12384 13688 12436
rect 13912 12384 13964 12436
rect 9036 12316 9088 12368
rect 9496 12316 9548 12368
rect 14188 12316 14240 12368
rect 9956 12248 10008 12300
rect 10876 12248 10928 12300
rect 12624 12291 12676 12300
rect 12624 12257 12633 12291
rect 12633 12257 12667 12291
rect 12667 12257 12676 12291
rect 12624 12248 12676 12257
rect 1860 12112 1912 12164
rect 5724 12180 5776 12232
rect 8668 12180 8720 12232
rect 13360 12248 13412 12300
rect 14556 12316 14608 12368
rect 14648 12291 14700 12300
rect 14648 12257 14657 12291
rect 14657 12257 14691 12291
rect 14691 12257 14700 12291
rect 14648 12248 14700 12257
rect 13912 12180 13964 12232
rect 14740 12180 14792 12232
rect 15660 12180 15712 12232
rect 5448 12112 5500 12164
rect 5816 12112 5868 12164
rect 9496 12112 9548 12164
rect 12072 12112 12124 12164
rect 12624 12112 12676 12164
rect 13820 12112 13872 12164
rect 2136 12044 2188 12096
rect 3976 12044 4028 12096
rect 4436 12087 4488 12096
rect 4436 12053 4445 12087
rect 4445 12053 4479 12087
rect 4479 12053 4488 12087
rect 4436 12044 4488 12053
rect 5540 12044 5592 12096
rect 11244 12044 11296 12096
rect 14464 12087 14516 12096
rect 14464 12053 14473 12087
rect 14473 12053 14507 12087
rect 14507 12053 14516 12087
rect 14464 12044 14516 12053
rect 15660 12087 15712 12096
rect 15660 12053 15669 12087
rect 15669 12053 15703 12087
rect 15703 12053 15712 12087
rect 15660 12044 15712 12053
rect 4698 11942 4750 11994
rect 4762 11942 4814 11994
rect 4826 11942 4878 11994
rect 4890 11942 4942 11994
rect 4954 11942 5006 11994
rect 8446 11942 8498 11994
rect 8510 11942 8562 11994
rect 8574 11942 8626 11994
rect 8638 11942 8690 11994
rect 8702 11942 8754 11994
rect 12194 11942 12246 11994
rect 12258 11942 12310 11994
rect 12322 11942 12374 11994
rect 12386 11942 12438 11994
rect 12450 11942 12502 11994
rect 5724 11840 5776 11892
rect 1676 11747 1728 11756
rect 1676 11713 1685 11747
rect 1685 11713 1719 11747
rect 1719 11713 1728 11747
rect 1676 11704 1728 11713
rect 5264 11704 5316 11756
rect 2596 11636 2648 11688
rect 3884 11636 3936 11688
rect 7012 11840 7064 11892
rect 9680 11840 9732 11892
rect 10324 11840 10376 11892
rect 11520 11883 11572 11892
rect 9220 11772 9272 11824
rect 9864 11772 9916 11824
rect 10508 11772 10560 11824
rect 11520 11849 11529 11883
rect 11529 11849 11563 11883
rect 11563 11849 11572 11883
rect 11520 11840 11572 11849
rect 11980 11883 12032 11892
rect 11980 11849 11989 11883
rect 11989 11849 12023 11883
rect 12023 11849 12032 11883
rect 11980 11840 12032 11849
rect 14188 11883 14240 11892
rect 14188 11849 14197 11883
rect 14197 11849 14231 11883
rect 14231 11849 14240 11883
rect 14188 11840 14240 11849
rect 15476 11883 15528 11892
rect 15476 11849 15485 11883
rect 15485 11849 15519 11883
rect 15519 11849 15528 11883
rect 15476 11840 15528 11849
rect 16028 11840 16080 11892
rect 10876 11772 10928 11824
rect 6368 11747 6420 11756
rect 6368 11713 6377 11747
rect 6377 11713 6411 11747
rect 6411 11713 6420 11747
rect 6368 11704 6420 11713
rect 7472 11704 7524 11756
rect 11336 11772 11388 11824
rect 12256 11772 12308 11824
rect 9496 11636 9548 11688
rect 11980 11704 12032 11756
rect 13268 11772 13320 11824
rect 12992 11704 13044 11756
rect 14648 11704 14700 11756
rect 12348 11679 12400 11688
rect 12348 11645 12357 11679
rect 12357 11645 12391 11679
rect 12391 11645 12400 11679
rect 12348 11636 12400 11645
rect 1492 11543 1544 11552
rect 1492 11509 1501 11543
rect 1501 11509 1535 11543
rect 1535 11509 1544 11543
rect 1492 11500 1544 11509
rect 4160 11500 4212 11552
rect 4620 11500 4672 11552
rect 5632 11543 5684 11552
rect 5632 11509 5641 11543
rect 5641 11509 5675 11543
rect 5675 11509 5684 11543
rect 5632 11500 5684 11509
rect 7840 11568 7892 11620
rect 11520 11568 11572 11620
rect 7288 11500 7340 11552
rect 7564 11500 7616 11552
rect 10784 11500 10836 11552
rect 12072 11500 12124 11552
rect 14740 11679 14792 11688
rect 14740 11645 14749 11679
rect 14749 11645 14783 11679
rect 14783 11645 14792 11679
rect 14740 11636 14792 11645
rect 13636 11500 13688 11552
rect 15292 11543 15344 11552
rect 15292 11509 15301 11543
rect 15301 11509 15335 11543
rect 15335 11509 15344 11543
rect 15292 11500 15344 11509
rect 2824 11398 2876 11450
rect 2888 11398 2940 11450
rect 2952 11398 3004 11450
rect 3016 11398 3068 11450
rect 3080 11398 3132 11450
rect 6572 11398 6624 11450
rect 6636 11398 6688 11450
rect 6700 11398 6752 11450
rect 6764 11398 6816 11450
rect 6828 11398 6880 11450
rect 10320 11398 10372 11450
rect 10384 11398 10436 11450
rect 10448 11398 10500 11450
rect 10512 11398 10564 11450
rect 10576 11398 10628 11450
rect 14068 11398 14120 11450
rect 14132 11398 14184 11450
rect 14196 11398 14248 11450
rect 14260 11398 14312 11450
rect 14324 11398 14376 11450
rect 1584 11296 1636 11348
rect 2504 11296 2556 11348
rect 3884 11296 3936 11348
rect 5540 11228 5592 11280
rect 10324 11296 10376 11348
rect 11428 11296 11480 11348
rect 11888 11296 11940 11348
rect 13544 11296 13596 11348
rect 9220 11271 9272 11280
rect 3240 11092 3292 11144
rect 4712 11092 4764 11144
rect 7012 11092 7064 11144
rect 7380 11135 7432 11144
rect 7380 11101 7389 11135
rect 7389 11101 7423 11135
rect 7423 11101 7432 11135
rect 9220 11237 9229 11271
rect 9229 11237 9263 11271
rect 9263 11237 9272 11271
rect 9220 11228 9272 11237
rect 12256 11228 12308 11280
rect 10692 11203 10744 11212
rect 10692 11169 10701 11203
rect 10701 11169 10735 11203
rect 10735 11169 10744 11203
rect 10692 11160 10744 11169
rect 11888 11203 11940 11212
rect 11888 11169 11897 11203
rect 11897 11169 11931 11203
rect 11931 11169 11940 11203
rect 11888 11160 11940 11169
rect 12072 11160 12124 11212
rect 7380 11092 7432 11101
rect 12348 11092 12400 11144
rect 13360 11228 13412 11280
rect 13636 11203 13688 11212
rect 13636 11169 13645 11203
rect 13645 11169 13679 11203
rect 13679 11169 13688 11203
rect 13636 11160 13688 11169
rect 13912 11160 13964 11212
rect 15752 11160 15804 11212
rect 14372 11135 14424 11144
rect 14372 11101 14381 11135
rect 14381 11101 14415 11135
rect 14415 11101 14424 11135
rect 14372 11092 14424 11101
rect 14648 11092 14700 11144
rect 7656 11067 7708 11076
rect 7656 11033 7690 11067
rect 7690 11033 7708 11067
rect 7656 11024 7708 11033
rect 7840 11024 7892 11076
rect 1400 10956 1452 11008
rect 2872 10956 2924 11008
rect 5264 10956 5316 11008
rect 9220 10956 9272 11008
rect 10784 11024 10836 11076
rect 11428 11024 11480 11076
rect 15752 11024 15804 11076
rect 10232 10956 10284 11008
rect 14924 10956 14976 11008
rect 15844 10956 15896 11008
rect 4698 10854 4750 10906
rect 4762 10854 4814 10906
rect 4826 10854 4878 10906
rect 4890 10854 4942 10906
rect 4954 10854 5006 10906
rect 8446 10854 8498 10906
rect 8510 10854 8562 10906
rect 8574 10854 8626 10906
rect 8638 10854 8690 10906
rect 8702 10854 8754 10906
rect 12194 10854 12246 10906
rect 12258 10854 12310 10906
rect 12322 10854 12374 10906
rect 12386 10854 12438 10906
rect 12450 10854 12502 10906
rect 3148 10795 3200 10804
rect 3148 10761 3157 10795
rect 3157 10761 3191 10795
rect 3191 10761 3200 10795
rect 3148 10752 3200 10761
rect 3700 10752 3752 10804
rect 3884 10752 3936 10804
rect 6368 10752 6420 10804
rect 5632 10684 5684 10736
rect 2044 10616 2096 10668
rect 3884 10659 3936 10668
rect 2136 10523 2188 10532
rect 2136 10489 2145 10523
rect 2145 10489 2179 10523
rect 2179 10489 2188 10523
rect 2136 10480 2188 10489
rect 3884 10625 3893 10659
rect 3893 10625 3927 10659
rect 3927 10625 3936 10659
rect 3884 10616 3936 10625
rect 4160 10659 4212 10668
rect 4160 10625 4194 10659
rect 4194 10625 4212 10659
rect 7380 10752 7432 10804
rect 13268 10752 13320 10804
rect 15292 10752 15344 10804
rect 4160 10616 4212 10625
rect 2872 10591 2924 10600
rect 2872 10557 2881 10591
rect 2881 10557 2915 10591
rect 2915 10557 2924 10591
rect 2872 10548 2924 10557
rect 5724 10548 5776 10600
rect 6000 10548 6052 10600
rect 9864 10684 9916 10736
rect 14464 10727 14516 10736
rect 7748 10616 7800 10668
rect 9220 10616 9272 10668
rect 13360 10659 13412 10668
rect 13360 10625 13369 10659
rect 13369 10625 13403 10659
rect 13403 10625 13412 10659
rect 13360 10616 13412 10625
rect 12900 10591 12952 10600
rect 12900 10557 12909 10591
rect 12909 10557 12943 10591
rect 12943 10557 12952 10591
rect 12900 10548 12952 10557
rect 14464 10693 14473 10727
rect 14473 10693 14507 10727
rect 14507 10693 14516 10727
rect 14464 10684 14516 10693
rect 15016 10684 15068 10736
rect 14832 10616 14884 10668
rect 13912 10548 13964 10600
rect 14924 10548 14976 10600
rect 12992 10523 13044 10532
rect 3148 10412 3200 10464
rect 4160 10412 4212 10464
rect 8208 10412 8260 10464
rect 9496 10412 9548 10464
rect 12992 10489 13001 10523
rect 13001 10489 13035 10523
rect 13035 10489 13044 10523
rect 12992 10480 13044 10489
rect 13728 10480 13780 10532
rect 14648 10480 14700 10532
rect 11152 10412 11204 10464
rect 11704 10412 11756 10464
rect 13268 10412 13320 10464
rect 13544 10412 13596 10464
rect 14740 10412 14792 10464
rect 15476 10412 15528 10464
rect 2824 10310 2876 10362
rect 2888 10310 2940 10362
rect 2952 10310 3004 10362
rect 3016 10310 3068 10362
rect 3080 10310 3132 10362
rect 6572 10310 6624 10362
rect 6636 10310 6688 10362
rect 6700 10310 6752 10362
rect 6764 10310 6816 10362
rect 6828 10310 6880 10362
rect 10320 10310 10372 10362
rect 10384 10310 10436 10362
rect 10448 10310 10500 10362
rect 10512 10310 10564 10362
rect 10576 10310 10628 10362
rect 14068 10310 14120 10362
rect 14132 10310 14184 10362
rect 14196 10310 14248 10362
rect 14260 10310 14312 10362
rect 14324 10310 14376 10362
rect 1492 10251 1544 10260
rect 1492 10217 1501 10251
rect 1501 10217 1535 10251
rect 1535 10217 1544 10251
rect 1492 10208 1544 10217
rect 7656 10208 7708 10260
rect 7472 10140 7524 10192
rect 10968 10208 11020 10260
rect 12624 10208 12676 10260
rect 12992 10208 13044 10260
rect 13360 10208 13412 10260
rect 14648 10208 14700 10260
rect 14924 10251 14976 10260
rect 14924 10217 14933 10251
rect 14933 10217 14967 10251
rect 14967 10217 14976 10251
rect 14924 10208 14976 10217
rect 10692 10072 10744 10124
rect 12072 10072 12124 10124
rect 12716 10115 12768 10124
rect 12716 10081 12725 10115
rect 12725 10081 12759 10115
rect 12759 10081 12768 10115
rect 12716 10072 12768 10081
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 5448 9936 5500 9988
rect 5724 9936 5776 9988
rect 8852 10004 8904 10056
rect 9772 10004 9824 10056
rect 7932 9936 7984 9988
rect 11244 9936 11296 9988
rect 11704 9979 11756 9988
rect 11704 9945 11722 9979
rect 11722 9945 11756 9979
rect 11704 9936 11756 9945
rect 2228 9868 2280 9920
rect 11152 9868 11204 9920
rect 12624 10004 12676 10056
rect 13268 10072 13320 10124
rect 13820 10115 13872 10124
rect 13820 10081 13829 10115
rect 13829 10081 13863 10115
rect 13863 10081 13872 10115
rect 13820 10072 13872 10081
rect 14004 10072 14056 10124
rect 14556 10072 14608 10124
rect 14648 10072 14700 10124
rect 15384 10115 15436 10124
rect 15384 10081 15393 10115
rect 15393 10081 15427 10115
rect 15427 10081 15436 10115
rect 15384 10072 15436 10081
rect 15476 10115 15528 10124
rect 15476 10081 15485 10115
rect 15485 10081 15519 10115
rect 15519 10081 15528 10115
rect 15476 10072 15528 10081
rect 15660 10004 15712 10056
rect 13820 9936 13872 9988
rect 13452 9868 13504 9920
rect 13636 9911 13688 9920
rect 13636 9877 13645 9911
rect 13645 9877 13679 9911
rect 13679 9877 13688 9911
rect 13636 9868 13688 9877
rect 14464 9911 14516 9920
rect 14464 9877 14473 9911
rect 14473 9877 14507 9911
rect 14507 9877 14516 9911
rect 14464 9868 14516 9877
rect 4698 9766 4750 9818
rect 4762 9766 4814 9818
rect 4826 9766 4878 9818
rect 4890 9766 4942 9818
rect 4954 9766 5006 9818
rect 8446 9766 8498 9818
rect 8510 9766 8562 9818
rect 8574 9766 8626 9818
rect 8638 9766 8690 9818
rect 8702 9766 8754 9818
rect 12194 9766 12246 9818
rect 12258 9766 12310 9818
rect 12322 9766 12374 9818
rect 12386 9766 12438 9818
rect 12450 9766 12502 9818
rect 1676 9664 1728 9716
rect 2320 9664 2372 9716
rect 5724 9664 5776 9716
rect 7564 9664 7616 9716
rect 5448 9596 5500 9648
rect 1768 9528 1820 9580
rect 2136 9528 2188 9580
rect 3976 9528 4028 9580
rect 5356 9528 5408 9580
rect 9496 9664 9548 9716
rect 10692 9707 10744 9716
rect 7472 9571 7524 9580
rect 7472 9537 7490 9571
rect 7490 9537 7524 9571
rect 7472 9528 7524 9537
rect 8668 9596 8720 9648
rect 8852 9596 8904 9648
rect 9864 9596 9916 9648
rect 10692 9673 10701 9707
rect 10701 9673 10735 9707
rect 10735 9673 10744 9707
rect 10692 9664 10744 9673
rect 11704 9664 11756 9716
rect 12624 9664 12676 9716
rect 12900 9664 12952 9716
rect 14464 9664 14516 9716
rect 7840 9528 7892 9580
rect 1492 9435 1544 9444
rect 1492 9401 1501 9435
rect 1501 9401 1535 9435
rect 1535 9401 1544 9435
rect 1492 9392 1544 9401
rect 4344 9435 4396 9444
rect 4344 9401 4353 9435
rect 4353 9401 4387 9435
rect 4387 9401 4396 9435
rect 4344 9392 4396 9401
rect 3148 9324 3200 9376
rect 3976 9324 4028 9376
rect 5540 9324 5592 9376
rect 8852 9460 8904 9512
rect 11796 9596 11848 9648
rect 12624 9528 12676 9580
rect 12808 9528 12860 9580
rect 11612 9435 11664 9444
rect 9128 9367 9180 9376
rect 9128 9333 9137 9367
rect 9137 9333 9171 9367
rect 9171 9333 9180 9367
rect 9128 9324 9180 9333
rect 11612 9401 11621 9435
rect 11621 9401 11655 9435
rect 11655 9401 11664 9435
rect 11612 9392 11664 9401
rect 12164 9503 12216 9512
rect 12164 9469 12173 9503
rect 12173 9469 12207 9503
rect 12207 9469 12216 9503
rect 12164 9460 12216 9469
rect 13084 9460 13136 9512
rect 13176 9460 13228 9512
rect 13636 9596 13688 9648
rect 15292 9596 15344 9648
rect 13912 9528 13964 9580
rect 14464 9528 14516 9580
rect 15568 9528 15620 9580
rect 15476 9503 15528 9512
rect 15476 9469 15485 9503
rect 15485 9469 15519 9503
rect 15519 9469 15528 9503
rect 15476 9460 15528 9469
rect 12808 9435 12860 9444
rect 12808 9401 12817 9435
rect 12817 9401 12851 9435
rect 12851 9401 12860 9435
rect 12808 9392 12860 9401
rect 11796 9324 11848 9376
rect 12624 9367 12676 9376
rect 12624 9333 12633 9367
rect 12633 9333 12667 9367
rect 12667 9333 12676 9367
rect 12624 9324 12676 9333
rect 13636 9367 13688 9376
rect 13636 9333 13645 9367
rect 13645 9333 13679 9367
rect 13679 9333 13688 9367
rect 13636 9324 13688 9333
rect 15476 9324 15528 9376
rect 2824 9222 2876 9274
rect 2888 9222 2940 9274
rect 2952 9222 3004 9274
rect 3016 9222 3068 9274
rect 3080 9222 3132 9274
rect 6572 9222 6624 9274
rect 6636 9222 6688 9274
rect 6700 9222 6752 9274
rect 6764 9222 6816 9274
rect 6828 9222 6880 9274
rect 10320 9222 10372 9274
rect 10384 9222 10436 9274
rect 10448 9222 10500 9274
rect 10512 9222 10564 9274
rect 10576 9222 10628 9274
rect 14068 9222 14120 9274
rect 14132 9222 14184 9274
rect 14196 9222 14248 9274
rect 14260 9222 14312 9274
rect 14324 9222 14376 9274
rect 1768 9163 1820 9172
rect 1768 9129 1777 9163
rect 1777 9129 1811 9163
rect 1811 9129 1820 9163
rect 1768 9120 1820 9129
rect 3148 9120 3200 9172
rect 3516 9052 3568 9104
rect 3792 9052 3844 9104
rect 7380 9120 7432 9172
rect 8852 9120 8904 9172
rect 9312 9120 9364 9172
rect 9588 9120 9640 9172
rect 15200 9120 15252 9172
rect 5356 9052 5408 9104
rect 7472 9052 7524 9104
rect 5448 9027 5500 9036
rect 1768 8916 1820 8968
rect 1952 8959 2004 8968
rect 1952 8925 1961 8959
rect 1961 8925 1995 8959
rect 1995 8925 2004 8959
rect 1952 8916 2004 8925
rect 2044 8848 2096 8900
rect 2228 8848 2280 8900
rect 1492 8823 1544 8832
rect 1492 8789 1501 8823
rect 1501 8789 1535 8823
rect 1535 8789 1544 8823
rect 1492 8780 1544 8789
rect 2320 8780 2372 8832
rect 3976 8916 4028 8968
rect 5448 8993 5457 9027
rect 5457 8993 5491 9027
rect 5491 8993 5500 9027
rect 5448 8984 5500 8993
rect 9036 9052 9088 9104
rect 9496 9052 9548 9104
rect 11612 9052 11664 9104
rect 11888 9052 11940 9104
rect 12164 9052 12216 9104
rect 12532 9095 12584 9104
rect 12532 9061 12541 9095
rect 12541 9061 12575 9095
rect 12575 9061 12584 9095
rect 12532 9052 12584 9061
rect 13084 9052 13136 9104
rect 14924 9095 14976 9104
rect 11980 8984 12032 9036
rect 14924 9061 14933 9095
rect 14933 9061 14967 9095
rect 14967 9061 14976 9095
rect 14924 9052 14976 9061
rect 15108 9052 15160 9104
rect 14740 8984 14792 9036
rect 15292 9027 15344 9036
rect 15292 8993 15301 9027
rect 15301 8993 15335 9027
rect 15335 8993 15344 9027
rect 15292 8984 15344 8993
rect 9036 8916 9088 8968
rect 10692 8916 10744 8968
rect 13268 8959 13320 8968
rect 13268 8925 13277 8959
rect 13277 8925 13311 8959
rect 13311 8925 13320 8959
rect 13268 8916 13320 8925
rect 14556 8916 14608 8968
rect 15108 8916 15160 8968
rect 15476 8916 15528 8968
rect 3700 8848 3752 8900
rect 3792 8780 3844 8832
rect 4344 8848 4396 8900
rect 6092 8848 6144 8900
rect 6460 8848 6512 8900
rect 8300 8848 8352 8900
rect 9220 8848 9272 8900
rect 10324 8848 10376 8900
rect 11336 8848 11388 8900
rect 10692 8780 10744 8832
rect 12072 8780 12124 8832
rect 12992 8848 13044 8900
rect 14280 8848 14332 8900
rect 16396 8848 16448 8900
rect 12532 8780 12584 8832
rect 12900 8823 12952 8832
rect 12900 8789 12909 8823
rect 12909 8789 12943 8823
rect 12943 8789 12952 8823
rect 12900 8780 12952 8789
rect 13176 8780 13228 8832
rect 13636 8780 13688 8832
rect 14096 8823 14148 8832
rect 14096 8789 14105 8823
rect 14105 8789 14139 8823
rect 14139 8789 14148 8823
rect 14096 8780 14148 8789
rect 14464 8823 14516 8832
rect 14464 8789 14473 8823
rect 14473 8789 14507 8823
rect 14507 8789 14516 8823
rect 14464 8780 14516 8789
rect 4698 8678 4750 8730
rect 4762 8678 4814 8730
rect 4826 8678 4878 8730
rect 4890 8678 4942 8730
rect 4954 8678 5006 8730
rect 8446 8678 8498 8730
rect 8510 8678 8562 8730
rect 8574 8678 8626 8730
rect 8638 8678 8690 8730
rect 8702 8678 8754 8730
rect 12194 8678 12246 8730
rect 12258 8678 12310 8730
rect 12322 8678 12374 8730
rect 12386 8678 12438 8730
rect 12450 8678 12502 8730
rect 1860 8619 1912 8628
rect 1860 8585 1869 8619
rect 1869 8585 1903 8619
rect 1903 8585 1912 8619
rect 1860 8576 1912 8585
rect 1952 8576 2004 8628
rect 5264 8576 5316 8628
rect 6736 8508 6788 8560
rect 7932 8576 7984 8628
rect 9036 8619 9088 8628
rect 9036 8585 9045 8619
rect 9045 8585 9079 8619
rect 9079 8585 9088 8619
rect 9036 8576 9088 8585
rect 9680 8576 9732 8628
rect 10324 8576 10376 8628
rect 10876 8576 10928 8628
rect 13544 8619 13596 8628
rect 3700 8483 3752 8492
rect 3700 8449 3718 8483
rect 3718 8449 3752 8483
rect 3976 8483 4028 8492
rect 3700 8440 3752 8449
rect 3976 8449 3985 8483
rect 3985 8449 4019 8483
rect 4019 8449 4028 8483
rect 3976 8440 4028 8449
rect 4620 8440 4672 8492
rect 2412 8236 2464 8288
rect 5540 8304 5592 8356
rect 5356 8236 5408 8288
rect 7656 8236 7708 8288
rect 9128 8508 9180 8560
rect 11612 8508 11664 8560
rect 11704 8508 11756 8560
rect 7932 8372 7984 8424
rect 11060 8440 11112 8492
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 11704 8372 11756 8424
rect 11980 8415 12032 8424
rect 11980 8381 11989 8415
rect 11989 8381 12023 8415
rect 12023 8381 12032 8415
rect 11980 8372 12032 8381
rect 13544 8585 13553 8619
rect 13553 8585 13587 8619
rect 13587 8585 13596 8619
rect 13544 8576 13596 8585
rect 13912 8576 13964 8628
rect 12808 8508 12860 8560
rect 13452 8508 13504 8560
rect 14280 8508 14332 8560
rect 14648 8508 14700 8560
rect 14924 8576 14976 8628
rect 15108 8508 15160 8560
rect 12808 8415 12860 8424
rect 10600 8304 10652 8356
rect 11888 8304 11940 8356
rect 12348 8347 12400 8356
rect 12348 8313 12357 8347
rect 12357 8313 12391 8347
rect 12391 8313 12400 8347
rect 12348 8304 12400 8313
rect 12808 8381 12817 8415
rect 12817 8381 12851 8415
rect 12851 8381 12860 8415
rect 12808 8372 12860 8381
rect 14188 8440 14240 8492
rect 14464 8440 14516 8492
rect 14924 8440 14976 8492
rect 13636 8372 13688 8424
rect 15108 8415 15160 8424
rect 15108 8381 15117 8415
rect 15117 8381 15151 8415
rect 15151 8381 15160 8415
rect 15108 8372 15160 8381
rect 15660 8304 15712 8356
rect 9404 8236 9456 8288
rect 11336 8236 11388 8288
rect 13820 8236 13872 8288
rect 14372 8236 14424 8288
rect 14648 8236 14700 8288
rect 2824 8134 2876 8186
rect 2888 8134 2940 8186
rect 2952 8134 3004 8186
rect 3016 8134 3068 8186
rect 3080 8134 3132 8186
rect 6572 8134 6624 8186
rect 6636 8134 6688 8186
rect 6700 8134 6752 8186
rect 6764 8134 6816 8186
rect 6828 8134 6880 8186
rect 10320 8134 10372 8186
rect 10384 8134 10436 8186
rect 10448 8134 10500 8186
rect 10512 8134 10564 8186
rect 10576 8134 10628 8186
rect 14068 8134 14120 8186
rect 14132 8134 14184 8186
rect 14196 8134 14248 8186
rect 14260 8134 14312 8186
rect 14324 8134 14376 8186
rect 2136 8075 2188 8084
rect 2136 8041 2145 8075
rect 2145 8041 2179 8075
rect 2179 8041 2188 8075
rect 2136 8032 2188 8041
rect 3884 7964 3936 8016
rect 2495 7871 2547 7880
rect 2495 7837 2504 7871
rect 2504 7837 2538 7871
rect 2538 7837 2547 7871
rect 2495 7828 2547 7837
rect 9036 8032 9088 8084
rect 9220 8075 9272 8084
rect 9220 8041 9229 8075
rect 9229 8041 9263 8075
rect 9263 8041 9272 8075
rect 9220 8032 9272 8041
rect 9680 7964 9732 8016
rect 4620 7871 4672 7880
rect 4620 7837 4629 7871
rect 4629 7837 4663 7871
rect 4663 7837 4672 7871
rect 4620 7828 4672 7837
rect 7656 7939 7708 7948
rect 7656 7905 7665 7939
rect 7665 7905 7699 7939
rect 7699 7905 7708 7939
rect 7656 7896 7708 7905
rect 9036 7896 9088 7948
rect 12716 8032 12768 8084
rect 14464 8032 14516 8084
rect 14740 8032 14792 8084
rect 11336 7964 11388 8016
rect 12072 8007 12124 8016
rect 12072 7973 12081 8007
rect 12081 7973 12115 8007
rect 12115 7973 12124 8007
rect 12072 7964 12124 7973
rect 13820 7964 13872 8016
rect 7748 7828 7800 7880
rect 1676 7735 1728 7744
rect 1676 7701 1685 7735
rect 1685 7701 1719 7735
rect 1719 7701 1728 7735
rect 1676 7692 1728 7701
rect 5356 7760 5408 7812
rect 6276 7692 6328 7744
rect 7380 7803 7432 7812
rect 7380 7769 7398 7803
rect 7398 7769 7432 7803
rect 7380 7760 7432 7769
rect 8300 7692 8352 7744
rect 8852 7692 8904 7744
rect 10140 7828 10192 7880
rect 10968 7828 11020 7880
rect 11796 7896 11848 7948
rect 12164 7939 12216 7948
rect 12164 7905 12173 7939
rect 12173 7905 12207 7939
rect 12207 7905 12216 7939
rect 12164 7896 12216 7905
rect 12900 7896 12952 7948
rect 13176 7939 13228 7948
rect 13176 7905 13185 7939
rect 13185 7905 13219 7939
rect 13219 7905 13228 7939
rect 13176 7896 13228 7905
rect 13544 7896 13596 7948
rect 13912 7896 13964 7948
rect 14556 7896 14608 7948
rect 11520 7828 11572 7880
rect 14096 7828 14148 7880
rect 14372 7828 14424 7880
rect 15108 7871 15160 7880
rect 10416 7760 10468 7812
rect 10692 7760 10744 7812
rect 10876 7760 10928 7812
rect 15108 7837 15117 7871
rect 15117 7837 15151 7871
rect 15151 7837 15160 7871
rect 15108 7828 15160 7837
rect 9588 7692 9640 7744
rect 11428 7735 11480 7744
rect 11428 7701 11437 7735
rect 11437 7701 11471 7735
rect 11471 7701 11480 7735
rect 11428 7692 11480 7701
rect 11612 7692 11664 7744
rect 12532 7692 12584 7744
rect 13452 7735 13504 7744
rect 13452 7701 13461 7735
rect 13461 7701 13495 7735
rect 13495 7701 13504 7735
rect 13452 7692 13504 7701
rect 13912 7692 13964 7744
rect 14372 7692 14424 7744
rect 4698 7590 4750 7642
rect 4762 7590 4814 7642
rect 4826 7590 4878 7642
rect 4890 7590 4942 7642
rect 4954 7590 5006 7642
rect 8446 7590 8498 7642
rect 8510 7590 8562 7642
rect 8574 7590 8626 7642
rect 8638 7590 8690 7642
rect 8702 7590 8754 7642
rect 12194 7590 12246 7642
rect 12258 7590 12310 7642
rect 12322 7590 12374 7642
rect 12386 7590 12438 7642
rect 12450 7590 12502 7642
rect 1492 7531 1544 7540
rect 1492 7497 1501 7531
rect 1501 7497 1535 7531
rect 1535 7497 1544 7531
rect 1492 7488 1544 7497
rect 1768 7531 1820 7540
rect 1768 7497 1777 7531
rect 1777 7497 1811 7531
rect 1811 7497 1820 7531
rect 1768 7488 1820 7497
rect 1768 7352 1820 7404
rect 1952 7395 2004 7404
rect 1952 7361 1961 7395
rect 1961 7361 1995 7395
rect 1995 7361 2004 7395
rect 1952 7352 2004 7361
rect 3976 7352 4028 7404
rect 5540 7420 5592 7472
rect 4620 7352 4672 7404
rect 7656 7488 7708 7540
rect 9220 7531 9272 7540
rect 9220 7497 9229 7531
rect 9229 7497 9263 7531
rect 9263 7497 9272 7531
rect 9220 7488 9272 7497
rect 9404 7488 9456 7540
rect 9956 7488 10008 7540
rect 10968 7488 11020 7540
rect 11060 7488 11112 7540
rect 11796 7488 11848 7540
rect 12164 7488 12216 7540
rect 12348 7488 12400 7540
rect 7196 7352 7248 7404
rect 8484 7352 8536 7404
rect 6460 7284 6512 7336
rect 7840 7284 7892 7336
rect 10416 7463 10468 7472
rect 10416 7429 10434 7463
rect 10434 7429 10468 7463
rect 12900 7463 12952 7472
rect 10416 7420 10468 7429
rect 9312 7284 9364 7336
rect 7932 7216 7984 7268
rect 10692 7216 10744 7268
rect 11244 7352 11296 7404
rect 11060 7284 11112 7336
rect 11520 7284 11572 7336
rect 12900 7429 12909 7463
rect 12909 7429 12943 7463
rect 12943 7429 12952 7463
rect 12900 7420 12952 7429
rect 13084 7420 13136 7472
rect 14372 7420 14424 7472
rect 12716 7352 12768 7404
rect 12992 7352 13044 7404
rect 13544 7352 13596 7404
rect 3148 7191 3200 7200
rect 3148 7157 3157 7191
rect 3157 7157 3191 7191
rect 3191 7157 3200 7191
rect 3148 7148 3200 7157
rect 6368 7148 6420 7200
rect 12624 7216 12676 7268
rect 12900 7216 12952 7268
rect 13452 7216 13504 7268
rect 14464 7352 14516 7404
rect 14556 7399 14608 7404
rect 14556 7365 14565 7399
rect 14565 7365 14599 7399
rect 14599 7365 14608 7399
rect 16764 7420 16816 7472
rect 14556 7352 14608 7365
rect 14096 7327 14148 7336
rect 14096 7293 14105 7327
rect 14105 7293 14139 7327
rect 14139 7293 14148 7327
rect 15292 7352 15344 7404
rect 15568 7352 15620 7404
rect 14096 7284 14148 7293
rect 14556 7216 14608 7268
rect 11336 7191 11388 7200
rect 11336 7157 11345 7191
rect 11345 7157 11379 7191
rect 11379 7157 11388 7191
rect 11336 7148 11388 7157
rect 11520 7191 11572 7200
rect 11520 7157 11529 7191
rect 11529 7157 11563 7191
rect 11563 7157 11572 7191
rect 11520 7148 11572 7157
rect 13084 7191 13136 7200
rect 13084 7157 13093 7191
rect 13093 7157 13127 7191
rect 13127 7157 13136 7191
rect 13084 7148 13136 7157
rect 13544 7191 13596 7200
rect 13544 7157 13553 7191
rect 13553 7157 13587 7191
rect 13587 7157 13596 7191
rect 13544 7148 13596 7157
rect 14372 7191 14424 7200
rect 14372 7157 14381 7191
rect 14381 7157 14415 7191
rect 14415 7157 14424 7191
rect 14372 7148 14424 7157
rect 14648 7191 14700 7200
rect 14648 7157 14657 7191
rect 14657 7157 14691 7191
rect 14691 7157 14700 7191
rect 14648 7148 14700 7157
rect 15108 7216 15160 7268
rect 2824 7046 2876 7098
rect 2888 7046 2940 7098
rect 2952 7046 3004 7098
rect 3016 7046 3068 7098
rect 3080 7046 3132 7098
rect 6572 7046 6624 7098
rect 6636 7046 6688 7098
rect 6700 7046 6752 7098
rect 6764 7046 6816 7098
rect 6828 7046 6880 7098
rect 10320 7046 10372 7098
rect 10384 7046 10436 7098
rect 10448 7046 10500 7098
rect 10512 7046 10564 7098
rect 10576 7046 10628 7098
rect 14068 7046 14120 7098
rect 14132 7046 14184 7098
rect 14196 7046 14248 7098
rect 14260 7046 14312 7098
rect 14324 7046 14376 7098
rect 4620 6944 4672 6996
rect 2596 6876 2648 6928
rect 3424 6876 3476 6928
rect 1952 6851 2004 6860
rect 1952 6817 1961 6851
rect 1961 6817 1995 6851
rect 1995 6817 2004 6851
rect 1952 6808 2004 6817
rect 7564 6944 7616 6996
rect 7656 6876 7708 6928
rect 8392 6987 8444 6996
rect 8392 6953 8401 6987
rect 8401 6953 8435 6987
rect 8435 6953 8444 6987
rect 8392 6944 8444 6953
rect 9220 6944 9272 6996
rect 10968 6944 11020 6996
rect 11428 6944 11480 6996
rect 11796 6944 11848 6996
rect 13820 6944 13872 6996
rect 14188 6944 14240 6996
rect 7564 6808 7616 6860
rect 7932 6808 7984 6860
rect 3424 6740 3476 6792
rect 6644 6740 6696 6792
rect 9680 6876 9732 6928
rect 10232 6876 10284 6928
rect 2228 6715 2280 6724
rect 2228 6681 2237 6715
rect 2237 6681 2271 6715
rect 2271 6681 2280 6715
rect 2228 6672 2280 6681
rect 5448 6672 5500 6724
rect 9128 6808 9180 6860
rect 9496 6851 9548 6860
rect 9496 6817 9505 6851
rect 9505 6817 9539 6851
rect 9539 6817 9548 6851
rect 9864 6851 9916 6860
rect 9496 6808 9548 6817
rect 9864 6817 9873 6851
rect 9873 6817 9907 6851
rect 9907 6817 9916 6851
rect 9864 6808 9916 6817
rect 8484 6740 8536 6792
rect 1492 6647 1544 6656
rect 1492 6613 1501 6647
rect 1501 6613 1535 6647
rect 1535 6613 1544 6647
rect 1492 6604 1544 6613
rect 2504 6604 2556 6656
rect 2688 6604 2740 6656
rect 3608 6604 3660 6656
rect 5632 6604 5684 6656
rect 6920 6604 6972 6656
rect 7196 6604 7248 6656
rect 8760 6604 8812 6656
rect 11336 6808 11388 6860
rect 11888 6876 11940 6928
rect 11796 6808 11848 6860
rect 13176 6808 13228 6860
rect 14004 6808 14056 6860
rect 15108 6944 15160 6996
rect 14372 6876 14424 6928
rect 14740 6876 14792 6928
rect 15844 6808 15896 6860
rect 9220 6740 9272 6792
rect 10692 6740 10744 6792
rect 10876 6740 10928 6792
rect 11520 6783 11572 6792
rect 11520 6749 11529 6783
rect 11529 6749 11563 6783
rect 11563 6749 11572 6783
rect 11520 6740 11572 6749
rect 13544 6740 13596 6792
rect 13820 6740 13872 6792
rect 12992 6672 13044 6724
rect 14096 6740 14148 6792
rect 14280 6740 14332 6792
rect 9128 6604 9180 6656
rect 9404 6604 9456 6656
rect 9588 6604 9640 6656
rect 10140 6647 10192 6656
rect 10140 6613 10149 6647
rect 10149 6613 10183 6647
rect 10183 6613 10192 6647
rect 10140 6604 10192 6613
rect 10232 6604 10284 6656
rect 10692 6604 10744 6656
rect 11796 6604 11848 6656
rect 11888 6604 11940 6656
rect 12624 6604 12676 6656
rect 12808 6647 12860 6656
rect 12808 6613 12817 6647
rect 12817 6613 12851 6647
rect 12851 6613 12860 6647
rect 12808 6604 12860 6613
rect 13636 6604 13688 6656
rect 13820 6604 13872 6656
rect 14740 6740 14792 6792
rect 15108 6783 15160 6792
rect 15108 6749 15117 6783
rect 15117 6749 15151 6783
rect 15151 6749 15160 6783
rect 15108 6740 15160 6749
rect 15752 6604 15804 6656
rect 4698 6502 4750 6554
rect 4762 6502 4814 6554
rect 4826 6502 4878 6554
rect 4890 6502 4942 6554
rect 4954 6502 5006 6554
rect 8446 6502 8498 6554
rect 8510 6502 8562 6554
rect 8574 6502 8626 6554
rect 8638 6502 8690 6554
rect 8702 6502 8754 6554
rect 12194 6502 12246 6554
rect 12258 6502 12310 6554
rect 12322 6502 12374 6554
rect 12386 6502 12438 6554
rect 12450 6502 12502 6554
rect 1676 6400 1728 6452
rect 4252 6400 4304 6452
rect 4620 6400 4672 6452
rect 4712 6400 4764 6452
rect 5172 6400 5224 6452
rect 5632 6443 5684 6452
rect 5632 6409 5641 6443
rect 5641 6409 5675 6443
rect 5675 6409 5684 6443
rect 5632 6400 5684 6409
rect 5908 6400 5960 6452
rect 6460 6400 6512 6452
rect 7748 6400 7800 6452
rect 9036 6400 9088 6452
rect 10048 6400 10100 6452
rect 3516 6332 3568 6384
rect 4988 6375 5040 6384
rect 4988 6341 4997 6375
rect 4997 6341 5031 6375
rect 5031 6341 5040 6375
rect 4988 6332 5040 6341
rect 5448 6332 5500 6384
rect 6920 6332 6972 6384
rect 7840 6375 7892 6384
rect 7840 6341 7849 6375
rect 7849 6341 7883 6375
rect 7883 6341 7892 6375
rect 7840 6332 7892 6341
rect 8208 6375 8260 6384
rect 8208 6341 8242 6375
rect 8242 6341 8260 6375
rect 8208 6332 8260 6341
rect 8852 6332 8904 6384
rect 9772 6375 9824 6384
rect 9772 6341 9781 6375
rect 9781 6341 9815 6375
rect 9815 6341 9824 6375
rect 9772 6332 9824 6341
rect 10324 6332 10376 6384
rect 11244 6400 11296 6452
rect 12072 6400 12124 6452
rect 12624 6443 12676 6452
rect 12624 6409 12633 6443
rect 12633 6409 12667 6443
rect 12667 6409 12676 6443
rect 12624 6400 12676 6409
rect 12992 6400 13044 6452
rect 13820 6443 13872 6452
rect 13820 6409 13829 6443
rect 13829 6409 13863 6443
rect 13863 6409 13872 6443
rect 13820 6400 13872 6409
rect 14096 6400 14148 6452
rect 14648 6400 14700 6452
rect 14924 6443 14976 6452
rect 14924 6409 14933 6443
rect 14933 6409 14967 6443
rect 14967 6409 14976 6443
rect 14924 6400 14976 6409
rect 15292 6443 15344 6452
rect 15292 6409 15301 6443
rect 15301 6409 15335 6443
rect 15335 6409 15344 6443
rect 15292 6400 15344 6409
rect 3884 6264 3936 6316
rect 4068 6264 4120 6316
rect 5540 6307 5592 6316
rect 5540 6273 5549 6307
rect 5549 6273 5583 6307
rect 5583 6273 5592 6307
rect 5540 6264 5592 6273
rect 7012 6264 7064 6316
rect 7104 6307 7156 6316
rect 7104 6273 7113 6307
rect 7113 6273 7147 6307
rect 7147 6273 7156 6307
rect 7104 6264 7156 6273
rect 7380 6264 7432 6316
rect 2044 6239 2096 6248
rect 2044 6205 2053 6239
rect 2053 6205 2087 6239
rect 2087 6205 2096 6239
rect 2044 6196 2096 6205
rect 2320 6196 2372 6248
rect 3148 6128 3200 6180
rect 4528 6196 4580 6248
rect 5448 6196 5500 6248
rect 5816 6239 5868 6248
rect 5816 6205 5825 6239
rect 5825 6205 5859 6239
rect 5859 6205 5868 6239
rect 5816 6196 5868 6205
rect 6828 6239 6880 6248
rect 6828 6205 6837 6239
rect 6837 6205 6871 6239
rect 6871 6205 6880 6239
rect 6828 6196 6880 6205
rect 4344 6128 4396 6180
rect 1400 6103 1452 6112
rect 1400 6069 1409 6103
rect 1409 6069 1443 6103
rect 1443 6069 1452 6103
rect 1400 6060 1452 6069
rect 3700 6060 3752 6112
rect 4620 6103 4672 6112
rect 4620 6069 4629 6103
rect 4629 6069 4663 6103
rect 4663 6069 4672 6103
rect 4620 6060 4672 6069
rect 5172 6103 5224 6112
rect 5172 6069 5181 6103
rect 5181 6069 5215 6103
rect 5215 6069 5224 6103
rect 5172 6060 5224 6069
rect 6460 6060 6512 6112
rect 7104 6060 7156 6112
rect 7564 6128 7616 6180
rect 7472 6103 7524 6112
rect 7472 6069 7481 6103
rect 7481 6069 7515 6103
rect 7515 6069 7524 6103
rect 7472 6060 7524 6069
rect 7840 6060 7892 6112
rect 8668 6060 8720 6112
rect 9036 6264 9088 6316
rect 9312 6171 9364 6180
rect 9312 6137 9321 6171
rect 9321 6137 9355 6171
rect 9355 6137 9364 6171
rect 9312 6128 9364 6137
rect 10140 6264 10192 6316
rect 11428 6332 11480 6384
rect 15108 6332 15160 6384
rect 11796 6264 11848 6316
rect 12164 6307 12216 6316
rect 12164 6273 12173 6307
rect 12173 6273 12207 6307
rect 12207 6273 12216 6307
rect 12164 6264 12216 6273
rect 12716 6264 12768 6316
rect 9588 6196 9640 6248
rect 10600 6196 10652 6248
rect 12624 6196 12676 6248
rect 12900 6196 12952 6248
rect 13728 6264 13780 6316
rect 13912 6264 13964 6316
rect 15568 6307 15620 6316
rect 14372 6196 14424 6248
rect 15568 6273 15577 6307
rect 15577 6273 15611 6307
rect 15611 6273 15620 6307
rect 15568 6264 15620 6273
rect 16580 6264 16632 6316
rect 10140 6060 10192 6112
rect 10968 6060 11020 6112
rect 11244 6103 11296 6112
rect 11244 6069 11253 6103
rect 11253 6069 11287 6103
rect 11287 6069 11296 6103
rect 11244 6060 11296 6069
rect 11336 6060 11388 6112
rect 11980 6060 12032 6112
rect 12348 6060 12400 6112
rect 13820 6060 13872 6112
rect 14004 6060 14056 6112
rect 14188 6060 14240 6112
rect 14648 6060 14700 6112
rect 15108 6196 15160 6248
rect 15384 6103 15436 6112
rect 15384 6069 15393 6103
rect 15393 6069 15427 6103
rect 15427 6069 15436 6103
rect 15384 6060 15436 6069
rect 2824 5958 2876 6010
rect 2888 5958 2940 6010
rect 2952 5958 3004 6010
rect 3016 5958 3068 6010
rect 3080 5958 3132 6010
rect 6572 5958 6624 6010
rect 6636 5958 6688 6010
rect 6700 5958 6752 6010
rect 6764 5958 6816 6010
rect 6828 5958 6880 6010
rect 10320 5958 10372 6010
rect 10384 5958 10436 6010
rect 10448 5958 10500 6010
rect 10512 5958 10564 6010
rect 10576 5958 10628 6010
rect 14068 5958 14120 6010
rect 14132 5958 14184 6010
rect 14196 5958 14248 6010
rect 14260 5958 14312 6010
rect 14324 5958 14376 6010
rect 1768 5899 1820 5908
rect 1768 5865 1777 5899
rect 1777 5865 1811 5899
rect 1811 5865 1820 5899
rect 1768 5856 1820 5865
rect 2044 5856 2096 5908
rect 5264 5856 5316 5908
rect 5816 5856 5868 5908
rect 6276 5856 6328 5908
rect 6736 5856 6788 5908
rect 12624 5856 12676 5908
rect 14004 5856 14056 5908
rect 15568 5856 15620 5908
rect 2136 5720 2188 5772
rect 3148 5788 3200 5840
rect 3424 5831 3476 5840
rect 3424 5797 3433 5831
rect 3433 5797 3467 5831
rect 3467 5797 3476 5831
rect 3424 5788 3476 5797
rect 2320 5652 2372 5704
rect 4344 5720 4396 5772
rect 5080 5788 5132 5840
rect 5540 5788 5592 5840
rect 7840 5788 7892 5840
rect 7932 5831 7984 5840
rect 7932 5797 7941 5831
rect 7941 5797 7975 5831
rect 7975 5797 7984 5831
rect 7932 5788 7984 5797
rect 5264 5763 5316 5772
rect 5264 5729 5273 5763
rect 5273 5729 5307 5763
rect 5307 5729 5316 5763
rect 5264 5720 5316 5729
rect 5448 5720 5500 5772
rect 6000 5720 6052 5772
rect 6460 5720 6512 5772
rect 6736 5763 6788 5772
rect 6736 5729 6745 5763
rect 6745 5729 6779 5763
rect 6779 5729 6788 5763
rect 6736 5720 6788 5729
rect 7104 5763 7156 5772
rect 7104 5729 7113 5763
rect 7113 5729 7147 5763
rect 7147 5729 7156 5763
rect 7104 5720 7156 5729
rect 7196 5720 7248 5772
rect 9036 5788 9088 5840
rect 9312 5788 9364 5840
rect 9496 5788 9548 5840
rect 9772 5788 9824 5840
rect 10416 5788 10468 5840
rect 10968 5788 11020 5840
rect 4712 5652 4764 5704
rect 5080 5652 5132 5704
rect 2228 5627 2280 5636
rect 2228 5593 2237 5627
rect 2237 5593 2271 5627
rect 2271 5593 2280 5627
rect 2228 5584 2280 5593
rect 2596 5584 2648 5636
rect 6276 5652 6328 5704
rect 8392 5720 8444 5772
rect 9128 5720 9180 5772
rect 9588 5720 9640 5772
rect 10140 5720 10192 5772
rect 11796 5788 11848 5840
rect 14740 5788 14792 5840
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 7380 5584 7432 5636
rect 8300 5652 8352 5704
rect 8852 5652 8904 5704
rect 9036 5695 9088 5704
rect 9036 5661 9045 5695
rect 9045 5661 9079 5695
rect 9079 5661 9088 5695
rect 9036 5652 9088 5661
rect 7840 5584 7892 5636
rect 8576 5584 8628 5636
rect 8668 5584 8720 5636
rect 9588 5584 9640 5636
rect 10048 5652 10100 5704
rect 10968 5652 11020 5704
rect 11152 5695 11204 5704
rect 11152 5661 11161 5695
rect 11161 5661 11195 5695
rect 11195 5661 11204 5695
rect 11152 5652 11204 5661
rect 11244 5652 11296 5704
rect 12440 5763 12492 5772
rect 12440 5729 12449 5763
rect 12449 5729 12483 5763
rect 12483 5729 12492 5763
rect 13360 5763 13412 5772
rect 12440 5720 12492 5729
rect 13360 5729 13369 5763
rect 13369 5729 13403 5763
rect 13403 5729 13412 5763
rect 13360 5720 13412 5729
rect 14280 5720 14332 5772
rect 11980 5652 12032 5704
rect 14096 5695 14148 5704
rect 14096 5661 14105 5695
rect 14105 5661 14139 5695
rect 14139 5661 14148 5695
rect 14096 5652 14148 5661
rect 14648 5652 14700 5704
rect 14832 5695 14884 5704
rect 14832 5661 14841 5695
rect 14841 5661 14875 5695
rect 14875 5661 14884 5695
rect 14832 5652 14884 5661
rect 3516 5516 3568 5568
rect 4160 5516 4212 5568
rect 4252 5559 4304 5568
rect 4252 5525 4261 5559
rect 4261 5525 4295 5559
rect 4295 5525 4304 5559
rect 4252 5516 4304 5525
rect 5264 5516 5316 5568
rect 5448 5516 5500 5568
rect 8208 5516 8260 5568
rect 9036 5516 9088 5568
rect 9772 5559 9824 5568
rect 9772 5525 9781 5559
rect 9781 5525 9815 5559
rect 9815 5525 9824 5559
rect 9772 5516 9824 5525
rect 10232 5559 10284 5568
rect 10232 5525 10241 5559
rect 10241 5525 10275 5559
rect 10275 5525 10284 5559
rect 10232 5516 10284 5525
rect 10692 5559 10744 5568
rect 10692 5525 10701 5559
rect 10701 5525 10735 5559
rect 10735 5525 10744 5559
rect 10692 5516 10744 5525
rect 11428 5516 11480 5568
rect 11796 5559 11848 5568
rect 11796 5525 11805 5559
rect 11805 5525 11839 5559
rect 11839 5525 11848 5559
rect 11796 5516 11848 5525
rect 12348 5516 12400 5568
rect 14188 5584 14240 5636
rect 13728 5516 13780 5568
rect 14372 5559 14424 5568
rect 14372 5525 14381 5559
rect 14381 5525 14415 5559
rect 14415 5525 14424 5559
rect 14372 5516 14424 5525
rect 15016 5516 15068 5568
rect 4698 5414 4750 5466
rect 4762 5414 4814 5466
rect 4826 5414 4878 5466
rect 4890 5414 4942 5466
rect 4954 5414 5006 5466
rect 8446 5414 8498 5466
rect 8510 5414 8562 5466
rect 8574 5414 8626 5466
rect 8638 5414 8690 5466
rect 8702 5414 8754 5466
rect 12194 5414 12246 5466
rect 12258 5414 12310 5466
rect 12322 5414 12374 5466
rect 12386 5414 12438 5466
rect 12450 5414 12502 5466
rect 3516 5312 3568 5364
rect 3976 5312 4028 5364
rect 1676 5219 1728 5228
rect 1676 5185 1685 5219
rect 1685 5185 1719 5219
rect 1719 5185 1728 5219
rect 1676 5176 1728 5185
rect 2504 5176 2556 5228
rect 2688 5244 2740 5296
rect 4160 5244 4212 5296
rect 3792 5176 3844 5228
rect 3976 5219 4028 5228
rect 3976 5185 3985 5219
rect 3985 5185 4019 5219
rect 4019 5185 4028 5219
rect 3976 5176 4028 5185
rect 1952 5151 2004 5160
rect 1952 5117 1961 5151
rect 1961 5117 1995 5151
rect 1995 5117 2004 5151
rect 1952 5108 2004 5117
rect 3424 5108 3476 5160
rect 3608 5108 3660 5160
rect 4988 5312 5040 5364
rect 5356 5312 5408 5364
rect 5448 5312 5500 5364
rect 5264 5244 5316 5296
rect 7656 5312 7708 5364
rect 7748 5312 7800 5364
rect 9772 5312 9824 5364
rect 10232 5312 10284 5364
rect 10968 5355 11020 5364
rect 10968 5321 10977 5355
rect 10977 5321 11011 5355
rect 11011 5321 11020 5355
rect 10968 5312 11020 5321
rect 11888 5312 11940 5364
rect 12256 5355 12308 5364
rect 12256 5321 12265 5355
rect 12265 5321 12299 5355
rect 12299 5321 12308 5355
rect 12256 5312 12308 5321
rect 12348 5312 12400 5364
rect 13820 5312 13872 5364
rect 14096 5355 14148 5364
rect 14096 5321 14105 5355
rect 14105 5321 14139 5355
rect 14139 5321 14148 5355
rect 14096 5312 14148 5321
rect 14464 5312 14516 5364
rect 14740 5312 14792 5364
rect 15476 5355 15528 5364
rect 15476 5321 15485 5355
rect 15485 5321 15519 5355
rect 15519 5321 15528 5355
rect 15476 5312 15528 5321
rect 5908 5287 5960 5296
rect 5908 5253 5917 5287
rect 5917 5253 5951 5287
rect 5951 5253 5960 5287
rect 5908 5244 5960 5253
rect 6184 5244 6236 5296
rect 6460 5244 6512 5296
rect 6736 5244 6788 5296
rect 6920 5244 6972 5296
rect 5540 5176 5592 5228
rect 5816 5176 5868 5228
rect 7196 5176 7248 5228
rect 7288 5176 7340 5228
rect 11336 5244 11388 5296
rect 9036 5219 9088 5228
rect 2320 5040 2372 5092
rect 1492 5015 1544 5024
rect 1492 4981 1501 5015
rect 1501 4981 1535 5015
rect 1535 4981 1544 5015
rect 1492 4972 1544 4981
rect 1860 4972 1912 5024
rect 3148 4972 3200 5024
rect 3700 4972 3752 5024
rect 4068 4972 4120 5024
rect 4896 5015 4948 5024
rect 4896 4981 4905 5015
rect 4905 4981 4939 5015
rect 4939 4981 4948 5015
rect 4896 4972 4948 4981
rect 7104 5108 7156 5160
rect 7840 5151 7892 5160
rect 7840 5117 7849 5151
rect 7849 5117 7883 5151
rect 7883 5117 7892 5151
rect 7840 5108 7892 5117
rect 5448 5040 5500 5092
rect 6000 4972 6052 5024
rect 6368 5015 6420 5024
rect 6368 4981 6377 5015
rect 6377 4981 6411 5015
rect 6411 4981 6420 5015
rect 6368 4972 6420 4981
rect 7104 4972 7156 5024
rect 7380 4972 7432 5024
rect 8484 5108 8536 5160
rect 9036 5185 9045 5219
rect 9045 5185 9079 5219
rect 9079 5185 9088 5219
rect 9036 5176 9088 5185
rect 10048 5176 10100 5228
rect 10232 5176 10284 5228
rect 10600 5176 10652 5228
rect 12440 5244 12492 5296
rect 13544 5287 13596 5296
rect 9128 5151 9180 5160
rect 8208 5040 8260 5092
rect 8392 5040 8444 5092
rect 8760 4972 8812 5024
rect 9128 5117 9137 5151
rect 9137 5117 9171 5151
rect 9171 5117 9180 5151
rect 9128 5108 9180 5117
rect 9864 5151 9916 5160
rect 9864 5117 9873 5151
rect 9873 5117 9907 5151
rect 9907 5117 9916 5151
rect 9864 5108 9916 5117
rect 9956 5108 10008 5160
rect 10508 5108 10560 5160
rect 10692 5151 10744 5160
rect 10692 5117 10701 5151
rect 10701 5117 10735 5151
rect 10735 5117 10744 5151
rect 10692 5108 10744 5117
rect 11428 5108 11480 5160
rect 12716 5219 12768 5228
rect 12716 5185 12725 5219
rect 12725 5185 12759 5219
rect 12759 5185 12768 5219
rect 12716 5176 12768 5185
rect 12900 5176 12952 5228
rect 13084 5176 13136 5228
rect 13544 5253 13553 5287
rect 13553 5253 13587 5287
rect 13587 5253 13596 5287
rect 13544 5244 13596 5253
rect 14280 5244 14332 5296
rect 12808 5151 12860 5160
rect 12808 5117 12817 5151
rect 12817 5117 12851 5151
rect 12851 5117 12860 5151
rect 12808 5108 12860 5117
rect 13544 5108 13596 5160
rect 14096 5108 14148 5160
rect 14648 5108 14700 5160
rect 15292 5176 15344 5228
rect 9496 5040 9548 5092
rect 10324 4972 10376 5024
rect 11336 5015 11388 5024
rect 11336 4981 11345 5015
rect 11345 4981 11379 5015
rect 11379 4981 11388 5015
rect 11336 4972 11388 4981
rect 12348 5015 12400 5024
rect 12348 4981 12357 5015
rect 12357 4981 12391 5015
rect 12391 4981 12400 5015
rect 12348 4972 12400 4981
rect 12440 4972 12492 5024
rect 14464 5015 14516 5024
rect 14464 4981 14473 5015
rect 14473 4981 14507 5015
rect 14507 4981 14516 5015
rect 14464 4972 14516 4981
rect 15108 5040 15160 5092
rect 15844 5244 15896 5296
rect 15660 5219 15712 5228
rect 15660 5185 15669 5219
rect 15669 5185 15703 5219
rect 15703 5185 15712 5219
rect 15660 5176 15712 5185
rect 2824 4870 2876 4922
rect 2888 4870 2940 4922
rect 2952 4870 3004 4922
rect 3016 4870 3068 4922
rect 3080 4870 3132 4922
rect 6572 4870 6624 4922
rect 6636 4870 6688 4922
rect 6700 4870 6752 4922
rect 6764 4870 6816 4922
rect 6828 4870 6880 4922
rect 10320 4870 10372 4922
rect 10384 4870 10436 4922
rect 10448 4870 10500 4922
rect 10512 4870 10564 4922
rect 10576 4870 10628 4922
rect 14068 4870 14120 4922
rect 14132 4870 14184 4922
rect 14196 4870 14248 4922
rect 14260 4870 14312 4922
rect 14324 4870 14376 4922
rect 1676 4811 1728 4820
rect 1676 4777 1685 4811
rect 1685 4777 1719 4811
rect 1719 4777 1728 4811
rect 1676 4768 1728 4777
rect 2412 4811 2464 4820
rect 2412 4777 2421 4811
rect 2421 4777 2455 4811
rect 2455 4777 2464 4811
rect 2412 4768 2464 4777
rect 2596 4768 2648 4820
rect 4528 4768 4580 4820
rect 5448 4768 5500 4820
rect 6276 4768 6328 4820
rect 6368 4768 6420 4820
rect 6552 4768 6604 4820
rect 7288 4768 7340 4820
rect 9036 4768 9088 4820
rect 9772 4768 9824 4820
rect 10968 4768 11020 4820
rect 11060 4768 11112 4820
rect 11336 4768 11388 4820
rect 1584 4743 1636 4752
rect 1584 4709 1593 4743
rect 1593 4709 1627 4743
rect 1627 4709 1636 4743
rect 1584 4700 1636 4709
rect 3332 4700 3384 4752
rect 3608 4700 3660 4752
rect 1400 4607 1452 4616
rect 1400 4573 1409 4607
rect 1409 4573 1443 4607
rect 1443 4573 1452 4607
rect 1400 4564 1452 4573
rect 2596 4632 2648 4684
rect 6828 4700 6880 4752
rect 8760 4700 8812 4752
rect 4436 4675 4488 4684
rect 4436 4641 4445 4675
rect 4445 4641 4479 4675
rect 4479 4641 4488 4675
rect 4436 4632 4488 4641
rect 4988 4675 5040 4684
rect 4988 4641 4997 4675
rect 4997 4641 5031 4675
rect 5031 4641 5040 4675
rect 4988 4632 5040 4641
rect 5816 4632 5868 4684
rect 6276 4675 6328 4684
rect 6276 4641 6285 4675
rect 6285 4641 6319 4675
rect 6319 4641 6328 4675
rect 6276 4632 6328 4641
rect 6460 4675 6512 4684
rect 6460 4641 6469 4675
rect 6469 4641 6503 4675
rect 6503 4641 6512 4675
rect 6460 4632 6512 4641
rect 7104 4675 7156 4684
rect 7104 4641 7113 4675
rect 7113 4641 7147 4675
rect 7147 4641 7156 4675
rect 7104 4632 7156 4641
rect 7288 4675 7340 4684
rect 7288 4641 7297 4675
rect 7297 4641 7331 4675
rect 7331 4641 7340 4675
rect 7288 4632 7340 4641
rect 7932 4675 7984 4684
rect 7932 4641 7941 4675
rect 7941 4641 7975 4675
rect 7975 4641 7984 4675
rect 7932 4632 7984 4641
rect 8024 4675 8076 4684
rect 8024 4641 8033 4675
rect 8033 4641 8067 4675
rect 8067 4641 8076 4675
rect 8944 4700 8996 4752
rect 9496 4700 9548 4752
rect 9864 4675 9916 4684
rect 8024 4632 8076 4641
rect 9864 4641 9873 4675
rect 9873 4641 9907 4675
rect 9907 4641 9916 4675
rect 9864 4632 9916 4641
rect 10692 4632 10744 4684
rect 10784 4632 10836 4684
rect 2228 4607 2280 4616
rect 2228 4573 2237 4607
rect 2237 4573 2271 4607
rect 2271 4573 2280 4607
rect 2228 4564 2280 4573
rect 5724 4564 5776 4616
rect 5908 4564 5960 4616
rect 6920 4564 6972 4616
rect 7472 4564 7524 4616
rect 2412 4496 2464 4548
rect 2688 4496 2740 4548
rect 2044 4428 2096 4480
rect 2504 4428 2556 4480
rect 3240 4496 3292 4548
rect 3516 4496 3568 4548
rect 5540 4496 5592 4548
rect 7932 4540 7984 4592
rect 3056 4471 3108 4480
rect 3056 4437 3065 4471
rect 3065 4437 3099 4471
rect 3099 4437 3108 4471
rect 3056 4428 3108 4437
rect 3792 4428 3844 4480
rect 4160 4471 4212 4480
rect 4160 4437 4169 4471
rect 4169 4437 4203 4471
rect 4203 4437 4212 4471
rect 4160 4428 4212 4437
rect 5448 4428 5500 4480
rect 5908 4428 5960 4480
rect 8300 4496 8352 4548
rect 8576 4583 8628 4592
rect 8576 4549 8585 4583
rect 8585 4549 8619 4583
rect 8619 4549 8628 4583
rect 8760 4564 8812 4616
rect 8576 4540 8628 4549
rect 7104 4428 7156 4480
rect 7288 4428 7340 4480
rect 7748 4428 7800 4480
rect 8392 4428 8444 4480
rect 9588 4564 9640 4616
rect 12348 4768 12400 4820
rect 12716 4811 12768 4820
rect 12716 4777 12725 4811
rect 12725 4777 12759 4811
rect 12759 4777 12768 4811
rect 12716 4768 12768 4777
rect 13912 4811 13964 4820
rect 13912 4777 13921 4811
rect 13921 4777 13955 4811
rect 13955 4777 13964 4811
rect 13912 4768 13964 4777
rect 14556 4811 14608 4820
rect 14556 4777 14565 4811
rect 14565 4777 14599 4811
rect 14599 4777 14608 4811
rect 14556 4768 14608 4777
rect 14648 4768 14700 4820
rect 15476 4768 15528 4820
rect 12072 4700 12124 4752
rect 12900 4632 12952 4684
rect 13176 4632 13228 4684
rect 13360 4675 13412 4684
rect 13360 4641 13369 4675
rect 13369 4641 13403 4675
rect 13403 4641 13412 4675
rect 13360 4632 13412 4641
rect 13452 4632 13504 4684
rect 13728 4632 13780 4684
rect 15016 4675 15068 4684
rect 15016 4641 15025 4675
rect 15025 4641 15059 4675
rect 15059 4641 15068 4675
rect 15016 4632 15068 4641
rect 15108 4675 15160 4684
rect 15108 4641 15117 4675
rect 15117 4641 15151 4675
rect 15151 4641 15160 4675
rect 15108 4632 15160 4641
rect 12072 4564 12124 4616
rect 12256 4564 12308 4616
rect 14096 4564 14148 4616
rect 9864 4496 9916 4548
rect 11060 4539 11112 4548
rect 10600 4471 10652 4480
rect 10600 4437 10609 4471
rect 10609 4437 10643 4471
rect 10643 4437 10652 4471
rect 10600 4428 10652 4437
rect 11060 4505 11069 4539
rect 11069 4505 11103 4539
rect 11103 4505 11112 4539
rect 11060 4496 11112 4505
rect 12164 4496 12216 4548
rect 12716 4496 12768 4548
rect 13728 4496 13780 4548
rect 14832 4496 14884 4548
rect 11336 4428 11388 4480
rect 11980 4428 12032 4480
rect 12992 4428 13044 4480
rect 15108 4428 15160 4480
rect 4698 4326 4750 4378
rect 4762 4326 4814 4378
rect 4826 4326 4878 4378
rect 4890 4326 4942 4378
rect 4954 4326 5006 4378
rect 8446 4326 8498 4378
rect 8510 4326 8562 4378
rect 8574 4326 8626 4378
rect 8638 4326 8690 4378
rect 8702 4326 8754 4378
rect 12194 4326 12246 4378
rect 12258 4326 12310 4378
rect 12322 4326 12374 4378
rect 12386 4326 12438 4378
rect 12450 4326 12502 4378
rect 1860 4267 1912 4276
rect 1860 4233 1869 4267
rect 1869 4233 1903 4267
rect 1903 4233 1912 4267
rect 1860 4224 1912 4233
rect 1952 4224 2004 4276
rect 2320 4224 2372 4276
rect 3056 4224 3108 4276
rect 3700 4224 3752 4276
rect 4344 4224 4396 4276
rect 4528 4224 4580 4276
rect 5540 4224 5592 4276
rect 1952 4131 2004 4140
rect 1952 4097 1961 4131
rect 1961 4097 1995 4131
rect 1995 4097 2004 4131
rect 1952 4088 2004 4097
rect 1768 4063 1820 4072
rect 1768 4029 1777 4063
rect 1777 4029 1811 4063
rect 1811 4029 1820 4063
rect 1768 4020 1820 4029
rect 2872 4131 2924 4140
rect 2872 4097 2881 4131
rect 2881 4097 2915 4131
rect 2915 4097 2924 4131
rect 2872 4088 2924 4097
rect 3240 4088 3292 4140
rect 3332 4088 3384 4140
rect 3976 4156 4028 4208
rect 4160 4156 4212 4208
rect 5724 4156 5776 4208
rect 8852 4224 8904 4276
rect 10048 4224 10100 4276
rect 12900 4224 12952 4276
rect 13452 4224 13504 4276
rect 13912 4224 13964 4276
rect 14832 4224 14884 4276
rect 7564 4156 7616 4208
rect 3792 4063 3844 4072
rect 3792 4029 3801 4063
rect 3801 4029 3835 4063
rect 3835 4029 3844 4063
rect 3792 4020 3844 4029
rect 3332 3952 3384 4004
rect 4068 4088 4120 4140
rect 5264 4088 5316 4140
rect 6368 4088 6420 4140
rect 7380 4131 7432 4140
rect 7380 4097 7389 4131
rect 7389 4097 7423 4131
rect 7423 4097 7432 4131
rect 7380 4088 7432 4097
rect 7472 4088 7524 4140
rect 8116 4131 8168 4140
rect 8116 4097 8125 4131
rect 8125 4097 8159 4131
rect 8159 4097 8168 4131
rect 8116 4088 8168 4097
rect 8208 4112 8260 4164
rect 10600 4156 10652 4208
rect 4252 3995 4304 4004
rect 4252 3961 4261 3995
rect 4261 3961 4295 3995
rect 4295 3961 4304 3995
rect 4252 3952 4304 3961
rect 5356 3952 5408 4004
rect 6092 3952 6144 4004
rect 1676 3884 1728 3936
rect 2596 3884 2648 3936
rect 3240 3927 3292 3936
rect 3240 3893 3249 3927
rect 3249 3893 3283 3927
rect 3283 3893 3292 3927
rect 3240 3884 3292 3893
rect 3884 3884 3936 3936
rect 4436 3884 4488 3936
rect 4528 3884 4580 3936
rect 5264 3884 5316 3936
rect 6276 3884 6328 3936
rect 6460 3884 6512 3936
rect 6644 3884 6696 3936
rect 7196 4020 7248 4072
rect 7840 4063 7892 4072
rect 7840 4029 7849 4063
rect 7849 4029 7883 4063
rect 7883 4029 7892 4063
rect 7840 4020 7892 4029
rect 8208 4020 8260 4072
rect 7104 3952 7156 4004
rect 8668 4020 8720 4072
rect 9036 4063 9088 4072
rect 9036 4029 9045 4063
rect 9045 4029 9079 4063
rect 9079 4029 9088 4063
rect 9036 4020 9088 4029
rect 9404 4088 9456 4140
rect 9772 4088 9824 4140
rect 10968 4131 11020 4140
rect 10968 4097 10977 4131
rect 10977 4097 11011 4131
rect 11011 4097 11020 4131
rect 10968 4088 11020 4097
rect 11336 4088 11388 4140
rect 12256 4088 12308 4140
rect 9220 3952 9272 4004
rect 7196 3927 7248 3936
rect 7196 3893 7205 3927
rect 7205 3893 7239 3927
rect 7239 3893 7248 3927
rect 7196 3884 7248 3893
rect 7380 3884 7432 3936
rect 7840 3884 7892 3936
rect 8944 3884 8996 3936
rect 10324 4020 10376 4072
rect 10784 4020 10836 4072
rect 11428 4020 11480 4072
rect 12164 4063 12216 4072
rect 12164 4029 12173 4063
rect 12173 4029 12207 4063
rect 12207 4029 12216 4063
rect 12164 4020 12216 4029
rect 13084 4156 13136 4208
rect 12992 4088 13044 4140
rect 13176 4088 13228 4140
rect 13820 4088 13872 4140
rect 10600 3927 10652 3936
rect 10600 3893 10609 3927
rect 10609 3893 10643 3927
rect 10643 3893 10652 3927
rect 10600 3884 10652 3893
rect 11520 3927 11572 3936
rect 11520 3893 11529 3927
rect 11529 3893 11563 3927
rect 11563 3893 11572 3927
rect 11520 3884 11572 3893
rect 13268 3952 13320 4004
rect 13360 3952 13412 4004
rect 13820 3952 13872 4004
rect 15292 4156 15344 4208
rect 14648 4063 14700 4072
rect 14648 4029 14657 4063
rect 14657 4029 14691 4063
rect 14691 4029 14700 4063
rect 14648 4020 14700 4029
rect 14832 4063 14884 4072
rect 14832 4029 14841 4063
rect 14841 4029 14875 4063
rect 14875 4029 14884 4063
rect 14832 4020 14884 4029
rect 16120 4088 16172 4140
rect 16396 4020 16448 4072
rect 15016 3952 15068 4004
rect 14096 3884 14148 3936
rect 14648 3884 14700 3936
rect 15292 3927 15344 3936
rect 15292 3893 15301 3927
rect 15301 3893 15335 3927
rect 15335 3893 15344 3927
rect 15292 3884 15344 3893
rect 15568 3927 15620 3936
rect 15568 3893 15577 3927
rect 15577 3893 15611 3927
rect 15611 3893 15620 3927
rect 15568 3884 15620 3893
rect 2824 3782 2876 3834
rect 2888 3782 2940 3834
rect 2952 3782 3004 3834
rect 3016 3782 3068 3834
rect 3080 3782 3132 3834
rect 6572 3782 6624 3834
rect 6636 3782 6688 3834
rect 6700 3782 6752 3834
rect 6764 3782 6816 3834
rect 6828 3782 6880 3834
rect 10320 3782 10372 3834
rect 10384 3782 10436 3834
rect 10448 3782 10500 3834
rect 10512 3782 10564 3834
rect 10576 3782 10628 3834
rect 14068 3782 14120 3834
rect 14132 3782 14184 3834
rect 14196 3782 14248 3834
rect 14260 3782 14312 3834
rect 14324 3782 14376 3834
rect 1492 3723 1544 3732
rect 1492 3689 1501 3723
rect 1501 3689 1535 3723
rect 1535 3689 1544 3723
rect 1492 3680 1544 3689
rect 2504 3680 2556 3732
rect 3976 3680 4028 3732
rect 4068 3680 4120 3732
rect 6368 3680 6420 3732
rect 7104 3680 7156 3732
rect 8024 3680 8076 3732
rect 8576 3680 8628 3732
rect 8944 3723 8996 3732
rect 8944 3689 8953 3723
rect 8953 3689 8987 3723
rect 8987 3689 8996 3723
rect 8944 3680 8996 3689
rect 9036 3680 9088 3732
rect 11060 3723 11112 3732
rect 11060 3689 11069 3723
rect 11069 3689 11103 3723
rect 11103 3689 11112 3723
rect 11060 3680 11112 3689
rect 11152 3680 11204 3732
rect 12716 3680 12768 3732
rect 13544 3680 13596 3732
rect 14464 3680 14516 3732
rect 3056 3612 3108 3664
rect 2688 3544 2740 3596
rect 1676 3519 1728 3528
rect 1676 3485 1685 3519
rect 1685 3485 1719 3519
rect 1719 3485 1728 3519
rect 1676 3476 1728 3485
rect 2044 3519 2096 3528
rect 2044 3485 2053 3519
rect 2053 3485 2087 3519
rect 2087 3485 2096 3519
rect 2044 3476 2096 3485
rect 2136 3476 2188 3528
rect 2872 3519 2924 3528
rect 2872 3485 2881 3519
rect 2881 3485 2915 3519
rect 2915 3485 2924 3519
rect 2872 3476 2924 3485
rect 3148 3519 3200 3528
rect 3148 3485 3157 3519
rect 3157 3485 3191 3519
rect 3191 3485 3200 3519
rect 3148 3476 3200 3485
rect 3700 3544 3752 3596
rect 4528 3544 4580 3596
rect 5080 3612 5132 3664
rect 5724 3544 5776 3596
rect 4436 3519 4488 3528
rect 4436 3485 4445 3519
rect 4445 3485 4479 3519
rect 4479 3485 4488 3519
rect 4436 3476 4488 3485
rect 5356 3476 5408 3528
rect 6828 3544 6880 3596
rect 7288 3587 7340 3596
rect 7288 3553 7297 3587
rect 7297 3553 7331 3587
rect 7331 3553 7340 3587
rect 7288 3544 7340 3553
rect 6276 3476 6328 3528
rect 6644 3476 6696 3528
rect 1860 3383 1912 3392
rect 1860 3349 1869 3383
rect 1869 3349 1903 3383
rect 1903 3349 1912 3383
rect 1860 3340 1912 3349
rect 1952 3340 2004 3392
rect 2228 3340 2280 3392
rect 2504 3340 2556 3392
rect 2964 3383 3016 3392
rect 2964 3349 2973 3383
rect 2973 3349 3007 3383
rect 3007 3349 3016 3383
rect 2964 3340 3016 3349
rect 5448 3408 5500 3460
rect 5540 3408 5592 3460
rect 8024 3544 8076 3596
rect 8208 3476 8260 3528
rect 8392 3544 8444 3596
rect 10416 3612 10468 3664
rect 9496 3544 9548 3596
rect 7288 3408 7340 3460
rect 7472 3408 7524 3460
rect 7748 3408 7800 3460
rect 4160 3340 4212 3392
rect 4620 3340 4672 3392
rect 5080 3340 5132 3392
rect 5816 3340 5868 3392
rect 6368 3340 6420 3392
rect 6828 3340 6880 3392
rect 9220 3476 9272 3528
rect 10048 3544 10100 3596
rect 11336 3612 11388 3664
rect 11428 3612 11480 3664
rect 10600 3544 10652 3596
rect 10784 3476 10836 3528
rect 10968 3544 11020 3596
rect 11980 3544 12032 3596
rect 12624 3544 12676 3596
rect 11888 3476 11940 3528
rect 10232 3408 10284 3460
rect 11980 3408 12032 3460
rect 13084 3544 13136 3596
rect 13176 3476 13228 3528
rect 13912 3544 13964 3596
rect 14556 3544 14608 3596
rect 14924 3544 14976 3596
rect 15476 3587 15528 3596
rect 15476 3553 15485 3587
rect 15485 3553 15519 3587
rect 15519 3553 15528 3587
rect 15476 3544 15528 3553
rect 13084 3408 13136 3460
rect 13452 3408 13504 3460
rect 13636 3485 13645 3504
rect 13645 3485 13679 3504
rect 13679 3485 13688 3504
rect 13636 3452 13688 3485
rect 14004 3476 14056 3528
rect 14832 3476 14884 3528
rect 15292 3519 15344 3528
rect 15292 3485 15301 3519
rect 15301 3485 15335 3519
rect 15335 3485 15344 3519
rect 15292 3476 15344 3485
rect 8668 3340 8720 3392
rect 9128 3340 9180 3392
rect 9496 3383 9548 3392
rect 9496 3349 9505 3383
rect 9505 3349 9539 3383
rect 9539 3349 9548 3383
rect 9496 3340 9548 3349
rect 10416 3383 10468 3392
rect 10416 3349 10425 3383
rect 10425 3349 10459 3383
rect 10459 3349 10468 3383
rect 10784 3383 10836 3392
rect 10416 3340 10468 3349
rect 10784 3349 10793 3383
rect 10793 3349 10827 3383
rect 10827 3349 10836 3383
rect 10784 3340 10836 3349
rect 11888 3340 11940 3392
rect 12624 3340 12676 3392
rect 14372 3383 14424 3392
rect 14372 3349 14381 3383
rect 14381 3349 14415 3383
rect 14415 3349 14424 3383
rect 14372 3340 14424 3349
rect 14464 3383 14516 3392
rect 14464 3349 14473 3383
rect 14473 3349 14507 3383
rect 14507 3349 14516 3383
rect 14832 3383 14884 3392
rect 14464 3340 14516 3349
rect 14832 3349 14841 3383
rect 14841 3349 14875 3383
rect 14875 3349 14884 3383
rect 14832 3340 14884 3349
rect 15292 3340 15344 3392
rect 4698 3238 4750 3290
rect 4762 3238 4814 3290
rect 4826 3238 4878 3290
rect 4890 3238 4942 3290
rect 4954 3238 5006 3290
rect 8446 3238 8498 3290
rect 8510 3238 8562 3290
rect 8574 3238 8626 3290
rect 8638 3238 8690 3290
rect 8702 3238 8754 3290
rect 12194 3238 12246 3290
rect 12258 3238 12310 3290
rect 12322 3238 12374 3290
rect 12386 3238 12438 3290
rect 12450 3238 12502 3290
rect 3884 3136 3936 3188
rect 3976 3136 4028 3188
rect 1952 3000 2004 3052
rect 2964 3043 3016 3052
rect 2596 2932 2648 2984
rect 2964 3009 2973 3043
rect 2973 3009 3007 3043
rect 3007 3009 3016 3043
rect 2964 3000 3016 3009
rect 3240 2932 3292 2984
rect 3976 3000 4028 3052
rect 4252 3068 4304 3120
rect 4620 3136 4672 3188
rect 5908 3179 5960 3188
rect 5908 3145 5917 3179
rect 5917 3145 5951 3179
rect 5951 3145 5960 3179
rect 5908 3136 5960 3145
rect 6460 3136 6512 3188
rect 5264 3068 5316 3120
rect 6092 3068 6144 3120
rect 6552 3068 6604 3120
rect 7564 3136 7616 3188
rect 3700 2864 3752 2916
rect 4160 2932 4212 2984
rect 4528 2932 4580 2984
rect 5448 2932 5500 2984
rect 5264 2864 5316 2916
rect 5540 2864 5592 2916
rect 5816 2932 5868 2984
rect 6460 3000 6512 3052
rect 7012 3000 7064 3052
rect 7288 3000 7340 3052
rect 8208 3068 8260 3120
rect 7840 3000 7892 3052
rect 7932 3000 7984 3052
rect 8116 3043 8168 3052
rect 8116 3009 8125 3043
rect 8125 3009 8159 3043
rect 8159 3009 8168 3043
rect 8116 3000 8168 3009
rect 8392 3000 8444 3052
rect 8852 3000 8904 3052
rect 1492 2839 1544 2848
rect 1492 2805 1501 2839
rect 1501 2805 1535 2839
rect 1535 2805 1544 2839
rect 1492 2796 1544 2805
rect 1768 2796 1820 2848
rect 2044 2796 2096 2848
rect 2688 2796 2740 2848
rect 4252 2796 4304 2848
rect 6184 2796 6236 2848
rect 6828 2864 6880 2916
rect 8760 2975 8812 2984
rect 8760 2941 8769 2975
rect 8769 2941 8803 2975
rect 8803 2941 8812 2975
rect 8760 2932 8812 2941
rect 9496 3136 9548 3188
rect 10784 3136 10836 3188
rect 10968 3179 11020 3188
rect 10968 3145 10977 3179
rect 10977 3145 11011 3179
rect 11011 3145 11020 3179
rect 10968 3136 11020 3145
rect 11796 3136 11848 3188
rect 14740 3136 14792 3188
rect 9220 3000 9272 3052
rect 10692 3068 10744 3120
rect 10876 3068 10928 3120
rect 10048 3000 10100 3052
rect 12532 3068 12584 3120
rect 10508 2975 10560 2984
rect 9680 2907 9732 2916
rect 9680 2873 9689 2907
rect 9689 2873 9723 2907
rect 9723 2873 9732 2907
rect 10508 2941 10517 2975
rect 10517 2941 10551 2975
rect 10551 2941 10560 2975
rect 10508 2932 10560 2941
rect 11704 3000 11756 3052
rect 11152 2932 11204 2984
rect 12256 3000 12308 3052
rect 12900 3000 12952 3052
rect 12992 3000 13044 3052
rect 13176 2932 13228 2984
rect 13820 3000 13872 3052
rect 14096 3000 14148 3052
rect 14924 3000 14976 3052
rect 15200 3000 15252 3052
rect 9680 2864 9732 2873
rect 8208 2796 8260 2848
rect 8300 2796 8352 2848
rect 11336 2796 11388 2848
rect 11704 2796 11756 2848
rect 12256 2796 12308 2848
rect 12532 2864 12584 2916
rect 12808 2864 12860 2916
rect 13452 2864 13504 2916
rect 15476 2932 15528 2984
rect 13728 2796 13780 2848
rect 15660 2796 15712 2848
rect 2824 2694 2876 2746
rect 2888 2694 2940 2746
rect 2952 2694 3004 2746
rect 3016 2694 3068 2746
rect 3080 2694 3132 2746
rect 6572 2694 6624 2746
rect 6636 2694 6688 2746
rect 6700 2694 6752 2746
rect 6764 2694 6816 2746
rect 6828 2694 6880 2746
rect 10320 2694 10372 2746
rect 10384 2694 10436 2746
rect 10448 2694 10500 2746
rect 10512 2694 10564 2746
rect 10576 2694 10628 2746
rect 14068 2694 14120 2746
rect 14132 2694 14184 2746
rect 14196 2694 14248 2746
rect 14260 2694 14312 2746
rect 14324 2694 14376 2746
rect 3424 2592 3476 2644
rect 3792 2592 3844 2644
rect 6000 2592 6052 2644
rect 7196 2592 7248 2644
rect 7840 2592 7892 2644
rect 8300 2592 8352 2644
rect 9772 2592 9824 2644
rect 2596 2524 2648 2576
rect 3976 2524 4028 2576
rect 4068 2524 4120 2576
rect 4160 2524 4212 2576
rect 4712 2524 4764 2576
rect 5632 2524 5684 2576
rect 6460 2524 6512 2576
rect 7472 2524 7524 2576
rect 8208 2524 8260 2576
rect 8668 2524 8720 2576
rect 3332 2456 3384 2508
rect 2228 2388 2280 2440
rect 2504 2431 2556 2440
rect 2504 2397 2513 2431
rect 2513 2397 2547 2431
rect 2547 2397 2556 2431
rect 2504 2388 2556 2397
rect 2964 2388 3016 2440
rect 5264 2456 5316 2508
rect 12624 2592 12676 2644
rect 9956 2524 10008 2576
rect 10600 2524 10652 2576
rect 10784 2499 10836 2508
rect 3884 2388 3936 2440
rect 4068 2431 4120 2440
rect 4068 2397 4077 2431
rect 4077 2397 4111 2431
rect 4111 2397 4120 2431
rect 4068 2388 4120 2397
rect 4436 2431 4488 2440
rect 4436 2397 4445 2431
rect 4445 2397 4479 2431
rect 4479 2397 4488 2431
rect 4436 2388 4488 2397
rect 4896 2431 4948 2440
rect 4896 2397 4905 2431
rect 4905 2397 4939 2431
rect 4939 2397 4948 2431
rect 4896 2388 4948 2397
rect 5172 2388 5224 2440
rect 5816 2431 5868 2440
rect 5816 2397 5825 2431
rect 5825 2397 5859 2431
rect 5859 2397 5868 2431
rect 5816 2388 5868 2397
rect 2228 2252 2280 2304
rect 4344 2320 4396 2372
rect 3792 2252 3844 2304
rect 5264 2320 5316 2372
rect 6276 2388 6328 2440
rect 6828 2388 6880 2440
rect 7288 2431 7340 2440
rect 7288 2397 7297 2431
rect 7297 2397 7331 2431
rect 7331 2397 7340 2431
rect 7288 2388 7340 2397
rect 8300 2431 8352 2440
rect 7472 2320 7524 2372
rect 7656 2320 7708 2372
rect 7748 2320 7800 2372
rect 5448 2295 5500 2304
rect 5448 2261 5457 2295
rect 5457 2261 5491 2295
rect 5491 2261 5500 2295
rect 5448 2252 5500 2261
rect 5908 2252 5960 2304
rect 6460 2252 6512 2304
rect 6736 2295 6788 2304
rect 6736 2261 6745 2295
rect 6745 2261 6779 2295
rect 6779 2261 6788 2295
rect 6736 2252 6788 2261
rect 7012 2252 7064 2304
rect 7932 2295 7984 2304
rect 7932 2261 7941 2295
rect 7941 2261 7975 2295
rect 7975 2261 7984 2295
rect 7932 2252 7984 2261
rect 8300 2397 8309 2431
rect 8309 2397 8343 2431
rect 8343 2397 8352 2431
rect 8300 2388 8352 2397
rect 8944 2388 8996 2440
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 9404 2431 9456 2440
rect 9404 2397 9413 2431
rect 9413 2397 9447 2431
rect 9447 2397 9456 2431
rect 9404 2388 9456 2397
rect 9588 2431 9640 2440
rect 9588 2397 9597 2431
rect 9597 2397 9631 2431
rect 9631 2397 9640 2431
rect 9588 2388 9640 2397
rect 9864 2431 9916 2440
rect 9864 2397 9873 2431
rect 9873 2397 9907 2431
rect 9907 2397 9916 2431
rect 9864 2388 9916 2397
rect 10784 2465 10793 2499
rect 10793 2465 10827 2499
rect 10827 2465 10836 2499
rect 10784 2456 10836 2465
rect 11796 2499 11848 2508
rect 11796 2465 11805 2499
rect 11805 2465 11839 2499
rect 11839 2465 11848 2499
rect 11796 2456 11848 2465
rect 11888 2456 11940 2508
rect 13728 2592 13780 2644
rect 13820 2524 13872 2576
rect 14464 2524 14516 2576
rect 13176 2456 13228 2508
rect 14372 2499 14424 2508
rect 14372 2465 14381 2499
rect 14381 2465 14415 2499
rect 14415 2465 14424 2499
rect 14372 2456 14424 2465
rect 8208 2320 8260 2372
rect 8668 2363 8720 2372
rect 8668 2329 8677 2363
rect 8677 2329 8711 2363
rect 8711 2329 8720 2363
rect 8668 2320 8720 2329
rect 10140 2320 10192 2372
rect 10324 2320 10376 2372
rect 11244 2388 11296 2440
rect 11612 2388 11664 2440
rect 10784 2320 10836 2372
rect 12072 2320 12124 2372
rect 12808 2388 12860 2440
rect 13636 2388 13688 2440
rect 15016 2431 15068 2440
rect 15016 2397 15025 2431
rect 15025 2397 15059 2431
rect 15059 2397 15068 2431
rect 15016 2388 15068 2397
rect 15384 2431 15436 2440
rect 15384 2397 15393 2431
rect 15393 2397 15427 2431
rect 15427 2397 15436 2431
rect 15384 2388 15436 2397
rect 9680 2252 9732 2304
rect 14556 2320 14608 2372
rect 13728 2295 13780 2304
rect 13728 2261 13737 2295
rect 13737 2261 13771 2295
rect 13771 2261 13780 2295
rect 13728 2252 13780 2261
rect 14188 2252 14240 2304
rect 4698 2150 4750 2202
rect 4762 2150 4814 2202
rect 4826 2150 4878 2202
rect 4890 2150 4942 2202
rect 4954 2150 5006 2202
rect 8446 2150 8498 2202
rect 8510 2150 8562 2202
rect 8574 2150 8626 2202
rect 8638 2150 8690 2202
rect 8702 2150 8754 2202
rect 12194 2150 12246 2202
rect 12258 2150 12310 2202
rect 12322 2150 12374 2202
rect 12386 2150 12438 2202
rect 12450 2150 12502 2202
rect 3792 2048 3844 2100
rect 5172 2048 5224 2100
rect 6276 2048 6328 2100
rect 4068 1980 4120 2032
rect 7104 1980 7156 2032
rect 4160 1912 4212 1964
rect 5632 1912 5684 1964
rect 6000 1912 6052 1964
rect 9404 1980 9456 2032
rect 9588 1980 9640 2032
rect 13728 1980 13780 2032
rect 7288 1912 7340 1964
rect 16028 1912 16080 1964
rect 4436 1844 4488 1896
rect 9312 1844 9364 1896
rect 12256 1844 12308 1896
rect 13176 1844 13228 1896
rect 2964 1776 3016 1828
rect 7380 1776 7432 1828
rect 5540 1708 5592 1760
rect 7932 1708 7984 1760
rect 11152 1708 11204 1760
rect 11612 1708 11664 1760
rect 3516 1640 3568 1692
rect 8208 1640 8260 1692
rect 5448 1572 5500 1624
rect 9220 1572 9272 1624
rect 6920 1300 6972 1352
rect 7840 1300 7892 1352
<< metal2 >>
rect 294 19200 350 20000
rect 662 19200 718 20000
rect 1030 19200 1086 20000
rect 1136 19230 1348 19258
rect 308 16590 336 19200
rect 296 16584 348 16590
rect 296 16526 348 16532
rect 676 16046 704 19200
rect 1044 19122 1072 19200
rect 1136 19122 1164 19230
rect 1044 19094 1164 19122
rect 1320 17320 1348 19230
rect 1398 19200 1454 20000
rect 1766 19200 1822 20000
rect 2134 19200 2190 20000
rect 2502 19200 2558 20000
rect 2870 19200 2926 20000
rect 3238 19200 3294 20000
rect 3606 19200 3662 20000
rect 3974 19200 4030 20000
rect 4342 19200 4398 20000
rect 4710 19200 4766 20000
rect 5078 19200 5134 20000
rect 5446 19200 5502 20000
rect 5814 19200 5870 20000
rect 6182 19200 6238 20000
rect 6550 19200 6606 20000
rect 6918 19200 6974 20000
rect 7286 19200 7342 20000
rect 7654 19200 7710 20000
rect 8022 19200 8078 20000
rect 8390 19200 8446 20000
rect 8758 19200 8814 20000
rect 9126 19200 9182 20000
rect 9494 19200 9550 20000
rect 9862 19200 9918 20000
rect 9968 19230 10180 19258
rect 1412 19122 1440 19200
rect 1412 19094 1624 19122
rect 1490 19000 1546 19009
rect 1490 18935 1546 18944
rect 1400 17332 1452 17338
rect 1320 17292 1400 17320
rect 1400 17274 1452 17280
rect 1504 16590 1532 18935
rect 1492 16584 1544 16590
rect 1492 16526 1544 16532
rect 1596 16454 1624 19094
rect 1780 17184 1808 19200
rect 1858 18048 1914 18057
rect 1858 17983 1914 17992
rect 1688 17156 1808 17184
rect 1688 17066 1716 17156
rect 1676 17060 1728 17066
rect 1676 17002 1728 17008
rect 1768 16720 1820 16726
rect 1768 16662 1820 16668
rect 1780 16590 1808 16662
rect 1768 16584 1820 16590
rect 1768 16526 1820 16532
rect 1584 16448 1636 16454
rect 1584 16390 1636 16396
rect 1872 16250 1900 17983
rect 2044 17196 2096 17202
rect 2044 17138 2096 17144
rect 2056 17105 2084 17138
rect 2042 17096 2098 17105
rect 2042 17031 2098 17040
rect 2148 16998 2176 19200
rect 2516 17320 2544 19200
rect 2424 17292 2544 17320
rect 2320 17264 2372 17270
rect 2320 17206 2372 17212
rect 2136 16992 2188 16998
rect 2136 16934 2188 16940
rect 2134 16552 2190 16561
rect 2044 16516 2096 16522
rect 2134 16487 2190 16496
rect 2044 16458 2096 16464
rect 1492 16244 1544 16250
rect 1492 16186 1544 16192
rect 1860 16244 1912 16250
rect 1860 16186 1912 16192
rect 1504 16153 1532 16186
rect 1490 16144 1546 16153
rect 1490 16079 1546 16088
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 664 16040 716 16046
rect 664 15982 716 15988
rect 1492 15360 1544 15366
rect 1492 15302 1544 15308
rect 1504 15201 1532 15302
rect 1490 15192 1546 15201
rect 1490 15127 1546 15136
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 1676 14952 1728 14958
rect 1676 14894 1728 14900
rect 1412 11014 1440 14894
rect 1492 14272 1544 14278
rect 1490 14240 1492 14249
rect 1544 14240 1546 14249
rect 1490 14175 1546 14184
rect 1688 14074 1716 14894
rect 1780 14618 1808 16050
rect 2056 15042 2084 16458
rect 2148 16114 2176 16487
rect 2332 16250 2360 17206
rect 2424 16998 2452 17292
rect 2504 17196 2556 17202
rect 2504 17138 2556 17144
rect 2412 16992 2464 16998
rect 2412 16934 2464 16940
rect 2412 16584 2464 16590
rect 2412 16526 2464 16532
rect 2320 16244 2372 16250
rect 2320 16186 2372 16192
rect 2136 16108 2188 16114
rect 2136 16050 2188 16056
rect 2148 15162 2176 16050
rect 2320 15904 2372 15910
rect 2320 15846 2372 15852
rect 2332 15434 2360 15846
rect 2320 15428 2372 15434
rect 2320 15370 2372 15376
rect 2228 15360 2280 15366
rect 2226 15328 2228 15337
rect 2424 15337 2452 16526
rect 2280 15328 2282 15337
rect 2410 15328 2466 15337
rect 2282 15286 2360 15314
rect 2226 15263 2282 15272
rect 2136 15156 2188 15162
rect 2136 15098 2188 15104
rect 2056 15014 2268 15042
rect 1860 14884 1912 14890
rect 1860 14826 1912 14832
rect 1768 14612 1820 14618
rect 1768 14554 1820 14560
rect 1768 14408 1820 14414
rect 1768 14350 1820 14356
rect 1780 14074 1808 14350
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 1768 14068 1820 14074
rect 1768 14010 1820 14016
rect 1872 13326 1900 14826
rect 2044 14816 2096 14822
rect 2044 14758 2096 14764
rect 1950 14512 2006 14521
rect 1950 14447 2006 14456
rect 1964 14414 1992 14447
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 1860 13320 1912 13326
rect 1490 13288 1546 13297
rect 1490 13223 1546 13232
rect 1766 13288 1822 13297
rect 1860 13262 1912 13268
rect 1766 13223 1822 13232
rect 1504 13190 1532 13223
rect 1492 13184 1544 13190
rect 1492 13126 1544 13132
rect 1584 12844 1636 12850
rect 1584 12786 1636 12792
rect 1492 12640 1544 12646
rect 1492 12582 1544 12588
rect 1504 12345 1532 12582
rect 1490 12336 1546 12345
rect 1490 12271 1546 12280
rect 1492 11552 1544 11558
rect 1492 11494 1544 11500
rect 1504 11393 1532 11494
rect 1490 11384 1546 11393
rect 1596 11354 1624 12786
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1688 11762 1716 12582
rect 1780 12238 1808 13223
rect 1952 12844 2004 12850
rect 1952 12786 2004 12792
rect 1964 12442 1992 12786
rect 1952 12436 2004 12442
rect 1952 12378 2004 12384
rect 1768 12232 1820 12238
rect 1768 12174 1820 12180
rect 1860 12164 1912 12170
rect 1860 12106 1912 12112
rect 1676 11756 1728 11762
rect 1676 11698 1728 11704
rect 1490 11319 1546 11328
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 1400 11008 1452 11014
rect 1400 10950 1452 10956
rect 1490 10432 1546 10441
rect 1490 10367 1546 10376
rect 1504 10266 1532 10367
rect 1492 10260 1544 10266
rect 1492 10202 1544 10208
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1688 9722 1716 9998
rect 1676 9716 1728 9722
rect 1676 9658 1728 9664
rect 1768 9580 1820 9586
rect 1768 9522 1820 9528
rect 1490 9480 1546 9489
rect 1490 9415 1492 9424
rect 1544 9415 1546 9424
rect 1492 9386 1544 9392
rect 1780 9178 1808 9522
rect 1768 9172 1820 9178
rect 1768 9114 1820 9120
rect 1872 9058 1900 12106
rect 2056 10674 2084 14758
rect 2240 14414 2268 15014
rect 2228 14408 2280 14414
rect 2228 14350 2280 14356
rect 2240 13530 2268 14350
rect 2332 14006 2360 15286
rect 2410 15263 2466 15272
rect 2516 15162 2544 17138
rect 2596 17128 2648 17134
rect 2596 17070 2648 17076
rect 2504 15156 2556 15162
rect 2504 15098 2556 15104
rect 2410 15056 2466 15065
rect 2410 14991 2412 15000
rect 2464 14991 2466 15000
rect 2504 15020 2556 15026
rect 2412 14962 2464 14968
rect 2504 14962 2556 14968
rect 2320 14000 2372 14006
rect 2320 13942 2372 13948
rect 2410 13968 2466 13977
rect 2410 13903 2412 13912
rect 2464 13903 2466 13912
rect 2412 13874 2464 13880
rect 2320 13728 2372 13734
rect 2516 13716 2544 14962
rect 2608 14074 2636 17070
rect 2884 16998 2912 19200
rect 3252 17066 3280 19200
rect 3332 17196 3384 17202
rect 3332 17138 3384 17144
rect 3240 17060 3292 17066
rect 3240 17002 3292 17008
rect 2872 16992 2924 16998
rect 2872 16934 2924 16940
rect 2824 16892 3132 16901
rect 2824 16890 2830 16892
rect 2886 16890 2910 16892
rect 2966 16890 2990 16892
rect 3046 16890 3070 16892
rect 3126 16890 3132 16892
rect 2886 16838 2888 16890
rect 3068 16838 3070 16890
rect 2824 16836 2830 16838
rect 2886 16836 2910 16838
rect 2966 16836 2990 16838
rect 3046 16836 3070 16838
rect 3126 16836 3132 16838
rect 2824 16827 3132 16836
rect 3056 16584 3108 16590
rect 3056 16526 3108 16532
rect 3148 16584 3200 16590
rect 3148 16526 3200 16532
rect 2688 16516 2740 16522
rect 2688 16458 2740 16464
rect 2700 15609 2728 16458
rect 2872 16448 2924 16454
rect 2872 16390 2924 16396
rect 2884 16046 2912 16390
rect 3068 16153 3096 16526
rect 3054 16144 3110 16153
rect 3054 16079 3110 16088
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 2824 15804 3132 15813
rect 2824 15802 2830 15804
rect 2886 15802 2910 15804
rect 2966 15802 2990 15804
rect 3046 15802 3070 15804
rect 3126 15802 3132 15804
rect 2886 15750 2888 15802
rect 3068 15750 3070 15802
rect 2824 15748 2830 15750
rect 2886 15748 2910 15750
rect 2966 15748 2990 15750
rect 3046 15748 3070 15750
rect 3126 15748 3132 15750
rect 2824 15739 3132 15748
rect 2686 15600 2742 15609
rect 2686 15535 2742 15544
rect 3160 15434 3188 16526
rect 3344 16250 3372 17138
rect 3424 17128 3476 17134
rect 3424 17070 3476 17076
rect 3332 16244 3384 16250
rect 3332 16186 3384 16192
rect 3240 16108 3292 16114
rect 3240 16050 3292 16056
rect 2780 15428 2832 15434
rect 2780 15370 2832 15376
rect 3148 15428 3200 15434
rect 3148 15370 3200 15376
rect 2792 15026 2820 15370
rect 2780 15020 2832 15026
rect 2700 14980 2780 15008
rect 2700 14464 2728 14980
rect 2780 14962 2832 14968
rect 2824 14716 3132 14725
rect 2824 14714 2830 14716
rect 2886 14714 2910 14716
rect 2966 14714 2990 14716
rect 3046 14714 3070 14716
rect 3126 14714 3132 14716
rect 2886 14662 2888 14714
rect 3068 14662 3070 14714
rect 2824 14660 2830 14662
rect 2886 14660 2910 14662
rect 2966 14660 2990 14662
rect 3046 14660 3070 14662
rect 3126 14660 3132 14662
rect 2824 14651 3132 14660
rect 2872 14476 2924 14482
rect 2700 14436 2872 14464
rect 2872 14418 2924 14424
rect 3148 14476 3200 14482
rect 3148 14418 3200 14424
rect 2780 14340 2832 14346
rect 2780 14282 2832 14288
rect 2596 14068 2648 14074
rect 2596 14010 2648 14016
rect 2792 13870 2820 14282
rect 2870 14240 2926 14249
rect 2870 14175 2926 14184
rect 2884 14074 2912 14175
rect 3160 14074 3188 14418
rect 3252 14278 3280 16050
rect 3436 15978 3464 17070
rect 3620 17066 3648 19200
rect 3792 17196 3844 17202
rect 3792 17138 3844 17144
rect 3884 17196 3936 17202
rect 3884 17138 3936 17144
rect 3608 17060 3660 17066
rect 3608 17002 3660 17008
rect 3804 16726 3832 17138
rect 3792 16720 3844 16726
rect 3792 16662 3844 16668
rect 3792 16584 3844 16590
rect 3792 16526 3844 16532
rect 3608 16108 3660 16114
rect 3608 16050 3660 16056
rect 3424 15972 3476 15978
rect 3424 15914 3476 15920
rect 3620 15910 3648 16050
rect 3700 16040 3752 16046
rect 3700 15982 3752 15988
rect 3608 15904 3660 15910
rect 3608 15846 3660 15852
rect 3516 15428 3568 15434
rect 3516 15370 3568 15376
rect 3424 14816 3476 14822
rect 3344 14776 3424 14804
rect 3240 14272 3292 14278
rect 3240 14214 3292 14220
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 3148 14068 3200 14074
rect 3148 14010 3200 14016
rect 2884 13938 2912 14010
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2372 13688 2544 13716
rect 2320 13670 2372 13676
rect 2228 13524 2280 13530
rect 2228 13466 2280 13472
rect 2136 12096 2188 12102
rect 2136 12038 2188 12044
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 2148 10538 2176 12038
rect 2136 10532 2188 10538
rect 2136 10474 2188 10480
rect 2228 9920 2280 9926
rect 2228 9862 2280 9868
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 1596 9030 1900 9058
rect 1492 8832 1544 8838
rect 1492 8774 1544 8780
rect 1504 8537 1532 8774
rect 1490 8528 1546 8537
rect 1490 8463 1546 8472
rect 1490 7576 1546 7585
rect 1490 7511 1492 7520
rect 1544 7511 1546 7520
rect 1492 7482 1544 7488
rect 1492 6656 1544 6662
rect 1490 6624 1492 6633
rect 1544 6624 1546 6633
rect 1490 6559 1546 6568
rect 1400 6112 1452 6118
rect 1400 6054 1452 6060
rect 1412 4622 1440 6054
rect 1490 5672 1546 5681
rect 1490 5607 1546 5616
rect 1504 5574 1532 5607
rect 1492 5568 1544 5574
rect 1492 5510 1544 5516
rect 1492 5024 1544 5030
rect 1492 4966 1544 4972
rect 1504 4729 1532 4966
rect 1596 4758 1624 9030
rect 1768 8968 1820 8974
rect 1952 8968 2004 8974
rect 1768 8910 1820 8916
rect 1858 8936 1914 8945
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 1688 6458 1716 7686
rect 1780 7546 1808 8910
rect 1952 8910 2004 8916
rect 1858 8871 1914 8880
rect 1872 8634 1900 8871
rect 1964 8634 1992 8910
rect 2044 8900 2096 8906
rect 2044 8842 2096 8848
rect 1860 8628 1912 8634
rect 1860 8570 1912 8576
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 1950 8392 2006 8401
rect 1950 8327 2006 8336
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 1964 7410 1992 8327
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1780 5914 1808 7346
rect 1952 6860 2004 6866
rect 2056 6848 2084 8842
rect 2148 8090 2176 9522
rect 2240 8906 2268 9862
rect 2332 9722 2360 13670
rect 2824 13628 3132 13637
rect 2824 13626 2830 13628
rect 2886 13626 2910 13628
rect 2966 13626 2990 13628
rect 3046 13626 3070 13628
rect 3126 13626 3132 13628
rect 2886 13574 2888 13626
rect 3068 13574 3070 13626
rect 2824 13572 2830 13574
rect 2886 13572 2910 13574
rect 2966 13572 2990 13574
rect 3046 13572 3070 13574
rect 3126 13572 3132 13574
rect 2824 13563 3132 13572
rect 3160 12986 3188 14010
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 2824 12540 3132 12549
rect 2824 12538 2830 12540
rect 2886 12538 2910 12540
rect 2966 12538 2990 12540
rect 3046 12538 3070 12540
rect 3126 12538 3132 12540
rect 2886 12486 2888 12538
rect 3068 12486 3070 12538
rect 2824 12484 2830 12486
rect 2886 12484 2910 12486
rect 2966 12484 2990 12486
rect 3046 12484 3070 12486
rect 3126 12484 3132 12486
rect 2824 12475 3132 12484
rect 3160 12442 3188 12922
rect 3252 12442 3280 14214
rect 2596 12436 2648 12442
rect 2596 12378 2648 12384
rect 3148 12436 3200 12442
rect 3148 12378 3200 12384
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 2608 11694 2636 12378
rect 2596 11688 2648 11694
rect 2516 11648 2596 11676
rect 2516 11354 2544 11648
rect 2596 11630 2648 11636
rect 2824 11452 3132 11461
rect 2824 11450 2830 11452
rect 2886 11450 2910 11452
rect 2966 11450 2990 11452
rect 3046 11450 3070 11452
rect 3126 11450 3132 11452
rect 2886 11398 2888 11450
rect 3068 11398 3070 11450
rect 2824 11396 2830 11398
rect 2886 11396 2910 11398
rect 2966 11396 2990 11398
rect 3046 11396 3070 11398
rect 3126 11396 3132 11398
rect 2824 11387 3132 11396
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 2872 11008 2924 11014
rect 2872 10950 2924 10956
rect 2884 10606 2912 10950
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 3160 10470 3188 10746
rect 3252 10577 3280 11086
rect 3238 10568 3294 10577
rect 3238 10503 3294 10512
rect 3148 10464 3200 10470
rect 3200 10424 3280 10452
rect 3148 10406 3200 10412
rect 2824 10364 3132 10373
rect 2824 10362 2830 10364
rect 2886 10362 2910 10364
rect 2966 10362 2990 10364
rect 3046 10362 3070 10364
rect 3126 10362 3132 10364
rect 2886 10310 2888 10362
rect 3068 10310 3070 10362
rect 2824 10308 2830 10310
rect 2886 10308 2910 10310
rect 2966 10308 2990 10310
rect 3046 10308 3070 10310
rect 3126 10308 3132 10310
rect 2824 10299 3132 10308
rect 2320 9716 2372 9722
rect 2320 9658 2372 9664
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 2824 9276 3132 9285
rect 2824 9274 2830 9276
rect 2886 9274 2910 9276
rect 2966 9274 2990 9276
rect 3046 9274 3070 9276
rect 3126 9274 3132 9276
rect 2886 9222 2888 9274
rect 3068 9222 3070 9274
rect 2824 9220 2830 9222
rect 2886 9220 2910 9222
rect 2966 9220 2990 9222
rect 3046 9220 3070 9222
rect 3126 9220 3132 9222
rect 2824 9211 3132 9220
rect 3160 9178 3188 9318
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 2228 8900 2280 8906
rect 2228 8842 2280 8848
rect 2320 8832 2372 8838
rect 2320 8774 2372 8780
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 2004 6820 2084 6848
rect 1952 6802 2004 6808
rect 1768 5908 1820 5914
rect 1768 5850 1820 5856
rect 1676 5228 1728 5234
rect 1676 5170 1728 5176
rect 1688 4826 1716 5170
rect 1964 5166 1992 6802
rect 2226 6760 2282 6769
rect 2226 6695 2228 6704
rect 2280 6695 2282 6704
rect 2228 6666 2280 6672
rect 2332 6254 2360 8774
rect 2412 8288 2464 8294
rect 2412 8230 2464 8236
rect 2424 7868 2452 8230
rect 2824 8188 3132 8197
rect 2824 8186 2830 8188
rect 2886 8186 2910 8188
rect 2966 8186 2990 8188
rect 3046 8186 3070 8188
rect 3126 8186 3132 8188
rect 2886 8134 2888 8186
rect 3068 8134 3070 8186
rect 2824 8132 2830 8134
rect 2886 8132 2910 8134
rect 2966 8132 2990 8134
rect 3046 8132 3070 8134
rect 3126 8132 3132 8134
rect 2824 8123 3132 8132
rect 2495 7880 2547 7886
rect 2424 7840 2495 7868
rect 2044 6248 2096 6254
rect 2044 6190 2096 6196
rect 2320 6248 2372 6254
rect 2320 6190 2372 6196
rect 2056 5914 2084 6190
rect 2044 5908 2096 5914
rect 2044 5850 2096 5856
rect 2226 5808 2282 5817
rect 2136 5772 2188 5778
rect 2226 5743 2282 5752
rect 2136 5714 2188 5720
rect 1952 5160 2004 5166
rect 1952 5102 2004 5108
rect 1860 5024 1912 5030
rect 1860 4966 1912 4972
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1584 4752 1636 4758
rect 1490 4720 1546 4729
rect 1584 4694 1636 4700
rect 1490 4655 1546 4664
rect 1400 4616 1452 4622
rect 1400 4558 1452 4564
rect 1412 921 1440 4558
rect 1872 4282 1900 4966
rect 1964 4282 1992 5102
rect 2044 4480 2096 4486
rect 2044 4422 2096 4428
rect 1860 4276 1912 4282
rect 1860 4218 1912 4224
rect 1952 4276 2004 4282
rect 1952 4218 2004 4224
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 1768 4072 1820 4078
rect 1766 4040 1768 4049
rect 1820 4040 1822 4049
rect 1766 3975 1822 3984
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 1490 3768 1546 3777
rect 1490 3703 1492 3712
rect 1544 3703 1546 3712
rect 1492 3674 1544 3680
rect 1688 3534 1716 3878
rect 1676 3528 1728 3534
rect 1964 3505 1992 4082
rect 2056 3534 2084 4422
rect 2148 3534 2176 5714
rect 2240 5642 2268 5743
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 2228 5636 2280 5642
rect 2228 5578 2280 5584
rect 2226 5128 2282 5137
rect 2332 5098 2360 5646
rect 2226 5063 2282 5072
rect 2320 5092 2372 5098
rect 2240 4622 2268 5063
rect 2320 5034 2372 5040
rect 2424 4978 2452 7840
rect 2495 7822 2547 7828
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 2824 7100 3132 7109
rect 2824 7098 2830 7100
rect 2886 7098 2910 7100
rect 2966 7098 2990 7100
rect 3046 7098 3070 7100
rect 3126 7098 3132 7100
rect 2886 7046 2888 7098
rect 3068 7046 3070 7098
rect 2824 7044 2830 7046
rect 2886 7044 2910 7046
rect 2966 7044 2990 7046
rect 3046 7044 3070 7046
rect 3126 7044 3132 7046
rect 2824 7035 3132 7044
rect 2596 6928 2648 6934
rect 2596 6870 2648 6876
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2516 5386 2544 6598
rect 2608 5642 2636 6870
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2596 5636 2648 5642
rect 2596 5578 2648 5584
rect 2516 5358 2636 5386
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 2332 4950 2452 4978
rect 2332 4729 2360 4950
rect 2410 4856 2466 4865
rect 2410 4791 2412 4800
rect 2464 4791 2466 4800
rect 2412 4762 2464 4768
rect 2318 4720 2374 4729
rect 2318 4655 2374 4664
rect 2228 4616 2280 4622
rect 2228 4558 2280 4564
rect 2412 4548 2464 4554
rect 2412 4490 2464 4496
rect 2320 4276 2372 4282
rect 2320 4218 2372 4224
rect 2044 3528 2096 3534
rect 1676 3470 1728 3476
rect 1950 3496 2006 3505
rect 2044 3470 2096 3476
rect 2136 3528 2188 3534
rect 2136 3470 2188 3476
rect 1950 3431 2006 3440
rect 1860 3392 1912 3398
rect 1860 3334 1912 3340
rect 1952 3392 2004 3398
rect 1952 3334 2004 3340
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 1492 2848 1544 2854
rect 1490 2816 1492 2825
rect 1768 2848 1820 2854
rect 1544 2816 1546 2825
rect 1768 2790 1820 2796
rect 1490 2751 1546 2760
rect 1398 912 1454 921
rect 1398 847 1454 856
rect 1780 800 1808 2790
rect 1872 1873 1900 3334
rect 1964 3058 1992 3334
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 2044 2848 2096 2854
rect 2044 2790 2096 2796
rect 1858 1864 1914 1873
rect 1858 1799 1914 1808
rect 2056 800 2084 2790
rect 2240 2446 2268 3334
rect 2332 2961 2360 4218
rect 2318 2952 2374 2961
rect 2318 2887 2374 2896
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 2228 2304 2280 2310
rect 2280 2264 2360 2292
rect 2228 2246 2280 2252
rect 2332 800 2360 2264
rect 2424 2009 2452 4490
rect 2516 4486 2544 5170
rect 2608 4826 2636 5358
rect 2700 5302 2728 6598
rect 3160 6186 3188 7142
rect 3148 6180 3200 6186
rect 3148 6122 3200 6128
rect 2824 6012 3132 6021
rect 2824 6010 2830 6012
rect 2886 6010 2910 6012
rect 2966 6010 2990 6012
rect 3046 6010 3070 6012
rect 3126 6010 3132 6012
rect 2886 5958 2888 6010
rect 3068 5958 3070 6010
rect 2824 5956 2830 5958
rect 2886 5956 2910 5958
rect 2966 5956 2990 5958
rect 3046 5956 3070 5958
rect 3126 5956 3132 5958
rect 2824 5947 3132 5956
rect 3160 5846 3188 6122
rect 3148 5840 3200 5846
rect 3148 5782 3200 5788
rect 2688 5296 2740 5302
rect 2688 5238 2740 5244
rect 3148 5024 3200 5030
rect 3148 4966 3200 4972
rect 2824 4924 3132 4933
rect 2824 4922 2830 4924
rect 2886 4922 2910 4924
rect 2966 4922 2990 4924
rect 3046 4922 3070 4924
rect 3126 4922 3132 4924
rect 2886 4870 2888 4922
rect 3068 4870 3070 4922
rect 2824 4868 2830 4870
rect 2886 4868 2910 4870
rect 2966 4868 2990 4870
rect 3046 4868 3070 4870
rect 3126 4868 3132 4870
rect 2824 4859 3132 4868
rect 2596 4820 2648 4826
rect 2596 4762 2648 4768
rect 2596 4684 2648 4690
rect 2596 4626 2648 4632
rect 2504 4480 2556 4486
rect 2504 4422 2556 4428
rect 2608 4026 2636 4626
rect 2688 4548 2740 4554
rect 2688 4490 2740 4496
rect 2516 3998 2636 4026
rect 2516 3738 2544 3998
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 2516 2446 2544 3334
rect 2608 2990 2636 3878
rect 2700 3602 2728 4490
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 3068 4282 3096 4422
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 2870 4176 2926 4185
rect 2870 4111 2872 4120
rect 2924 4111 2926 4120
rect 2872 4082 2924 4088
rect 2824 3836 3132 3845
rect 2824 3834 2830 3836
rect 2886 3834 2910 3836
rect 2966 3834 2990 3836
rect 3046 3834 3070 3836
rect 3126 3834 3132 3836
rect 2886 3782 2888 3834
rect 3068 3782 3070 3834
rect 2824 3780 2830 3782
rect 2886 3780 2910 3782
rect 2966 3780 2990 3782
rect 3046 3780 3070 3782
rect 3126 3780 3132 3782
rect 2824 3771 3132 3780
rect 3056 3664 3108 3670
rect 2870 3632 2926 3641
rect 2688 3596 2740 3602
rect 3056 3606 3108 3612
rect 2870 3567 2926 3576
rect 2688 3538 2740 3544
rect 2884 3534 2912 3567
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 2976 3058 3004 3334
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 2688 2848 2740 2854
rect 3068 2836 3096 3606
rect 3160 3534 3188 4966
rect 3252 4554 3280 10424
rect 3344 4758 3372 14776
rect 3424 14758 3476 14764
rect 3424 12436 3476 12442
rect 3424 12378 3476 12384
rect 3436 6934 3464 12378
rect 3528 9110 3556 15370
rect 3620 13394 3648 15846
rect 3608 13388 3660 13394
rect 3608 13330 3660 13336
rect 3712 12434 3740 15982
rect 3804 14550 3832 16526
rect 3896 16454 3924 17138
rect 3988 17066 4016 19200
rect 4356 17354 4384 19200
rect 4724 17524 4752 19200
rect 4632 17496 4752 17524
rect 4356 17326 4476 17354
rect 4344 17196 4396 17202
rect 4344 17138 4396 17144
rect 3976 17060 4028 17066
rect 3976 17002 4028 17008
rect 4356 16726 4384 17138
rect 4344 16720 4396 16726
rect 4344 16662 4396 16668
rect 4068 16584 4120 16590
rect 4252 16584 4304 16590
rect 4120 16544 4200 16572
rect 4068 16526 4120 16532
rect 3884 16448 3936 16454
rect 3884 16390 3936 16396
rect 4068 16176 4120 16182
rect 4068 16118 4120 16124
rect 3884 15904 3936 15910
rect 3882 15872 3884 15881
rect 3936 15872 3938 15881
rect 3882 15807 3938 15816
rect 3976 15564 4028 15570
rect 3976 15506 4028 15512
rect 3884 15360 3936 15366
rect 3884 15302 3936 15308
rect 3792 14544 3844 14550
rect 3792 14486 3844 14492
rect 3804 12646 3832 14486
rect 3896 14006 3924 15302
rect 3884 14000 3936 14006
rect 3884 13942 3936 13948
rect 3792 12640 3844 12646
rect 3792 12582 3844 12588
rect 3620 12406 3740 12434
rect 3516 9104 3568 9110
rect 3516 9046 3568 9052
rect 3424 6928 3476 6934
rect 3476 6888 3556 6916
rect 3424 6870 3476 6876
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 3436 5846 3464 6734
rect 3528 6390 3556 6888
rect 3620 6662 3648 12406
rect 3804 11234 3832 12582
rect 3896 12434 3924 13942
rect 3988 13938 4016 15506
rect 4080 14278 4108 16118
rect 4172 15094 4200 16544
rect 4252 16526 4304 16532
rect 4264 16250 4292 16526
rect 4448 16454 4476 17326
rect 4632 17066 4660 17496
rect 4698 17436 5006 17445
rect 4698 17434 4704 17436
rect 4760 17434 4784 17436
rect 4840 17434 4864 17436
rect 4920 17434 4944 17436
rect 5000 17434 5006 17436
rect 4760 17382 4762 17434
rect 4942 17382 4944 17434
rect 4698 17380 4704 17382
rect 4760 17380 4784 17382
rect 4840 17380 4864 17382
rect 4920 17380 4944 17382
rect 5000 17380 5006 17382
rect 4698 17371 5006 17380
rect 4620 17060 4672 17066
rect 4620 17002 4672 17008
rect 5092 16454 5120 19200
rect 5460 17270 5488 19200
rect 5448 17264 5500 17270
rect 5448 17206 5500 17212
rect 5630 17232 5686 17241
rect 5172 17196 5224 17202
rect 5630 17167 5632 17176
rect 5172 17138 5224 17144
rect 5684 17167 5686 17176
rect 5632 17138 5684 17144
rect 4344 16448 4396 16454
rect 4344 16390 4396 16396
rect 4436 16448 4488 16454
rect 4712 16448 4764 16454
rect 4436 16390 4488 16396
rect 4632 16408 4712 16436
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 4160 15088 4212 15094
rect 4160 15030 4212 15036
rect 4252 15020 4304 15026
rect 4252 14962 4304 14968
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 4068 14272 4120 14278
rect 4066 14240 4068 14249
rect 4120 14240 4122 14249
rect 4066 14175 4122 14184
rect 3976 13932 4028 13938
rect 3976 13874 4028 13880
rect 4172 13530 4200 14418
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4160 13388 4212 13394
rect 4160 13330 4212 13336
rect 4172 12458 4200 13330
rect 4264 13190 4292 14962
rect 4356 14822 4384 16390
rect 4632 16182 4660 16408
rect 4712 16390 4764 16396
rect 5080 16448 5132 16454
rect 5080 16390 5132 16396
rect 4698 16348 5006 16357
rect 4698 16346 4704 16348
rect 4760 16346 4784 16348
rect 4840 16346 4864 16348
rect 4920 16346 4944 16348
rect 5000 16346 5006 16348
rect 4760 16294 4762 16346
rect 4942 16294 4944 16346
rect 4698 16292 4704 16294
rect 4760 16292 4784 16294
rect 4840 16292 4864 16294
rect 4920 16292 4944 16294
rect 5000 16292 5006 16294
rect 4698 16283 5006 16292
rect 5184 16250 5212 17138
rect 5264 16992 5316 16998
rect 5264 16934 5316 16940
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5172 16244 5224 16250
rect 5172 16186 5224 16192
rect 4620 16176 4672 16182
rect 4620 16118 4672 16124
rect 4528 16108 4580 16114
rect 4528 16050 4580 16056
rect 4344 14816 4396 14822
rect 4344 14758 4396 14764
rect 4252 13184 4304 13190
rect 4252 13126 4304 13132
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 4252 12640 4304 12646
rect 4250 12608 4252 12617
rect 4304 12608 4306 12617
rect 4250 12543 4306 12552
rect 3896 12406 4108 12434
rect 3884 12368 3936 12374
rect 3884 12310 3936 12316
rect 3896 11694 3924 12310
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 3896 11354 3924 11630
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3712 11206 3832 11234
rect 3712 10810 3740 11206
rect 3896 10810 3924 11290
rect 3700 10804 3752 10810
rect 3700 10746 3752 10752
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 3896 10674 3924 10746
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 3988 9586 4016 12038
rect 3976 9580 4028 9586
rect 3976 9522 4028 9528
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3792 9104 3844 9110
rect 3792 9046 3844 9052
rect 3700 8900 3752 8906
rect 3700 8842 3752 8848
rect 3712 8498 3740 8842
rect 3804 8838 3832 9046
rect 3988 8974 4016 9318
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 3516 6384 3568 6390
rect 3516 6326 3568 6332
rect 3424 5840 3476 5846
rect 3424 5782 3476 5788
rect 3516 5568 3568 5574
rect 3516 5510 3568 5516
rect 3528 5370 3556 5510
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 3620 5166 3648 6598
rect 3700 6112 3752 6118
rect 3700 6054 3752 6060
rect 3712 5273 3740 6054
rect 3698 5264 3754 5273
rect 3804 5234 3832 8774
rect 3988 8498 4016 8910
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 3884 8016 3936 8022
rect 3884 7958 3936 7964
rect 3896 7313 3924 7958
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3882 7304 3938 7313
rect 3882 7239 3938 7248
rect 3882 6352 3938 6361
rect 3882 6287 3884 6296
rect 3936 6287 3938 6296
rect 3884 6258 3936 6264
rect 3698 5199 3754 5208
rect 3792 5228 3844 5234
rect 3424 5160 3476 5166
rect 3424 5102 3476 5108
rect 3608 5160 3660 5166
rect 3608 5102 3660 5108
rect 3332 4752 3384 4758
rect 3332 4694 3384 4700
rect 3240 4548 3292 4554
rect 3240 4490 3292 4496
rect 3330 4448 3386 4457
rect 3330 4383 3386 4392
rect 3238 4312 3294 4321
rect 3238 4247 3294 4256
rect 3252 4146 3280 4247
rect 3344 4146 3372 4383
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3436 4049 3464 5102
rect 3712 5030 3740 5199
rect 3792 5170 3844 5176
rect 3700 5024 3752 5030
rect 3700 4966 3752 4972
rect 3698 4856 3754 4865
rect 3698 4791 3754 4800
rect 3608 4752 3660 4758
rect 3608 4694 3660 4700
rect 3516 4548 3568 4554
rect 3516 4490 3568 4496
rect 3422 4040 3478 4049
rect 3332 4004 3384 4010
rect 3422 3975 3478 3984
rect 3332 3946 3384 3952
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 3148 3528 3200 3534
rect 3148 3470 3200 3476
rect 3252 2990 3280 3878
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 3068 2808 3188 2836
rect 2688 2790 2740 2796
rect 2596 2576 2648 2582
rect 2596 2518 2648 2524
rect 2700 2530 2728 2790
rect 2824 2748 3132 2757
rect 2824 2746 2830 2748
rect 2886 2746 2910 2748
rect 2966 2746 2990 2748
rect 3046 2746 3070 2748
rect 3126 2746 3132 2748
rect 2886 2694 2888 2746
rect 3068 2694 3070 2746
rect 2824 2692 2830 2694
rect 2886 2692 2910 2694
rect 2966 2692 2990 2694
rect 3046 2692 3070 2694
rect 3126 2692 3132 2694
rect 2824 2683 3132 2692
rect 2504 2440 2556 2446
rect 2504 2382 2556 2388
rect 2410 2000 2466 2009
rect 2410 1935 2466 1944
rect 2608 800 2636 2518
rect 2700 2502 2912 2530
rect 2884 800 2912 2502
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 2976 1834 3004 2382
rect 2964 1828 3016 1834
rect 2964 1770 3016 1776
rect 3160 800 3188 2808
rect 3344 2514 3372 3946
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3332 2508 3384 2514
rect 3332 2450 3384 2456
rect 3436 800 3464 2586
rect 3528 1698 3556 4490
rect 3620 1873 3648 4694
rect 3712 4282 3740 4791
rect 3790 4584 3846 4593
rect 3790 4519 3846 4528
rect 3804 4486 3832 4519
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 3700 4276 3752 4282
rect 3700 4218 3752 4224
rect 3712 3602 3740 4218
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 3896 4026 3924 6258
rect 3988 5370 4016 7346
rect 4080 6497 4108 12406
rect 4163 12430 4200 12458
rect 4163 12356 4191 12430
rect 4344 12368 4396 12374
rect 4163 12328 4292 12356
rect 4158 11792 4214 11801
rect 4158 11727 4214 11736
rect 4172 11558 4200 11727
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4172 10674 4200 11494
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4160 10464 4212 10470
rect 4160 10406 4212 10412
rect 4066 6488 4122 6497
rect 4066 6423 4122 6432
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 3976 5228 4028 5234
rect 4080 5216 4108 6258
rect 4172 5574 4200 10406
rect 4264 6458 4292 12328
rect 4344 12310 4396 12316
rect 4356 9450 4384 12310
rect 4448 12102 4476 12718
rect 4540 12442 4568 16050
rect 4632 15502 4660 16118
rect 5276 15706 5304 16934
rect 5552 16572 5580 16934
rect 5632 16584 5684 16590
rect 5552 16544 5632 16572
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4632 14958 4660 15438
rect 5172 15428 5224 15434
rect 5172 15370 5224 15376
rect 4698 15260 5006 15269
rect 4698 15258 4704 15260
rect 4760 15258 4784 15260
rect 4840 15258 4864 15260
rect 4920 15258 4944 15260
rect 5000 15258 5006 15260
rect 4760 15206 4762 15258
rect 4942 15206 4944 15258
rect 4698 15204 4704 15206
rect 4760 15204 4784 15206
rect 4840 15204 4864 15206
rect 4920 15204 4944 15206
rect 5000 15204 5006 15206
rect 4698 15195 5006 15204
rect 4804 15088 4856 15094
rect 4804 15030 4856 15036
rect 4620 14952 4672 14958
rect 4620 14894 4672 14900
rect 4632 14482 4660 14894
rect 4816 14822 4844 15030
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 5184 14278 5212 15370
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5172 14272 5224 14278
rect 5172 14214 5224 14220
rect 4698 14172 5006 14181
rect 4698 14170 4704 14172
rect 4760 14170 4784 14172
rect 4840 14170 4864 14172
rect 4920 14170 4944 14172
rect 5000 14170 5006 14172
rect 4760 14118 4762 14170
rect 4942 14118 4944 14170
rect 4698 14116 4704 14118
rect 4760 14116 4784 14118
rect 4840 14116 4864 14118
rect 4920 14116 4944 14118
rect 5000 14116 5006 14118
rect 4698 14107 5006 14116
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 4528 12436 4580 12442
rect 4528 12378 4580 12384
rect 4436 12096 4488 12102
rect 4436 12038 4488 12044
rect 4448 9489 4476 12038
rect 4434 9480 4490 9489
rect 4344 9444 4396 9450
rect 4434 9415 4490 9424
rect 4344 9386 4396 9392
rect 4540 9058 4568 12378
rect 4632 11744 4660 14010
rect 4712 13796 4764 13802
rect 4712 13738 4764 13744
rect 4724 13394 4752 13738
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 4698 13084 5006 13093
rect 4698 13082 4704 13084
rect 4760 13082 4784 13084
rect 4840 13082 4864 13084
rect 4920 13082 4944 13084
rect 5000 13082 5006 13084
rect 4760 13030 4762 13082
rect 4942 13030 4944 13082
rect 4698 13028 4704 13030
rect 4760 13028 4784 13030
rect 4840 13028 4864 13030
rect 4920 13028 4944 13030
rect 5000 13028 5006 13030
rect 4698 13019 5006 13028
rect 5092 12918 5120 13126
rect 5080 12912 5132 12918
rect 5080 12854 5132 12860
rect 5184 12434 5212 14214
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 5276 12753 5304 12786
rect 5262 12744 5318 12753
rect 5262 12679 5318 12688
rect 5368 12434 5396 14758
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 5460 14074 5488 14418
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 5448 13252 5500 13258
rect 5448 13194 5500 13200
rect 5092 12406 5212 12434
rect 5276 12406 5396 12434
rect 4698 11996 5006 12005
rect 4698 11994 4704 11996
rect 4760 11994 4784 11996
rect 4840 11994 4864 11996
rect 4920 11994 4944 11996
rect 5000 11994 5006 11996
rect 4760 11942 4762 11994
rect 4942 11942 4944 11994
rect 4698 11940 4704 11942
rect 4760 11940 4784 11942
rect 4840 11940 4864 11942
rect 4920 11940 4944 11942
rect 5000 11940 5006 11942
rect 4698 11931 5006 11940
rect 4632 11716 4752 11744
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4448 9030 4568 9058
rect 4344 8900 4396 8906
rect 4344 8842 4396 8848
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4356 6186 4384 8842
rect 4344 6180 4396 6186
rect 4344 6122 4396 6128
rect 4342 5808 4398 5817
rect 4342 5743 4344 5752
rect 4396 5743 4398 5752
rect 4344 5714 4396 5720
rect 4448 5658 4476 9030
rect 4632 8498 4660 11494
rect 4724 11150 4752 11716
rect 4712 11144 4764 11150
rect 4710 11112 4712 11121
rect 4764 11112 4766 11121
rect 4710 11047 4766 11056
rect 4698 10908 5006 10917
rect 4698 10906 4704 10908
rect 4760 10906 4784 10908
rect 4840 10906 4864 10908
rect 4920 10906 4944 10908
rect 5000 10906 5006 10908
rect 4760 10854 4762 10906
rect 4942 10854 4944 10906
rect 4698 10852 4704 10854
rect 4760 10852 4784 10854
rect 4840 10852 4864 10854
rect 4920 10852 4944 10854
rect 5000 10852 5006 10854
rect 4698 10843 5006 10852
rect 4698 9820 5006 9829
rect 4698 9818 4704 9820
rect 4760 9818 4784 9820
rect 4840 9818 4864 9820
rect 4920 9818 4944 9820
rect 5000 9818 5006 9820
rect 4760 9766 4762 9818
rect 4942 9766 4944 9818
rect 4698 9764 4704 9766
rect 4760 9764 4784 9766
rect 4840 9764 4864 9766
rect 4920 9764 4944 9766
rect 5000 9764 5006 9766
rect 4698 9755 5006 9764
rect 4698 8732 5006 8741
rect 4698 8730 4704 8732
rect 4760 8730 4784 8732
rect 4840 8730 4864 8732
rect 4920 8730 4944 8732
rect 5000 8730 5006 8732
rect 4760 8678 4762 8730
rect 4942 8678 4944 8730
rect 4698 8676 4704 8678
rect 4760 8676 4784 8678
rect 4840 8676 4864 8678
rect 4920 8676 4944 8678
rect 5000 8676 5006 8678
rect 4698 8667 5006 8676
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4632 7410 4660 7822
rect 4698 7644 5006 7653
rect 4698 7642 4704 7644
rect 4760 7642 4784 7644
rect 4840 7642 4864 7644
rect 4920 7642 4944 7644
rect 5000 7642 5006 7644
rect 4760 7590 4762 7642
rect 4942 7590 4944 7642
rect 4698 7588 4704 7590
rect 4760 7588 4784 7590
rect 4840 7588 4864 7590
rect 4920 7588 4944 7590
rect 5000 7588 5006 7590
rect 4698 7579 5006 7588
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4632 7002 4660 7346
rect 4620 6996 4672 7002
rect 4620 6938 4672 6944
rect 4698 6556 5006 6565
rect 4698 6554 4704 6556
rect 4760 6554 4784 6556
rect 4840 6554 4864 6556
rect 4920 6554 4944 6556
rect 5000 6554 5006 6556
rect 4760 6502 4762 6554
rect 4942 6502 4944 6554
rect 4698 6500 4704 6502
rect 4760 6500 4784 6502
rect 4840 6500 4864 6502
rect 4920 6500 4944 6502
rect 5000 6500 5006 6502
rect 4698 6491 5006 6500
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4528 6248 4580 6254
rect 4528 6190 4580 6196
rect 4356 5630 4476 5658
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 4172 5302 4200 5510
rect 4160 5296 4212 5302
rect 4160 5238 4212 5244
rect 4028 5188 4108 5216
rect 3976 5170 4028 5176
rect 3988 4214 4016 5170
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4080 4865 4108 4966
rect 4066 4856 4122 4865
rect 4066 4791 4122 4800
rect 4172 4570 4200 5238
rect 4080 4542 4200 4570
rect 4080 4321 4108 4542
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 4066 4312 4122 4321
rect 4066 4247 4122 4256
rect 3976 4208 4028 4214
rect 3976 4150 4028 4156
rect 4080 4146 4108 4247
rect 4172 4214 4200 4422
rect 4160 4208 4212 4214
rect 4158 4176 4160 4185
rect 4212 4176 4214 4185
rect 4068 4140 4120 4146
rect 4158 4111 4214 4120
rect 4068 4082 4120 4088
rect 3700 3596 3752 3602
rect 3700 3538 3752 3544
rect 3700 2916 3752 2922
rect 3700 2858 3752 2864
rect 3606 1864 3662 1873
rect 3606 1799 3662 1808
rect 3516 1692 3568 1698
rect 3516 1634 3568 1640
rect 3712 800 3740 2858
rect 3804 2650 3832 4014
rect 3896 3998 4200 4026
rect 4264 4010 4292 5510
rect 4356 4570 4384 5630
rect 4434 4856 4490 4865
rect 4540 4826 4568 6190
rect 4632 6118 4660 6394
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4434 4791 4490 4800
rect 4528 4820 4580 4826
rect 4448 4690 4476 4791
rect 4528 4762 4580 4768
rect 4632 4706 4660 6054
rect 4724 5710 4752 6394
rect 4988 6384 5040 6390
rect 4988 6326 5040 6332
rect 4712 5704 4764 5710
rect 5000 5681 5028 6326
rect 5092 5846 5120 12406
rect 5276 11914 5304 12406
rect 5460 12170 5488 13194
rect 5552 12866 5580 16544
rect 5632 16526 5684 16532
rect 5828 16250 5856 19200
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 6012 16794 6040 17138
rect 6196 17066 6224 19200
rect 6276 17264 6328 17270
rect 6276 17206 6328 17212
rect 6184 17060 6236 17066
rect 6184 17002 6236 17008
rect 6288 16794 6316 17206
rect 6564 16980 6592 19200
rect 6932 17338 6960 19200
rect 7300 17338 7328 19200
rect 7668 17338 7696 19200
rect 8036 17338 8064 19200
rect 8404 17524 8432 19200
rect 8312 17496 8432 17524
rect 8772 17524 8800 19200
rect 8772 17496 8892 17524
rect 8312 17338 8340 17496
rect 8446 17436 8754 17445
rect 8446 17434 8452 17436
rect 8508 17434 8532 17436
rect 8588 17434 8612 17436
rect 8668 17434 8692 17436
rect 8748 17434 8754 17436
rect 8508 17382 8510 17434
rect 8690 17382 8692 17434
rect 8446 17380 8452 17382
rect 8508 17380 8532 17382
rect 8588 17380 8612 17382
rect 8668 17380 8692 17382
rect 8748 17380 8754 17382
rect 8446 17371 8754 17380
rect 8864 17338 8892 17496
rect 9140 17338 9168 19200
rect 9220 17740 9272 17746
rect 9220 17682 9272 17688
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 7288 17332 7340 17338
rect 7288 17274 7340 17280
rect 7656 17332 7708 17338
rect 7656 17274 7708 17280
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 9128 17332 9180 17338
rect 9128 17274 9180 17280
rect 9232 17202 9260 17682
rect 9508 17338 9536 19200
rect 9876 19122 9904 19200
rect 9968 19122 9996 19230
rect 9876 19094 9996 19122
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9496 17332 9548 17338
rect 9496 17274 9548 17280
rect 9312 17264 9364 17270
rect 9312 17206 9364 17212
rect 7288 17196 7340 17202
rect 7288 17138 7340 17144
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 8392 17196 8444 17202
rect 8392 17138 8444 17144
rect 9220 17196 9272 17202
rect 9220 17138 9272 17144
rect 6472 16952 6592 16980
rect 6000 16788 6052 16794
rect 6000 16730 6052 16736
rect 6276 16788 6328 16794
rect 6276 16730 6328 16736
rect 6472 16250 6500 16952
rect 6572 16892 6880 16901
rect 6572 16890 6578 16892
rect 6634 16890 6658 16892
rect 6714 16890 6738 16892
rect 6794 16890 6818 16892
rect 6874 16890 6880 16892
rect 6634 16838 6636 16890
rect 6816 16838 6818 16890
rect 6572 16836 6578 16838
rect 6634 16836 6658 16838
rect 6714 16836 6738 16838
rect 6794 16836 6818 16838
rect 6874 16836 6880 16838
rect 6572 16827 6880 16836
rect 7300 16794 7328 17138
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 7472 16652 7524 16658
rect 7472 16594 7524 16600
rect 7286 16552 7342 16561
rect 7286 16487 7342 16496
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 5816 16244 5868 16250
rect 5816 16186 5868 16192
rect 6460 16244 6512 16250
rect 6460 16186 6512 16192
rect 5632 16108 5684 16114
rect 5632 16050 5684 16056
rect 5644 16017 5672 16050
rect 5630 16008 5686 16017
rect 5630 15943 5686 15952
rect 5644 14822 5672 15943
rect 6366 15872 6422 15881
rect 6366 15807 6422 15816
rect 5908 15360 5960 15366
rect 5908 15302 5960 15308
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5644 12986 5672 14758
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5724 14068 5776 14074
rect 5724 14010 5776 14016
rect 5736 13394 5764 14010
rect 5724 13388 5776 13394
rect 5724 13330 5776 13336
rect 5632 12980 5684 12986
rect 5632 12922 5684 12928
rect 5552 12838 5672 12866
rect 5736 12850 5764 13330
rect 5644 12628 5672 12838
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5552 12600 5672 12628
rect 5448 12164 5500 12170
rect 5448 12106 5500 12112
rect 5552 12102 5580 12600
rect 5630 12472 5686 12481
rect 5630 12407 5686 12416
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5184 11886 5304 11914
rect 5184 7857 5212 11886
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5276 11014 5304 11698
rect 5552 11286 5580 12038
rect 5644 11558 5672 12407
rect 5736 12238 5764 12786
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 5736 11898 5764 12174
rect 5828 12170 5856 14214
rect 5920 13938 5948 15302
rect 6092 15020 6144 15026
rect 6092 14962 6144 14968
rect 6000 14884 6052 14890
rect 6000 14826 6052 14832
rect 5908 13932 5960 13938
rect 5908 13874 5960 13880
rect 5920 13190 5948 13874
rect 6012 13240 6040 14826
rect 6104 14346 6132 14962
rect 6380 14346 6408 15807
rect 6572 15804 6880 15813
rect 6572 15802 6578 15804
rect 6634 15802 6658 15804
rect 6714 15802 6738 15804
rect 6794 15802 6818 15804
rect 6874 15802 6880 15804
rect 6634 15750 6636 15802
rect 6816 15750 6818 15802
rect 6572 15748 6578 15750
rect 6634 15748 6658 15750
rect 6714 15748 6738 15750
rect 6794 15748 6818 15750
rect 6874 15748 6880 15750
rect 6572 15739 6880 15748
rect 6920 15428 6972 15434
rect 6920 15370 6972 15376
rect 6828 15360 6880 15366
rect 6826 15328 6828 15337
rect 6880 15328 6882 15337
rect 6826 15263 6882 15272
rect 6932 15026 6960 15370
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6472 14414 6500 14758
rect 6572 14716 6880 14725
rect 6572 14714 6578 14716
rect 6634 14714 6658 14716
rect 6714 14714 6738 14716
rect 6794 14714 6818 14716
rect 6874 14714 6880 14716
rect 6634 14662 6636 14714
rect 6816 14662 6818 14714
rect 6572 14660 6578 14662
rect 6634 14660 6658 14662
rect 6714 14660 6738 14662
rect 6794 14660 6818 14662
rect 6874 14660 6880 14662
rect 6572 14651 6880 14660
rect 6460 14408 6512 14414
rect 6460 14350 6512 14356
rect 6092 14340 6144 14346
rect 6092 14282 6144 14288
rect 6368 14340 6420 14346
rect 6368 14282 6420 14288
rect 6472 14074 6500 14350
rect 6644 14340 6696 14346
rect 6644 14282 6696 14288
rect 6460 14068 6512 14074
rect 6460 14010 6512 14016
rect 6092 14000 6144 14006
rect 6092 13942 6144 13948
rect 6104 13258 6132 13942
rect 6460 13864 6512 13870
rect 6656 13841 6684 14282
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 6932 13938 6960 14010
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 6460 13806 6512 13812
rect 6642 13832 6698 13841
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 6196 13530 6224 13670
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6092 13252 6144 13258
rect 6012 13212 6049 13240
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 6021 13002 6049 13212
rect 6092 13194 6144 13200
rect 6368 13252 6420 13258
rect 6368 13194 6420 13200
rect 6184 13184 6236 13190
rect 6184 13126 6236 13132
rect 6012 12974 6049 13002
rect 6092 12980 6144 12986
rect 5816 12164 5868 12170
rect 5816 12106 5868 12112
rect 5724 11892 5776 11898
rect 5724 11834 5776 11840
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5540 11280 5592 11286
rect 5540 11222 5592 11228
rect 5264 11008 5316 11014
rect 5264 10950 5316 10956
rect 5276 8634 5304 10950
rect 5644 10742 5672 11494
rect 5632 10736 5684 10742
rect 5632 10678 5684 10684
rect 5724 10600 5776 10606
rect 5724 10542 5776 10548
rect 5736 9994 5764 10542
rect 5448 9988 5500 9994
rect 5448 9930 5500 9936
rect 5724 9988 5776 9994
rect 5724 9930 5776 9936
rect 5460 9654 5488 9930
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 5448 9648 5500 9654
rect 5448 9590 5500 9596
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5368 9110 5396 9522
rect 5356 9104 5408 9110
rect 5356 9046 5408 9052
rect 5460 9042 5488 9590
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5552 8362 5580 9318
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5170 7848 5226 7857
rect 5368 7818 5396 8230
rect 5170 7783 5226 7792
rect 5356 7812 5408 7818
rect 5356 7754 5408 7760
rect 5170 6488 5226 6497
rect 5170 6423 5172 6432
rect 5224 6423 5226 6432
rect 5172 6394 5224 6400
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 5080 5840 5132 5846
rect 5080 5782 5132 5788
rect 5080 5704 5132 5710
rect 4712 5646 4764 5652
rect 4986 5672 5042 5681
rect 5080 5646 5132 5652
rect 4986 5607 5042 5616
rect 4698 5468 5006 5477
rect 4698 5466 4704 5468
rect 4760 5466 4784 5468
rect 4840 5466 4864 5468
rect 4920 5466 4944 5468
rect 5000 5466 5006 5468
rect 4760 5414 4762 5466
rect 4942 5414 4944 5466
rect 4698 5412 4704 5414
rect 4760 5412 4784 5414
rect 4840 5412 4864 5414
rect 4920 5412 4944 5414
rect 5000 5412 5006 5414
rect 4698 5403 5006 5412
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 4896 5024 4948 5030
rect 4894 4992 4896 5001
rect 4948 4992 4950 5001
rect 4894 4927 4950 4936
rect 4436 4684 4488 4690
rect 4436 4626 4488 4632
rect 4540 4678 4660 4706
rect 5000 4690 5028 5306
rect 4988 4684 5040 4690
rect 4356 4542 4476 4570
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3896 3194 3924 3878
rect 3974 3768 4030 3777
rect 3974 3703 3976 3712
rect 4028 3703 4030 3712
rect 4068 3732 4120 3738
rect 3976 3674 4028 3680
rect 4068 3674 4120 3680
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 3988 3058 4016 3130
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 4080 2582 4108 3674
rect 4172 3398 4200 3998
rect 4252 4004 4304 4010
rect 4252 3946 4304 3952
rect 4356 3890 4384 4218
rect 4448 4026 4476 4542
rect 4540 4282 4568 4678
rect 4988 4626 5040 4632
rect 5000 4593 5028 4626
rect 4986 4584 5042 4593
rect 4986 4519 5042 4528
rect 4698 4380 5006 4389
rect 4698 4378 4704 4380
rect 4760 4378 4784 4380
rect 4840 4378 4864 4380
rect 4920 4378 4944 4380
rect 5000 4378 5006 4380
rect 4760 4326 4762 4378
rect 4942 4326 4944 4378
rect 4698 4324 4704 4326
rect 4760 4324 4784 4326
rect 4840 4324 4864 4326
rect 4920 4324 4944 4326
rect 5000 4324 5006 4326
rect 4698 4315 5006 4324
rect 4528 4276 4580 4282
rect 4528 4218 4580 4224
rect 4618 4176 4674 4185
rect 4618 4111 4674 4120
rect 4632 4026 4660 4111
rect 4448 3998 4660 4026
rect 4264 3862 4384 3890
rect 4436 3936 4488 3942
rect 4436 3878 4488 3884
rect 4528 3936 4580 3942
rect 4528 3878 4580 3884
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 4172 2990 4200 3334
rect 4264 3126 4292 3862
rect 4448 3534 4476 3878
rect 4540 3602 4568 3878
rect 4528 3596 4580 3602
rect 4528 3538 4580 3544
rect 4436 3528 4488 3534
rect 4632 3482 4660 3998
rect 5092 3670 5120 5646
rect 5080 3664 5132 3670
rect 5080 3606 5132 3612
rect 4436 3470 4488 3476
rect 4540 3454 4660 3482
rect 4252 3120 4304 3126
rect 4252 3062 4304 3068
rect 4160 2984 4212 2990
rect 4264 2972 4292 3062
rect 4540 2990 4568 3454
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 5080 3392 5132 3398
rect 5080 3334 5132 3340
rect 4632 3194 4660 3334
rect 4698 3292 5006 3301
rect 4698 3290 4704 3292
rect 4760 3290 4784 3292
rect 4840 3290 4864 3292
rect 4920 3290 4944 3292
rect 5000 3290 5006 3292
rect 4760 3238 4762 3290
rect 4942 3238 4944 3290
rect 4698 3236 4704 3238
rect 4760 3236 4784 3238
rect 4840 3236 4864 3238
rect 4920 3236 4944 3238
rect 5000 3236 5006 3238
rect 4698 3227 5006 3236
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4528 2984 4580 2990
rect 4264 2944 4384 2972
rect 4160 2926 4212 2932
rect 4252 2848 4304 2854
rect 4356 2825 4384 2944
rect 4580 2944 4752 2972
rect 4528 2926 4580 2932
rect 4252 2790 4304 2796
rect 4342 2816 4398 2825
rect 3976 2576 4028 2582
rect 3976 2518 4028 2524
rect 4068 2576 4120 2582
rect 4068 2518 4120 2524
rect 4160 2576 4212 2582
rect 4160 2518 4212 2524
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 3792 2304 3844 2310
rect 3792 2246 3844 2252
rect 3804 2106 3832 2246
rect 3792 2100 3844 2106
rect 3792 2042 3844 2048
rect 3896 1737 3924 2382
rect 3882 1728 3938 1737
rect 3882 1663 3938 1672
rect 3988 800 4016 2518
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 4080 2038 4108 2382
rect 4068 2032 4120 2038
rect 4068 1974 4120 1980
rect 4172 1970 4200 2518
rect 4160 1964 4212 1970
rect 4160 1906 4212 1912
rect 4264 800 4292 2790
rect 4342 2751 4398 2760
rect 4724 2582 4752 2944
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 4894 2544 4950 2553
rect 4894 2479 4950 2488
rect 4908 2446 4936 2479
rect 4436 2440 4488 2446
rect 4436 2382 4488 2388
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 4344 2372 4396 2378
rect 4344 2314 4396 2320
rect 4356 1170 4384 2314
rect 4448 1902 4476 2382
rect 4698 2204 5006 2213
rect 4698 2202 4704 2204
rect 4760 2202 4784 2204
rect 4840 2202 4864 2204
rect 4920 2202 4944 2204
rect 5000 2202 5006 2204
rect 4760 2150 4762 2202
rect 4942 2150 4944 2202
rect 4698 2148 4704 2150
rect 4760 2148 4784 2150
rect 4840 2148 4864 2150
rect 4920 2148 4944 2150
rect 5000 2148 5006 2150
rect 4698 2139 5006 2148
rect 4436 1896 4488 1902
rect 4436 1838 4488 1844
rect 5092 1442 5120 3334
rect 5184 2446 5212 6054
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5276 5778 5304 5850
rect 5264 5772 5316 5778
rect 5264 5714 5316 5720
rect 5264 5568 5316 5574
rect 5262 5536 5264 5545
rect 5316 5536 5318 5545
rect 5262 5471 5318 5480
rect 5368 5370 5396 7754
rect 5552 7478 5580 8298
rect 5540 7472 5592 7478
rect 5540 7414 5592 7420
rect 5448 6724 5500 6730
rect 5448 6666 5500 6672
rect 5460 6390 5488 6666
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5644 6458 5672 6598
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5448 6384 5500 6390
rect 5448 6326 5500 6332
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5460 5778 5488 6190
rect 5552 5846 5580 6258
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 5448 5772 5500 5778
rect 5448 5714 5500 5720
rect 5538 5672 5594 5681
rect 5538 5607 5594 5616
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5460 5370 5488 5510
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 5264 5296 5316 5302
rect 5446 5264 5502 5273
rect 5316 5244 5396 5250
rect 5264 5238 5396 5244
rect 5276 5222 5396 5238
rect 5368 4978 5396 5222
rect 5552 5234 5580 5607
rect 5446 5199 5502 5208
rect 5540 5228 5592 5234
rect 5460 5098 5488 5199
rect 5540 5170 5592 5176
rect 5448 5092 5500 5098
rect 5448 5034 5500 5040
rect 5276 4950 5396 4978
rect 5276 4146 5304 4950
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5460 4486 5488 4762
rect 5540 4548 5592 4554
rect 5540 4490 5592 4496
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 5446 4312 5502 4321
rect 5552 4282 5580 4490
rect 5446 4247 5502 4256
rect 5540 4276 5592 4282
rect 5264 4140 5316 4146
rect 5460 4128 5488 4247
rect 5540 4218 5592 4224
rect 5264 4082 5316 4088
rect 5368 4100 5488 4128
rect 5368 4010 5396 4100
rect 5356 4004 5408 4010
rect 5356 3946 5408 3952
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 5276 3126 5304 3878
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 5264 3120 5316 3126
rect 5264 3062 5316 3068
rect 5264 2916 5316 2922
rect 5264 2858 5316 2864
rect 5276 2514 5304 2858
rect 5264 2508 5316 2514
rect 5264 2450 5316 2456
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5264 2372 5316 2378
rect 5264 2314 5316 2320
rect 5172 2100 5224 2106
rect 5172 2042 5224 2048
rect 4816 1414 5120 1442
rect 4356 1142 4568 1170
rect 4540 800 4568 1142
rect 4816 800 4844 1414
rect 5184 1170 5212 2042
rect 5092 1142 5212 1170
rect 5276 1170 5304 2314
rect 5368 1601 5396 3470
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 5540 3460 5592 3466
rect 5540 3402 5592 3408
rect 5460 3369 5488 3402
rect 5446 3360 5502 3369
rect 5446 3295 5502 3304
rect 5446 3224 5502 3233
rect 5446 3159 5502 3168
rect 5460 2990 5488 3159
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5552 2922 5580 3402
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 5644 2582 5672 6394
rect 5736 4622 5764 9658
rect 5828 6254 5856 12106
rect 6012 10606 6040 12974
rect 6092 12922 6144 12928
rect 6000 10600 6052 10606
rect 6000 10542 6052 10548
rect 6104 9058 6132 12922
rect 6012 9030 6132 9058
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 5920 5953 5948 6394
rect 5906 5944 5962 5953
rect 5816 5908 5868 5914
rect 5906 5879 5962 5888
rect 5816 5850 5868 5856
rect 5828 5234 5856 5850
rect 6012 5778 6040 9030
rect 6092 8900 6144 8906
rect 6092 8842 6144 8848
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 5906 5400 5962 5409
rect 5906 5335 5962 5344
rect 5920 5302 5948 5335
rect 5908 5296 5960 5302
rect 6104 5273 6132 8842
rect 6196 5302 6224 13126
rect 6380 12617 6408 13194
rect 6366 12608 6422 12617
rect 6366 12543 6422 12552
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6380 10810 6408 11698
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6472 8906 6500 13806
rect 6642 13767 6698 13776
rect 6572 13628 6880 13637
rect 6572 13626 6578 13628
rect 6634 13626 6658 13628
rect 6714 13626 6738 13628
rect 6794 13626 6818 13628
rect 6874 13626 6880 13628
rect 6634 13574 6636 13626
rect 6816 13574 6818 13626
rect 6572 13572 6578 13574
rect 6634 13572 6658 13574
rect 6714 13572 6738 13574
rect 6794 13572 6818 13574
rect 6874 13572 6880 13574
rect 6572 13563 6880 13572
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 6932 12714 6960 12922
rect 6920 12708 6972 12714
rect 6920 12650 6972 12656
rect 6572 12540 6880 12549
rect 6572 12538 6578 12540
rect 6634 12538 6658 12540
rect 6714 12538 6738 12540
rect 6794 12538 6818 12540
rect 6874 12538 6880 12540
rect 6634 12486 6636 12538
rect 6816 12486 6818 12538
rect 6572 12484 6578 12486
rect 6634 12484 6658 12486
rect 6714 12484 6738 12486
rect 6794 12484 6818 12486
rect 6874 12484 6880 12486
rect 6572 12475 6880 12484
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 6572 11452 6880 11461
rect 6572 11450 6578 11452
rect 6634 11450 6658 11452
rect 6714 11450 6738 11452
rect 6794 11450 6818 11452
rect 6874 11450 6880 11452
rect 6634 11398 6636 11450
rect 6816 11398 6818 11450
rect 6572 11396 6578 11398
rect 6634 11396 6658 11398
rect 6714 11396 6738 11398
rect 6794 11396 6818 11398
rect 6874 11396 6880 11398
rect 6572 11387 6880 11396
rect 6572 10364 6880 10373
rect 6572 10362 6578 10364
rect 6634 10362 6658 10364
rect 6714 10362 6738 10364
rect 6794 10362 6818 10364
rect 6874 10362 6880 10364
rect 6634 10310 6636 10362
rect 6816 10310 6818 10362
rect 6572 10308 6578 10310
rect 6634 10308 6658 10310
rect 6714 10308 6738 10310
rect 6794 10308 6818 10310
rect 6874 10308 6880 10310
rect 6572 10299 6880 10308
rect 6572 9276 6880 9285
rect 6572 9274 6578 9276
rect 6634 9274 6658 9276
rect 6714 9274 6738 9276
rect 6794 9274 6818 9276
rect 6874 9274 6880 9276
rect 6634 9222 6636 9274
rect 6816 9222 6818 9274
rect 6572 9220 6578 9222
rect 6634 9220 6658 9222
rect 6714 9220 6738 9222
rect 6794 9220 6818 9222
rect 6874 9220 6880 9222
rect 6572 9211 6880 9220
rect 6460 8900 6512 8906
rect 6460 8842 6512 8848
rect 6736 8560 6788 8566
rect 6734 8528 6736 8537
rect 6788 8528 6790 8537
rect 6734 8463 6790 8472
rect 6572 8188 6880 8197
rect 6572 8186 6578 8188
rect 6634 8186 6658 8188
rect 6714 8186 6738 8188
rect 6794 8186 6818 8188
rect 6874 8186 6880 8188
rect 6634 8134 6636 8186
rect 6816 8134 6818 8186
rect 6572 8132 6578 8134
rect 6634 8132 6658 8134
rect 6714 8132 6738 8134
rect 6794 8132 6818 8134
rect 6874 8132 6880 8134
rect 6572 8123 6880 8132
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6288 5914 6316 7686
rect 6460 7336 6512 7342
rect 6460 7278 6512 7284
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6380 6905 6408 7142
rect 6366 6896 6422 6905
rect 6366 6831 6422 6840
rect 6472 6458 6500 7278
rect 6572 7100 6880 7109
rect 6572 7098 6578 7100
rect 6634 7098 6658 7100
rect 6714 7098 6738 7100
rect 6794 7098 6818 7100
rect 6874 7098 6880 7100
rect 6634 7046 6636 7098
rect 6816 7046 6818 7098
rect 6572 7044 6578 7046
rect 6634 7044 6658 7046
rect 6714 7044 6738 7046
rect 6794 7044 6818 7046
rect 6874 7044 6880 7046
rect 6572 7035 6880 7044
rect 6642 6896 6698 6905
rect 6642 6831 6698 6840
rect 6656 6798 6684 6831
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6932 6662 6960 12378
rect 7024 11898 7052 16390
rect 7104 16176 7156 16182
rect 7104 16118 7156 16124
rect 7116 15994 7144 16118
rect 7116 15966 7236 15994
rect 7104 15904 7156 15910
rect 7104 15846 7156 15852
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 7024 11150 7052 11834
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 7024 7993 7052 11086
rect 7010 7984 7066 7993
rect 7010 7919 7066 7928
rect 7116 6914 7144 15846
rect 7208 14278 7236 15966
rect 7196 14272 7248 14278
rect 7196 14214 7248 14220
rect 7300 14074 7328 16487
rect 7380 15700 7432 15706
rect 7380 15642 7432 15648
rect 7392 15094 7420 15642
rect 7484 15502 7512 16594
rect 7576 16250 7604 17070
rect 7668 16250 7696 17138
rect 8300 17128 8352 17134
rect 8300 17070 8352 17076
rect 7932 16720 7984 16726
rect 7932 16662 7984 16668
rect 7840 16584 7892 16590
rect 7840 16526 7892 16532
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 7656 16244 7708 16250
rect 7656 16186 7708 16192
rect 7656 16108 7708 16114
rect 7708 16068 7788 16096
rect 7656 16050 7708 16056
rect 7564 16040 7616 16046
rect 7564 15982 7616 15988
rect 7472 15496 7524 15502
rect 7472 15438 7524 15444
rect 7380 15088 7432 15094
rect 7380 15030 7432 15036
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7196 13932 7248 13938
rect 7196 13874 7248 13880
rect 7208 12442 7236 13874
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 7300 12442 7328 13126
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7484 11762 7512 15438
rect 7576 15094 7604 15982
rect 7656 15972 7708 15978
rect 7656 15914 7708 15920
rect 7668 15638 7696 15914
rect 7656 15632 7708 15638
rect 7656 15574 7708 15580
rect 7668 15162 7696 15574
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 7564 15088 7616 15094
rect 7564 15030 7616 15036
rect 7656 14340 7708 14346
rect 7656 14282 7708 14288
rect 7668 14249 7696 14282
rect 7654 14240 7710 14249
rect 7654 14175 7710 14184
rect 7654 12880 7710 12889
rect 7654 12815 7710 12824
rect 7564 12436 7616 12442
rect 7564 12378 7616 12384
rect 7576 12345 7604 12378
rect 7562 12336 7618 12345
rect 7562 12271 7618 12280
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7024 6886 7144 6914
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6932 6474 6960 6598
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6840 6446 6960 6474
rect 6840 6254 6868 6446
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6460 6112 6512 6118
rect 6460 6054 6512 6060
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6472 5778 6500 6054
rect 6572 6012 6880 6021
rect 6572 6010 6578 6012
rect 6634 6010 6658 6012
rect 6714 6010 6738 6012
rect 6794 6010 6818 6012
rect 6874 6010 6880 6012
rect 6634 5958 6636 6010
rect 6816 5958 6818 6010
rect 6572 5956 6578 5958
rect 6634 5956 6658 5958
rect 6714 5956 6738 5958
rect 6794 5956 6818 5958
rect 6874 5956 6880 5958
rect 6572 5947 6880 5956
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6748 5778 6776 5850
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6184 5296 6236 5302
rect 5908 5238 5960 5244
rect 6090 5264 6146 5273
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5828 4690 5856 5170
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5920 4622 5948 5238
rect 6184 5238 6236 5244
rect 6090 5199 6146 5208
rect 6000 5024 6052 5030
rect 6104 5001 6132 5199
rect 6000 4966 6052 4972
rect 6090 4992 6146 5001
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 5736 4214 5764 4558
rect 5908 4480 5960 4486
rect 5908 4422 5960 4428
rect 5724 4208 5776 4214
rect 5724 4150 5776 4156
rect 5736 3720 5764 4150
rect 5736 3692 5856 3720
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 5736 2972 5764 3538
rect 5828 3505 5856 3692
rect 5814 3496 5870 3505
rect 5814 3431 5870 3440
rect 5816 3392 5868 3398
rect 5816 3334 5868 3340
rect 5828 3074 5856 3334
rect 5920 3194 5948 4422
rect 6012 4128 6040 4966
rect 6090 4927 6146 4936
rect 6104 4706 6132 4927
rect 6288 4826 6316 5646
rect 6932 5545 6960 6326
rect 7024 6322 7052 6886
rect 7208 6746 7236 7346
rect 7116 6718 7236 6746
rect 7116 6497 7144 6718
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7102 6488 7158 6497
rect 7102 6423 7158 6432
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 6918 5536 6974 5545
rect 6918 5471 6974 5480
rect 6932 5386 6960 5471
rect 6748 5358 6960 5386
rect 6748 5302 6776 5358
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 6736 5296 6788 5302
rect 6736 5238 6788 5244
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6380 4826 6408 4966
rect 6276 4820 6328 4826
rect 6276 4762 6328 4768
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6104 4690 6316 4706
rect 6472 4690 6500 5238
rect 6572 4924 6880 4933
rect 6572 4922 6578 4924
rect 6634 4922 6658 4924
rect 6714 4922 6738 4924
rect 6794 4922 6818 4924
rect 6874 4922 6880 4924
rect 6634 4870 6636 4922
rect 6816 4870 6818 4922
rect 6572 4868 6578 4870
rect 6634 4868 6658 4870
rect 6714 4868 6738 4870
rect 6794 4868 6818 4870
rect 6874 4868 6880 4870
rect 6572 4859 6880 4868
rect 6552 4820 6604 4826
rect 6552 4762 6604 4768
rect 6104 4684 6328 4690
rect 6104 4678 6276 4684
rect 6276 4626 6328 4632
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6472 4457 6500 4626
rect 6458 4448 6514 4457
rect 6458 4383 6514 4392
rect 6368 4140 6420 4146
rect 6012 4100 6368 4128
rect 6092 4004 6144 4010
rect 6012 3964 6092 3992
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 5828 3046 5948 3074
rect 5816 2984 5868 2990
rect 5736 2944 5816 2972
rect 5816 2926 5868 2932
rect 5814 2680 5870 2689
rect 5814 2615 5870 2624
rect 5632 2576 5684 2582
rect 5538 2544 5594 2553
rect 5632 2518 5684 2524
rect 5538 2479 5594 2488
rect 5448 2304 5500 2310
rect 5448 2246 5500 2252
rect 5460 1630 5488 2246
rect 5552 1766 5580 2479
rect 5828 2446 5856 2615
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 5920 2394 5948 3046
rect 6012 2650 6040 3964
rect 6092 3946 6144 3952
rect 6092 3120 6144 3126
rect 6196 3097 6224 4100
rect 6368 4082 6420 4088
rect 6564 4049 6592 4762
rect 6828 4752 6880 4758
rect 6828 4694 6880 4700
rect 6642 4176 6698 4185
rect 6642 4111 6698 4120
rect 6550 4040 6606 4049
rect 6550 3975 6606 3984
rect 6656 3942 6684 4111
rect 6276 3936 6328 3942
rect 6274 3904 6276 3913
rect 6460 3936 6512 3942
rect 6328 3904 6330 3913
rect 6460 3878 6512 3884
rect 6644 3936 6696 3942
rect 6840 3924 6868 4694
rect 6932 4622 6960 5238
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6840 3896 6960 3924
rect 6644 3878 6696 3884
rect 6274 3839 6330 3848
rect 6366 3768 6422 3777
rect 6366 3703 6368 3712
rect 6420 3703 6422 3712
rect 6368 3674 6420 3680
rect 6274 3632 6330 3641
rect 6274 3567 6330 3576
rect 6288 3534 6316 3567
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 6368 3392 6420 3398
rect 6368 3334 6420 3340
rect 6472 3346 6500 3878
rect 6572 3836 6880 3845
rect 6572 3834 6578 3836
rect 6634 3834 6658 3836
rect 6714 3834 6738 3836
rect 6794 3834 6818 3836
rect 6874 3834 6880 3836
rect 6634 3782 6636 3834
rect 6816 3782 6818 3834
rect 6572 3780 6578 3782
rect 6634 3780 6658 3782
rect 6714 3780 6738 3782
rect 6794 3780 6818 3782
rect 6874 3780 6880 3782
rect 6572 3771 6880 3780
rect 6642 3632 6698 3641
rect 6826 3632 6882 3641
rect 6698 3590 6776 3618
rect 6642 3567 6698 3576
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6092 3062 6144 3068
rect 6182 3088 6238 3097
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 5920 2366 6040 2394
rect 5908 2304 5960 2310
rect 5908 2246 5960 2252
rect 5632 1964 5684 1970
rect 5632 1906 5684 1912
rect 5540 1760 5592 1766
rect 5540 1702 5592 1708
rect 5448 1624 5500 1630
rect 5354 1592 5410 1601
rect 5448 1566 5500 1572
rect 5354 1527 5410 1536
rect 5276 1142 5396 1170
rect 5092 800 5120 1142
rect 5368 800 5396 1142
rect 5644 800 5672 1906
rect 5920 800 5948 2246
rect 6012 1970 6040 2366
rect 6000 1964 6052 1970
rect 6000 1906 6052 1912
rect 6104 1873 6132 3062
rect 6182 3023 6238 3032
rect 6184 2848 6236 2854
rect 6184 2790 6236 2796
rect 6090 1864 6146 1873
rect 6090 1799 6146 1808
rect 6196 800 6224 2790
rect 6276 2440 6328 2446
rect 6276 2382 6328 2388
rect 6288 2106 6316 2382
rect 6276 2100 6328 2106
rect 6276 2042 6328 2048
rect 6380 2009 6408 3334
rect 6472 3318 6592 3346
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6472 3058 6500 3130
rect 6564 3126 6592 3318
rect 6552 3120 6604 3126
rect 6552 3062 6604 3068
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6656 2938 6684 3470
rect 6748 3380 6776 3590
rect 6826 3567 6828 3576
rect 6880 3567 6882 3576
rect 6828 3538 6880 3544
rect 6828 3392 6880 3398
rect 6748 3352 6828 3380
rect 6828 3334 6880 3340
rect 6472 2910 6684 2938
rect 6826 2952 6882 2961
rect 6472 2582 6500 2910
rect 6826 2887 6828 2896
rect 6880 2887 6882 2896
rect 6828 2858 6880 2864
rect 6572 2748 6880 2757
rect 6572 2746 6578 2748
rect 6634 2746 6658 2748
rect 6714 2746 6738 2748
rect 6794 2746 6818 2748
rect 6874 2746 6880 2748
rect 6634 2694 6636 2746
rect 6816 2694 6818 2746
rect 6572 2692 6578 2694
rect 6634 2692 6658 2694
rect 6714 2692 6738 2694
rect 6794 2692 6818 2694
rect 6874 2692 6880 2694
rect 6572 2683 6880 2692
rect 6460 2576 6512 2582
rect 6460 2518 6512 2524
rect 6828 2440 6880 2446
rect 6932 2428 6960 3896
rect 7024 3058 7052 6258
rect 7116 6118 7144 6258
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 7102 5944 7158 5953
rect 7102 5879 7158 5888
rect 7116 5778 7144 5879
rect 7208 5778 7236 6598
rect 7104 5772 7156 5778
rect 7104 5714 7156 5720
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7116 5166 7144 5714
rect 7300 5234 7328 11494
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7392 10810 7420 11086
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 7484 10198 7512 11698
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7472 10192 7524 10198
rect 7472 10134 7524 10140
rect 7576 9722 7604 11494
rect 7668 11234 7696 12815
rect 7760 11665 7788 16068
rect 7852 15366 7880 16526
rect 7840 15360 7892 15366
rect 7840 15302 7892 15308
rect 7746 11656 7802 11665
rect 7746 11591 7802 11600
rect 7840 11620 7892 11626
rect 7840 11562 7892 11568
rect 7668 11206 7788 11234
rect 7656 11076 7708 11082
rect 7656 11018 7708 11024
rect 7668 10266 7696 11018
rect 7760 10674 7788 11206
rect 7852 11082 7880 11562
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7472 9580 7524 9586
rect 7576 9568 7604 9658
rect 7524 9540 7604 9568
rect 7472 9522 7524 9528
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7392 7818 7420 9114
rect 7472 9104 7524 9110
rect 7472 9046 7524 9052
rect 7380 7812 7432 7818
rect 7380 7754 7432 7760
rect 7392 6905 7420 7754
rect 7378 6896 7434 6905
rect 7378 6831 7434 6840
rect 7484 6769 7512 9046
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7668 7954 7696 8230
rect 7656 7948 7708 7954
rect 7656 7890 7708 7896
rect 7668 7546 7696 7890
rect 7760 7886 7788 10610
rect 7944 9994 7972 16662
rect 8312 16250 8340 17070
rect 8404 16794 8432 17138
rect 9220 16992 9272 16998
rect 9220 16934 9272 16940
rect 8392 16788 8444 16794
rect 8392 16730 8444 16736
rect 8390 16552 8446 16561
rect 8390 16487 8446 16496
rect 8404 16454 8432 16487
rect 8392 16448 8444 16454
rect 8392 16390 8444 16396
rect 8446 16348 8754 16357
rect 8446 16346 8452 16348
rect 8508 16346 8532 16348
rect 8588 16346 8612 16348
rect 8668 16346 8692 16348
rect 8748 16346 8754 16348
rect 8508 16294 8510 16346
rect 8690 16294 8692 16346
rect 8446 16292 8452 16294
rect 8508 16292 8532 16294
rect 8588 16292 8612 16294
rect 8668 16292 8692 16294
rect 8748 16292 8754 16294
rect 8446 16283 8754 16292
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8576 16244 8628 16250
rect 8576 16186 8628 16192
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 8116 16040 8168 16046
rect 8116 15982 8168 15988
rect 8128 15434 8156 15982
rect 8220 15910 8248 16050
rect 8588 16017 8616 16186
rect 9128 16176 9180 16182
rect 9128 16118 9180 16124
rect 8574 16008 8630 16017
rect 8574 15943 8630 15952
rect 8944 15972 8996 15978
rect 8944 15914 8996 15920
rect 8208 15904 8260 15910
rect 8208 15846 8260 15852
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 8116 15428 8168 15434
rect 8116 15370 8168 15376
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 7932 9988 7984 9994
rect 7932 9930 7984 9936
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 7656 7540 7708 7546
rect 7576 7500 7656 7528
rect 7576 7002 7604 7500
rect 7656 7482 7708 7488
rect 7852 7342 7880 9522
rect 7944 8634 7972 9930
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 7840 7336 7892 7342
rect 7760 7296 7840 7324
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7656 6928 7708 6934
rect 7656 6870 7708 6876
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 7470 6760 7526 6769
rect 7470 6695 7526 6704
rect 7576 6610 7604 6802
rect 7392 6582 7604 6610
rect 7392 6322 7420 6582
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7564 6180 7616 6186
rect 7564 6122 7616 6128
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 7380 5636 7432 5642
rect 7380 5578 7432 5584
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 7104 5024 7156 5030
rect 7208 5001 7236 5170
rect 7392 5114 7420 5578
rect 7300 5086 7420 5114
rect 7104 4966 7156 4972
rect 7194 4992 7250 5001
rect 7116 4690 7144 4966
rect 7194 4927 7250 4936
rect 7300 4826 7328 5086
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7300 4593 7328 4626
rect 7286 4584 7342 4593
rect 7286 4519 7342 4528
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7116 4010 7144 4422
rect 7194 4312 7250 4321
rect 7194 4247 7250 4256
rect 7208 4078 7236 4247
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 7104 4004 7156 4010
rect 7104 3946 7156 3952
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 7116 3505 7144 3674
rect 7102 3496 7158 3505
rect 7102 3431 7158 3440
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 6880 2400 6960 2428
rect 7024 2417 7052 2994
rect 7208 2904 7236 3878
rect 7300 3602 7328 4422
rect 7392 4146 7420 4966
rect 7484 4622 7512 6054
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7576 4321 7604 6122
rect 7668 5370 7696 6870
rect 7760 6633 7788 7296
rect 7840 7278 7892 7284
rect 7944 7274 7972 8366
rect 7932 7268 7984 7274
rect 7932 7210 7984 7216
rect 7838 7168 7894 7177
rect 8036 7154 8064 14010
rect 8128 13802 8156 14894
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8116 13796 8168 13802
rect 8116 13738 8168 13744
rect 7894 7126 8064 7154
rect 7838 7103 7894 7112
rect 7746 6624 7802 6633
rect 7746 6559 7802 6568
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7760 5370 7788 6394
rect 7852 6390 7880 7103
rect 7930 7032 7986 7041
rect 8128 7018 8156 13738
rect 8220 10470 8248 14350
rect 8312 14346 8340 15846
rect 8760 15632 8812 15638
rect 8680 15580 8760 15586
rect 8680 15574 8812 15580
rect 8680 15558 8800 15574
rect 8680 15434 8708 15558
rect 8956 15502 8984 15914
rect 9036 15632 9088 15638
rect 9036 15574 9088 15580
rect 8944 15496 8996 15502
rect 8944 15438 8996 15444
rect 8668 15428 8720 15434
rect 8668 15370 8720 15376
rect 8852 15360 8904 15366
rect 8852 15302 8904 15308
rect 8446 15260 8754 15269
rect 8446 15258 8452 15260
rect 8508 15258 8532 15260
rect 8588 15258 8612 15260
rect 8668 15258 8692 15260
rect 8748 15258 8754 15260
rect 8508 15206 8510 15258
rect 8690 15206 8692 15258
rect 8446 15204 8452 15206
rect 8508 15204 8532 15206
rect 8588 15204 8612 15206
rect 8668 15204 8692 15206
rect 8748 15204 8754 15206
rect 8446 15195 8754 15204
rect 8300 14340 8352 14346
rect 8300 14282 8352 14288
rect 8446 14172 8754 14181
rect 8446 14170 8452 14172
rect 8508 14170 8532 14172
rect 8588 14170 8612 14172
rect 8668 14170 8692 14172
rect 8748 14170 8754 14172
rect 8508 14118 8510 14170
rect 8690 14118 8692 14170
rect 8446 14116 8452 14118
rect 8508 14116 8532 14118
rect 8588 14116 8612 14118
rect 8668 14116 8692 14118
rect 8748 14116 8754 14118
rect 8446 14107 8754 14116
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8312 12782 8340 13874
rect 8446 13084 8754 13093
rect 8446 13082 8452 13084
rect 8508 13082 8532 13084
rect 8588 13082 8612 13084
rect 8668 13082 8692 13084
rect 8748 13082 8754 13084
rect 8508 13030 8510 13082
rect 8690 13030 8692 13082
rect 8446 13028 8452 13030
rect 8508 13028 8532 13030
rect 8588 13028 8612 13030
rect 8668 13028 8692 13030
rect 8748 13028 8754 13030
rect 8446 13019 8754 13028
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8680 12238 8708 12582
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8446 11996 8754 12005
rect 8446 11994 8452 11996
rect 8508 11994 8532 11996
rect 8588 11994 8612 11996
rect 8668 11994 8692 11996
rect 8748 11994 8754 11996
rect 8508 11942 8510 11994
rect 8690 11942 8692 11994
rect 8446 11940 8452 11942
rect 8508 11940 8532 11942
rect 8588 11940 8612 11942
rect 8668 11940 8692 11942
rect 8748 11940 8754 11942
rect 8446 11931 8754 11940
rect 8446 10908 8754 10917
rect 8446 10906 8452 10908
rect 8508 10906 8532 10908
rect 8588 10906 8612 10908
rect 8668 10906 8692 10908
rect 8748 10906 8754 10908
rect 8508 10854 8510 10906
rect 8690 10854 8692 10906
rect 8446 10852 8452 10854
rect 8508 10852 8532 10854
rect 8588 10852 8612 10854
rect 8668 10852 8692 10854
rect 8748 10852 8754 10854
rect 8446 10843 8754 10852
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 7930 6967 7986 6976
rect 8036 6990 8156 7018
rect 7944 6866 7972 6967
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 7840 6384 7892 6390
rect 7840 6326 7892 6332
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7852 5846 7880 6054
rect 7840 5840 7892 5846
rect 7840 5782 7892 5788
rect 7932 5840 7984 5846
rect 7932 5782 7984 5788
rect 7840 5636 7892 5642
rect 7840 5578 7892 5584
rect 7656 5364 7708 5370
rect 7656 5306 7708 5312
rect 7748 5364 7800 5370
rect 7748 5306 7800 5312
rect 7852 5250 7880 5578
rect 7668 5222 7880 5250
rect 7562 4312 7618 4321
rect 7562 4247 7618 4256
rect 7564 4208 7616 4214
rect 7470 4176 7526 4185
rect 7380 4140 7432 4146
rect 7564 4150 7616 4156
rect 7470 4111 7472 4120
rect 7380 4082 7432 4088
rect 7524 4111 7526 4120
rect 7472 4082 7524 4088
rect 7470 4040 7526 4049
rect 7470 3975 7526 3984
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 7392 3777 7420 3878
rect 7378 3768 7434 3777
rect 7378 3703 7434 3712
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 7286 3496 7342 3505
rect 7484 3466 7512 3975
rect 7286 3431 7288 3440
rect 7340 3431 7342 3440
rect 7472 3460 7524 3466
rect 7288 3402 7340 3408
rect 7472 3402 7524 3408
rect 7576 3194 7604 4150
rect 7668 3777 7696 5222
rect 7840 5160 7892 5166
rect 7840 5102 7892 5108
rect 7748 4480 7800 4486
rect 7748 4422 7800 4428
rect 7654 3768 7710 3777
rect 7654 3703 7710 3712
rect 7760 3466 7788 4422
rect 7852 4078 7880 5102
rect 7944 4690 7972 5782
rect 8036 4690 8064 6990
rect 8220 6882 8248 10406
rect 8864 10146 8892 15302
rect 8956 15162 8984 15438
rect 8944 15156 8996 15162
rect 8944 15098 8996 15104
rect 9048 14346 9076 15574
rect 9140 14958 9168 16118
rect 9232 15638 9260 16934
rect 9324 16454 9352 17206
rect 9496 16516 9548 16522
rect 9416 16476 9496 16504
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9220 15632 9272 15638
rect 9220 15574 9272 15580
rect 9128 14952 9180 14958
rect 9128 14894 9180 14900
rect 9128 14816 9180 14822
rect 9128 14758 9180 14764
rect 9036 14340 9088 14346
rect 9036 14282 9088 14288
rect 9048 13938 9076 14282
rect 9036 13932 9088 13938
rect 9036 13874 9088 13880
rect 9036 13320 9088 13326
rect 9036 13262 9088 13268
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 8312 10118 8892 10146
rect 8312 9217 8340 10118
rect 8852 10056 8904 10062
rect 8852 9998 8904 10004
rect 8446 9820 8754 9829
rect 8446 9818 8452 9820
rect 8508 9818 8532 9820
rect 8588 9818 8612 9820
rect 8668 9818 8692 9820
rect 8748 9818 8754 9820
rect 8508 9766 8510 9818
rect 8690 9766 8692 9818
rect 8446 9764 8452 9766
rect 8508 9764 8532 9766
rect 8588 9764 8612 9766
rect 8668 9764 8692 9766
rect 8748 9764 8754 9766
rect 8446 9755 8754 9764
rect 8864 9654 8892 9998
rect 8668 9648 8720 9654
rect 8668 9590 8720 9596
rect 8852 9648 8904 9654
rect 8852 9590 8904 9596
rect 8298 9208 8354 9217
rect 8298 9143 8354 9152
rect 8300 8900 8352 8906
rect 8300 8842 8352 8848
rect 8312 8809 8340 8842
rect 8680 8820 8708 9590
rect 8864 9518 8892 9590
rect 8852 9512 8904 9518
rect 8852 9454 8904 9460
rect 8864 9178 8892 9454
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 8298 8800 8354 8809
rect 8680 8792 8892 8820
rect 8298 8735 8354 8744
rect 8446 8732 8754 8741
rect 8446 8730 8452 8732
rect 8508 8730 8532 8732
rect 8588 8730 8612 8732
rect 8668 8730 8692 8732
rect 8748 8730 8754 8732
rect 8508 8678 8510 8730
rect 8690 8678 8692 8730
rect 8446 8676 8452 8678
rect 8508 8676 8532 8678
rect 8588 8676 8612 8678
rect 8668 8676 8692 8678
rect 8748 8676 8754 8678
rect 8446 8667 8754 8676
rect 8864 8673 8892 8792
rect 8850 8664 8906 8673
rect 8850 8599 8906 8608
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8852 7744 8904 7750
rect 8852 7686 8904 7692
rect 8312 7177 8340 7686
rect 8446 7644 8754 7653
rect 8446 7642 8452 7644
rect 8508 7642 8532 7644
rect 8588 7642 8612 7644
rect 8668 7642 8692 7644
rect 8748 7642 8754 7644
rect 8508 7590 8510 7642
rect 8690 7590 8692 7642
rect 8446 7588 8452 7590
rect 8508 7588 8532 7590
rect 8588 7588 8612 7590
rect 8668 7588 8692 7590
rect 8748 7588 8754 7590
rect 8446 7579 8754 7588
rect 8864 7585 8892 7686
rect 8850 7576 8906 7585
rect 8850 7511 8906 7520
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 8298 7168 8354 7177
rect 8298 7103 8354 7112
rect 8390 7032 8446 7041
rect 8390 6967 8392 6976
rect 8444 6967 8446 6976
rect 8392 6938 8444 6944
rect 8220 6854 8294 6882
rect 8266 6712 8294 6854
rect 8496 6798 8524 7346
rect 8956 7041 8984 13126
rect 9048 12986 9076 13262
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 9036 12368 9088 12374
rect 9036 12310 9088 12316
rect 9048 9110 9076 12310
rect 9140 9674 9168 14758
rect 9232 12918 9260 15574
rect 9324 13705 9352 16390
rect 9310 13696 9366 13705
rect 9310 13631 9366 13640
rect 9312 13524 9364 13530
rect 9312 13466 9364 13472
rect 9220 12912 9272 12918
rect 9220 12854 9272 12860
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 9232 12442 9260 12718
rect 9220 12436 9272 12442
rect 9220 12378 9272 12384
rect 9220 11824 9272 11830
rect 9220 11766 9272 11772
rect 9232 11286 9260 11766
rect 9220 11280 9272 11286
rect 9220 11222 9272 11228
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9232 10674 9260 10950
rect 9220 10668 9272 10674
rect 9220 10610 9272 10616
rect 9140 9646 9260 9674
rect 9128 9376 9180 9382
rect 9128 9318 9180 9324
rect 9036 9104 9088 9110
rect 9140 9081 9168 9318
rect 9036 9046 9088 9052
rect 9126 9072 9182 9081
rect 9126 9007 9182 9016
rect 9036 8968 9088 8974
rect 9036 8910 9088 8916
rect 9048 8634 9076 8910
rect 9232 8906 9260 9646
rect 9324 9178 9352 13466
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9220 8900 9272 8906
rect 9220 8842 9272 8848
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 9048 8090 9076 8570
rect 9128 8560 9180 8566
rect 9128 8502 9180 8508
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 9048 7954 9076 8026
rect 9036 7948 9088 7954
rect 9036 7890 9088 7896
rect 8942 7032 8998 7041
rect 8942 6967 8998 6976
rect 9140 6866 9168 8502
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 9232 7546 9260 8026
rect 9220 7540 9272 7546
rect 9220 7482 9272 7488
rect 9232 7002 9260 7482
rect 9324 7342 9352 9114
rect 9416 8294 9444 16476
rect 9496 16458 9548 16464
rect 9588 16448 9640 16454
rect 9588 16390 9640 16396
rect 9600 16250 9628 16390
rect 9588 16244 9640 16250
rect 9588 16186 9640 16192
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9600 14929 9628 16050
rect 9586 14920 9642 14929
rect 9496 14884 9548 14890
rect 9586 14855 9642 14864
rect 9496 14826 9548 14832
rect 9508 13841 9536 14826
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9494 13832 9550 13841
rect 9494 13767 9550 13776
rect 9494 13696 9550 13705
rect 9494 13631 9550 13640
rect 9508 12374 9536 13631
rect 9496 12368 9548 12374
rect 9496 12310 9548 12316
rect 9496 12164 9548 12170
rect 9496 12106 9548 12112
rect 9508 11694 9536 12106
rect 9496 11688 9548 11694
rect 9496 11630 9548 11636
rect 9508 10470 9536 11630
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9494 9888 9550 9897
rect 9494 9823 9550 9832
rect 9508 9722 9536 9823
rect 9496 9716 9548 9722
rect 9496 9658 9548 9664
rect 9600 9178 9628 14554
rect 9692 14074 9720 17818
rect 10152 17252 10180 19230
rect 10230 19200 10286 20000
rect 10598 19200 10654 20000
rect 10966 19200 11022 20000
rect 11334 19200 11390 20000
rect 11702 19200 11758 20000
rect 12070 19200 12126 20000
rect 12438 19200 12494 20000
rect 12806 19200 12862 20000
rect 13174 19200 13230 20000
rect 13542 19200 13598 20000
rect 13910 19200 13966 20000
rect 14278 19200 14334 20000
rect 14646 19200 14702 20000
rect 15014 19200 15070 20000
rect 15382 19200 15438 20000
rect 15750 19200 15806 20000
rect 16118 19200 16174 20000
rect 16486 19200 16542 20000
rect 16854 19200 16910 20000
rect 10244 17882 10272 19200
rect 10232 17876 10284 17882
rect 10232 17818 10284 17824
rect 10152 17224 10272 17252
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9956 17128 10008 17134
rect 9956 17070 10008 17076
rect 9784 16402 9812 17070
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9876 16658 9904 16730
rect 9864 16652 9916 16658
rect 9864 16594 9916 16600
rect 9784 16374 9904 16402
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9784 15366 9812 16186
rect 9772 15360 9824 15366
rect 9772 15302 9824 15308
rect 9876 15314 9904 16374
rect 9968 15434 9996 17070
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 10060 16425 10088 16526
rect 10046 16416 10102 16425
rect 10046 16351 10102 16360
rect 10048 16176 10100 16182
rect 10048 16118 10100 16124
rect 9956 15428 10008 15434
rect 9956 15370 10008 15376
rect 9876 15286 9996 15314
rect 9770 15192 9826 15201
rect 9770 15127 9826 15136
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9678 13424 9734 13433
rect 9678 13359 9734 13368
rect 9692 13258 9720 13359
rect 9680 13252 9732 13258
rect 9680 13194 9732 13200
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9692 12782 9720 12922
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9692 12209 9720 12582
rect 9678 12200 9734 12209
rect 9678 12135 9734 12144
rect 9692 11898 9720 12135
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9678 11112 9734 11121
rect 9678 11047 9734 11056
rect 9692 9674 9720 11047
rect 9784 10062 9812 15127
rect 9864 15020 9916 15026
rect 9864 14962 9916 14968
rect 9876 12481 9904 14962
rect 9968 14414 9996 15286
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 9968 13161 9996 14350
rect 9954 13152 10010 13161
rect 9954 13087 10010 13096
rect 9862 12472 9918 12481
rect 10060 12442 10088 16118
rect 10152 15094 10180 16934
rect 10244 16794 10272 17224
rect 10612 17116 10640 19200
rect 10784 17128 10836 17134
rect 10612 17088 10732 17116
rect 10320 16892 10628 16901
rect 10320 16890 10326 16892
rect 10382 16890 10406 16892
rect 10462 16890 10486 16892
rect 10542 16890 10566 16892
rect 10622 16890 10628 16892
rect 10382 16838 10384 16890
rect 10564 16838 10566 16890
rect 10320 16836 10326 16838
rect 10382 16836 10406 16838
rect 10462 16836 10486 16838
rect 10542 16836 10566 16838
rect 10622 16836 10628 16838
rect 10320 16827 10628 16836
rect 10232 16788 10284 16794
rect 10232 16730 10284 16736
rect 10324 16788 10376 16794
rect 10324 16730 10376 16736
rect 10244 16114 10272 16730
rect 10336 16182 10364 16730
rect 10508 16720 10560 16726
rect 10506 16688 10508 16697
rect 10560 16688 10562 16697
rect 10506 16623 10562 16632
rect 10416 16516 10468 16522
rect 10416 16458 10468 16464
rect 10324 16176 10376 16182
rect 10324 16118 10376 16124
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 10232 15972 10284 15978
rect 10232 15914 10284 15920
rect 10140 15088 10192 15094
rect 10244 15065 10272 15914
rect 10428 15910 10456 16458
rect 10704 16182 10732 17088
rect 10784 17070 10836 17076
rect 10796 16561 10824 17070
rect 10782 16552 10838 16561
rect 10980 16538 11008 19200
rect 11348 17898 11376 19200
rect 11716 17950 11744 19200
rect 11704 17944 11756 17950
rect 11348 17870 11560 17898
rect 11704 17886 11756 17892
rect 11336 17604 11388 17610
rect 11336 17546 11388 17552
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 11164 16658 11192 17274
rect 11348 17202 11376 17546
rect 11532 17338 11560 17870
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 11336 17196 11388 17202
rect 11336 17138 11388 17144
rect 11532 17134 11560 17274
rect 12084 17202 12112 19200
rect 12452 17814 12480 19200
rect 12440 17808 12492 17814
rect 12440 17750 12492 17756
rect 12624 17672 12676 17678
rect 12624 17614 12676 17620
rect 12194 17436 12502 17445
rect 12194 17434 12200 17436
rect 12256 17434 12280 17436
rect 12336 17434 12360 17436
rect 12416 17434 12440 17436
rect 12496 17434 12502 17436
rect 12256 17382 12258 17434
rect 12438 17382 12440 17434
rect 12194 17380 12200 17382
rect 12256 17380 12280 17382
rect 12336 17380 12360 17382
rect 12416 17380 12440 17382
rect 12496 17380 12502 17382
rect 12194 17371 12502 17380
rect 12072 17196 12124 17202
rect 12072 17138 12124 17144
rect 11520 17128 11572 17134
rect 11520 17070 11572 17076
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11808 16726 11836 17070
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 12268 16726 12296 16934
rect 12440 16788 12492 16794
rect 12440 16730 12492 16736
rect 11796 16720 11848 16726
rect 11796 16662 11848 16668
rect 12256 16720 12308 16726
rect 12256 16662 12308 16668
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 11244 16584 11296 16590
rect 10980 16532 11244 16538
rect 12452 16561 12480 16730
rect 12636 16590 12664 17614
rect 12820 17542 12848 19200
rect 13084 17944 13136 17950
rect 13084 17886 13136 17892
rect 12808 17536 12860 17542
rect 12808 17478 12860 17484
rect 12716 17060 12768 17066
rect 12716 17002 12768 17008
rect 12728 16590 12756 17002
rect 12624 16584 12676 16590
rect 10980 16526 11296 16532
rect 12438 16552 12494 16561
rect 10980 16510 11284 16526
rect 10782 16487 10838 16496
rect 12624 16526 12676 16532
rect 12716 16584 12768 16590
rect 12716 16526 12768 16532
rect 12438 16487 12494 16496
rect 11152 16448 11204 16454
rect 12072 16448 12124 16454
rect 11152 16390 11204 16396
rect 11886 16416 11942 16425
rect 10692 16176 10744 16182
rect 10692 16118 10744 16124
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 10692 16040 10744 16046
rect 10692 15982 10744 15988
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10320 15804 10628 15813
rect 10320 15802 10326 15804
rect 10382 15802 10406 15804
rect 10462 15802 10486 15804
rect 10542 15802 10566 15804
rect 10622 15802 10628 15804
rect 10382 15750 10384 15802
rect 10564 15750 10566 15802
rect 10320 15748 10326 15750
rect 10382 15748 10406 15750
rect 10462 15748 10486 15750
rect 10542 15748 10566 15750
rect 10622 15748 10628 15750
rect 10320 15739 10628 15748
rect 10600 15496 10652 15502
rect 10704 15484 10732 15982
rect 10784 15972 10836 15978
rect 10784 15914 10836 15920
rect 10652 15456 10732 15484
rect 10600 15438 10652 15444
rect 10140 15030 10192 15036
rect 10230 15056 10286 15065
rect 10230 14991 10286 15000
rect 10612 14958 10640 15438
rect 10600 14952 10652 14958
rect 10652 14912 10732 14940
rect 10600 14894 10652 14900
rect 10140 14816 10192 14822
rect 10140 14758 10192 14764
rect 10152 13705 10180 14758
rect 10320 14716 10628 14725
rect 10320 14714 10326 14716
rect 10382 14714 10406 14716
rect 10462 14714 10486 14716
rect 10542 14714 10566 14716
rect 10622 14714 10628 14716
rect 10382 14662 10384 14714
rect 10564 14662 10566 14714
rect 10320 14660 10326 14662
rect 10382 14660 10406 14662
rect 10462 14660 10486 14662
rect 10542 14660 10566 14662
rect 10622 14660 10628 14662
rect 10320 14651 10628 14660
rect 10704 14362 10732 14912
rect 10612 14334 10732 14362
rect 10612 14006 10640 14334
rect 10692 14272 10744 14278
rect 10796 14249 10824 15914
rect 10888 15162 10916 15982
rect 10980 15706 11008 16050
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 11164 15450 11192 16390
rect 12072 16390 12124 16396
rect 12624 16448 12676 16454
rect 12624 16390 12676 16396
rect 11886 16351 11942 16360
rect 11900 16114 11928 16351
rect 12084 16250 12112 16390
rect 12194 16348 12502 16357
rect 12194 16346 12200 16348
rect 12256 16346 12280 16348
rect 12336 16346 12360 16348
rect 12416 16346 12440 16348
rect 12496 16346 12502 16348
rect 12256 16294 12258 16346
rect 12438 16294 12440 16346
rect 12194 16292 12200 16294
rect 12256 16292 12280 16294
rect 12336 16292 12360 16294
rect 12416 16292 12440 16294
rect 12496 16292 12502 16294
rect 12194 16283 12502 16292
rect 12072 16244 12124 16250
rect 12072 16186 12124 16192
rect 11888 16108 11940 16114
rect 11888 16050 11940 16056
rect 12164 16108 12216 16114
rect 12164 16050 12216 16056
rect 12532 16108 12584 16114
rect 12532 16050 12584 16056
rect 11980 16040 12032 16046
rect 11978 16008 11980 16017
rect 12072 16040 12124 16046
rect 12032 16008 12034 16017
rect 11336 15972 11388 15978
rect 12072 15982 12124 15988
rect 11978 15943 12034 15952
rect 11336 15914 11388 15920
rect 11348 15638 11376 15914
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 11336 15632 11388 15638
rect 11336 15574 11388 15580
rect 11440 15570 11468 15846
rect 12084 15688 12112 15982
rect 11900 15660 12112 15688
rect 11612 15632 11664 15638
rect 11612 15574 11664 15580
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 11520 15564 11572 15570
rect 11520 15506 11572 15512
rect 10968 15428 11020 15434
rect 11164 15422 11468 15450
rect 10968 15370 11020 15376
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 10874 14648 10930 14657
rect 10980 14618 11008 15370
rect 11336 15360 11388 15366
rect 11336 15302 11388 15308
rect 11060 15088 11112 15094
rect 11060 15030 11112 15036
rect 10874 14583 10930 14592
rect 10968 14612 11020 14618
rect 10692 14214 10744 14220
rect 10782 14240 10838 14249
rect 10704 14090 10732 14214
rect 10782 14175 10838 14184
rect 10704 14062 10824 14090
rect 10600 14000 10652 14006
rect 10652 13960 10732 13988
rect 10600 13942 10652 13948
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 10138 13696 10194 13705
rect 10138 13631 10194 13640
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 9862 12407 9918 12416
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 9864 11824 9916 11830
rect 9864 11766 9916 11772
rect 9876 10742 9904 11766
rect 9864 10736 9916 10742
rect 9864 10678 9916 10684
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9692 9646 9812 9674
rect 9876 9654 9904 10678
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9496 9104 9548 9110
rect 9496 9046 9548 9052
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9416 7546 9444 8230
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 9402 7032 9458 7041
rect 9220 6996 9272 7002
rect 9402 6967 9458 6976
rect 9508 6984 9536 9046
rect 9784 8809 9812 9646
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 9968 9500 9996 12242
rect 9876 9472 9996 9500
rect 9770 8800 9826 8809
rect 9770 8735 9826 8744
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9586 8528 9642 8537
rect 9586 8463 9642 8472
rect 9600 7750 9628 8463
rect 9692 8022 9720 8570
rect 9784 8129 9812 8735
rect 9770 8120 9826 8129
rect 9770 8055 9826 8064
rect 9680 8016 9732 8022
rect 9680 7958 9732 7964
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9770 7712 9826 7721
rect 9770 7647 9826 7656
rect 9220 6938 9272 6944
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 9220 6792 9272 6798
rect 9416 6746 9444 6967
rect 9508 6956 9628 6984
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9220 6734 9272 6740
rect 8128 6684 8294 6712
rect 8128 6372 8156 6684
rect 8760 6656 8812 6662
rect 9128 6656 9180 6662
rect 8812 6604 8820 6644
rect 8760 6598 8820 6604
rect 9128 6598 9180 6604
rect 8446 6556 8754 6565
rect 8446 6554 8452 6556
rect 8508 6554 8532 6556
rect 8588 6554 8612 6556
rect 8668 6554 8692 6556
rect 8748 6554 8754 6556
rect 8508 6502 8510 6554
rect 8690 6502 8692 6554
rect 8446 6500 8452 6502
rect 8508 6500 8532 6502
rect 8588 6500 8612 6502
rect 8668 6500 8692 6502
rect 8748 6500 8754 6502
rect 8446 6491 8754 6500
rect 8792 6474 8820 6598
rect 8792 6458 9076 6474
rect 8792 6452 9088 6458
rect 8792 6446 9036 6452
rect 8792 6440 8820 6446
rect 8680 6412 8820 6440
rect 8208 6384 8260 6390
rect 8128 6344 8208 6372
rect 8208 6326 8260 6332
rect 8680 6202 8708 6412
rect 9036 6394 9088 6400
rect 8852 6384 8904 6390
rect 8588 6174 8708 6202
rect 8772 6344 8852 6372
rect 8390 6080 8446 6089
rect 8390 6015 8446 6024
rect 8298 5808 8354 5817
rect 8404 5778 8432 6015
rect 8298 5743 8354 5752
rect 8392 5772 8444 5778
rect 8312 5710 8340 5743
rect 8392 5714 8444 5720
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8588 5642 8616 6174
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8680 5642 8708 6054
rect 8576 5636 8628 5642
rect 8576 5578 8628 5584
rect 8668 5636 8720 5642
rect 8668 5578 8720 5584
rect 8208 5568 8260 5574
rect 8772 5556 8800 6344
rect 8852 6326 8904 6332
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 8942 6216 8998 6225
rect 8942 6151 8998 6160
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8772 5528 8820 5556
rect 8864 5545 8892 5646
rect 8208 5510 8260 5516
rect 8220 5250 8248 5510
rect 8446 5468 8754 5477
rect 8446 5466 8452 5468
rect 8508 5466 8532 5468
rect 8588 5466 8612 5468
rect 8668 5466 8692 5468
rect 8748 5466 8754 5468
rect 8508 5414 8510 5466
rect 8690 5414 8692 5466
rect 8446 5412 8452 5414
rect 8508 5412 8532 5414
rect 8588 5412 8612 5414
rect 8668 5412 8692 5414
rect 8748 5412 8754 5414
rect 8446 5403 8754 5412
rect 8792 5352 8820 5528
rect 8850 5536 8906 5545
rect 8850 5471 8906 5480
rect 8772 5324 8820 5352
rect 8772 5284 8800 5324
rect 8482 5264 8538 5273
rect 8220 5222 8340 5250
rect 8206 5128 8262 5137
rect 8206 5063 8208 5072
rect 8260 5063 8262 5072
rect 8208 5034 8260 5040
rect 7932 4684 7984 4690
rect 7932 4626 7984 4632
rect 8024 4684 8076 4690
rect 8076 4644 8248 4672
rect 8024 4626 8076 4632
rect 7932 4592 7984 4598
rect 7932 4534 7984 4540
rect 7944 4152 7972 4534
rect 8220 4170 8248 4644
rect 8312 4554 8340 5222
rect 8404 5222 8482 5250
rect 8404 5098 8432 5222
rect 8482 5199 8538 5208
rect 8588 5256 8800 5284
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 8392 5092 8444 5098
rect 8392 5034 8444 5040
rect 8496 4842 8524 5102
rect 8588 5001 8616 5256
rect 8760 5024 8812 5030
rect 8574 4992 8630 5001
rect 8956 5012 8984 6151
rect 9048 5846 9076 6258
rect 9140 6225 9168 6598
rect 9126 6216 9182 6225
rect 9126 6151 9182 6160
rect 9036 5840 9088 5846
rect 9036 5782 9088 5788
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 9048 5574 9076 5646
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 9048 5137 9076 5170
rect 9140 5166 9168 5714
rect 9128 5160 9180 5166
rect 9034 5128 9090 5137
rect 9232 5137 9260 6734
rect 9324 6718 9444 6746
rect 9324 6186 9352 6718
rect 9404 6656 9456 6662
rect 9508 6633 9536 6802
rect 9600 6662 9628 6956
rect 9680 6928 9732 6934
rect 9680 6870 9732 6876
rect 9588 6656 9640 6662
rect 9404 6598 9456 6604
rect 9494 6624 9550 6633
rect 9312 6180 9364 6186
rect 9312 6122 9364 6128
rect 9310 5944 9366 5953
rect 9416 5930 9444 6598
rect 9588 6598 9640 6604
rect 9494 6559 9550 6568
rect 9692 6338 9720 6870
rect 9784 6390 9812 7647
rect 9876 7041 9904 9472
rect 9954 8528 10010 8537
rect 9954 8463 10010 8472
rect 9968 7546 9996 8463
rect 9956 7540 10008 7546
rect 9956 7482 10008 7488
rect 9862 7032 9918 7041
rect 9862 6967 9918 6976
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9366 5902 9444 5930
rect 9508 6310 9720 6338
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 9310 5879 9366 5888
rect 9324 5846 9352 5879
rect 9508 5846 9536 6310
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 9312 5840 9364 5846
rect 9496 5840 9548 5846
rect 9312 5782 9364 5788
rect 9402 5808 9458 5817
rect 9496 5782 9548 5788
rect 9402 5743 9458 5752
rect 9416 5692 9444 5743
rect 9324 5664 9444 5692
rect 9128 5102 9180 5108
rect 9218 5128 9274 5137
rect 9034 5063 9090 5072
rect 9218 5063 9274 5072
rect 8812 4984 8984 5012
rect 8760 4966 8812 4972
rect 8574 4927 8630 4936
rect 9048 4842 9076 5063
rect 9324 5012 9352 5664
rect 9402 5400 9458 5409
rect 9508 5386 9536 5782
rect 9600 5778 9628 6190
rect 9876 6168 9904 6802
rect 10060 6458 10088 12378
rect 10152 7886 10180 13466
rect 10244 12753 10272 13874
rect 10320 13628 10628 13637
rect 10320 13626 10326 13628
rect 10382 13626 10406 13628
rect 10462 13626 10486 13628
rect 10542 13626 10566 13628
rect 10622 13626 10628 13628
rect 10382 13574 10384 13626
rect 10564 13574 10566 13626
rect 10320 13572 10326 13574
rect 10382 13572 10406 13574
rect 10462 13572 10486 13574
rect 10542 13572 10566 13574
rect 10622 13572 10628 13574
rect 10320 13563 10628 13572
rect 10230 12744 10286 12753
rect 10230 12679 10286 12688
rect 10244 11234 10272 12679
rect 10704 12646 10732 13960
rect 10796 13410 10824 14062
rect 10888 13530 10916 14583
rect 10968 14554 11020 14560
rect 10968 14408 11020 14414
rect 10966 14376 10968 14385
rect 11020 14376 11022 14385
rect 10966 14311 11022 14320
rect 10966 14240 11022 14249
rect 10966 14175 11022 14184
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10796 13382 10916 13410
rect 10784 13252 10836 13258
rect 10784 13194 10836 13200
rect 10796 12986 10824 13194
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10320 12540 10628 12549
rect 10320 12538 10326 12540
rect 10382 12538 10406 12540
rect 10462 12538 10486 12540
rect 10542 12538 10566 12540
rect 10622 12538 10628 12540
rect 10382 12486 10384 12538
rect 10564 12486 10566 12538
rect 10320 12484 10326 12486
rect 10382 12484 10406 12486
rect 10462 12484 10486 12486
rect 10542 12484 10566 12486
rect 10622 12484 10628 12486
rect 10320 12475 10628 12484
rect 10704 11937 10732 12582
rect 10322 11928 10378 11937
rect 10690 11928 10746 11937
rect 10322 11863 10324 11872
rect 10376 11863 10378 11872
rect 10612 11886 10690 11914
rect 10324 11834 10376 11840
rect 10508 11824 10560 11830
rect 10612 11812 10640 11886
rect 10690 11863 10746 11872
rect 10560 11784 10640 11812
rect 10508 11766 10560 11772
rect 10320 11452 10628 11461
rect 10320 11450 10326 11452
rect 10382 11450 10406 11452
rect 10462 11450 10486 11452
rect 10542 11450 10566 11452
rect 10622 11450 10628 11452
rect 10382 11398 10384 11450
rect 10564 11398 10566 11450
rect 10320 11396 10326 11398
rect 10382 11396 10406 11398
rect 10462 11396 10486 11398
rect 10542 11396 10566 11398
rect 10622 11396 10628 11398
rect 10320 11387 10628 11396
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10336 11234 10364 11290
rect 10244 11206 10364 11234
rect 10704 11218 10732 11863
rect 10796 11642 10824 12786
rect 10888 12306 10916 13382
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10874 11928 10930 11937
rect 10874 11863 10930 11872
rect 10888 11830 10916 11863
rect 10876 11824 10928 11830
rect 10876 11766 10928 11772
rect 10796 11614 10916 11642
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 10244 9874 10272 10950
rect 10320 10364 10628 10373
rect 10320 10362 10326 10364
rect 10382 10362 10406 10364
rect 10462 10362 10486 10364
rect 10542 10362 10566 10364
rect 10622 10362 10628 10364
rect 10382 10310 10384 10362
rect 10564 10310 10566 10362
rect 10320 10308 10326 10310
rect 10382 10308 10406 10310
rect 10462 10308 10486 10310
rect 10542 10308 10566 10310
rect 10622 10308 10628 10310
rect 10320 10299 10628 10308
rect 10704 10130 10732 11154
rect 10796 11082 10824 11494
rect 10784 11076 10836 11082
rect 10784 11018 10836 11024
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10244 9846 10364 9874
rect 10336 9674 10364 9846
rect 10704 9722 10732 10066
rect 10244 9646 10364 9674
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10244 7936 10272 9646
rect 10320 9276 10628 9285
rect 10320 9274 10326 9276
rect 10382 9274 10406 9276
rect 10462 9274 10486 9276
rect 10542 9274 10566 9276
rect 10622 9274 10628 9276
rect 10382 9222 10384 9274
rect 10564 9222 10566 9274
rect 10320 9220 10326 9222
rect 10382 9220 10406 9222
rect 10462 9220 10486 9222
rect 10542 9220 10566 9222
rect 10622 9220 10628 9222
rect 10320 9211 10628 9220
rect 10704 8974 10732 9658
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10324 8900 10376 8906
rect 10324 8842 10376 8848
rect 10336 8634 10364 8842
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10598 8664 10654 8673
rect 10324 8628 10376 8634
rect 10598 8599 10654 8608
rect 10324 8570 10376 8576
rect 10612 8362 10640 8599
rect 10600 8356 10652 8362
rect 10600 8298 10652 8304
rect 10320 8188 10628 8197
rect 10320 8186 10326 8188
rect 10382 8186 10406 8188
rect 10462 8186 10486 8188
rect 10542 8186 10566 8188
rect 10622 8186 10628 8188
rect 10382 8134 10384 8186
rect 10564 8134 10566 8186
rect 10320 8132 10326 8134
rect 10382 8132 10406 8134
rect 10462 8132 10486 8134
rect 10542 8132 10566 8134
rect 10622 8132 10628 8134
rect 10320 8123 10628 8132
rect 10244 7908 10364 7936
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10336 7324 10364 7908
rect 10704 7818 10732 8774
rect 10416 7812 10468 7818
rect 10416 7754 10468 7760
rect 10692 7812 10744 7818
rect 10692 7754 10744 7760
rect 10428 7478 10456 7754
rect 10416 7472 10468 7478
rect 10416 7414 10468 7420
rect 10244 7296 10364 7324
rect 10138 7168 10194 7177
rect 10138 7103 10194 7112
rect 10152 6769 10180 7103
rect 10244 6934 10272 7296
rect 10692 7268 10744 7274
rect 10692 7210 10744 7216
rect 10320 7100 10628 7109
rect 10320 7098 10326 7100
rect 10382 7098 10406 7100
rect 10462 7098 10486 7100
rect 10542 7098 10566 7100
rect 10622 7098 10628 7100
rect 10382 7046 10384 7098
rect 10564 7046 10566 7098
rect 10320 7044 10326 7046
rect 10382 7044 10406 7046
rect 10462 7044 10486 7046
rect 10542 7044 10566 7046
rect 10622 7044 10628 7046
rect 10320 7035 10628 7044
rect 10704 6984 10732 7210
rect 10336 6956 10732 6984
rect 10232 6928 10284 6934
rect 10232 6870 10284 6876
rect 10138 6760 10194 6769
rect 10138 6695 10194 6704
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10046 6352 10102 6361
rect 10152 6322 10180 6598
rect 10244 6361 10272 6598
rect 10336 6390 10364 6956
rect 10692 6792 10744 6798
rect 10612 6752 10692 6780
rect 10324 6384 10376 6390
rect 10230 6352 10286 6361
rect 10046 6287 10102 6296
rect 10140 6316 10192 6322
rect 10060 6236 10088 6287
rect 10324 6326 10376 6332
rect 10230 6287 10286 6296
rect 10140 6258 10192 6264
rect 9784 6140 9904 6168
rect 9968 6208 10088 6236
rect 9784 5930 9812 6140
rect 9692 5902 9812 5930
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 9588 5636 9640 5642
rect 9588 5578 9640 5584
rect 9600 5545 9628 5578
rect 9586 5536 9642 5545
rect 9586 5471 9642 5480
rect 9586 5400 9642 5409
rect 9508 5358 9586 5386
rect 9402 5335 9458 5344
rect 9586 5335 9642 5344
rect 8496 4814 8708 4842
rect 8680 4604 8708 4814
rect 8864 4826 9076 4842
rect 9140 4984 9352 5012
rect 8864 4820 9088 4826
rect 8864 4814 9036 4820
rect 8760 4752 8812 4758
rect 8758 4720 8760 4729
rect 8812 4720 8814 4729
rect 8758 4655 8814 4664
rect 8760 4616 8812 4622
rect 8404 4598 8616 4604
rect 8404 4592 8628 4598
rect 8404 4576 8576 4592
rect 8300 4548 8352 4554
rect 8300 4490 8352 4496
rect 8208 4164 8260 4170
rect 7944 4124 8064 4152
rect 7840 4072 7892 4078
rect 8036 4026 8064 4124
rect 8116 4140 8168 4146
rect 8208 4106 8260 4112
rect 8116 4082 8168 4088
rect 7840 4014 7892 4020
rect 7944 3998 8064 4026
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 7852 3505 7880 3878
rect 7838 3496 7894 3505
rect 7748 3460 7800 3466
rect 7838 3431 7894 3440
rect 7748 3402 7800 3408
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 7286 3088 7342 3097
rect 7286 3023 7288 3032
rect 7340 3023 7342 3032
rect 7288 2994 7340 3000
rect 7760 2972 7788 3402
rect 7944 3058 7972 3998
rect 8128 3924 8156 4082
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 8036 3913 8156 3924
rect 8220 3913 8248 4014
rect 8022 3904 8156 3913
rect 8078 3896 8156 3904
rect 8206 3904 8262 3913
rect 8022 3839 8078 3848
rect 8206 3839 8262 3848
rect 8036 3738 8064 3839
rect 8220 3754 8248 3839
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 8128 3726 8248 3754
rect 8024 3596 8076 3602
rect 8024 3538 8076 3544
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 7116 2876 7236 2904
rect 7576 2944 7788 2972
rect 6828 2382 6880 2388
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 6736 2304 6788 2310
rect 6736 2246 6788 2252
rect 6366 2000 6422 2009
rect 6366 1935 6422 1944
rect 6472 800 6500 2246
rect 6748 800 6776 2246
rect 6932 1358 6960 2400
rect 7010 2408 7066 2417
rect 7010 2343 7066 2352
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 6920 1352 6972 1358
rect 6920 1294 6972 1300
rect 7024 800 7052 2246
rect 7116 2038 7144 2876
rect 7194 2680 7250 2689
rect 7194 2615 7196 2624
rect 7248 2615 7250 2624
rect 7378 2680 7434 2689
rect 7378 2615 7434 2624
rect 7196 2586 7248 2592
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 7104 2032 7156 2038
rect 7104 1974 7156 1980
rect 7300 1970 7328 2382
rect 7288 1964 7340 1970
rect 7288 1906 7340 1912
rect 7392 1834 7420 2615
rect 7472 2576 7524 2582
rect 7470 2544 7472 2553
rect 7524 2544 7526 2553
rect 7470 2479 7526 2488
rect 7472 2372 7524 2378
rect 7472 2314 7524 2320
rect 7484 2281 7512 2314
rect 7470 2272 7526 2281
rect 7470 2207 7526 2216
rect 7380 1828 7432 1834
rect 7380 1770 7432 1776
rect 7576 1714 7604 2944
rect 7852 2650 7880 2994
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 7656 2372 7708 2378
rect 7656 2314 7708 2320
rect 7748 2372 7800 2378
rect 7748 2314 7800 2320
rect 7300 1686 7604 1714
rect 7300 800 7328 1686
rect 7668 1612 7696 2314
rect 7760 2145 7788 2314
rect 7932 2304 7984 2310
rect 8036 2292 8064 3538
rect 8128 3369 8156 3726
rect 8208 3528 8260 3534
rect 8312 3516 8340 4490
rect 8404 4486 8432 4576
rect 8680 4576 8760 4604
rect 8760 4558 8812 4564
rect 8576 4534 8628 4540
rect 8392 4480 8444 4486
rect 8864 4434 8892 4814
rect 9036 4762 9088 4768
rect 8944 4752 8996 4758
rect 8944 4694 8996 4700
rect 8392 4422 8444 4428
rect 8792 4406 8892 4434
rect 8446 4380 8754 4389
rect 8446 4378 8452 4380
rect 8508 4378 8532 4380
rect 8588 4378 8612 4380
rect 8668 4378 8692 4380
rect 8748 4378 8754 4380
rect 8508 4326 8510 4378
rect 8690 4326 8692 4378
rect 8446 4324 8452 4326
rect 8508 4324 8532 4326
rect 8588 4324 8612 4326
rect 8668 4324 8692 4326
rect 8748 4324 8754 4326
rect 8446 4315 8754 4324
rect 8792 4264 8820 4406
rect 8956 4321 8984 4694
rect 8942 4312 8998 4321
rect 8772 4236 8820 4264
rect 8852 4276 8904 4282
rect 8482 4176 8538 4185
rect 8666 4176 8722 4185
rect 8482 4111 8538 4120
rect 8588 4134 8666 4162
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 8260 3488 8340 3516
rect 8208 3470 8260 3476
rect 8404 3380 8432 3538
rect 8496 3505 8524 4111
rect 8588 3738 8616 4134
rect 8666 4111 8722 4120
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8482 3496 8538 3505
rect 8482 3431 8538 3440
rect 8680 3398 8708 4014
rect 8114 3360 8170 3369
rect 8114 3295 8170 3304
rect 8220 3352 8432 3380
rect 8668 3392 8720 3398
rect 8220 3126 8248 3352
rect 8772 3380 8800 4236
rect 8942 4247 8998 4256
rect 8852 4218 8904 4224
rect 8772 3352 8820 3380
rect 8668 3334 8720 3340
rect 8446 3292 8754 3301
rect 8446 3290 8452 3292
rect 8508 3290 8532 3292
rect 8588 3290 8612 3292
rect 8668 3290 8692 3292
rect 8748 3290 8754 3292
rect 8508 3238 8510 3290
rect 8690 3238 8692 3290
rect 8446 3236 8452 3238
rect 8508 3236 8532 3238
rect 8588 3236 8612 3238
rect 8668 3236 8692 3238
rect 8748 3236 8754 3238
rect 8446 3227 8754 3236
rect 8792 3176 8820 3352
rect 8772 3148 8820 3176
rect 8208 3120 8260 3126
rect 8114 3088 8170 3097
rect 8208 3062 8260 3068
rect 8114 3023 8116 3032
rect 8168 3023 8170 3032
rect 8392 3052 8444 3058
rect 8116 2994 8168 3000
rect 8392 2994 8444 3000
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 8220 2582 8248 2790
rect 8312 2650 8340 2790
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8208 2576 8260 2582
rect 8208 2518 8260 2524
rect 8298 2544 8354 2553
rect 8298 2479 8354 2488
rect 8312 2446 8340 2479
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 8208 2372 8260 2378
rect 8208 2314 8260 2320
rect 7984 2264 8064 2292
rect 7932 2246 7984 2252
rect 7746 2136 7802 2145
rect 7746 2071 7802 2080
rect 7944 1766 7972 2246
rect 8114 2136 8170 2145
rect 8114 2071 8170 2080
rect 7932 1760 7984 1766
rect 7932 1702 7984 1708
rect 7576 1584 7696 1612
rect 7576 800 7604 1584
rect 7840 1352 7892 1358
rect 7840 1294 7892 1300
rect 7852 800 7880 1294
rect 8128 800 8156 2071
rect 8220 1698 8248 2314
rect 8404 2292 8432 2994
rect 8772 2990 8800 3148
rect 8864 3058 8892 4218
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8956 3738 8984 3878
rect 9048 3738 9076 4014
rect 9140 3913 9168 4984
rect 9218 4720 9274 4729
rect 9218 4655 9274 4664
rect 9232 4010 9260 4655
rect 9416 4593 9444 5335
rect 9586 5264 9642 5273
rect 9586 5199 9642 5208
rect 9496 5092 9548 5098
rect 9496 5034 9548 5040
rect 9508 4865 9536 5034
rect 9494 4856 9550 4865
rect 9494 4791 9550 4800
rect 9496 4752 9548 4758
rect 9496 4694 9548 4700
rect 9402 4584 9458 4593
rect 9402 4519 9458 4528
rect 9310 4312 9366 4321
rect 9310 4247 9366 4256
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 9126 3904 9182 3913
rect 9126 3839 9182 3848
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 9218 3632 9274 3641
rect 9218 3567 9274 3576
rect 9232 3534 9260 3567
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 8668 2576 8720 2582
rect 8668 2518 8720 2524
rect 8850 2544 8906 2553
rect 8680 2378 8708 2518
rect 8850 2479 8906 2488
rect 8668 2372 8720 2378
rect 8668 2314 8720 2320
rect 8312 2264 8432 2292
rect 8312 2088 8340 2264
rect 8446 2204 8754 2213
rect 8446 2202 8452 2204
rect 8508 2202 8532 2204
rect 8588 2202 8612 2204
rect 8668 2202 8692 2204
rect 8748 2202 8754 2204
rect 8508 2150 8510 2202
rect 8690 2150 8692 2202
rect 8446 2148 8452 2150
rect 8508 2148 8532 2150
rect 8588 2148 8612 2150
rect 8668 2148 8692 2150
rect 8748 2148 8754 2150
rect 8446 2139 8754 2148
rect 8864 2088 8892 2479
rect 9140 2446 9168 3334
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 8944 2440 8996 2446
rect 8944 2382 8996 2388
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 8312 2060 8432 2088
rect 8208 1692 8260 1698
rect 8208 1634 8260 1640
rect 8404 800 8432 2060
rect 8680 2060 8892 2088
rect 8680 800 8708 2060
rect 8956 800 8984 2382
rect 9140 2281 9168 2382
rect 9126 2272 9182 2281
rect 9126 2207 9182 2216
rect 9232 1630 9260 2994
rect 9324 1902 9352 4247
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9416 2961 9444 4082
rect 9508 3602 9536 4694
rect 9600 4622 9628 5199
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 9508 3194 9536 3334
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9692 3040 9720 5902
rect 9772 5840 9824 5846
rect 9770 5808 9772 5817
rect 9824 5808 9826 5817
rect 9770 5743 9826 5752
rect 9772 5568 9824 5574
rect 9770 5536 9772 5545
rect 9824 5536 9826 5545
rect 9770 5471 9826 5480
rect 9772 5364 9824 5370
rect 9968 5352 9996 6208
rect 10140 6112 10192 6118
rect 10336 6100 10364 6326
rect 10612 6254 10640 6752
rect 10692 6734 10744 6740
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 10140 6054 10192 6060
rect 10244 6072 10364 6100
rect 10046 5944 10102 5953
rect 10046 5879 10102 5888
rect 10060 5710 10088 5879
rect 10152 5778 10180 6054
rect 10140 5772 10192 5778
rect 10140 5714 10192 5720
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 10244 5658 10272 6072
rect 10320 6012 10628 6021
rect 10320 6010 10326 6012
rect 10382 6010 10406 6012
rect 10462 6010 10486 6012
rect 10542 6010 10566 6012
rect 10622 6010 10628 6012
rect 10382 5958 10384 6010
rect 10564 5958 10566 6010
rect 10320 5956 10326 5958
rect 10382 5956 10406 5958
rect 10462 5956 10486 5958
rect 10542 5956 10566 5958
rect 10622 5956 10628 5958
rect 10320 5947 10628 5956
rect 10704 5896 10732 6598
rect 10520 5868 10732 5896
rect 10416 5840 10468 5846
rect 10416 5782 10468 5788
rect 10244 5630 10364 5658
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10244 5370 10272 5510
rect 10232 5364 10284 5370
rect 9968 5324 10180 5352
rect 9772 5306 9824 5312
rect 9784 4865 9812 5306
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 9956 5160 10008 5166
rect 9956 5102 10008 5108
rect 9770 4856 9826 4865
rect 9770 4791 9772 4800
rect 9824 4791 9826 4800
rect 9772 4762 9824 4768
rect 9876 4729 9904 5102
rect 9862 4720 9918 4729
rect 9862 4655 9864 4664
rect 9916 4655 9918 4664
rect 9864 4626 9916 4632
rect 9864 4548 9916 4554
rect 9864 4490 9916 4496
rect 9770 4312 9826 4321
rect 9770 4247 9826 4256
rect 9784 4146 9812 4247
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9600 3012 9720 3040
rect 9402 2952 9458 2961
rect 9402 2887 9458 2896
rect 9600 2446 9628 3012
rect 9680 2916 9732 2922
rect 9680 2858 9732 2864
rect 9404 2440 9456 2446
rect 9588 2440 9640 2446
rect 9404 2382 9456 2388
rect 9508 2400 9588 2428
rect 9416 2038 9444 2382
rect 9404 2032 9456 2038
rect 9404 1974 9456 1980
rect 9312 1896 9364 1902
rect 9312 1838 9364 1844
rect 9220 1624 9272 1630
rect 9220 1566 9272 1572
rect 9232 800 9260 1566
rect 9508 800 9536 2400
rect 9588 2382 9640 2388
rect 9692 2310 9720 2858
rect 9772 2644 9824 2650
rect 9876 2632 9904 4490
rect 9824 2604 9904 2632
rect 9772 2586 9824 2592
rect 9968 2582 9996 5102
rect 10060 4282 10088 5170
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 10046 3768 10102 3777
rect 10046 3703 10102 3712
rect 10060 3602 10088 3703
rect 10048 3596 10100 3602
rect 10048 3538 10100 3544
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 9956 2576 10008 2582
rect 9956 2518 10008 2524
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9588 2032 9640 2038
rect 9588 1974 9640 1980
rect 9600 1714 9628 1974
rect 9876 1873 9904 2382
rect 9862 1864 9918 1873
rect 9862 1799 9918 1808
rect 9600 1686 9812 1714
rect 9784 800 9812 1686
rect 10060 800 10088 2994
rect 10152 2378 10180 5324
rect 10232 5306 10284 5312
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 10244 3466 10272 5170
rect 10336 5030 10364 5630
rect 10428 5409 10456 5782
rect 10414 5400 10470 5409
rect 10414 5335 10470 5344
rect 10520 5166 10548 5868
rect 10598 5808 10654 5817
rect 10598 5743 10654 5752
rect 10612 5234 10640 5743
rect 10690 5672 10746 5681
rect 10690 5607 10746 5616
rect 10704 5574 10732 5607
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 10690 5264 10746 5273
rect 10600 5228 10652 5234
rect 10690 5199 10746 5208
rect 10600 5170 10652 5176
rect 10508 5160 10560 5166
rect 10508 5102 10560 5108
rect 10324 5024 10376 5030
rect 10612 5012 10640 5170
rect 10704 5166 10732 5199
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 10612 4984 10732 5012
rect 10324 4966 10376 4972
rect 10320 4924 10628 4933
rect 10320 4922 10326 4924
rect 10382 4922 10406 4924
rect 10462 4922 10486 4924
rect 10542 4922 10566 4924
rect 10622 4922 10628 4924
rect 10382 4870 10384 4922
rect 10564 4870 10566 4922
rect 10320 4868 10326 4870
rect 10382 4868 10406 4870
rect 10462 4868 10486 4870
rect 10542 4868 10566 4870
rect 10622 4868 10628 4870
rect 10320 4859 10628 4868
rect 10704 4690 10732 4984
rect 10796 4690 10824 11018
rect 10888 8634 10916 11614
rect 10980 10266 11008 14175
rect 11072 13938 11100 15030
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 11058 13288 11114 13297
rect 11058 13223 11114 13232
rect 11072 13190 11100 13223
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10980 7886 11008 10202
rect 11072 8498 11100 12854
rect 11164 10470 11192 14758
rect 11256 12714 11284 14894
rect 11348 14618 11376 15302
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 11440 14362 11468 15422
rect 11532 14822 11560 15506
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11520 14544 11572 14550
rect 11520 14486 11572 14492
rect 11348 14334 11468 14362
rect 11244 12708 11296 12714
rect 11244 12650 11296 12656
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 11256 10656 11284 12038
rect 11348 11830 11376 14334
rect 11532 14278 11560 14486
rect 11428 14272 11480 14278
rect 11428 14214 11480 14220
rect 11520 14272 11572 14278
rect 11520 14214 11572 14220
rect 11440 13705 11468 14214
rect 11624 14074 11652 15574
rect 11796 15360 11848 15366
rect 11796 15302 11848 15308
rect 11702 14784 11758 14793
rect 11702 14719 11758 14728
rect 11716 14414 11744 14719
rect 11808 14521 11836 15302
rect 11900 15162 11928 15660
rect 12072 15564 12124 15570
rect 12072 15506 12124 15512
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11888 14884 11940 14890
rect 11888 14826 11940 14832
rect 11794 14512 11850 14521
rect 11794 14447 11850 14456
rect 11704 14408 11756 14414
rect 11704 14350 11756 14356
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11520 13932 11572 13938
rect 11520 13874 11572 13880
rect 11426 13696 11482 13705
rect 11426 13631 11482 13640
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 11336 11824 11388 11830
rect 11336 11766 11388 11772
rect 11440 11354 11468 13126
rect 11532 12918 11560 13874
rect 11716 13802 11744 14214
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11704 13796 11756 13802
rect 11704 13738 11756 13744
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 11624 13530 11652 13670
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 11520 12912 11572 12918
rect 11520 12854 11572 12860
rect 11518 11928 11574 11937
rect 11518 11863 11520 11872
rect 11572 11863 11574 11872
rect 11520 11834 11572 11840
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11428 11348 11480 11354
rect 11428 11290 11480 11296
rect 11428 11076 11480 11082
rect 11428 11018 11480 11024
rect 11256 10628 11376 10656
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 11242 10024 11298 10033
rect 11242 9959 11244 9968
rect 11296 9959 11298 9968
rect 11244 9930 11296 9936
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 11058 7848 11114 7857
rect 10876 7812 10928 7818
rect 11058 7783 11114 7792
rect 10876 7754 10928 7760
rect 10888 6882 10916 7754
rect 11072 7546 11100 7783
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 10980 7002 11008 7482
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 10888 6854 11008 6882
rect 10876 6792 10928 6798
rect 10876 6734 10928 6740
rect 10692 4684 10744 4690
rect 10692 4626 10744 4632
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10598 4584 10654 4593
rect 10598 4519 10654 4528
rect 10612 4486 10640 4519
rect 10600 4480 10652 4486
rect 10600 4422 10652 4428
rect 10322 4312 10378 4321
rect 10322 4247 10378 4256
rect 10336 4078 10364 4247
rect 10600 4208 10652 4214
rect 10600 4150 10652 4156
rect 10324 4072 10376 4078
rect 10324 4014 10376 4020
rect 10612 3942 10640 4150
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10600 3936 10652 3942
rect 10796 3913 10824 4014
rect 10782 3904 10838 3913
rect 10600 3878 10652 3884
rect 10704 3862 10782 3890
rect 10320 3836 10628 3845
rect 10320 3834 10326 3836
rect 10382 3834 10406 3836
rect 10462 3834 10486 3836
rect 10542 3834 10566 3836
rect 10622 3834 10628 3836
rect 10382 3782 10384 3834
rect 10564 3782 10566 3834
rect 10320 3780 10326 3782
rect 10382 3780 10406 3782
rect 10462 3780 10486 3782
rect 10542 3780 10566 3782
rect 10622 3780 10628 3782
rect 10320 3771 10628 3780
rect 10428 3670 10456 3701
rect 10416 3664 10468 3670
rect 10414 3632 10416 3641
rect 10468 3632 10470 3641
rect 10414 3567 10470 3576
rect 10600 3596 10652 3602
rect 10232 3460 10284 3466
rect 10232 3402 10284 3408
rect 10428 3398 10456 3567
rect 10600 3538 10652 3544
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 10506 3088 10562 3097
rect 10506 3023 10562 3032
rect 10520 2990 10548 3023
rect 10508 2984 10560 2990
rect 10508 2926 10560 2932
rect 10612 2836 10640 3538
rect 10704 3126 10732 3862
rect 10782 3839 10838 3848
rect 10782 3768 10838 3777
rect 10782 3703 10838 3712
rect 10796 3534 10824 3703
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 10784 3392 10836 3398
rect 10784 3334 10836 3340
rect 10796 3194 10824 3334
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 10888 3126 10916 6734
rect 10980 6118 11008 6854
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10966 5944 11022 5953
rect 10966 5879 11022 5888
rect 10980 5846 11008 5879
rect 10968 5840 11020 5846
rect 10968 5782 11020 5788
rect 10968 5704 11020 5710
rect 10966 5672 10968 5681
rect 11020 5672 11022 5681
rect 10966 5607 11022 5616
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 10980 4826 11008 5306
rect 11072 5114 11100 7278
rect 11164 5710 11192 9862
rect 11348 8906 11376 10628
rect 11336 8900 11388 8906
rect 11336 8842 11388 8848
rect 11440 8378 11468 11018
rect 11256 8350 11468 8378
rect 11256 7410 11284 8350
rect 11532 8294 11560 11562
rect 11624 9450 11652 13126
rect 11716 11801 11744 13738
rect 11808 13530 11836 13806
rect 11796 13524 11848 13530
rect 11796 13466 11848 13472
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11808 12918 11836 13330
rect 11796 12912 11848 12918
rect 11796 12854 11848 12860
rect 11702 11792 11758 11801
rect 11702 11727 11758 11736
rect 11900 11354 11928 14826
rect 11992 13734 12020 15302
rect 12084 15065 12112 15506
rect 12176 15502 12204 16050
rect 12544 15706 12572 16050
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12194 15260 12502 15269
rect 12194 15258 12200 15260
rect 12256 15258 12280 15260
rect 12336 15258 12360 15260
rect 12416 15258 12440 15260
rect 12496 15258 12502 15260
rect 12256 15206 12258 15258
rect 12438 15206 12440 15258
rect 12194 15204 12200 15206
rect 12256 15204 12280 15206
rect 12336 15204 12360 15206
rect 12416 15204 12440 15206
rect 12496 15204 12502 15206
rect 12194 15195 12502 15204
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 12070 15056 12126 15065
rect 12070 14991 12126 15000
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 12084 13802 12112 14758
rect 12176 14550 12204 15098
rect 12636 15042 12664 16390
rect 12716 16040 12768 16046
rect 12716 15982 12768 15988
rect 12728 15178 12756 15982
rect 12820 15434 12848 17478
rect 12900 17128 12952 17134
rect 12900 17070 12952 17076
rect 12992 17128 13044 17134
rect 12992 17070 13044 17076
rect 12912 16794 12940 17070
rect 12900 16788 12952 16794
rect 12900 16730 12952 16736
rect 13004 16697 13032 17070
rect 13096 17066 13124 17886
rect 13084 17060 13136 17066
rect 13084 17002 13136 17008
rect 13096 16833 13124 17002
rect 13082 16824 13138 16833
rect 13082 16759 13138 16768
rect 12990 16688 13046 16697
rect 12990 16623 13046 16632
rect 12992 16584 13044 16590
rect 12992 16526 13044 16532
rect 13084 16584 13136 16590
rect 13084 16526 13136 16532
rect 12900 16516 12952 16522
rect 12900 16458 12952 16464
rect 12912 16114 12940 16458
rect 12900 16108 12952 16114
rect 12900 16050 12952 16056
rect 12900 15972 12952 15978
rect 12900 15914 12952 15920
rect 12912 15570 12940 15914
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 12808 15428 12860 15434
rect 12808 15370 12860 15376
rect 12728 15150 12848 15178
rect 12360 15014 12664 15042
rect 12714 15056 12770 15065
rect 12256 14884 12308 14890
rect 12256 14826 12308 14832
rect 12268 14657 12296 14826
rect 12254 14648 12310 14657
rect 12254 14583 12310 14592
rect 12164 14544 12216 14550
rect 12162 14512 12164 14521
rect 12216 14512 12218 14521
rect 12162 14447 12218 14456
rect 12360 14385 12388 15014
rect 12714 14991 12770 15000
rect 12728 14958 12756 14991
rect 12716 14952 12768 14958
rect 12716 14894 12768 14900
rect 12532 14816 12584 14822
rect 12532 14758 12584 14764
rect 12346 14376 12402 14385
rect 12346 14311 12402 14320
rect 12256 14272 12308 14278
rect 12440 14272 12492 14278
rect 12308 14232 12440 14260
rect 12256 14214 12308 14220
rect 12440 14214 12492 14220
rect 12194 14172 12502 14181
rect 12194 14170 12200 14172
rect 12256 14170 12280 14172
rect 12336 14170 12360 14172
rect 12416 14170 12440 14172
rect 12496 14170 12502 14172
rect 12256 14118 12258 14170
rect 12438 14118 12440 14170
rect 12194 14116 12200 14118
rect 12256 14116 12280 14118
rect 12336 14116 12360 14118
rect 12416 14116 12440 14118
rect 12496 14116 12502 14118
rect 12194 14107 12502 14116
rect 12440 14000 12492 14006
rect 12544 13977 12572 14758
rect 12624 14544 12676 14550
rect 12622 14512 12624 14521
rect 12676 14512 12678 14521
rect 12622 14447 12678 14456
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12636 14074 12664 14214
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12440 13942 12492 13948
rect 12530 13968 12586 13977
rect 12072 13796 12124 13802
rect 12072 13738 12124 13744
rect 11980 13728 12032 13734
rect 12452 13705 12480 13942
rect 12530 13903 12586 13912
rect 12728 13841 12756 14894
rect 12820 14482 12848 15150
rect 12808 14476 12860 14482
rect 12808 14418 12860 14424
rect 12714 13832 12770 13841
rect 12714 13767 12770 13776
rect 11980 13670 12032 13676
rect 12438 13696 12494 13705
rect 12820 13682 12848 14418
rect 12912 13870 12940 15506
rect 13004 15450 13032 16526
rect 13096 16289 13124 16526
rect 13082 16280 13138 16289
rect 13188 16250 13216 19200
rect 13360 17808 13412 17814
rect 13360 17750 13412 17756
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 13280 16522 13308 17138
rect 13372 16658 13400 17750
rect 13452 17740 13504 17746
rect 13452 17682 13504 17688
rect 13360 16652 13412 16658
rect 13360 16594 13412 16600
rect 13268 16516 13320 16522
rect 13268 16458 13320 16464
rect 13082 16215 13138 16224
rect 13176 16244 13228 16250
rect 13176 16186 13228 16192
rect 13188 15722 13216 16186
rect 13266 16008 13322 16017
rect 13266 15943 13322 15952
rect 13280 15910 13308 15943
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 13096 15694 13216 15722
rect 13096 15638 13124 15694
rect 13084 15632 13136 15638
rect 13084 15574 13136 15580
rect 13268 15496 13320 15502
rect 13004 15422 13216 15450
rect 13268 15438 13320 15444
rect 12992 15360 13044 15366
rect 12992 15302 13044 15308
rect 13084 15360 13136 15366
rect 13084 15302 13136 15308
rect 13004 14822 13032 15302
rect 12992 14816 13044 14822
rect 12992 14758 13044 14764
rect 12992 14476 13044 14482
rect 12992 14418 13044 14424
rect 12900 13864 12952 13870
rect 12900 13806 12952 13812
rect 12438 13631 12494 13640
rect 12636 13654 12848 13682
rect 12636 13546 12664 13654
rect 13004 13546 13032 14418
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 12544 13518 12664 13546
rect 12728 13518 13032 13546
rect 11980 13456 12032 13462
rect 11980 13398 12032 13404
rect 11992 11898 12020 13398
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 12084 12170 12112 13330
rect 12268 13258 12296 13466
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 12194 13084 12502 13093
rect 12194 13082 12200 13084
rect 12256 13082 12280 13084
rect 12336 13082 12360 13084
rect 12416 13082 12440 13084
rect 12496 13082 12502 13084
rect 12256 13030 12258 13082
rect 12438 13030 12440 13082
rect 12194 13028 12200 13030
rect 12256 13028 12280 13030
rect 12336 13028 12360 13030
rect 12416 13028 12440 13030
rect 12496 13028 12502 13030
rect 12194 13019 12502 13028
rect 12544 12900 12572 13518
rect 12360 12872 12572 12900
rect 12360 12345 12388 12872
rect 12346 12336 12402 12345
rect 12346 12271 12402 12280
rect 12530 12336 12586 12345
rect 12530 12271 12586 12280
rect 12624 12300 12676 12306
rect 12072 12164 12124 12170
rect 12072 12106 12124 12112
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 11716 9994 11744 10406
rect 11704 9988 11756 9994
rect 11704 9930 11756 9936
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11612 9444 11664 9450
rect 11612 9386 11664 9392
rect 11612 9104 11664 9110
rect 11612 9046 11664 9052
rect 11624 8566 11652 9046
rect 11716 8566 11744 9658
rect 11796 9648 11848 9654
rect 11796 9590 11848 9596
rect 11808 9382 11836 9590
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11612 8560 11664 8566
rect 11612 8502 11664 8508
rect 11704 8560 11756 8566
rect 11704 8502 11756 8508
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11440 8266 11560 8294
rect 11348 8022 11376 8230
rect 11336 8016 11388 8022
rect 11336 7958 11388 7964
rect 11440 7868 11468 8266
rect 11348 7840 11468 7868
rect 11520 7880 11572 7886
rect 11348 7721 11376 7840
rect 11520 7822 11572 7828
rect 11428 7744 11480 7750
rect 11334 7712 11390 7721
rect 11428 7686 11480 7692
rect 11334 7647 11390 7656
rect 11244 7404 11296 7410
rect 11244 7346 11296 7352
rect 11348 7313 11376 7647
rect 11334 7304 11390 7313
rect 11334 7239 11390 7248
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11348 7041 11376 7142
rect 11334 7032 11390 7041
rect 11440 7002 11468 7686
rect 11532 7342 11560 7822
rect 11612 7744 11664 7750
rect 11612 7686 11664 7692
rect 11520 7336 11572 7342
rect 11520 7278 11572 7284
rect 11520 7200 11572 7206
rect 11520 7142 11572 7148
rect 11334 6967 11390 6976
rect 11428 6996 11480 7002
rect 11428 6938 11480 6944
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11242 6624 11298 6633
rect 11242 6559 11298 6568
rect 11256 6458 11284 6559
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 11348 6225 11376 6802
rect 11532 6798 11560 7142
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11518 6624 11574 6633
rect 11518 6559 11574 6568
rect 11428 6384 11480 6390
rect 11428 6326 11480 6332
rect 11334 6216 11390 6225
rect 11334 6151 11390 6160
rect 11244 6112 11296 6118
rect 11244 6054 11296 6060
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11256 5710 11284 6054
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 11072 5086 11192 5114
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 11072 4554 11100 4762
rect 11060 4548 11112 4554
rect 11060 4490 11112 4496
rect 11058 4176 11114 4185
rect 10968 4140 11020 4146
rect 11058 4111 11114 4120
rect 10968 4082 11020 4088
rect 10980 3602 11008 4082
rect 11072 3913 11100 4111
rect 11058 3904 11114 3913
rect 11058 3839 11114 3848
rect 11072 3738 11100 3839
rect 11164 3738 11192 5086
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10966 3496 11022 3505
rect 10966 3431 11022 3440
rect 10980 3194 11008 3431
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 10692 3120 10744 3126
rect 10876 3120 10928 3126
rect 10692 3062 10744 3068
rect 10782 3088 10838 3097
rect 10876 3062 10928 3068
rect 10782 3023 10838 3032
rect 10612 2808 10732 2836
rect 10320 2748 10628 2757
rect 10320 2746 10326 2748
rect 10382 2746 10406 2748
rect 10462 2746 10486 2748
rect 10542 2746 10566 2748
rect 10622 2746 10628 2748
rect 10382 2694 10384 2746
rect 10564 2694 10566 2746
rect 10320 2692 10326 2694
rect 10382 2692 10406 2694
rect 10462 2692 10486 2694
rect 10542 2692 10566 2694
rect 10622 2692 10628 2694
rect 10320 2683 10628 2692
rect 10600 2576 10652 2582
rect 10600 2518 10652 2524
rect 10140 2372 10192 2378
rect 10140 2314 10192 2320
rect 10324 2372 10376 2378
rect 10324 2314 10376 2320
rect 10336 800 10364 2314
rect 10612 800 10640 2518
rect 10704 1737 10732 2808
rect 10796 2514 10824 3023
rect 10784 2508 10836 2514
rect 10784 2450 10836 2456
rect 10782 2408 10838 2417
rect 10782 2343 10784 2352
rect 10836 2343 10838 2352
rect 10784 2314 10836 2320
rect 10690 1728 10746 1737
rect 10690 1663 10746 1672
rect 10888 800 10916 3062
rect 11072 2972 11100 3674
rect 11152 2984 11204 2990
rect 11072 2944 11152 2972
rect 11152 2926 11204 2932
rect 11256 2446 11284 5646
rect 11348 5302 11376 6054
rect 11440 5574 11468 6326
rect 11428 5568 11480 5574
rect 11428 5510 11480 5516
rect 11426 5400 11482 5409
rect 11426 5335 11482 5344
rect 11336 5296 11388 5302
rect 11336 5238 11388 5244
rect 11440 5166 11468 5335
rect 11428 5160 11480 5166
rect 11428 5102 11480 5108
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 11348 4826 11376 4966
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 11348 4146 11376 4422
rect 11440 4185 11468 5102
rect 11532 4321 11560 6559
rect 11518 4312 11574 4321
rect 11518 4247 11574 4256
rect 11426 4176 11482 4185
rect 11336 4140 11388 4146
rect 11426 4111 11482 4120
rect 11336 4082 11388 4088
rect 11348 4049 11376 4082
rect 11428 4072 11480 4078
rect 11334 4040 11390 4049
rect 11428 4014 11480 4020
rect 11334 3975 11390 3984
rect 11440 3924 11468 4014
rect 11348 3896 11468 3924
rect 11520 3936 11572 3942
rect 11348 3670 11376 3896
rect 11520 3878 11572 3884
rect 11336 3664 11388 3670
rect 11336 3606 11388 3612
rect 11428 3664 11480 3670
rect 11428 3606 11480 3612
rect 11336 2848 11388 2854
rect 11334 2816 11336 2825
rect 11388 2816 11390 2825
rect 11334 2751 11390 2760
rect 11440 2689 11468 3606
rect 11426 2680 11482 2689
rect 11426 2615 11482 2624
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 11152 1760 11204 1766
rect 11152 1702 11204 1708
rect 11164 800 11192 1702
rect 11440 800 11468 2615
rect 11532 1465 11560 3878
rect 11624 2446 11652 7686
rect 11716 3058 11744 8366
rect 11808 7954 11836 9318
rect 11900 9110 11928 11154
rect 11992 9489 12020 11698
rect 12084 11558 12112 12106
rect 12194 11996 12502 12005
rect 12194 11994 12200 11996
rect 12256 11994 12280 11996
rect 12336 11994 12360 11996
rect 12416 11994 12440 11996
rect 12496 11994 12502 11996
rect 12256 11942 12258 11994
rect 12438 11942 12440 11994
rect 12194 11940 12200 11942
rect 12256 11940 12280 11942
rect 12336 11940 12360 11942
rect 12416 11940 12440 11942
rect 12496 11940 12502 11942
rect 12194 11931 12502 11940
rect 12256 11824 12308 11830
rect 12256 11766 12308 11772
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 12084 11218 12112 11494
rect 12268 11286 12296 11766
rect 12348 11688 12400 11694
rect 12348 11630 12400 11636
rect 12256 11280 12308 11286
rect 12256 11222 12308 11228
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 12360 11150 12388 11630
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12194 10908 12502 10917
rect 12194 10906 12200 10908
rect 12256 10906 12280 10908
rect 12336 10906 12360 10908
rect 12416 10906 12440 10908
rect 12496 10906 12502 10908
rect 12256 10854 12258 10906
rect 12438 10854 12440 10906
rect 12194 10852 12200 10854
rect 12256 10852 12280 10854
rect 12336 10852 12360 10854
rect 12416 10852 12440 10854
rect 12496 10852 12502 10854
rect 12194 10843 12502 10852
rect 12070 10296 12126 10305
rect 12070 10231 12126 10240
rect 12084 10130 12112 10231
rect 12072 10124 12124 10130
rect 12072 10066 12124 10072
rect 11978 9480 12034 9489
rect 11978 9415 12034 9424
rect 12084 9353 12112 10066
rect 12194 9820 12502 9829
rect 12194 9818 12200 9820
rect 12256 9818 12280 9820
rect 12336 9818 12360 9820
rect 12416 9818 12440 9820
rect 12496 9818 12502 9820
rect 12256 9766 12258 9818
rect 12438 9766 12440 9818
rect 12194 9764 12200 9766
rect 12256 9764 12280 9766
rect 12336 9764 12360 9766
rect 12416 9764 12440 9766
rect 12496 9764 12502 9766
rect 12194 9755 12502 9764
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 12070 9344 12126 9353
rect 12070 9279 12126 9288
rect 12176 9110 12204 9454
rect 12544 9110 12572 12271
rect 12624 12242 12676 12248
rect 12636 12170 12664 12242
rect 12624 12164 12676 12170
rect 12624 12106 12676 12112
rect 12728 10962 12756 13518
rect 12992 13456 13044 13462
rect 12992 13398 13044 13404
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12636 10934 12756 10962
rect 12636 10266 12664 10934
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12716 10124 12768 10130
rect 12716 10066 12768 10072
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12636 9722 12664 9998
rect 12728 9897 12756 10066
rect 12820 10033 12848 13330
rect 13004 12866 13032 13398
rect 13096 12986 13124 15302
rect 13188 14482 13216 15422
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 13176 14340 13228 14346
rect 13176 14282 13228 14288
rect 13188 14074 13216 14282
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13176 13456 13228 13462
rect 13176 13398 13228 13404
rect 13188 13002 13216 13398
rect 13280 13258 13308 15438
rect 13372 15162 13400 16594
rect 13464 15638 13492 17682
rect 13556 16182 13584 19200
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13636 17536 13688 17542
rect 13636 17478 13688 17484
rect 13648 17134 13676 17478
rect 13740 17202 13768 17818
rect 13924 17202 13952 19200
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 13912 17196 13964 17202
rect 13912 17138 13964 17144
rect 13636 17128 13688 17134
rect 13636 17070 13688 17076
rect 13910 17096 13966 17105
rect 14292 17082 14320 19200
rect 14292 17054 14504 17082
rect 13910 17031 13966 17040
rect 13728 16992 13780 16998
rect 13728 16934 13780 16940
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13544 16176 13596 16182
rect 13544 16118 13596 16124
rect 13452 15632 13504 15638
rect 13452 15574 13504 15580
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 13360 15156 13412 15162
rect 13360 15098 13412 15104
rect 13360 14952 13412 14958
rect 13360 14894 13412 14900
rect 13268 13252 13320 13258
rect 13268 13194 13320 13200
rect 13280 13161 13308 13194
rect 13266 13152 13322 13161
rect 13266 13087 13322 13096
rect 13084 12980 13136 12986
rect 13188 12974 13308 13002
rect 13084 12922 13136 12928
rect 13280 12918 13308 12974
rect 13268 12912 13320 12918
rect 13004 12838 13124 12866
rect 13372 12889 13400 14894
rect 13464 14074 13492 15302
rect 13556 15042 13584 16118
rect 13648 15978 13676 16526
rect 13636 15972 13688 15978
rect 13636 15914 13688 15920
rect 13648 15366 13676 15914
rect 13636 15360 13688 15366
rect 13636 15302 13688 15308
rect 13556 15014 13676 15042
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13556 14618 13584 14758
rect 13648 14618 13676 15014
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13636 14612 13688 14618
rect 13636 14554 13688 14560
rect 13544 14340 13596 14346
rect 13544 14282 13596 14288
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13452 13796 13504 13802
rect 13452 13738 13504 13744
rect 13464 13190 13492 13738
rect 13556 13705 13584 14282
rect 13636 13728 13688 13734
rect 13542 13696 13598 13705
rect 13636 13670 13688 13676
rect 13542 13631 13598 13640
rect 13542 13560 13598 13569
rect 13542 13495 13544 13504
rect 13596 13495 13598 13504
rect 13544 13466 13596 13472
rect 13452 13184 13504 13190
rect 13452 13126 13504 13132
rect 13452 12912 13504 12918
rect 13268 12854 13320 12860
rect 13358 12880 13414 12889
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 13004 11762 13032 12378
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12990 10568 13046 10577
rect 12806 10024 12862 10033
rect 12806 9959 12862 9968
rect 12714 9888 12770 9897
rect 12714 9823 12770 9832
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12820 9586 12848 9959
rect 12912 9722 12940 10542
rect 12990 10503 12992 10512
rect 13044 10503 13046 10512
rect 12992 10474 13044 10480
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 12900 9716 12952 9722
rect 12900 9658 12952 9664
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12636 9382 12664 9522
rect 12806 9480 12862 9489
rect 12806 9415 12808 9424
rect 12860 9415 12862 9424
rect 12808 9386 12860 9392
rect 12624 9376 12676 9382
rect 13004 9364 13032 10202
rect 13096 9518 13124 12838
rect 13176 12844 13228 12850
rect 13452 12854 13504 12860
rect 13358 12815 13414 12824
rect 13176 12786 13228 12792
rect 13188 10010 13216 12786
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 13280 11830 13308 12582
rect 13372 12306 13400 12718
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 13268 11824 13320 11830
rect 13268 11766 13320 11772
rect 13358 11792 13414 11801
rect 13358 11727 13414 11736
rect 13372 11286 13400 11727
rect 13360 11280 13412 11286
rect 13360 11222 13412 11228
rect 13268 10804 13320 10810
rect 13268 10746 13320 10752
rect 13280 10470 13308 10746
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13268 10464 13320 10470
rect 13268 10406 13320 10412
rect 13372 10266 13400 10610
rect 13464 10554 13492 12854
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 13556 11354 13584 12718
rect 13648 12442 13676 13670
rect 13740 13530 13768 16934
rect 13820 16516 13872 16522
rect 13820 16458 13872 16464
rect 13832 15434 13860 16458
rect 13924 15706 13952 17031
rect 14068 16892 14376 16901
rect 14068 16890 14074 16892
rect 14130 16890 14154 16892
rect 14210 16890 14234 16892
rect 14290 16890 14314 16892
rect 14370 16890 14376 16892
rect 14130 16838 14132 16890
rect 14312 16838 14314 16890
rect 14068 16836 14074 16838
rect 14130 16836 14154 16838
rect 14210 16836 14234 16838
rect 14290 16836 14314 16838
rect 14370 16836 14376 16838
rect 14068 16827 14376 16836
rect 14096 16652 14148 16658
rect 14096 16594 14148 16600
rect 14108 16250 14136 16594
rect 14096 16244 14148 16250
rect 14096 16186 14148 16192
rect 14476 16130 14504 17054
rect 14476 16114 14596 16130
rect 14464 16108 14596 16114
rect 14516 16102 14596 16108
rect 14464 16050 14516 16056
rect 14004 16040 14056 16046
rect 14002 16008 14004 16017
rect 14056 16008 14058 16017
rect 14002 15943 14058 15952
rect 14068 15804 14376 15813
rect 14068 15802 14074 15804
rect 14130 15802 14154 15804
rect 14210 15802 14234 15804
rect 14290 15802 14314 15804
rect 14370 15802 14376 15804
rect 14130 15750 14132 15802
rect 14312 15750 14314 15802
rect 14068 15748 14074 15750
rect 14130 15748 14154 15750
rect 14210 15748 14234 15750
rect 14290 15748 14314 15750
rect 14370 15748 14376 15750
rect 14068 15739 14376 15748
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 14464 15632 14516 15638
rect 14462 15600 14464 15609
rect 14516 15600 14518 15609
rect 13912 15564 13964 15570
rect 14462 15535 14518 15544
rect 13912 15506 13964 15512
rect 13820 15428 13872 15434
rect 13820 15370 13872 15376
rect 13820 15088 13872 15094
rect 13820 15030 13872 15036
rect 13832 14074 13860 15030
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13924 13954 13952 15506
rect 14004 15428 14056 15434
rect 14004 15370 14056 15376
rect 14016 15026 14044 15370
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 14068 14716 14376 14725
rect 14068 14714 14074 14716
rect 14130 14714 14154 14716
rect 14210 14714 14234 14716
rect 14290 14714 14314 14716
rect 14370 14714 14376 14716
rect 14130 14662 14132 14714
rect 14312 14662 14314 14714
rect 14068 14660 14074 14662
rect 14130 14660 14154 14662
rect 14210 14660 14234 14662
rect 14290 14660 14314 14662
rect 14370 14660 14376 14662
rect 14068 14651 14376 14660
rect 14004 14476 14056 14482
rect 14004 14418 14056 14424
rect 13832 13926 13952 13954
rect 13832 13870 13860 13926
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13912 13864 13964 13870
rect 13912 13806 13964 13812
rect 13818 13560 13874 13569
rect 13728 13524 13780 13530
rect 13818 13495 13820 13504
rect 13728 13466 13780 13472
rect 13872 13495 13874 13504
rect 13820 13466 13872 13472
rect 13832 13258 13860 13466
rect 13820 13252 13872 13258
rect 13820 13194 13872 13200
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13648 11218 13676 11494
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13464 10526 13676 10554
rect 13740 10538 13768 12922
rect 13832 12170 13860 12922
rect 13924 12442 13952 13806
rect 14016 13802 14044 14418
rect 14096 14272 14148 14278
rect 14096 14214 14148 14220
rect 14004 13796 14056 13802
rect 14004 13738 14056 13744
rect 14108 13734 14136 14214
rect 14096 13728 14148 13734
rect 14096 13670 14148 13676
rect 14464 13728 14516 13734
rect 14464 13670 14516 13676
rect 14068 13628 14376 13637
rect 14068 13626 14074 13628
rect 14130 13626 14154 13628
rect 14210 13626 14234 13628
rect 14290 13626 14314 13628
rect 14370 13626 14376 13628
rect 14130 13574 14132 13626
rect 14312 13574 14314 13626
rect 14068 13572 14074 13574
rect 14130 13572 14154 13574
rect 14210 13572 14234 13574
rect 14290 13572 14314 13574
rect 14370 13572 14376 13574
rect 14068 13563 14376 13572
rect 14476 13433 14504 13670
rect 14568 13530 14596 16102
rect 14660 15638 14688 19200
rect 14832 16652 14884 16658
rect 14832 16594 14884 16600
rect 14740 16176 14792 16182
rect 14740 16118 14792 16124
rect 14648 15632 14700 15638
rect 14648 15574 14700 15580
rect 14648 15496 14700 15502
rect 14648 15438 14700 15444
rect 14660 15337 14688 15438
rect 14646 15328 14702 15337
rect 14646 15263 14702 15272
rect 14752 14906 14780 16118
rect 14660 14878 14780 14906
rect 14660 14618 14688 14878
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 14648 13932 14700 13938
rect 14648 13874 14700 13880
rect 14660 13530 14688 13874
rect 14556 13524 14608 13530
rect 14556 13466 14608 13472
rect 14648 13524 14700 13530
rect 14648 13466 14700 13472
rect 14462 13424 14518 13433
rect 14462 13359 14518 13368
rect 14556 13388 14608 13394
rect 14556 13330 14608 13336
rect 14004 13184 14056 13190
rect 14280 13184 14332 13190
rect 14004 13126 14056 13132
rect 14278 13152 14280 13161
rect 14332 13152 14334 13161
rect 14016 12782 14044 13126
rect 14278 13087 14334 13096
rect 14464 12980 14516 12986
rect 14464 12922 14516 12928
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 14068 12540 14376 12549
rect 14068 12538 14074 12540
rect 14130 12538 14154 12540
rect 14210 12538 14234 12540
rect 14290 12538 14314 12540
rect 14370 12538 14376 12540
rect 14130 12486 14132 12538
rect 14312 12486 14314 12538
rect 14068 12484 14074 12486
rect 14130 12484 14154 12486
rect 14210 12484 14234 12486
rect 14290 12484 14314 12486
rect 14370 12484 14376 12486
rect 14068 12475 14376 12484
rect 13912 12436 13964 12442
rect 13912 12378 13964 12384
rect 14188 12368 14240 12374
rect 14188 12310 14240 12316
rect 13912 12232 13964 12238
rect 13912 12174 13964 12180
rect 13820 12164 13872 12170
rect 13820 12106 13872 12112
rect 13924 11218 13952 12174
rect 14200 11898 14228 12310
rect 14476 12186 14504 12922
rect 14568 12374 14596 13330
rect 14646 13288 14702 13297
rect 14646 13223 14702 13232
rect 14660 12782 14688 13223
rect 14648 12776 14700 12782
rect 14648 12718 14700 12724
rect 14556 12368 14608 12374
rect 14556 12310 14608 12316
rect 14660 12306 14688 12718
rect 14648 12300 14700 12306
rect 14648 12242 14700 12248
rect 14752 12238 14780 14758
rect 14844 12986 14872 16594
rect 15028 16538 15056 19200
rect 15200 16992 15252 16998
rect 15200 16934 15252 16940
rect 14936 16510 15056 16538
rect 14936 15094 14964 16510
rect 15016 16448 15068 16454
rect 15016 16390 15068 16396
rect 15028 16153 15056 16390
rect 15014 16144 15070 16153
rect 15014 16079 15070 16088
rect 15212 15162 15240 16934
rect 15396 16114 15424 19200
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15568 16448 15620 16454
rect 15568 16390 15620 16396
rect 15384 16108 15436 16114
rect 15384 16050 15436 16056
rect 15396 15994 15424 16050
rect 15396 15966 15516 15994
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15200 15156 15252 15162
rect 15200 15098 15252 15104
rect 14924 15088 14976 15094
rect 14976 15036 15056 15042
rect 14924 15030 15056 15036
rect 14936 15014 15056 15030
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 14832 12980 14884 12986
rect 14832 12922 14884 12928
rect 14832 12708 14884 12714
rect 14832 12650 14884 12656
rect 14740 12232 14792 12238
rect 14476 12158 14596 12186
rect 14740 12174 14792 12180
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14068 11452 14376 11461
rect 14068 11450 14074 11452
rect 14130 11450 14154 11452
rect 14210 11450 14234 11452
rect 14290 11450 14314 11452
rect 14370 11450 14376 11452
rect 14130 11398 14132 11450
rect 14312 11398 14314 11450
rect 14068 11396 14074 11398
rect 14130 11396 14154 11398
rect 14210 11396 14234 11398
rect 14290 11396 14314 11398
rect 14370 11396 14376 11398
rect 14068 11387 14376 11396
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 13924 10606 13952 11154
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 13912 10600 13964 10606
rect 13912 10542 13964 10548
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 13266 10160 13322 10169
rect 13266 10095 13268 10104
rect 13320 10095 13322 10104
rect 13268 10066 13320 10072
rect 13450 10024 13506 10033
rect 13188 9982 13308 10010
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 13188 9364 13216 9454
rect 13004 9336 13216 9364
rect 12624 9318 12676 9324
rect 11888 9104 11940 9110
rect 11888 9046 11940 9052
rect 12164 9104 12216 9110
rect 12164 9046 12216 9052
rect 12532 9104 12584 9110
rect 12532 9046 12584 9052
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 11992 8809 12020 8978
rect 12072 8832 12124 8838
rect 11978 8800 12034 8809
rect 12072 8774 12124 8780
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 11978 8735 12034 8744
rect 12084 8537 12112 8774
rect 12194 8732 12502 8741
rect 12194 8730 12200 8732
rect 12256 8730 12280 8732
rect 12336 8730 12360 8732
rect 12416 8730 12440 8732
rect 12496 8730 12502 8732
rect 12256 8678 12258 8730
rect 12438 8678 12440 8730
rect 12194 8676 12200 8678
rect 12256 8676 12280 8678
rect 12336 8676 12360 8678
rect 12416 8676 12440 8678
rect 12496 8676 12502 8678
rect 12194 8667 12502 8676
rect 11886 8528 11942 8537
rect 11886 8463 11888 8472
rect 11940 8463 11942 8472
rect 12070 8528 12126 8537
rect 12070 8463 12126 8472
rect 11888 8434 11940 8440
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 12346 8392 12402 8401
rect 11888 8356 11940 8362
rect 11888 8298 11940 8304
rect 11796 7948 11848 7954
rect 11796 7890 11848 7896
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 11808 7002 11836 7482
rect 11796 6996 11848 7002
rect 11796 6938 11848 6944
rect 11900 6934 11928 8298
rect 11888 6928 11940 6934
rect 11794 6896 11850 6905
rect 11888 6870 11940 6876
rect 11794 6831 11796 6840
rect 11848 6831 11850 6840
rect 11796 6802 11848 6808
rect 11886 6760 11942 6769
rect 11886 6695 11942 6704
rect 11900 6662 11928 6695
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11808 6322 11836 6598
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11992 6118 12020 8366
rect 12346 8327 12348 8336
rect 12400 8327 12402 8336
rect 12348 8298 12400 8304
rect 12072 8016 12124 8022
rect 12072 7958 12124 7964
rect 12162 7984 12218 7993
rect 12084 7041 12112 7958
rect 12162 7919 12164 7928
rect 12216 7919 12218 7928
rect 12164 7890 12216 7896
rect 12544 7857 12572 8774
rect 12530 7848 12586 7857
rect 12530 7783 12586 7792
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12194 7644 12502 7653
rect 12194 7642 12200 7644
rect 12256 7642 12280 7644
rect 12336 7642 12360 7644
rect 12416 7642 12440 7644
rect 12496 7642 12502 7644
rect 12256 7590 12258 7642
rect 12438 7590 12440 7642
rect 12194 7588 12200 7590
rect 12256 7588 12280 7590
rect 12336 7588 12360 7590
rect 12416 7588 12440 7590
rect 12496 7588 12502 7590
rect 12194 7579 12502 7588
rect 12164 7540 12216 7546
rect 12164 7482 12216 7488
rect 12348 7540 12400 7546
rect 12348 7482 12400 7488
rect 12176 7313 12204 7482
rect 12360 7449 12388 7482
rect 12346 7440 12402 7449
rect 12346 7375 12402 7384
rect 12162 7304 12218 7313
rect 12162 7239 12218 7248
rect 12162 7168 12218 7177
rect 12162 7103 12218 7112
rect 12070 7032 12126 7041
rect 12070 6967 12126 6976
rect 12176 6644 12204 7103
rect 12084 6616 12204 6644
rect 12084 6458 12112 6616
rect 12194 6556 12502 6565
rect 12194 6554 12200 6556
rect 12256 6554 12280 6556
rect 12336 6554 12360 6556
rect 12416 6554 12440 6556
rect 12496 6554 12502 6556
rect 12256 6502 12258 6554
rect 12438 6502 12440 6554
rect 12194 6500 12200 6502
rect 12256 6500 12280 6502
rect 12336 6500 12360 6502
rect 12416 6500 12440 6502
rect 12496 6500 12502 6502
rect 12194 6491 12502 6500
rect 12072 6452 12124 6458
rect 12072 6394 12124 6400
rect 12164 6316 12216 6322
rect 12084 6276 12164 6304
rect 11980 6112 12032 6118
rect 11886 6080 11942 6089
rect 11980 6054 12032 6060
rect 11886 6015 11942 6024
rect 11796 5840 11848 5846
rect 11796 5782 11848 5788
rect 11808 5681 11836 5782
rect 11794 5672 11850 5681
rect 11794 5607 11850 5616
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11808 3194 11836 5510
rect 11900 5370 11928 6015
rect 11980 5704 12032 5710
rect 11978 5672 11980 5681
rect 12032 5672 12034 5681
rect 11978 5607 12034 5616
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 11978 4992 12034 5001
rect 11978 4927 12034 4936
rect 11992 4604 12020 4927
rect 12084 4758 12112 6276
rect 12164 6258 12216 6264
rect 12438 6216 12494 6225
rect 12438 6151 12494 6160
rect 12348 6112 12400 6118
rect 12348 6054 12400 6060
rect 12360 5574 12388 6054
rect 12452 5778 12480 6151
rect 12440 5772 12492 5778
rect 12544 5760 12572 7686
rect 12636 7274 12664 9318
rect 13084 9104 13136 9110
rect 13084 9046 13136 9052
rect 12992 8900 13044 8906
rect 12992 8842 13044 8848
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12808 8560 12860 8566
rect 12728 8508 12808 8514
rect 12728 8502 12860 8508
rect 12728 8486 12848 8502
rect 12728 8090 12756 8486
rect 12808 8424 12860 8430
rect 12808 8366 12860 8372
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12624 7268 12676 7274
rect 12624 7210 12676 7216
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12636 6458 12664 6598
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12728 6361 12756 7346
rect 12820 6662 12848 8366
rect 12912 7954 12940 8774
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 12900 7472 12952 7478
rect 12898 7440 12900 7449
rect 12952 7440 12954 7449
rect 13004 7410 13032 8842
rect 13096 7478 13124 9046
rect 13188 8838 13216 9336
rect 13280 8974 13308 9982
rect 13450 9959 13506 9968
rect 13464 9926 13492 9959
rect 13452 9920 13504 9926
rect 13358 9888 13414 9897
rect 13452 9862 13504 9868
rect 13358 9823 13414 9832
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 13176 7948 13228 7954
rect 13176 7890 13228 7896
rect 13084 7472 13136 7478
rect 13084 7414 13136 7420
rect 12898 7375 12954 7384
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 12900 7268 12952 7274
rect 12900 7210 12952 7216
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12714 6352 12770 6361
rect 12912 6338 12940 7210
rect 13084 7200 13136 7206
rect 13084 7142 13136 7148
rect 12992 6724 13044 6730
rect 12992 6666 13044 6672
rect 13004 6458 13032 6666
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 12912 6310 13032 6338
rect 12714 6287 12716 6296
rect 12768 6287 12770 6296
rect 12716 6258 12768 6264
rect 12624 6248 12676 6254
rect 12622 6216 12624 6225
rect 12728 6227 12756 6258
rect 12900 6248 12952 6254
rect 12676 6216 12678 6225
rect 12900 6190 12952 6196
rect 12622 6151 12678 6160
rect 12636 5914 12664 6151
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12912 5817 12940 6190
rect 12898 5808 12954 5817
rect 12544 5732 12664 5760
rect 12898 5743 12954 5752
rect 12440 5714 12492 5720
rect 12530 5672 12586 5681
rect 12530 5607 12586 5616
rect 12348 5568 12400 5574
rect 12348 5510 12400 5516
rect 12194 5468 12502 5477
rect 12194 5466 12200 5468
rect 12256 5466 12280 5468
rect 12336 5466 12360 5468
rect 12416 5466 12440 5468
rect 12496 5466 12502 5468
rect 12256 5414 12258 5466
rect 12438 5414 12440 5466
rect 12194 5412 12200 5414
rect 12256 5412 12280 5414
rect 12336 5412 12360 5414
rect 12416 5412 12440 5414
rect 12496 5412 12502 5414
rect 12194 5403 12502 5412
rect 12256 5364 12308 5370
rect 12256 5306 12308 5312
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12162 4856 12218 4865
rect 12162 4791 12218 4800
rect 12072 4752 12124 4758
rect 12072 4694 12124 4700
rect 12072 4616 12124 4622
rect 11992 4576 12072 4604
rect 12072 4558 12124 4564
rect 11980 4480 12032 4486
rect 11900 4440 11980 4468
rect 11900 3534 11928 4440
rect 11980 4422 12032 4428
rect 11978 4040 12034 4049
rect 11978 3975 12034 3984
rect 11992 3602 12020 3975
rect 11980 3596 12032 3602
rect 11980 3538 12032 3544
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11980 3460 12032 3466
rect 11980 3402 12032 3408
rect 11888 3392 11940 3398
rect 11888 3334 11940 3340
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11794 3088 11850 3097
rect 11704 3052 11756 3058
rect 11794 3023 11850 3032
rect 11704 2994 11756 3000
rect 11704 2848 11756 2854
rect 11704 2790 11756 2796
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 11624 1766 11652 2382
rect 11612 1760 11664 1766
rect 11612 1702 11664 1708
rect 11518 1456 11574 1465
rect 11518 1391 11574 1400
rect 11716 800 11744 2790
rect 11808 2514 11836 3023
rect 11900 2514 11928 3334
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 11888 2508 11940 2514
rect 11888 2450 11940 2456
rect 11992 800 12020 3402
rect 12084 2378 12112 4558
rect 12176 4554 12204 4791
rect 12268 4622 12296 5306
rect 12360 5137 12388 5306
rect 12440 5296 12492 5302
rect 12440 5238 12492 5244
rect 12346 5128 12402 5137
rect 12346 5063 12402 5072
rect 12452 5030 12480 5238
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12360 4826 12388 4966
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12256 4616 12308 4622
rect 12256 4558 12308 4564
rect 12164 4548 12216 4554
rect 12164 4490 12216 4496
rect 12194 4380 12502 4389
rect 12194 4378 12200 4380
rect 12256 4378 12280 4380
rect 12336 4378 12360 4380
rect 12416 4378 12440 4380
rect 12496 4378 12502 4380
rect 12256 4326 12258 4378
rect 12438 4326 12440 4378
rect 12194 4324 12200 4326
rect 12256 4324 12280 4326
rect 12336 4324 12360 4326
rect 12416 4324 12440 4326
rect 12496 4324 12502 4326
rect 12194 4315 12502 4324
rect 12256 4140 12308 4146
rect 12256 4082 12308 4088
rect 12164 4072 12216 4078
rect 12268 4049 12296 4082
rect 12164 4014 12216 4020
rect 12254 4040 12310 4049
rect 12176 3641 12204 4014
rect 12254 3975 12310 3984
rect 12162 3632 12218 3641
rect 12162 3567 12218 3576
rect 12194 3292 12502 3301
rect 12194 3290 12200 3292
rect 12256 3290 12280 3292
rect 12336 3290 12360 3292
rect 12416 3290 12440 3292
rect 12496 3290 12502 3292
rect 12256 3238 12258 3290
rect 12438 3238 12440 3290
rect 12194 3236 12200 3238
rect 12256 3236 12280 3238
rect 12336 3236 12360 3238
rect 12416 3236 12440 3238
rect 12496 3236 12502 3238
rect 12194 3227 12502 3236
rect 12544 3126 12572 5607
rect 12636 3602 12664 5732
rect 12898 5264 12954 5273
rect 12716 5228 12768 5234
rect 12898 5199 12900 5208
rect 12716 5170 12768 5176
rect 12952 5199 12954 5208
rect 12900 5170 12952 5176
rect 12728 4826 12756 5170
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12716 4548 12768 4554
rect 12716 4490 12768 4496
rect 12728 4321 12756 4490
rect 12714 4312 12770 4321
rect 12714 4247 12770 4256
rect 12820 4264 12848 5102
rect 13004 5001 13032 6310
rect 13096 5234 13124 7142
rect 13188 6866 13216 7890
rect 13176 6860 13228 6866
rect 13176 6802 13228 6808
rect 13174 6488 13230 6497
rect 13174 6423 13230 6432
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 12990 4992 13046 5001
rect 12990 4927 13046 4936
rect 12990 4856 13046 4865
rect 12990 4791 13046 4800
rect 12900 4684 12952 4690
rect 12900 4626 12952 4632
rect 12912 4457 12940 4626
rect 13004 4486 13032 4791
rect 13188 4690 13216 6423
rect 13176 4684 13228 4690
rect 13176 4626 13228 4632
rect 13280 4570 13308 8910
rect 13372 5778 13400 9823
rect 13556 9330 13584 10406
rect 13648 10010 13676 10526
rect 13728 10532 13780 10538
rect 14384 10520 14412 11086
rect 14476 10742 14504 12038
rect 14464 10736 14516 10742
rect 14464 10678 14516 10684
rect 14384 10492 14504 10520
rect 13728 10474 13780 10480
rect 14068 10364 14376 10373
rect 14068 10362 14074 10364
rect 14130 10362 14154 10364
rect 14210 10362 14234 10364
rect 14290 10362 14314 10364
rect 14370 10362 14376 10364
rect 14130 10310 14132 10362
rect 14312 10310 14314 10362
rect 14068 10308 14074 10310
rect 14130 10308 14154 10310
rect 14210 10308 14234 10310
rect 14290 10308 14314 10310
rect 14370 10308 14376 10310
rect 13818 10296 13874 10305
rect 14068 10299 14376 10308
rect 13818 10231 13874 10240
rect 13832 10130 13860 10231
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 13648 9982 13768 10010
rect 13636 9920 13688 9926
rect 13636 9862 13688 9868
rect 13648 9654 13676 9862
rect 13636 9648 13688 9654
rect 13636 9590 13688 9596
rect 13464 9302 13584 9330
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13464 8566 13492 9302
rect 13542 9208 13598 9217
rect 13542 9143 13598 9152
rect 13556 8634 13584 9143
rect 13648 8945 13676 9318
rect 13634 8936 13690 8945
rect 13634 8871 13690 8880
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13452 8560 13504 8566
rect 13452 8502 13504 8508
rect 13648 8430 13676 8774
rect 13636 8424 13688 8430
rect 13636 8366 13688 8372
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 13452 7744 13504 7750
rect 13450 7712 13452 7721
rect 13504 7712 13506 7721
rect 13450 7647 13506 7656
rect 13556 7410 13584 7890
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13452 7268 13504 7274
rect 13452 7210 13504 7216
rect 13360 5772 13412 5778
rect 13360 5714 13412 5720
rect 13372 5001 13400 5714
rect 13464 5681 13492 7210
rect 13544 7200 13596 7206
rect 13544 7142 13596 7148
rect 13556 6798 13584 7142
rect 13544 6792 13596 6798
rect 13648 6769 13676 8366
rect 13544 6734 13596 6740
rect 13634 6760 13690 6769
rect 13634 6695 13690 6704
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13542 5808 13598 5817
rect 13542 5743 13598 5752
rect 13450 5672 13506 5681
rect 13450 5607 13506 5616
rect 13556 5302 13584 5743
rect 13544 5296 13596 5302
rect 13544 5238 13596 5244
rect 13544 5160 13596 5166
rect 13544 5102 13596 5108
rect 13358 4992 13414 5001
rect 13358 4927 13414 4936
rect 13358 4720 13414 4729
rect 13358 4655 13360 4664
rect 13412 4655 13414 4664
rect 13452 4684 13504 4690
rect 13360 4626 13412 4632
rect 13452 4626 13504 4632
rect 13096 4542 13308 4570
rect 12992 4480 13044 4486
rect 12898 4448 12954 4457
rect 12992 4422 13044 4428
rect 12898 4383 12954 4392
rect 13096 4298 13124 4542
rect 13266 4448 13322 4457
rect 13266 4383 13322 4392
rect 12900 4276 12952 4282
rect 12820 4236 12900 4264
rect 13096 4270 13216 4298
rect 12900 4218 12952 4224
rect 13084 4208 13136 4214
rect 13084 4150 13136 4156
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12532 3120 12584 3126
rect 12254 3088 12310 3097
rect 12532 3062 12584 3068
rect 12254 3023 12256 3032
rect 12308 3023 12310 3032
rect 12256 2994 12308 3000
rect 12268 2854 12296 2994
rect 12532 2916 12584 2922
rect 12532 2858 12584 2864
rect 12256 2848 12308 2854
rect 12256 2790 12308 2796
rect 12072 2372 12124 2378
rect 12072 2314 12124 2320
rect 12194 2204 12502 2213
rect 12194 2202 12200 2204
rect 12256 2202 12280 2204
rect 12336 2202 12360 2204
rect 12416 2202 12440 2204
rect 12496 2202 12502 2204
rect 12256 2150 12258 2202
rect 12438 2150 12440 2202
rect 12194 2148 12200 2150
rect 12256 2148 12280 2150
rect 12336 2148 12360 2150
rect 12416 2148 12440 2150
rect 12496 2148 12502 2150
rect 12194 2139 12502 2148
rect 12256 1896 12308 1902
rect 12256 1838 12308 1844
rect 12268 800 12296 1838
rect 12544 800 12572 2858
rect 12636 2650 12664 3334
rect 12624 2644 12676 2650
rect 12624 2586 12676 2592
rect 12728 2428 12756 3674
rect 12806 3496 12862 3505
rect 12806 3431 12862 3440
rect 12820 2922 12848 3431
rect 12898 3224 12954 3233
rect 12898 3159 12954 3168
rect 12912 3058 12940 3159
rect 13004 3058 13032 4082
rect 13096 3602 13124 4150
rect 13188 4146 13216 4270
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 13084 3596 13136 3602
rect 13084 3538 13136 3544
rect 13188 3534 13216 4082
rect 13280 4010 13308 4383
rect 13372 4010 13400 4626
rect 13464 4282 13492 4626
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13556 4060 13584 5102
rect 13464 4032 13584 4060
rect 13268 4004 13320 4010
rect 13268 3946 13320 3952
rect 13360 4004 13412 4010
rect 13360 3946 13412 3952
rect 13176 3528 13228 3534
rect 13176 3470 13228 3476
rect 13084 3460 13136 3466
rect 13084 3402 13136 3408
rect 12900 3052 12952 3058
rect 12900 2994 12952 3000
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 12808 2916 12860 2922
rect 12808 2858 12860 2864
rect 12808 2440 12860 2446
rect 12728 2400 12808 2428
rect 12808 2382 12860 2388
rect 12820 800 12848 2382
rect 13096 800 13124 3402
rect 13176 2984 13228 2990
rect 13176 2926 13228 2932
rect 13188 2514 13216 2926
rect 13280 2553 13308 3946
rect 13464 3466 13492 4032
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 13452 3460 13504 3466
rect 13452 3402 13504 3408
rect 13358 3088 13414 3097
rect 13358 3023 13414 3032
rect 13266 2544 13322 2553
rect 13176 2508 13228 2514
rect 13266 2479 13322 2488
rect 13176 2450 13228 2456
rect 13188 1902 13216 2450
rect 13176 1896 13228 1902
rect 13176 1838 13228 1844
rect 13372 800 13400 3023
rect 13452 2916 13504 2922
rect 13452 2858 13504 2864
rect 13464 2292 13492 2858
rect 13556 2689 13584 3674
rect 13648 3510 13676 6598
rect 13740 6322 13768 9982
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 13832 8294 13860 9930
rect 13912 9580 13964 9586
rect 13912 9522 13964 9528
rect 13924 8634 13952 9522
rect 14016 9489 14044 10066
rect 14476 10010 14504 10492
rect 14568 10130 14596 12158
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14660 11665 14688 11698
rect 14740 11688 14792 11694
rect 14646 11656 14702 11665
rect 14740 11630 14792 11636
rect 14646 11591 14702 11600
rect 14660 11150 14688 11591
rect 14648 11144 14700 11150
rect 14648 11086 14700 11092
rect 14648 10532 14700 10538
rect 14648 10474 14700 10480
rect 14660 10266 14688 10474
rect 14752 10470 14780 11630
rect 14844 10674 14872 12650
rect 14936 11014 14964 14758
rect 15028 12986 15056 15014
rect 15212 14074 15240 15098
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 15108 13796 15160 13802
rect 15108 13738 15160 13744
rect 15120 13462 15148 13738
rect 15212 13530 15240 14010
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15108 13456 15160 13462
rect 15304 13410 15332 15846
rect 15382 14920 15438 14929
rect 15382 14855 15438 14864
rect 15396 14414 15424 14855
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 15384 14068 15436 14074
rect 15384 14010 15436 14016
rect 15108 13398 15160 13404
rect 15212 13382 15332 13410
rect 15212 13258 15240 13382
rect 15200 13252 15252 13258
rect 15200 13194 15252 13200
rect 15016 12980 15068 12986
rect 15016 12922 15068 12928
rect 15212 12646 15240 13194
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 15304 12434 15332 13126
rect 15212 12406 15332 12434
rect 14924 11008 14976 11014
rect 14924 10950 14976 10956
rect 15016 10736 15068 10742
rect 15016 10678 15068 10684
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14648 10260 14700 10266
rect 14648 10202 14700 10208
rect 14660 10130 14688 10202
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 14648 10124 14700 10130
rect 14648 10066 14700 10072
rect 14738 10024 14794 10033
rect 14476 9982 14596 10010
rect 14464 9920 14516 9926
rect 14464 9862 14516 9868
rect 14476 9722 14504 9862
rect 14464 9716 14516 9722
rect 14464 9658 14516 9664
rect 14462 9616 14518 9625
rect 14462 9551 14464 9560
rect 14516 9551 14518 9560
rect 14464 9522 14516 9528
rect 14002 9480 14058 9489
rect 14002 9415 14058 9424
rect 14068 9276 14376 9285
rect 14068 9274 14074 9276
rect 14130 9274 14154 9276
rect 14210 9274 14234 9276
rect 14290 9274 14314 9276
rect 14370 9274 14376 9276
rect 14130 9222 14132 9274
rect 14312 9222 14314 9274
rect 14068 9220 14074 9222
rect 14130 9220 14154 9222
rect 14210 9220 14234 9222
rect 14290 9220 14314 9222
rect 14370 9220 14376 9222
rect 14068 9211 14376 9220
rect 14186 9072 14242 9081
rect 14186 9007 14242 9016
rect 14370 9072 14426 9081
rect 14370 9007 14426 9016
rect 14096 8832 14148 8838
rect 14094 8800 14096 8809
rect 14148 8800 14150 8809
rect 14094 8735 14150 8744
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 14200 8498 14228 9007
rect 14280 8900 14332 8906
rect 14280 8842 14332 8848
rect 14292 8566 14320 8842
rect 14280 8560 14332 8566
rect 14280 8502 14332 8508
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 14384 8294 14412 9007
rect 14476 8838 14504 9522
rect 14568 9081 14596 9982
rect 14738 9959 14794 9968
rect 14752 9194 14780 9959
rect 14660 9166 14780 9194
rect 14554 9072 14610 9081
rect 14554 9007 14610 9016
rect 14556 8968 14608 8974
rect 14660 8956 14688 9166
rect 14740 9036 14792 9042
rect 14740 8978 14792 8984
rect 14608 8928 14688 8956
rect 14556 8910 14608 8916
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14660 8566 14688 8928
rect 14648 8560 14700 8566
rect 14648 8502 14700 8508
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 14372 8288 14424 8294
rect 14372 8230 14424 8236
rect 14068 8188 14376 8197
rect 14068 8186 14074 8188
rect 14130 8186 14154 8188
rect 14210 8186 14234 8188
rect 14290 8186 14314 8188
rect 14370 8186 14376 8188
rect 14130 8134 14132 8186
rect 14312 8134 14314 8186
rect 14068 8132 14074 8134
rect 14130 8132 14154 8134
rect 14210 8132 14234 8134
rect 14290 8132 14314 8134
rect 14370 8132 14376 8134
rect 14068 8123 14376 8132
rect 14476 8090 14504 8434
rect 14752 8412 14780 8978
rect 14568 8384 14780 8412
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 13820 8016 13872 8022
rect 13820 7958 13872 7964
rect 13910 7984 13966 7993
rect 13832 7002 13860 7958
rect 14568 7954 14596 8384
rect 14648 8288 14700 8294
rect 14648 8230 14700 8236
rect 13910 7919 13912 7928
rect 13964 7919 13966 7928
rect 14556 7948 14608 7954
rect 13912 7890 13964 7896
rect 14556 7890 14608 7896
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 14372 7880 14424 7886
rect 14372 7822 14424 7828
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13820 6792 13872 6798
rect 13818 6760 13820 6769
rect 13872 6760 13874 6769
rect 13818 6695 13874 6704
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13832 6458 13860 6598
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13818 6352 13874 6361
rect 13728 6316 13780 6322
rect 13924 6322 13952 7686
rect 14108 7342 14136 7822
rect 14384 7750 14412 7822
rect 14372 7744 14424 7750
rect 14660 7721 14688 8230
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14372 7686 14424 7692
rect 14646 7712 14702 7721
rect 14384 7478 14412 7686
rect 14646 7647 14702 7656
rect 14554 7576 14610 7585
rect 14554 7511 14610 7520
rect 14372 7472 14424 7478
rect 14372 7414 14424 7420
rect 14568 7410 14596 7511
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 14370 7304 14426 7313
rect 14370 7239 14426 7248
rect 14384 7206 14412 7239
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14068 7100 14376 7109
rect 14068 7098 14074 7100
rect 14130 7098 14154 7100
rect 14210 7098 14234 7100
rect 14290 7098 14314 7100
rect 14370 7098 14376 7100
rect 14130 7046 14132 7098
rect 14312 7046 14314 7098
rect 14068 7044 14074 7046
rect 14130 7044 14154 7046
rect 14210 7044 14234 7046
rect 14290 7044 14314 7046
rect 14370 7044 14376 7046
rect 14068 7035 14376 7044
rect 14188 6996 14240 7002
rect 14188 6938 14240 6944
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 13818 6287 13874 6296
rect 13912 6316 13964 6322
rect 13728 6258 13780 6264
rect 13832 6202 13860 6287
rect 13912 6258 13964 6264
rect 13740 6174 13860 6202
rect 13740 5574 13768 6174
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13832 5953 13860 6054
rect 13818 5944 13874 5953
rect 13818 5879 13874 5888
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13740 4690 13768 5510
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13728 4684 13780 4690
rect 13728 4626 13780 4632
rect 13728 4548 13780 4554
rect 13728 4490 13780 4496
rect 13636 3504 13688 3510
rect 13636 3446 13688 3452
rect 13634 3360 13690 3369
rect 13634 3295 13690 3304
rect 13542 2680 13598 2689
rect 13542 2615 13598 2624
rect 13648 2446 13676 3295
rect 13740 2854 13768 4490
rect 13832 4146 13860 5306
rect 13924 5273 13952 6258
rect 14016 6118 14044 6802
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 14108 6633 14136 6734
rect 14094 6624 14150 6633
rect 14094 6559 14150 6568
rect 14094 6488 14150 6497
rect 14094 6423 14096 6432
rect 14148 6423 14150 6432
rect 14096 6394 14148 6400
rect 14200 6118 14228 6938
rect 14372 6928 14424 6934
rect 14372 6870 14424 6876
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14292 6225 14320 6734
rect 14384 6254 14412 6870
rect 14372 6248 14424 6254
rect 14278 6216 14334 6225
rect 14372 6190 14424 6196
rect 14278 6151 14334 6160
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 14068 6012 14376 6021
rect 14068 6010 14074 6012
rect 14130 6010 14154 6012
rect 14210 6010 14234 6012
rect 14290 6010 14314 6012
rect 14370 6010 14376 6012
rect 14130 5958 14132 6010
rect 14312 5958 14314 6010
rect 14068 5956 14074 5958
rect 14130 5956 14154 5958
rect 14210 5956 14234 5958
rect 14290 5956 14314 5958
rect 14370 5956 14376 5958
rect 14068 5947 14376 5956
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 13910 5264 13966 5273
rect 13910 5199 13966 5208
rect 14016 5148 14044 5850
rect 14186 5808 14242 5817
rect 14186 5743 14242 5752
rect 14280 5772 14332 5778
rect 14096 5704 14148 5710
rect 14094 5672 14096 5681
rect 14148 5672 14150 5681
rect 14200 5642 14228 5743
rect 14280 5714 14332 5720
rect 14094 5607 14150 5616
rect 14188 5636 14240 5642
rect 14188 5578 14240 5584
rect 14094 5400 14150 5409
rect 14094 5335 14096 5344
rect 14148 5335 14150 5344
rect 14096 5306 14148 5312
rect 14096 5160 14148 5166
rect 14016 5120 14096 5148
rect 14096 5102 14148 5108
rect 14200 5012 14228 5578
rect 14292 5302 14320 5714
rect 14372 5568 14424 5574
rect 14370 5536 14372 5545
rect 14424 5536 14426 5545
rect 14370 5471 14426 5480
rect 14476 5370 14504 7346
rect 14556 7268 14608 7274
rect 14556 7210 14608 7216
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 14280 5296 14332 5302
rect 14280 5238 14332 5244
rect 13924 4984 14228 5012
rect 14464 5024 14516 5030
rect 13924 4826 13952 4984
rect 14464 4966 14516 4972
rect 14068 4924 14376 4933
rect 14068 4922 14074 4924
rect 14130 4922 14154 4924
rect 14210 4922 14234 4924
rect 14290 4922 14314 4924
rect 14370 4922 14376 4924
rect 14130 4870 14132 4922
rect 14312 4870 14314 4922
rect 14068 4868 14074 4870
rect 14130 4868 14154 4870
rect 14210 4868 14234 4870
rect 14290 4868 14314 4870
rect 14370 4868 14376 4870
rect 14068 4859 14376 4868
rect 13912 4820 13964 4826
rect 13912 4762 13964 4768
rect 13924 4434 13952 4762
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 13924 4406 14044 4434
rect 13912 4276 13964 4282
rect 13912 4218 13964 4224
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 13832 3058 13860 3946
rect 13924 3602 13952 4218
rect 14016 4049 14044 4406
rect 14002 4040 14058 4049
rect 14002 3975 14058 3984
rect 14108 3942 14136 4558
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 14068 3836 14376 3845
rect 14068 3834 14074 3836
rect 14130 3834 14154 3836
rect 14210 3834 14234 3836
rect 14290 3834 14314 3836
rect 14370 3834 14376 3836
rect 14130 3782 14132 3834
rect 14312 3782 14314 3834
rect 14068 3780 14074 3782
rect 14130 3780 14154 3782
rect 14210 3780 14234 3782
rect 14290 3780 14314 3782
rect 14370 3780 14376 3782
rect 14068 3771 14376 3780
rect 14476 3738 14504 4966
rect 14568 4826 14596 7210
rect 14648 7200 14700 7206
rect 14648 7142 14700 7148
rect 14660 6769 14688 7142
rect 14752 6934 14780 8026
rect 14740 6928 14792 6934
rect 14740 6870 14792 6876
rect 14740 6792 14792 6798
rect 14646 6760 14702 6769
rect 14740 6734 14792 6740
rect 14646 6695 14702 6704
rect 14646 6488 14702 6497
rect 14646 6423 14648 6432
rect 14700 6423 14702 6432
rect 14648 6394 14700 6400
rect 14648 6112 14700 6118
rect 14646 6080 14648 6089
rect 14700 6080 14702 6089
rect 14646 6015 14702 6024
rect 14752 5846 14780 6734
rect 14740 5840 14792 5846
rect 14740 5782 14792 5788
rect 14648 5704 14700 5710
rect 14648 5646 14700 5652
rect 14660 5250 14688 5646
rect 14752 5370 14780 5782
rect 14844 5710 14872 10610
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 14936 10266 14964 10542
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 14924 9104 14976 9110
rect 14924 9046 14976 9052
rect 14936 8634 14964 9046
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 14936 6458 14964 8434
rect 14924 6452 14976 6458
rect 14924 6394 14976 6400
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 14740 5364 14792 5370
rect 14740 5306 14792 5312
rect 14660 5222 14780 5250
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 14660 4826 14688 5102
rect 14556 4820 14608 4826
rect 14556 4762 14608 4768
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14646 4176 14702 4185
rect 14646 4111 14702 4120
rect 14660 4078 14688 4111
rect 14648 4072 14700 4078
rect 14568 4032 14648 4060
rect 14464 3732 14516 3738
rect 14464 3674 14516 3680
rect 14094 3632 14150 3641
rect 13912 3596 13964 3602
rect 14568 3602 14596 4032
rect 14752 4060 14780 5222
rect 14844 4554 14872 5646
rect 14936 5545 14964 6394
rect 15028 5574 15056 10678
rect 15106 10024 15162 10033
rect 15106 9959 15162 9968
rect 15120 9110 15148 9959
rect 15212 9738 15240 12406
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15304 10810 15332 11494
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15396 10130 15424 14010
rect 15488 11898 15516 15966
rect 15580 13462 15608 16390
rect 15672 15026 15700 17614
rect 15764 16182 15792 19200
rect 16132 17678 16160 19200
rect 16120 17672 16172 17678
rect 16120 17614 16172 17620
rect 16500 17610 16528 19200
rect 16488 17604 16540 17610
rect 16488 17546 16540 17552
rect 16028 17196 16080 17202
rect 16028 17138 16080 17144
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15752 16176 15804 16182
rect 15752 16118 15804 16124
rect 15660 15020 15712 15026
rect 15856 15008 15884 16526
rect 15936 15428 15988 15434
rect 15936 15370 15988 15376
rect 15660 14962 15712 14968
rect 15764 14980 15884 15008
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15672 14074 15700 14418
rect 15660 14068 15712 14074
rect 15660 14010 15712 14016
rect 15568 13456 15620 13462
rect 15568 13398 15620 13404
rect 15764 13274 15792 14980
rect 15844 14884 15896 14890
rect 15844 14826 15896 14832
rect 15856 13870 15884 14826
rect 15844 13864 15896 13870
rect 15844 13806 15896 13812
rect 15672 13246 15792 13274
rect 15672 12918 15700 13246
rect 15752 13184 15804 13190
rect 15752 13126 15804 13132
rect 15660 12912 15712 12918
rect 15660 12854 15712 12860
rect 15660 12776 15712 12782
rect 15660 12718 15712 12724
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15476 10464 15528 10470
rect 15476 10406 15528 10412
rect 15488 10130 15516 10406
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15476 10124 15528 10130
rect 15476 10066 15528 10072
rect 15212 9710 15424 9738
rect 15292 9648 15344 9654
rect 15292 9590 15344 9596
rect 15200 9172 15252 9178
rect 15200 9114 15252 9120
rect 15108 9104 15160 9110
rect 15108 9046 15160 9052
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 15120 8566 15148 8910
rect 15108 8560 15160 8566
rect 15108 8502 15160 8508
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 15120 7886 15148 8366
rect 15108 7880 15160 7886
rect 15108 7822 15160 7828
rect 15106 7712 15162 7721
rect 15106 7647 15162 7656
rect 15120 7274 15148 7647
rect 15108 7268 15160 7274
rect 15108 7210 15160 7216
rect 15120 7002 15148 7210
rect 15108 6996 15160 7002
rect 15108 6938 15160 6944
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 15120 6390 15148 6734
rect 15108 6384 15160 6390
rect 15108 6326 15160 6332
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 15016 5568 15068 5574
rect 14922 5536 14978 5545
rect 15016 5510 15068 5516
rect 14922 5471 14978 5480
rect 15028 4690 15056 5510
rect 15120 5098 15148 6190
rect 15108 5092 15160 5098
rect 15108 5034 15160 5040
rect 15120 4690 15148 5034
rect 15016 4684 15068 4690
rect 15016 4626 15068 4632
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 14832 4548 14884 4554
rect 14832 4490 14884 4496
rect 14844 4282 14872 4490
rect 15108 4480 15160 4486
rect 15108 4422 15160 4428
rect 14922 4312 14978 4321
rect 14832 4276 14884 4282
rect 14922 4247 14978 4256
rect 14832 4218 14884 4224
rect 14832 4072 14884 4078
rect 14752 4032 14832 4060
rect 14648 4014 14700 4020
rect 14832 4014 14884 4020
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14094 3567 14150 3576
rect 14556 3596 14608 3602
rect 13912 3538 13964 3544
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 14016 2938 14044 3470
rect 14108 3058 14136 3567
rect 14556 3538 14608 3544
rect 14462 3496 14518 3505
rect 14462 3431 14518 3440
rect 14476 3398 14504 3431
rect 14372 3392 14424 3398
rect 14372 3334 14424 3340
rect 14464 3392 14516 3398
rect 14464 3334 14516 3340
rect 14554 3360 14610 3369
rect 14384 3210 14412 3334
rect 14554 3295 14610 3304
rect 14568 3210 14596 3295
rect 14384 3182 14596 3210
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 13832 2910 14044 2938
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 13832 2666 13860 2910
rect 13910 2816 13966 2825
rect 13910 2751 13966 2760
rect 13740 2650 13860 2666
rect 13728 2644 13860 2650
rect 13780 2638 13860 2644
rect 13728 2586 13780 2592
rect 13820 2576 13872 2582
rect 13820 2518 13872 2524
rect 13636 2440 13688 2446
rect 13636 2382 13688 2388
rect 13728 2304 13780 2310
rect 13464 2264 13676 2292
rect 13648 800 13676 2264
rect 13832 2281 13860 2518
rect 13728 2246 13780 2252
rect 13818 2272 13874 2281
rect 13740 2038 13768 2246
rect 13818 2207 13874 2216
rect 13728 2032 13780 2038
rect 13728 1974 13780 1980
rect 13924 800 13952 2751
rect 14068 2748 14376 2757
rect 14068 2746 14074 2748
rect 14130 2746 14154 2748
rect 14210 2746 14234 2748
rect 14290 2746 14314 2748
rect 14370 2746 14376 2748
rect 14130 2694 14132 2746
rect 14312 2694 14314 2746
rect 14068 2692 14074 2694
rect 14130 2692 14154 2694
rect 14210 2692 14234 2694
rect 14290 2692 14314 2694
rect 14370 2692 14376 2694
rect 14068 2683 14376 2692
rect 14464 2576 14516 2582
rect 14370 2544 14426 2553
rect 14464 2518 14516 2524
rect 14370 2479 14372 2488
rect 14424 2479 14426 2488
rect 14372 2450 14424 2456
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 14200 800 14228 2246
rect 14476 800 14504 2518
rect 14568 2378 14596 3182
rect 14556 2372 14608 2378
rect 14556 2314 14608 2320
rect 14660 1873 14688 3878
rect 14844 3534 14872 4014
rect 14936 3602 14964 4247
rect 15016 4004 15068 4010
rect 15016 3946 15068 3952
rect 14924 3596 14976 3602
rect 14924 3538 14976 3544
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 14832 3392 14884 3398
rect 14832 3334 14884 3340
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 14646 1864 14702 1873
rect 14646 1799 14702 1808
rect 14752 800 14780 3130
rect 14844 3040 14872 3334
rect 14924 3052 14976 3058
rect 14844 3012 14924 3040
rect 14924 2994 14976 3000
rect 15028 2446 15056 3946
rect 15016 2440 15068 2446
rect 15016 2382 15068 2388
rect 15120 2258 15148 4422
rect 15212 3058 15240 9114
rect 15304 9042 15332 9590
rect 15292 9036 15344 9042
rect 15292 8978 15344 8984
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 15304 6458 15332 7346
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 15396 6202 15424 9710
rect 15488 9518 15516 10066
rect 15580 9586 15608 12582
rect 15672 12238 15700 12718
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15672 10062 15700 12038
rect 15764 11218 15792 13126
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 15856 11098 15884 13806
rect 15764 11082 15884 11098
rect 15752 11076 15884 11082
rect 15804 11070 15884 11076
rect 15752 11018 15804 11024
rect 15660 10056 15712 10062
rect 15660 9998 15712 10004
rect 15568 9580 15620 9586
rect 15568 9522 15620 9528
rect 15476 9512 15528 9518
rect 15476 9454 15528 9460
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 15488 8974 15516 9318
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 15580 7410 15608 9522
rect 15660 8356 15712 8362
rect 15660 8298 15712 8304
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15568 6316 15620 6322
rect 15568 6258 15620 6264
rect 15304 6174 15424 6202
rect 15304 5234 15332 6174
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 15292 5228 15344 5234
rect 15292 5170 15344 5176
rect 15304 4214 15332 5170
rect 15292 4208 15344 4214
rect 15292 4150 15344 4156
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 15304 3534 15332 3878
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 15292 3392 15344 3398
rect 15292 3334 15344 3340
rect 15200 3052 15252 3058
rect 15200 2994 15252 3000
rect 15028 2230 15148 2258
rect 15028 800 15056 2230
rect 15304 800 15332 3334
rect 15396 2446 15424 6054
rect 15580 5914 15608 6258
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 15474 5400 15530 5409
rect 15474 5335 15476 5344
rect 15528 5335 15530 5344
rect 15476 5306 15528 5312
rect 15672 5234 15700 8298
rect 15764 6662 15792 11018
rect 15844 11008 15896 11014
rect 15844 10950 15896 10956
rect 15856 6866 15884 10950
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15856 5302 15884 6802
rect 15948 6497 15976 15370
rect 16040 11898 16068 17138
rect 16396 16992 16448 16998
rect 16396 16934 16448 16940
rect 16212 15496 16264 15502
rect 16212 15438 16264 15444
rect 16118 14376 16174 14385
rect 16118 14311 16174 14320
rect 16132 12782 16160 14311
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 16028 11892 16080 11898
rect 16028 11834 16080 11840
rect 16118 8664 16174 8673
rect 16118 8599 16174 8608
rect 16026 7304 16082 7313
rect 16026 7239 16082 7248
rect 15934 6488 15990 6497
rect 15934 6423 15990 6432
rect 15844 5296 15896 5302
rect 15844 5238 15896 5244
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 15476 4820 15528 4826
rect 15476 4762 15528 4768
rect 15488 3602 15516 4762
rect 15568 3936 15620 3942
rect 15568 3878 15620 3884
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15488 2990 15516 3538
rect 15580 3369 15608 3878
rect 15566 3360 15622 3369
rect 15566 3295 15622 3304
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 15672 2854 15700 5170
rect 15660 2848 15712 2854
rect 15660 2790 15712 2796
rect 15384 2440 15436 2446
rect 15384 2382 15436 2388
rect 16040 1970 16068 7239
rect 16132 4146 16160 8599
rect 16224 7993 16252 15438
rect 16408 8906 16436 16934
rect 16500 16794 16528 17546
rect 16580 17128 16632 17134
rect 16580 17070 16632 17076
rect 16488 16788 16540 16794
rect 16488 16730 16540 16736
rect 16592 16674 16620 17070
rect 16500 16646 16620 16674
rect 16396 8900 16448 8906
rect 16396 8842 16448 8848
rect 16210 7984 16266 7993
rect 16210 7919 16266 7928
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 16408 4078 16436 8842
rect 16500 5817 16528 16646
rect 16580 16516 16632 16522
rect 16580 16458 16632 16464
rect 16592 6322 16620 16458
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 16580 6316 16632 6322
rect 16580 6258 16632 6264
rect 16486 5808 16542 5817
rect 16486 5743 16542 5752
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16684 3097 16712 15302
rect 16868 14482 16896 19200
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16776 7478 16804 14350
rect 16854 12744 16910 12753
rect 16854 12679 16910 12688
rect 16764 7472 16816 7478
rect 16764 7414 16816 7420
rect 16868 3641 16896 12679
rect 16854 3632 16910 3641
rect 16854 3567 16910 3576
rect 16670 3088 16726 3097
rect 16670 3023 16726 3032
rect 16028 1964 16080 1970
rect 16028 1906 16080 1912
rect 1766 0 1822 800
rect 2042 0 2098 800
rect 2318 0 2374 800
rect 2594 0 2650 800
rect 2870 0 2926 800
rect 3146 0 3202 800
rect 3422 0 3478 800
rect 3698 0 3754 800
rect 3974 0 4030 800
rect 4250 0 4306 800
rect 4526 0 4582 800
rect 4802 0 4858 800
rect 5078 0 5134 800
rect 5354 0 5410 800
rect 5630 0 5686 800
rect 5906 0 5962 800
rect 6182 0 6238 800
rect 6458 0 6514 800
rect 6734 0 6790 800
rect 7010 0 7066 800
rect 7286 0 7342 800
rect 7562 0 7618 800
rect 7838 0 7894 800
rect 8114 0 8170 800
rect 8390 0 8446 800
rect 8666 0 8722 800
rect 8942 0 8998 800
rect 9218 0 9274 800
rect 9494 0 9550 800
rect 9770 0 9826 800
rect 10046 0 10102 800
rect 10322 0 10378 800
rect 10598 0 10654 800
rect 10874 0 10930 800
rect 11150 0 11206 800
rect 11426 0 11482 800
rect 11702 0 11758 800
rect 11978 0 12034 800
rect 12254 0 12310 800
rect 12530 0 12586 800
rect 12806 0 12862 800
rect 13082 0 13138 800
rect 13358 0 13414 800
rect 13634 0 13690 800
rect 13910 0 13966 800
rect 14186 0 14242 800
rect 14462 0 14518 800
rect 14738 0 14794 800
rect 15014 0 15070 800
rect 15290 0 15346 800
<< via2 >>
rect 1490 18944 1546 19000
rect 1858 17992 1914 18048
rect 2042 17040 2098 17096
rect 2134 16496 2190 16552
rect 1490 16088 1546 16144
rect 1490 15136 1546 15192
rect 1490 14220 1492 14240
rect 1492 14220 1544 14240
rect 1544 14220 1546 14240
rect 1490 14184 1546 14220
rect 2226 15308 2228 15328
rect 2228 15308 2280 15328
rect 2280 15308 2282 15328
rect 2226 15272 2282 15308
rect 1950 14456 2006 14512
rect 1490 13232 1546 13288
rect 1766 13232 1822 13288
rect 1490 12280 1546 12336
rect 1490 11328 1546 11384
rect 1490 10376 1546 10432
rect 1490 9444 1546 9480
rect 1490 9424 1492 9444
rect 1492 9424 1544 9444
rect 1544 9424 1546 9444
rect 2410 15272 2466 15328
rect 2410 15020 2466 15056
rect 2410 15000 2412 15020
rect 2412 15000 2464 15020
rect 2464 15000 2466 15020
rect 2410 13932 2466 13968
rect 2410 13912 2412 13932
rect 2412 13912 2464 13932
rect 2464 13912 2466 13932
rect 2830 16890 2886 16892
rect 2910 16890 2966 16892
rect 2990 16890 3046 16892
rect 3070 16890 3126 16892
rect 2830 16838 2876 16890
rect 2876 16838 2886 16890
rect 2910 16838 2940 16890
rect 2940 16838 2952 16890
rect 2952 16838 2966 16890
rect 2990 16838 3004 16890
rect 3004 16838 3016 16890
rect 3016 16838 3046 16890
rect 3070 16838 3080 16890
rect 3080 16838 3126 16890
rect 2830 16836 2886 16838
rect 2910 16836 2966 16838
rect 2990 16836 3046 16838
rect 3070 16836 3126 16838
rect 3054 16088 3110 16144
rect 2830 15802 2886 15804
rect 2910 15802 2966 15804
rect 2990 15802 3046 15804
rect 3070 15802 3126 15804
rect 2830 15750 2876 15802
rect 2876 15750 2886 15802
rect 2910 15750 2940 15802
rect 2940 15750 2952 15802
rect 2952 15750 2966 15802
rect 2990 15750 3004 15802
rect 3004 15750 3016 15802
rect 3016 15750 3046 15802
rect 3070 15750 3080 15802
rect 3080 15750 3126 15802
rect 2830 15748 2886 15750
rect 2910 15748 2966 15750
rect 2990 15748 3046 15750
rect 3070 15748 3126 15750
rect 2686 15544 2742 15600
rect 2830 14714 2886 14716
rect 2910 14714 2966 14716
rect 2990 14714 3046 14716
rect 3070 14714 3126 14716
rect 2830 14662 2876 14714
rect 2876 14662 2886 14714
rect 2910 14662 2940 14714
rect 2940 14662 2952 14714
rect 2952 14662 2966 14714
rect 2990 14662 3004 14714
rect 3004 14662 3016 14714
rect 3016 14662 3046 14714
rect 3070 14662 3080 14714
rect 3080 14662 3126 14714
rect 2830 14660 2886 14662
rect 2910 14660 2966 14662
rect 2990 14660 3046 14662
rect 3070 14660 3126 14662
rect 2870 14184 2926 14240
rect 1490 8472 1546 8528
rect 1490 7540 1546 7576
rect 1490 7520 1492 7540
rect 1492 7520 1544 7540
rect 1544 7520 1546 7540
rect 1490 6604 1492 6624
rect 1492 6604 1544 6624
rect 1544 6604 1546 6624
rect 1490 6568 1546 6604
rect 1490 5616 1546 5672
rect 1858 8880 1914 8936
rect 1950 8336 2006 8392
rect 2830 13626 2886 13628
rect 2910 13626 2966 13628
rect 2990 13626 3046 13628
rect 3070 13626 3126 13628
rect 2830 13574 2876 13626
rect 2876 13574 2886 13626
rect 2910 13574 2940 13626
rect 2940 13574 2952 13626
rect 2952 13574 2966 13626
rect 2990 13574 3004 13626
rect 3004 13574 3016 13626
rect 3016 13574 3046 13626
rect 3070 13574 3080 13626
rect 3080 13574 3126 13626
rect 2830 13572 2886 13574
rect 2910 13572 2966 13574
rect 2990 13572 3046 13574
rect 3070 13572 3126 13574
rect 2830 12538 2886 12540
rect 2910 12538 2966 12540
rect 2990 12538 3046 12540
rect 3070 12538 3126 12540
rect 2830 12486 2876 12538
rect 2876 12486 2886 12538
rect 2910 12486 2940 12538
rect 2940 12486 2952 12538
rect 2952 12486 2966 12538
rect 2990 12486 3004 12538
rect 3004 12486 3016 12538
rect 3016 12486 3046 12538
rect 3070 12486 3080 12538
rect 3080 12486 3126 12538
rect 2830 12484 2886 12486
rect 2910 12484 2966 12486
rect 2990 12484 3046 12486
rect 3070 12484 3126 12486
rect 2830 11450 2886 11452
rect 2910 11450 2966 11452
rect 2990 11450 3046 11452
rect 3070 11450 3126 11452
rect 2830 11398 2876 11450
rect 2876 11398 2886 11450
rect 2910 11398 2940 11450
rect 2940 11398 2952 11450
rect 2952 11398 2966 11450
rect 2990 11398 3004 11450
rect 3004 11398 3016 11450
rect 3016 11398 3046 11450
rect 3070 11398 3080 11450
rect 3080 11398 3126 11450
rect 2830 11396 2886 11398
rect 2910 11396 2966 11398
rect 2990 11396 3046 11398
rect 3070 11396 3126 11398
rect 3238 10512 3294 10568
rect 2830 10362 2886 10364
rect 2910 10362 2966 10364
rect 2990 10362 3046 10364
rect 3070 10362 3126 10364
rect 2830 10310 2876 10362
rect 2876 10310 2886 10362
rect 2910 10310 2940 10362
rect 2940 10310 2952 10362
rect 2952 10310 2966 10362
rect 2990 10310 3004 10362
rect 3004 10310 3016 10362
rect 3016 10310 3046 10362
rect 3070 10310 3080 10362
rect 3080 10310 3126 10362
rect 2830 10308 2886 10310
rect 2910 10308 2966 10310
rect 2990 10308 3046 10310
rect 3070 10308 3126 10310
rect 2830 9274 2886 9276
rect 2910 9274 2966 9276
rect 2990 9274 3046 9276
rect 3070 9274 3126 9276
rect 2830 9222 2876 9274
rect 2876 9222 2886 9274
rect 2910 9222 2940 9274
rect 2940 9222 2952 9274
rect 2952 9222 2966 9274
rect 2990 9222 3004 9274
rect 3004 9222 3016 9274
rect 3016 9222 3046 9274
rect 3070 9222 3080 9274
rect 3080 9222 3126 9274
rect 2830 9220 2886 9222
rect 2910 9220 2966 9222
rect 2990 9220 3046 9222
rect 3070 9220 3126 9222
rect 2226 6724 2282 6760
rect 2226 6704 2228 6724
rect 2228 6704 2280 6724
rect 2280 6704 2282 6724
rect 2830 8186 2886 8188
rect 2910 8186 2966 8188
rect 2990 8186 3046 8188
rect 3070 8186 3126 8188
rect 2830 8134 2876 8186
rect 2876 8134 2886 8186
rect 2910 8134 2940 8186
rect 2940 8134 2952 8186
rect 2952 8134 2966 8186
rect 2990 8134 3004 8186
rect 3004 8134 3016 8186
rect 3016 8134 3046 8186
rect 3070 8134 3080 8186
rect 3080 8134 3126 8186
rect 2830 8132 2886 8134
rect 2910 8132 2966 8134
rect 2990 8132 3046 8134
rect 3070 8132 3126 8134
rect 2226 5752 2282 5808
rect 1490 4664 1546 4720
rect 1766 4020 1768 4040
rect 1768 4020 1820 4040
rect 1820 4020 1822 4040
rect 1766 3984 1822 4020
rect 1490 3732 1546 3768
rect 1490 3712 1492 3732
rect 1492 3712 1544 3732
rect 1544 3712 1546 3732
rect 2226 5072 2282 5128
rect 2830 7098 2886 7100
rect 2910 7098 2966 7100
rect 2990 7098 3046 7100
rect 3070 7098 3126 7100
rect 2830 7046 2876 7098
rect 2876 7046 2886 7098
rect 2910 7046 2940 7098
rect 2940 7046 2952 7098
rect 2952 7046 2966 7098
rect 2990 7046 3004 7098
rect 3004 7046 3016 7098
rect 3016 7046 3046 7098
rect 3070 7046 3080 7098
rect 3080 7046 3126 7098
rect 2830 7044 2886 7046
rect 2910 7044 2966 7046
rect 2990 7044 3046 7046
rect 3070 7044 3126 7046
rect 2410 4820 2466 4856
rect 2410 4800 2412 4820
rect 2412 4800 2464 4820
rect 2464 4800 2466 4820
rect 2318 4664 2374 4720
rect 1950 3440 2006 3496
rect 1490 2796 1492 2816
rect 1492 2796 1544 2816
rect 1544 2796 1546 2816
rect 1490 2760 1546 2796
rect 1398 856 1454 912
rect 1858 1808 1914 1864
rect 2318 2896 2374 2952
rect 2830 6010 2886 6012
rect 2910 6010 2966 6012
rect 2990 6010 3046 6012
rect 3070 6010 3126 6012
rect 2830 5958 2876 6010
rect 2876 5958 2886 6010
rect 2910 5958 2940 6010
rect 2940 5958 2952 6010
rect 2952 5958 2966 6010
rect 2990 5958 3004 6010
rect 3004 5958 3016 6010
rect 3016 5958 3046 6010
rect 3070 5958 3080 6010
rect 3080 5958 3126 6010
rect 2830 5956 2886 5958
rect 2910 5956 2966 5958
rect 2990 5956 3046 5958
rect 3070 5956 3126 5958
rect 2830 4922 2886 4924
rect 2910 4922 2966 4924
rect 2990 4922 3046 4924
rect 3070 4922 3126 4924
rect 2830 4870 2876 4922
rect 2876 4870 2886 4922
rect 2910 4870 2940 4922
rect 2940 4870 2952 4922
rect 2952 4870 2966 4922
rect 2990 4870 3004 4922
rect 3004 4870 3016 4922
rect 3016 4870 3046 4922
rect 3070 4870 3080 4922
rect 3080 4870 3126 4922
rect 2830 4868 2886 4870
rect 2910 4868 2966 4870
rect 2990 4868 3046 4870
rect 3070 4868 3126 4870
rect 2870 4140 2926 4176
rect 2870 4120 2872 4140
rect 2872 4120 2924 4140
rect 2924 4120 2926 4140
rect 2830 3834 2886 3836
rect 2910 3834 2966 3836
rect 2990 3834 3046 3836
rect 3070 3834 3126 3836
rect 2830 3782 2876 3834
rect 2876 3782 2886 3834
rect 2910 3782 2940 3834
rect 2940 3782 2952 3834
rect 2952 3782 2966 3834
rect 2990 3782 3004 3834
rect 3004 3782 3016 3834
rect 3016 3782 3046 3834
rect 3070 3782 3080 3834
rect 3080 3782 3126 3834
rect 2830 3780 2886 3782
rect 2910 3780 2966 3782
rect 2990 3780 3046 3782
rect 3070 3780 3126 3782
rect 2870 3576 2926 3632
rect 3882 15852 3884 15872
rect 3884 15852 3936 15872
rect 3936 15852 3938 15872
rect 3882 15816 3938 15852
rect 4704 17434 4760 17436
rect 4784 17434 4840 17436
rect 4864 17434 4920 17436
rect 4944 17434 5000 17436
rect 4704 17382 4750 17434
rect 4750 17382 4760 17434
rect 4784 17382 4814 17434
rect 4814 17382 4826 17434
rect 4826 17382 4840 17434
rect 4864 17382 4878 17434
rect 4878 17382 4890 17434
rect 4890 17382 4920 17434
rect 4944 17382 4954 17434
rect 4954 17382 5000 17434
rect 4704 17380 4760 17382
rect 4784 17380 4840 17382
rect 4864 17380 4920 17382
rect 4944 17380 5000 17382
rect 5630 17196 5686 17232
rect 5630 17176 5632 17196
rect 5632 17176 5684 17196
rect 5684 17176 5686 17196
rect 4066 14220 4068 14240
rect 4068 14220 4120 14240
rect 4120 14220 4122 14240
rect 4066 14184 4122 14220
rect 4704 16346 4760 16348
rect 4784 16346 4840 16348
rect 4864 16346 4920 16348
rect 4944 16346 5000 16348
rect 4704 16294 4750 16346
rect 4750 16294 4760 16346
rect 4784 16294 4814 16346
rect 4814 16294 4826 16346
rect 4826 16294 4840 16346
rect 4864 16294 4878 16346
rect 4878 16294 4890 16346
rect 4890 16294 4920 16346
rect 4944 16294 4954 16346
rect 4954 16294 5000 16346
rect 4704 16292 4760 16294
rect 4784 16292 4840 16294
rect 4864 16292 4920 16294
rect 4944 16292 5000 16294
rect 4250 12588 4252 12608
rect 4252 12588 4304 12608
rect 4304 12588 4306 12608
rect 4250 12552 4306 12588
rect 3698 5208 3754 5264
rect 3882 7248 3938 7304
rect 3882 6316 3938 6352
rect 3882 6296 3884 6316
rect 3884 6296 3936 6316
rect 3936 6296 3938 6316
rect 3330 4392 3386 4448
rect 3238 4256 3294 4312
rect 3698 4800 3754 4856
rect 3422 3984 3478 4040
rect 2830 2746 2886 2748
rect 2910 2746 2966 2748
rect 2990 2746 3046 2748
rect 3070 2746 3126 2748
rect 2830 2694 2876 2746
rect 2876 2694 2886 2746
rect 2910 2694 2940 2746
rect 2940 2694 2952 2746
rect 2952 2694 2966 2746
rect 2990 2694 3004 2746
rect 3004 2694 3016 2746
rect 3016 2694 3046 2746
rect 3070 2694 3080 2746
rect 3080 2694 3126 2746
rect 2830 2692 2886 2694
rect 2910 2692 2966 2694
rect 2990 2692 3046 2694
rect 3070 2692 3126 2694
rect 2410 1944 2466 2000
rect 3790 4528 3846 4584
rect 4158 11736 4214 11792
rect 4066 6432 4122 6488
rect 4704 15258 4760 15260
rect 4784 15258 4840 15260
rect 4864 15258 4920 15260
rect 4944 15258 5000 15260
rect 4704 15206 4750 15258
rect 4750 15206 4760 15258
rect 4784 15206 4814 15258
rect 4814 15206 4826 15258
rect 4826 15206 4840 15258
rect 4864 15206 4878 15258
rect 4878 15206 4890 15258
rect 4890 15206 4920 15258
rect 4944 15206 4954 15258
rect 4954 15206 5000 15258
rect 4704 15204 4760 15206
rect 4784 15204 4840 15206
rect 4864 15204 4920 15206
rect 4944 15204 5000 15206
rect 4704 14170 4760 14172
rect 4784 14170 4840 14172
rect 4864 14170 4920 14172
rect 4944 14170 5000 14172
rect 4704 14118 4750 14170
rect 4750 14118 4760 14170
rect 4784 14118 4814 14170
rect 4814 14118 4826 14170
rect 4826 14118 4840 14170
rect 4864 14118 4878 14170
rect 4878 14118 4890 14170
rect 4890 14118 4920 14170
rect 4944 14118 4954 14170
rect 4954 14118 5000 14170
rect 4704 14116 4760 14118
rect 4784 14116 4840 14118
rect 4864 14116 4920 14118
rect 4944 14116 5000 14118
rect 4434 9424 4490 9480
rect 4704 13082 4760 13084
rect 4784 13082 4840 13084
rect 4864 13082 4920 13084
rect 4944 13082 5000 13084
rect 4704 13030 4750 13082
rect 4750 13030 4760 13082
rect 4784 13030 4814 13082
rect 4814 13030 4826 13082
rect 4826 13030 4840 13082
rect 4864 13030 4878 13082
rect 4878 13030 4890 13082
rect 4890 13030 4920 13082
rect 4944 13030 4954 13082
rect 4954 13030 5000 13082
rect 4704 13028 4760 13030
rect 4784 13028 4840 13030
rect 4864 13028 4920 13030
rect 4944 13028 5000 13030
rect 5262 12688 5318 12744
rect 4704 11994 4760 11996
rect 4784 11994 4840 11996
rect 4864 11994 4920 11996
rect 4944 11994 5000 11996
rect 4704 11942 4750 11994
rect 4750 11942 4760 11994
rect 4784 11942 4814 11994
rect 4814 11942 4826 11994
rect 4826 11942 4840 11994
rect 4864 11942 4878 11994
rect 4878 11942 4890 11994
rect 4890 11942 4920 11994
rect 4944 11942 4954 11994
rect 4954 11942 5000 11994
rect 4704 11940 4760 11942
rect 4784 11940 4840 11942
rect 4864 11940 4920 11942
rect 4944 11940 5000 11942
rect 4342 5772 4398 5808
rect 4342 5752 4344 5772
rect 4344 5752 4396 5772
rect 4396 5752 4398 5772
rect 4710 11092 4712 11112
rect 4712 11092 4764 11112
rect 4764 11092 4766 11112
rect 4710 11056 4766 11092
rect 4704 10906 4760 10908
rect 4784 10906 4840 10908
rect 4864 10906 4920 10908
rect 4944 10906 5000 10908
rect 4704 10854 4750 10906
rect 4750 10854 4760 10906
rect 4784 10854 4814 10906
rect 4814 10854 4826 10906
rect 4826 10854 4840 10906
rect 4864 10854 4878 10906
rect 4878 10854 4890 10906
rect 4890 10854 4920 10906
rect 4944 10854 4954 10906
rect 4954 10854 5000 10906
rect 4704 10852 4760 10854
rect 4784 10852 4840 10854
rect 4864 10852 4920 10854
rect 4944 10852 5000 10854
rect 4704 9818 4760 9820
rect 4784 9818 4840 9820
rect 4864 9818 4920 9820
rect 4944 9818 5000 9820
rect 4704 9766 4750 9818
rect 4750 9766 4760 9818
rect 4784 9766 4814 9818
rect 4814 9766 4826 9818
rect 4826 9766 4840 9818
rect 4864 9766 4878 9818
rect 4878 9766 4890 9818
rect 4890 9766 4920 9818
rect 4944 9766 4954 9818
rect 4954 9766 5000 9818
rect 4704 9764 4760 9766
rect 4784 9764 4840 9766
rect 4864 9764 4920 9766
rect 4944 9764 5000 9766
rect 4704 8730 4760 8732
rect 4784 8730 4840 8732
rect 4864 8730 4920 8732
rect 4944 8730 5000 8732
rect 4704 8678 4750 8730
rect 4750 8678 4760 8730
rect 4784 8678 4814 8730
rect 4814 8678 4826 8730
rect 4826 8678 4840 8730
rect 4864 8678 4878 8730
rect 4878 8678 4890 8730
rect 4890 8678 4920 8730
rect 4944 8678 4954 8730
rect 4954 8678 5000 8730
rect 4704 8676 4760 8678
rect 4784 8676 4840 8678
rect 4864 8676 4920 8678
rect 4944 8676 5000 8678
rect 4704 7642 4760 7644
rect 4784 7642 4840 7644
rect 4864 7642 4920 7644
rect 4944 7642 5000 7644
rect 4704 7590 4750 7642
rect 4750 7590 4760 7642
rect 4784 7590 4814 7642
rect 4814 7590 4826 7642
rect 4826 7590 4840 7642
rect 4864 7590 4878 7642
rect 4878 7590 4890 7642
rect 4890 7590 4920 7642
rect 4944 7590 4954 7642
rect 4954 7590 5000 7642
rect 4704 7588 4760 7590
rect 4784 7588 4840 7590
rect 4864 7588 4920 7590
rect 4944 7588 5000 7590
rect 4704 6554 4760 6556
rect 4784 6554 4840 6556
rect 4864 6554 4920 6556
rect 4944 6554 5000 6556
rect 4704 6502 4750 6554
rect 4750 6502 4760 6554
rect 4784 6502 4814 6554
rect 4814 6502 4826 6554
rect 4826 6502 4840 6554
rect 4864 6502 4878 6554
rect 4878 6502 4890 6554
rect 4890 6502 4920 6554
rect 4944 6502 4954 6554
rect 4954 6502 5000 6554
rect 4704 6500 4760 6502
rect 4784 6500 4840 6502
rect 4864 6500 4920 6502
rect 4944 6500 5000 6502
rect 4066 4800 4122 4856
rect 4066 4256 4122 4312
rect 4158 4156 4160 4176
rect 4160 4156 4212 4176
rect 4212 4156 4214 4176
rect 4158 4120 4214 4156
rect 3606 1808 3662 1864
rect 4434 4800 4490 4856
rect 8452 17434 8508 17436
rect 8532 17434 8588 17436
rect 8612 17434 8668 17436
rect 8692 17434 8748 17436
rect 8452 17382 8498 17434
rect 8498 17382 8508 17434
rect 8532 17382 8562 17434
rect 8562 17382 8574 17434
rect 8574 17382 8588 17434
rect 8612 17382 8626 17434
rect 8626 17382 8638 17434
rect 8638 17382 8668 17434
rect 8692 17382 8702 17434
rect 8702 17382 8748 17434
rect 8452 17380 8508 17382
rect 8532 17380 8588 17382
rect 8612 17380 8668 17382
rect 8692 17380 8748 17382
rect 6578 16890 6634 16892
rect 6658 16890 6714 16892
rect 6738 16890 6794 16892
rect 6818 16890 6874 16892
rect 6578 16838 6624 16890
rect 6624 16838 6634 16890
rect 6658 16838 6688 16890
rect 6688 16838 6700 16890
rect 6700 16838 6714 16890
rect 6738 16838 6752 16890
rect 6752 16838 6764 16890
rect 6764 16838 6794 16890
rect 6818 16838 6828 16890
rect 6828 16838 6874 16890
rect 6578 16836 6634 16838
rect 6658 16836 6714 16838
rect 6738 16836 6794 16838
rect 6818 16836 6874 16838
rect 7286 16496 7342 16552
rect 5630 15952 5686 16008
rect 6366 15816 6422 15872
rect 5630 12416 5686 12472
rect 6578 15802 6634 15804
rect 6658 15802 6714 15804
rect 6738 15802 6794 15804
rect 6818 15802 6874 15804
rect 6578 15750 6624 15802
rect 6624 15750 6634 15802
rect 6658 15750 6688 15802
rect 6688 15750 6700 15802
rect 6700 15750 6714 15802
rect 6738 15750 6752 15802
rect 6752 15750 6764 15802
rect 6764 15750 6794 15802
rect 6818 15750 6828 15802
rect 6828 15750 6874 15802
rect 6578 15748 6634 15750
rect 6658 15748 6714 15750
rect 6738 15748 6794 15750
rect 6818 15748 6874 15750
rect 6826 15308 6828 15328
rect 6828 15308 6880 15328
rect 6880 15308 6882 15328
rect 6826 15272 6882 15308
rect 6578 14714 6634 14716
rect 6658 14714 6714 14716
rect 6738 14714 6794 14716
rect 6818 14714 6874 14716
rect 6578 14662 6624 14714
rect 6624 14662 6634 14714
rect 6658 14662 6688 14714
rect 6688 14662 6700 14714
rect 6700 14662 6714 14714
rect 6738 14662 6752 14714
rect 6752 14662 6764 14714
rect 6764 14662 6794 14714
rect 6818 14662 6828 14714
rect 6828 14662 6874 14714
rect 6578 14660 6634 14662
rect 6658 14660 6714 14662
rect 6738 14660 6794 14662
rect 6818 14660 6874 14662
rect 5170 7792 5226 7848
rect 5170 6452 5226 6488
rect 5170 6432 5172 6452
rect 5172 6432 5224 6452
rect 5224 6432 5226 6452
rect 4986 5616 5042 5672
rect 4704 5466 4760 5468
rect 4784 5466 4840 5468
rect 4864 5466 4920 5468
rect 4944 5466 5000 5468
rect 4704 5414 4750 5466
rect 4750 5414 4760 5466
rect 4784 5414 4814 5466
rect 4814 5414 4826 5466
rect 4826 5414 4840 5466
rect 4864 5414 4878 5466
rect 4878 5414 4890 5466
rect 4890 5414 4920 5466
rect 4944 5414 4954 5466
rect 4954 5414 5000 5466
rect 4704 5412 4760 5414
rect 4784 5412 4840 5414
rect 4864 5412 4920 5414
rect 4944 5412 5000 5414
rect 4894 4972 4896 4992
rect 4896 4972 4948 4992
rect 4948 4972 4950 4992
rect 4894 4936 4950 4972
rect 3974 3732 4030 3768
rect 3974 3712 3976 3732
rect 3976 3712 4028 3732
rect 4028 3712 4030 3732
rect 4986 4528 5042 4584
rect 4704 4378 4760 4380
rect 4784 4378 4840 4380
rect 4864 4378 4920 4380
rect 4944 4378 5000 4380
rect 4704 4326 4750 4378
rect 4750 4326 4760 4378
rect 4784 4326 4814 4378
rect 4814 4326 4826 4378
rect 4826 4326 4840 4378
rect 4864 4326 4878 4378
rect 4878 4326 4890 4378
rect 4890 4326 4920 4378
rect 4944 4326 4954 4378
rect 4954 4326 5000 4378
rect 4704 4324 4760 4326
rect 4784 4324 4840 4326
rect 4864 4324 4920 4326
rect 4944 4324 5000 4326
rect 4618 4120 4674 4176
rect 4704 3290 4760 3292
rect 4784 3290 4840 3292
rect 4864 3290 4920 3292
rect 4944 3290 5000 3292
rect 4704 3238 4750 3290
rect 4750 3238 4760 3290
rect 4784 3238 4814 3290
rect 4814 3238 4826 3290
rect 4826 3238 4840 3290
rect 4864 3238 4878 3290
rect 4878 3238 4890 3290
rect 4890 3238 4920 3290
rect 4944 3238 4954 3290
rect 4954 3238 5000 3290
rect 4704 3236 4760 3238
rect 4784 3236 4840 3238
rect 4864 3236 4920 3238
rect 4944 3236 5000 3238
rect 3882 1672 3938 1728
rect 4342 2760 4398 2816
rect 4894 2488 4950 2544
rect 4704 2202 4760 2204
rect 4784 2202 4840 2204
rect 4864 2202 4920 2204
rect 4944 2202 5000 2204
rect 4704 2150 4750 2202
rect 4750 2150 4760 2202
rect 4784 2150 4814 2202
rect 4814 2150 4826 2202
rect 4826 2150 4840 2202
rect 4864 2150 4878 2202
rect 4878 2150 4890 2202
rect 4890 2150 4920 2202
rect 4944 2150 4954 2202
rect 4954 2150 5000 2202
rect 4704 2148 4760 2150
rect 4784 2148 4840 2150
rect 4864 2148 4920 2150
rect 4944 2148 5000 2150
rect 5262 5516 5264 5536
rect 5264 5516 5316 5536
rect 5316 5516 5318 5536
rect 5262 5480 5318 5516
rect 5538 5616 5594 5672
rect 5446 5208 5502 5264
rect 5446 4256 5502 4312
rect 5446 3304 5502 3360
rect 5446 3168 5502 3224
rect 5906 5888 5962 5944
rect 5906 5344 5962 5400
rect 6366 12552 6422 12608
rect 6642 13776 6698 13832
rect 6578 13626 6634 13628
rect 6658 13626 6714 13628
rect 6738 13626 6794 13628
rect 6818 13626 6874 13628
rect 6578 13574 6624 13626
rect 6624 13574 6634 13626
rect 6658 13574 6688 13626
rect 6688 13574 6700 13626
rect 6700 13574 6714 13626
rect 6738 13574 6752 13626
rect 6752 13574 6764 13626
rect 6764 13574 6794 13626
rect 6818 13574 6828 13626
rect 6828 13574 6874 13626
rect 6578 13572 6634 13574
rect 6658 13572 6714 13574
rect 6738 13572 6794 13574
rect 6818 13572 6874 13574
rect 6578 12538 6634 12540
rect 6658 12538 6714 12540
rect 6738 12538 6794 12540
rect 6818 12538 6874 12540
rect 6578 12486 6624 12538
rect 6624 12486 6634 12538
rect 6658 12486 6688 12538
rect 6688 12486 6700 12538
rect 6700 12486 6714 12538
rect 6738 12486 6752 12538
rect 6752 12486 6764 12538
rect 6764 12486 6794 12538
rect 6818 12486 6828 12538
rect 6828 12486 6874 12538
rect 6578 12484 6634 12486
rect 6658 12484 6714 12486
rect 6738 12484 6794 12486
rect 6818 12484 6874 12486
rect 6578 11450 6634 11452
rect 6658 11450 6714 11452
rect 6738 11450 6794 11452
rect 6818 11450 6874 11452
rect 6578 11398 6624 11450
rect 6624 11398 6634 11450
rect 6658 11398 6688 11450
rect 6688 11398 6700 11450
rect 6700 11398 6714 11450
rect 6738 11398 6752 11450
rect 6752 11398 6764 11450
rect 6764 11398 6794 11450
rect 6818 11398 6828 11450
rect 6828 11398 6874 11450
rect 6578 11396 6634 11398
rect 6658 11396 6714 11398
rect 6738 11396 6794 11398
rect 6818 11396 6874 11398
rect 6578 10362 6634 10364
rect 6658 10362 6714 10364
rect 6738 10362 6794 10364
rect 6818 10362 6874 10364
rect 6578 10310 6624 10362
rect 6624 10310 6634 10362
rect 6658 10310 6688 10362
rect 6688 10310 6700 10362
rect 6700 10310 6714 10362
rect 6738 10310 6752 10362
rect 6752 10310 6764 10362
rect 6764 10310 6794 10362
rect 6818 10310 6828 10362
rect 6828 10310 6874 10362
rect 6578 10308 6634 10310
rect 6658 10308 6714 10310
rect 6738 10308 6794 10310
rect 6818 10308 6874 10310
rect 6578 9274 6634 9276
rect 6658 9274 6714 9276
rect 6738 9274 6794 9276
rect 6818 9274 6874 9276
rect 6578 9222 6624 9274
rect 6624 9222 6634 9274
rect 6658 9222 6688 9274
rect 6688 9222 6700 9274
rect 6700 9222 6714 9274
rect 6738 9222 6752 9274
rect 6752 9222 6764 9274
rect 6764 9222 6794 9274
rect 6818 9222 6828 9274
rect 6828 9222 6874 9274
rect 6578 9220 6634 9222
rect 6658 9220 6714 9222
rect 6738 9220 6794 9222
rect 6818 9220 6874 9222
rect 6734 8508 6736 8528
rect 6736 8508 6788 8528
rect 6788 8508 6790 8528
rect 6734 8472 6790 8508
rect 6578 8186 6634 8188
rect 6658 8186 6714 8188
rect 6738 8186 6794 8188
rect 6818 8186 6874 8188
rect 6578 8134 6624 8186
rect 6624 8134 6634 8186
rect 6658 8134 6688 8186
rect 6688 8134 6700 8186
rect 6700 8134 6714 8186
rect 6738 8134 6752 8186
rect 6752 8134 6764 8186
rect 6764 8134 6794 8186
rect 6818 8134 6828 8186
rect 6828 8134 6874 8186
rect 6578 8132 6634 8134
rect 6658 8132 6714 8134
rect 6738 8132 6794 8134
rect 6818 8132 6874 8134
rect 6366 6840 6422 6896
rect 6578 7098 6634 7100
rect 6658 7098 6714 7100
rect 6738 7098 6794 7100
rect 6818 7098 6874 7100
rect 6578 7046 6624 7098
rect 6624 7046 6634 7098
rect 6658 7046 6688 7098
rect 6688 7046 6700 7098
rect 6700 7046 6714 7098
rect 6738 7046 6752 7098
rect 6752 7046 6764 7098
rect 6764 7046 6794 7098
rect 6818 7046 6828 7098
rect 6828 7046 6874 7098
rect 6578 7044 6634 7046
rect 6658 7044 6714 7046
rect 6738 7044 6794 7046
rect 6818 7044 6874 7046
rect 6642 6840 6698 6896
rect 7010 7928 7066 7984
rect 7654 14184 7710 14240
rect 7654 12824 7710 12880
rect 7562 12280 7618 12336
rect 6578 6010 6634 6012
rect 6658 6010 6714 6012
rect 6738 6010 6794 6012
rect 6818 6010 6874 6012
rect 6578 5958 6624 6010
rect 6624 5958 6634 6010
rect 6658 5958 6688 6010
rect 6688 5958 6700 6010
rect 6700 5958 6714 6010
rect 6738 5958 6752 6010
rect 6752 5958 6764 6010
rect 6764 5958 6794 6010
rect 6818 5958 6828 6010
rect 6828 5958 6874 6010
rect 6578 5956 6634 5958
rect 6658 5956 6714 5958
rect 6738 5956 6794 5958
rect 6818 5956 6874 5958
rect 6090 5208 6146 5264
rect 5814 3440 5870 3496
rect 6090 4936 6146 4992
rect 7102 6432 7158 6488
rect 6918 5480 6974 5536
rect 6578 4922 6634 4924
rect 6658 4922 6714 4924
rect 6738 4922 6794 4924
rect 6818 4922 6874 4924
rect 6578 4870 6624 4922
rect 6624 4870 6634 4922
rect 6658 4870 6688 4922
rect 6688 4870 6700 4922
rect 6700 4870 6714 4922
rect 6738 4870 6752 4922
rect 6752 4870 6764 4922
rect 6764 4870 6794 4922
rect 6818 4870 6828 4922
rect 6828 4870 6874 4922
rect 6578 4868 6634 4870
rect 6658 4868 6714 4870
rect 6738 4868 6794 4870
rect 6818 4868 6874 4870
rect 6458 4392 6514 4448
rect 5814 2624 5870 2680
rect 5538 2488 5594 2544
rect 6642 4120 6698 4176
rect 6550 3984 6606 4040
rect 6274 3884 6276 3904
rect 6276 3884 6328 3904
rect 6328 3884 6330 3904
rect 6274 3848 6330 3884
rect 6366 3732 6422 3768
rect 6366 3712 6368 3732
rect 6368 3712 6420 3732
rect 6420 3712 6422 3732
rect 6274 3576 6330 3632
rect 6578 3834 6634 3836
rect 6658 3834 6714 3836
rect 6738 3834 6794 3836
rect 6818 3834 6874 3836
rect 6578 3782 6624 3834
rect 6624 3782 6634 3834
rect 6658 3782 6688 3834
rect 6688 3782 6700 3834
rect 6700 3782 6714 3834
rect 6738 3782 6752 3834
rect 6752 3782 6764 3834
rect 6764 3782 6794 3834
rect 6818 3782 6828 3834
rect 6828 3782 6874 3834
rect 6578 3780 6634 3782
rect 6658 3780 6714 3782
rect 6738 3780 6794 3782
rect 6818 3780 6874 3782
rect 6642 3576 6698 3632
rect 5354 1536 5410 1592
rect 6182 3032 6238 3088
rect 6090 1808 6146 1864
rect 6826 3596 6882 3632
rect 6826 3576 6828 3596
rect 6828 3576 6880 3596
rect 6880 3576 6882 3596
rect 6826 2916 6882 2952
rect 6826 2896 6828 2916
rect 6828 2896 6880 2916
rect 6880 2896 6882 2916
rect 6578 2746 6634 2748
rect 6658 2746 6714 2748
rect 6738 2746 6794 2748
rect 6818 2746 6874 2748
rect 6578 2694 6624 2746
rect 6624 2694 6634 2746
rect 6658 2694 6688 2746
rect 6688 2694 6700 2746
rect 6700 2694 6714 2746
rect 6738 2694 6752 2746
rect 6752 2694 6764 2746
rect 6764 2694 6794 2746
rect 6818 2694 6828 2746
rect 6828 2694 6874 2746
rect 6578 2692 6634 2694
rect 6658 2692 6714 2694
rect 6738 2692 6794 2694
rect 6818 2692 6874 2694
rect 7102 5888 7158 5944
rect 7746 11600 7802 11656
rect 7378 6840 7434 6896
rect 8390 16496 8446 16552
rect 8452 16346 8508 16348
rect 8532 16346 8588 16348
rect 8612 16346 8668 16348
rect 8692 16346 8748 16348
rect 8452 16294 8498 16346
rect 8498 16294 8508 16346
rect 8532 16294 8562 16346
rect 8562 16294 8574 16346
rect 8574 16294 8588 16346
rect 8612 16294 8626 16346
rect 8626 16294 8638 16346
rect 8638 16294 8668 16346
rect 8692 16294 8702 16346
rect 8702 16294 8748 16346
rect 8452 16292 8508 16294
rect 8532 16292 8588 16294
rect 8612 16292 8668 16294
rect 8692 16292 8748 16294
rect 8574 15952 8630 16008
rect 7470 6704 7526 6760
rect 7194 4936 7250 4992
rect 7286 4528 7342 4584
rect 7194 4256 7250 4312
rect 7102 3440 7158 3496
rect 7838 7112 7894 7168
rect 7746 6568 7802 6624
rect 7930 6976 7986 7032
rect 8452 15258 8508 15260
rect 8532 15258 8588 15260
rect 8612 15258 8668 15260
rect 8692 15258 8748 15260
rect 8452 15206 8498 15258
rect 8498 15206 8508 15258
rect 8532 15206 8562 15258
rect 8562 15206 8574 15258
rect 8574 15206 8588 15258
rect 8612 15206 8626 15258
rect 8626 15206 8638 15258
rect 8638 15206 8668 15258
rect 8692 15206 8702 15258
rect 8702 15206 8748 15258
rect 8452 15204 8508 15206
rect 8532 15204 8588 15206
rect 8612 15204 8668 15206
rect 8692 15204 8748 15206
rect 8452 14170 8508 14172
rect 8532 14170 8588 14172
rect 8612 14170 8668 14172
rect 8692 14170 8748 14172
rect 8452 14118 8498 14170
rect 8498 14118 8508 14170
rect 8532 14118 8562 14170
rect 8562 14118 8574 14170
rect 8574 14118 8588 14170
rect 8612 14118 8626 14170
rect 8626 14118 8638 14170
rect 8638 14118 8668 14170
rect 8692 14118 8702 14170
rect 8702 14118 8748 14170
rect 8452 14116 8508 14118
rect 8532 14116 8588 14118
rect 8612 14116 8668 14118
rect 8692 14116 8748 14118
rect 8452 13082 8508 13084
rect 8532 13082 8588 13084
rect 8612 13082 8668 13084
rect 8692 13082 8748 13084
rect 8452 13030 8498 13082
rect 8498 13030 8508 13082
rect 8532 13030 8562 13082
rect 8562 13030 8574 13082
rect 8574 13030 8588 13082
rect 8612 13030 8626 13082
rect 8626 13030 8638 13082
rect 8638 13030 8668 13082
rect 8692 13030 8702 13082
rect 8702 13030 8748 13082
rect 8452 13028 8508 13030
rect 8532 13028 8588 13030
rect 8612 13028 8668 13030
rect 8692 13028 8748 13030
rect 8452 11994 8508 11996
rect 8532 11994 8588 11996
rect 8612 11994 8668 11996
rect 8692 11994 8748 11996
rect 8452 11942 8498 11994
rect 8498 11942 8508 11994
rect 8532 11942 8562 11994
rect 8562 11942 8574 11994
rect 8574 11942 8588 11994
rect 8612 11942 8626 11994
rect 8626 11942 8638 11994
rect 8638 11942 8668 11994
rect 8692 11942 8702 11994
rect 8702 11942 8748 11994
rect 8452 11940 8508 11942
rect 8532 11940 8588 11942
rect 8612 11940 8668 11942
rect 8692 11940 8748 11942
rect 8452 10906 8508 10908
rect 8532 10906 8588 10908
rect 8612 10906 8668 10908
rect 8692 10906 8748 10908
rect 8452 10854 8498 10906
rect 8498 10854 8508 10906
rect 8532 10854 8562 10906
rect 8562 10854 8574 10906
rect 8574 10854 8588 10906
rect 8612 10854 8626 10906
rect 8626 10854 8638 10906
rect 8638 10854 8668 10906
rect 8692 10854 8702 10906
rect 8702 10854 8748 10906
rect 8452 10852 8508 10854
rect 8532 10852 8588 10854
rect 8612 10852 8668 10854
rect 8692 10852 8748 10854
rect 7562 4256 7618 4312
rect 7470 4140 7526 4176
rect 7470 4120 7472 4140
rect 7472 4120 7524 4140
rect 7524 4120 7526 4140
rect 7470 3984 7526 4040
rect 7378 3712 7434 3768
rect 7286 3460 7342 3496
rect 7286 3440 7288 3460
rect 7288 3440 7340 3460
rect 7340 3440 7342 3460
rect 7654 3712 7710 3768
rect 8452 9818 8508 9820
rect 8532 9818 8588 9820
rect 8612 9818 8668 9820
rect 8692 9818 8748 9820
rect 8452 9766 8498 9818
rect 8498 9766 8508 9818
rect 8532 9766 8562 9818
rect 8562 9766 8574 9818
rect 8574 9766 8588 9818
rect 8612 9766 8626 9818
rect 8626 9766 8638 9818
rect 8638 9766 8668 9818
rect 8692 9766 8702 9818
rect 8702 9766 8748 9818
rect 8452 9764 8508 9766
rect 8532 9764 8588 9766
rect 8612 9764 8668 9766
rect 8692 9764 8748 9766
rect 8298 9152 8354 9208
rect 8298 8744 8354 8800
rect 8452 8730 8508 8732
rect 8532 8730 8588 8732
rect 8612 8730 8668 8732
rect 8692 8730 8748 8732
rect 8452 8678 8498 8730
rect 8498 8678 8508 8730
rect 8532 8678 8562 8730
rect 8562 8678 8574 8730
rect 8574 8678 8588 8730
rect 8612 8678 8626 8730
rect 8626 8678 8638 8730
rect 8638 8678 8668 8730
rect 8692 8678 8702 8730
rect 8702 8678 8748 8730
rect 8452 8676 8508 8678
rect 8532 8676 8588 8678
rect 8612 8676 8668 8678
rect 8692 8676 8748 8678
rect 8850 8608 8906 8664
rect 8452 7642 8508 7644
rect 8532 7642 8588 7644
rect 8612 7642 8668 7644
rect 8692 7642 8748 7644
rect 8452 7590 8498 7642
rect 8498 7590 8508 7642
rect 8532 7590 8562 7642
rect 8562 7590 8574 7642
rect 8574 7590 8588 7642
rect 8612 7590 8626 7642
rect 8626 7590 8638 7642
rect 8638 7590 8668 7642
rect 8692 7590 8702 7642
rect 8702 7590 8748 7642
rect 8452 7588 8508 7590
rect 8532 7588 8588 7590
rect 8612 7588 8668 7590
rect 8692 7588 8748 7590
rect 8850 7520 8906 7576
rect 8298 7112 8354 7168
rect 8390 6996 8446 7032
rect 8390 6976 8392 6996
rect 8392 6976 8444 6996
rect 8444 6976 8446 6996
rect 9310 13640 9366 13696
rect 9126 9016 9182 9072
rect 8942 6976 8998 7032
rect 9586 14864 9642 14920
rect 9494 13776 9550 13832
rect 9494 13640 9550 13696
rect 9494 9832 9550 9888
rect 10046 16360 10102 16416
rect 9770 15136 9826 15192
rect 9678 13368 9734 13424
rect 9678 12144 9734 12200
rect 9678 11056 9734 11112
rect 9954 13096 10010 13152
rect 9862 12416 9918 12472
rect 10326 16890 10382 16892
rect 10406 16890 10462 16892
rect 10486 16890 10542 16892
rect 10566 16890 10622 16892
rect 10326 16838 10372 16890
rect 10372 16838 10382 16890
rect 10406 16838 10436 16890
rect 10436 16838 10448 16890
rect 10448 16838 10462 16890
rect 10486 16838 10500 16890
rect 10500 16838 10512 16890
rect 10512 16838 10542 16890
rect 10566 16838 10576 16890
rect 10576 16838 10622 16890
rect 10326 16836 10382 16838
rect 10406 16836 10462 16838
rect 10486 16836 10542 16838
rect 10566 16836 10622 16838
rect 10506 16668 10508 16688
rect 10508 16668 10560 16688
rect 10560 16668 10562 16688
rect 10506 16632 10562 16668
rect 10782 16496 10838 16552
rect 12200 17434 12256 17436
rect 12280 17434 12336 17436
rect 12360 17434 12416 17436
rect 12440 17434 12496 17436
rect 12200 17382 12246 17434
rect 12246 17382 12256 17434
rect 12280 17382 12310 17434
rect 12310 17382 12322 17434
rect 12322 17382 12336 17434
rect 12360 17382 12374 17434
rect 12374 17382 12386 17434
rect 12386 17382 12416 17434
rect 12440 17382 12450 17434
rect 12450 17382 12496 17434
rect 12200 17380 12256 17382
rect 12280 17380 12336 17382
rect 12360 17380 12416 17382
rect 12440 17380 12496 17382
rect 12438 16496 12494 16552
rect 10326 15802 10382 15804
rect 10406 15802 10462 15804
rect 10486 15802 10542 15804
rect 10566 15802 10622 15804
rect 10326 15750 10372 15802
rect 10372 15750 10382 15802
rect 10406 15750 10436 15802
rect 10436 15750 10448 15802
rect 10448 15750 10462 15802
rect 10486 15750 10500 15802
rect 10500 15750 10512 15802
rect 10512 15750 10542 15802
rect 10566 15750 10576 15802
rect 10576 15750 10622 15802
rect 10326 15748 10382 15750
rect 10406 15748 10462 15750
rect 10486 15748 10542 15750
rect 10566 15748 10622 15750
rect 10230 15000 10286 15056
rect 10326 14714 10382 14716
rect 10406 14714 10462 14716
rect 10486 14714 10542 14716
rect 10566 14714 10622 14716
rect 10326 14662 10372 14714
rect 10372 14662 10382 14714
rect 10406 14662 10436 14714
rect 10436 14662 10448 14714
rect 10448 14662 10462 14714
rect 10486 14662 10500 14714
rect 10500 14662 10512 14714
rect 10512 14662 10542 14714
rect 10566 14662 10576 14714
rect 10576 14662 10622 14714
rect 10326 14660 10382 14662
rect 10406 14660 10462 14662
rect 10486 14660 10542 14662
rect 10566 14660 10622 14662
rect 11886 16360 11942 16416
rect 12200 16346 12256 16348
rect 12280 16346 12336 16348
rect 12360 16346 12416 16348
rect 12440 16346 12496 16348
rect 12200 16294 12246 16346
rect 12246 16294 12256 16346
rect 12280 16294 12310 16346
rect 12310 16294 12322 16346
rect 12322 16294 12336 16346
rect 12360 16294 12374 16346
rect 12374 16294 12386 16346
rect 12386 16294 12416 16346
rect 12440 16294 12450 16346
rect 12450 16294 12496 16346
rect 12200 16292 12256 16294
rect 12280 16292 12336 16294
rect 12360 16292 12416 16294
rect 12440 16292 12496 16294
rect 11978 15988 11980 16008
rect 11980 15988 12032 16008
rect 12032 15988 12034 16008
rect 11978 15952 12034 15988
rect 10874 14592 10930 14648
rect 10782 14184 10838 14240
rect 10138 13640 10194 13696
rect 9402 6976 9458 7032
rect 9770 8744 9826 8800
rect 9586 8472 9642 8528
rect 9770 8064 9826 8120
rect 9770 7656 9826 7712
rect 8452 6554 8508 6556
rect 8532 6554 8588 6556
rect 8612 6554 8668 6556
rect 8692 6554 8748 6556
rect 8452 6502 8498 6554
rect 8498 6502 8508 6554
rect 8532 6502 8562 6554
rect 8562 6502 8574 6554
rect 8574 6502 8588 6554
rect 8612 6502 8626 6554
rect 8626 6502 8638 6554
rect 8638 6502 8668 6554
rect 8692 6502 8702 6554
rect 8702 6502 8748 6554
rect 8452 6500 8508 6502
rect 8532 6500 8588 6502
rect 8612 6500 8668 6502
rect 8692 6500 8748 6502
rect 8390 6024 8446 6080
rect 8298 5752 8354 5808
rect 8942 6160 8998 6216
rect 8452 5466 8508 5468
rect 8532 5466 8588 5468
rect 8612 5466 8668 5468
rect 8692 5466 8748 5468
rect 8452 5414 8498 5466
rect 8498 5414 8508 5466
rect 8532 5414 8562 5466
rect 8562 5414 8574 5466
rect 8574 5414 8588 5466
rect 8612 5414 8626 5466
rect 8626 5414 8638 5466
rect 8638 5414 8668 5466
rect 8692 5414 8702 5466
rect 8702 5414 8748 5466
rect 8452 5412 8508 5414
rect 8532 5412 8588 5414
rect 8612 5412 8668 5414
rect 8692 5412 8748 5414
rect 8850 5480 8906 5536
rect 8206 5092 8262 5128
rect 8206 5072 8208 5092
rect 8208 5072 8260 5092
rect 8260 5072 8262 5092
rect 8482 5208 8538 5264
rect 8574 4936 8630 4992
rect 9126 6160 9182 6216
rect 9034 5072 9090 5128
rect 9310 5888 9366 5944
rect 9494 6568 9550 6624
rect 9954 8472 10010 8528
rect 9862 6976 9918 7032
rect 9402 5752 9458 5808
rect 9218 5072 9274 5128
rect 9402 5344 9458 5400
rect 10326 13626 10382 13628
rect 10406 13626 10462 13628
rect 10486 13626 10542 13628
rect 10566 13626 10622 13628
rect 10326 13574 10372 13626
rect 10372 13574 10382 13626
rect 10406 13574 10436 13626
rect 10436 13574 10448 13626
rect 10448 13574 10462 13626
rect 10486 13574 10500 13626
rect 10500 13574 10512 13626
rect 10512 13574 10542 13626
rect 10566 13574 10576 13626
rect 10576 13574 10622 13626
rect 10326 13572 10382 13574
rect 10406 13572 10462 13574
rect 10486 13572 10542 13574
rect 10566 13572 10622 13574
rect 10230 12688 10286 12744
rect 10966 14356 10968 14376
rect 10968 14356 11020 14376
rect 11020 14356 11022 14376
rect 10966 14320 11022 14356
rect 10966 14184 11022 14240
rect 10326 12538 10382 12540
rect 10406 12538 10462 12540
rect 10486 12538 10542 12540
rect 10566 12538 10622 12540
rect 10326 12486 10372 12538
rect 10372 12486 10382 12538
rect 10406 12486 10436 12538
rect 10436 12486 10448 12538
rect 10448 12486 10462 12538
rect 10486 12486 10500 12538
rect 10500 12486 10512 12538
rect 10512 12486 10542 12538
rect 10566 12486 10576 12538
rect 10576 12486 10622 12538
rect 10326 12484 10382 12486
rect 10406 12484 10462 12486
rect 10486 12484 10542 12486
rect 10566 12484 10622 12486
rect 10322 11892 10378 11928
rect 10322 11872 10324 11892
rect 10324 11872 10376 11892
rect 10376 11872 10378 11892
rect 10690 11872 10746 11928
rect 10326 11450 10382 11452
rect 10406 11450 10462 11452
rect 10486 11450 10542 11452
rect 10566 11450 10622 11452
rect 10326 11398 10372 11450
rect 10372 11398 10382 11450
rect 10406 11398 10436 11450
rect 10436 11398 10448 11450
rect 10448 11398 10462 11450
rect 10486 11398 10500 11450
rect 10500 11398 10512 11450
rect 10512 11398 10542 11450
rect 10566 11398 10576 11450
rect 10576 11398 10622 11450
rect 10326 11396 10382 11398
rect 10406 11396 10462 11398
rect 10486 11396 10542 11398
rect 10566 11396 10622 11398
rect 10874 11872 10930 11928
rect 10326 10362 10382 10364
rect 10406 10362 10462 10364
rect 10486 10362 10542 10364
rect 10566 10362 10622 10364
rect 10326 10310 10372 10362
rect 10372 10310 10382 10362
rect 10406 10310 10436 10362
rect 10436 10310 10448 10362
rect 10448 10310 10462 10362
rect 10486 10310 10500 10362
rect 10500 10310 10512 10362
rect 10512 10310 10542 10362
rect 10566 10310 10576 10362
rect 10576 10310 10622 10362
rect 10326 10308 10382 10310
rect 10406 10308 10462 10310
rect 10486 10308 10542 10310
rect 10566 10308 10622 10310
rect 10326 9274 10382 9276
rect 10406 9274 10462 9276
rect 10486 9274 10542 9276
rect 10566 9274 10622 9276
rect 10326 9222 10372 9274
rect 10372 9222 10382 9274
rect 10406 9222 10436 9274
rect 10436 9222 10448 9274
rect 10448 9222 10462 9274
rect 10486 9222 10500 9274
rect 10500 9222 10512 9274
rect 10512 9222 10542 9274
rect 10566 9222 10576 9274
rect 10576 9222 10622 9274
rect 10326 9220 10382 9222
rect 10406 9220 10462 9222
rect 10486 9220 10542 9222
rect 10566 9220 10622 9222
rect 10598 8608 10654 8664
rect 10326 8186 10382 8188
rect 10406 8186 10462 8188
rect 10486 8186 10542 8188
rect 10566 8186 10622 8188
rect 10326 8134 10372 8186
rect 10372 8134 10382 8186
rect 10406 8134 10436 8186
rect 10436 8134 10448 8186
rect 10448 8134 10462 8186
rect 10486 8134 10500 8186
rect 10500 8134 10512 8186
rect 10512 8134 10542 8186
rect 10566 8134 10576 8186
rect 10576 8134 10622 8186
rect 10326 8132 10382 8134
rect 10406 8132 10462 8134
rect 10486 8132 10542 8134
rect 10566 8132 10622 8134
rect 10138 7112 10194 7168
rect 10326 7098 10382 7100
rect 10406 7098 10462 7100
rect 10486 7098 10542 7100
rect 10566 7098 10622 7100
rect 10326 7046 10372 7098
rect 10372 7046 10382 7098
rect 10406 7046 10436 7098
rect 10436 7046 10448 7098
rect 10448 7046 10462 7098
rect 10486 7046 10500 7098
rect 10500 7046 10512 7098
rect 10512 7046 10542 7098
rect 10566 7046 10576 7098
rect 10576 7046 10622 7098
rect 10326 7044 10382 7046
rect 10406 7044 10462 7046
rect 10486 7044 10542 7046
rect 10566 7044 10622 7046
rect 10138 6704 10194 6760
rect 10046 6296 10102 6352
rect 10230 6296 10286 6352
rect 9586 5480 9642 5536
rect 9586 5344 9642 5400
rect 8758 4700 8760 4720
rect 8760 4700 8812 4720
rect 8812 4700 8814 4720
rect 8758 4664 8814 4700
rect 7838 3440 7894 3496
rect 7286 3052 7342 3088
rect 7286 3032 7288 3052
rect 7288 3032 7340 3052
rect 7340 3032 7342 3052
rect 8022 3848 8078 3904
rect 8206 3848 8262 3904
rect 6366 1944 6422 2000
rect 7010 2352 7066 2408
rect 7194 2644 7250 2680
rect 7194 2624 7196 2644
rect 7196 2624 7248 2644
rect 7248 2624 7250 2644
rect 7378 2624 7434 2680
rect 7470 2524 7472 2544
rect 7472 2524 7524 2544
rect 7524 2524 7526 2544
rect 7470 2488 7526 2524
rect 7470 2216 7526 2272
rect 8452 4378 8508 4380
rect 8532 4378 8588 4380
rect 8612 4378 8668 4380
rect 8692 4378 8748 4380
rect 8452 4326 8498 4378
rect 8498 4326 8508 4378
rect 8532 4326 8562 4378
rect 8562 4326 8574 4378
rect 8574 4326 8588 4378
rect 8612 4326 8626 4378
rect 8626 4326 8638 4378
rect 8638 4326 8668 4378
rect 8692 4326 8702 4378
rect 8702 4326 8748 4378
rect 8452 4324 8508 4326
rect 8532 4324 8588 4326
rect 8612 4324 8668 4326
rect 8692 4324 8748 4326
rect 8482 4120 8538 4176
rect 8666 4120 8722 4176
rect 8482 3440 8538 3496
rect 8114 3304 8170 3360
rect 8942 4256 8998 4312
rect 8452 3290 8508 3292
rect 8532 3290 8588 3292
rect 8612 3290 8668 3292
rect 8692 3290 8748 3292
rect 8452 3238 8498 3290
rect 8498 3238 8508 3290
rect 8532 3238 8562 3290
rect 8562 3238 8574 3290
rect 8574 3238 8588 3290
rect 8612 3238 8626 3290
rect 8626 3238 8638 3290
rect 8638 3238 8668 3290
rect 8692 3238 8702 3290
rect 8702 3238 8748 3290
rect 8452 3236 8508 3238
rect 8532 3236 8588 3238
rect 8612 3236 8668 3238
rect 8692 3236 8748 3238
rect 8114 3052 8170 3088
rect 8114 3032 8116 3052
rect 8116 3032 8168 3052
rect 8168 3032 8170 3052
rect 8298 2488 8354 2544
rect 7746 2080 7802 2136
rect 8114 2080 8170 2136
rect 9218 4664 9274 4720
rect 9586 5208 9642 5264
rect 9494 4800 9550 4856
rect 9402 4528 9458 4584
rect 9310 4256 9366 4312
rect 9126 3848 9182 3904
rect 9218 3576 9274 3632
rect 8850 2488 8906 2544
rect 8452 2202 8508 2204
rect 8532 2202 8588 2204
rect 8612 2202 8668 2204
rect 8692 2202 8748 2204
rect 8452 2150 8498 2202
rect 8498 2150 8508 2202
rect 8532 2150 8562 2202
rect 8562 2150 8574 2202
rect 8574 2150 8588 2202
rect 8612 2150 8626 2202
rect 8626 2150 8638 2202
rect 8638 2150 8668 2202
rect 8692 2150 8702 2202
rect 8702 2150 8748 2202
rect 8452 2148 8508 2150
rect 8532 2148 8588 2150
rect 8612 2148 8668 2150
rect 8692 2148 8748 2150
rect 9126 2216 9182 2272
rect 9770 5788 9772 5808
rect 9772 5788 9824 5808
rect 9824 5788 9826 5808
rect 9770 5752 9826 5788
rect 9770 5516 9772 5536
rect 9772 5516 9824 5536
rect 9824 5516 9826 5536
rect 9770 5480 9826 5516
rect 10046 5888 10102 5944
rect 10326 6010 10382 6012
rect 10406 6010 10462 6012
rect 10486 6010 10542 6012
rect 10566 6010 10622 6012
rect 10326 5958 10372 6010
rect 10372 5958 10382 6010
rect 10406 5958 10436 6010
rect 10436 5958 10448 6010
rect 10448 5958 10462 6010
rect 10486 5958 10500 6010
rect 10500 5958 10512 6010
rect 10512 5958 10542 6010
rect 10566 5958 10576 6010
rect 10576 5958 10622 6010
rect 10326 5956 10382 5958
rect 10406 5956 10462 5958
rect 10486 5956 10542 5958
rect 10566 5956 10622 5958
rect 9770 4820 9826 4856
rect 9770 4800 9772 4820
rect 9772 4800 9824 4820
rect 9824 4800 9826 4820
rect 9862 4684 9918 4720
rect 9862 4664 9864 4684
rect 9864 4664 9916 4684
rect 9916 4664 9918 4684
rect 9770 4256 9826 4312
rect 9402 2896 9458 2952
rect 10046 3712 10102 3768
rect 9862 1808 9918 1864
rect 10414 5344 10470 5400
rect 10598 5752 10654 5808
rect 10690 5616 10746 5672
rect 10690 5208 10746 5264
rect 10326 4922 10382 4924
rect 10406 4922 10462 4924
rect 10486 4922 10542 4924
rect 10566 4922 10622 4924
rect 10326 4870 10372 4922
rect 10372 4870 10382 4922
rect 10406 4870 10436 4922
rect 10436 4870 10448 4922
rect 10448 4870 10462 4922
rect 10486 4870 10500 4922
rect 10500 4870 10512 4922
rect 10512 4870 10542 4922
rect 10566 4870 10576 4922
rect 10576 4870 10622 4922
rect 10326 4868 10382 4870
rect 10406 4868 10462 4870
rect 10486 4868 10542 4870
rect 10566 4868 10622 4870
rect 11058 13232 11114 13288
rect 11702 14728 11758 14784
rect 11794 14456 11850 14512
rect 11426 13640 11482 13696
rect 11518 11892 11574 11928
rect 11518 11872 11520 11892
rect 11520 11872 11572 11892
rect 11572 11872 11574 11892
rect 11242 9988 11298 10024
rect 11242 9968 11244 9988
rect 11244 9968 11296 9988
rect 11296 9968 11298 9988
rect 11058 7792 11114 7848
rect 10598 4528 10654 4584
rect 10322 4256 10378 4312
rect 10326 3834 10382 3836
rect 10406 3834 10462 3836
rect 10486 3834 10542 3836
rect 10566 3834 10622 3836
rect 10326 3782 10372 3834
rect 10372 3782 10382 3834
rect 10406 3782 10436 3834
rect 10436 3782 10448 3834
rect 10448 3782 10462 3834
rect 10486 3782 10500 3834
rect 10500 3782 10512 3834
rect 10512 3782 10542 3834
rect 10566 3782 10576 3834
rect 10576 3782 10622 3834
rect 10326 3780 10382 3782
rect 10406 3780 10462 3782
rect 10486 3780 10542 3782
rect 10566 3780 10622 3782
rect 10414 3612 10416 3632
rect 10416 3612 10468 3632
rect 10468 3612 10470 3632
rect 10414 3576 10470 3612
rect 10506 3032 10562 3088
rect 10782 3848 10838 3904
rect 10782 3712 10838 3768
rect 10966 5888 11022 5944
rect 10966 5652 10968 5672
rect 10968 5652 11020 5672
rect 11020 5652 11022 5672
rect 10966 5616 11022 5652
rect 11702 11736 11758 11792
rect 12200 15258 12256 15260
rect 12280 15258 12336 15260
rect 12360 15258 12416 15260
rect 12440 15258 12496 15260
rect 12200 15206 12246 15258
rect 12246 15206 12256 15258
rect 12280 15206 12310 15258
rect 12310 15206 12322 15258
rect 12322 15206 12336 15258
rect 12360 15206 12374 15258
rect 12374 15206 12386 15258
rect 12386 15206 12416 15258
rect 12440 15206 12450 15258
rect 12450 15206 12496 15258
rect 12200 15204 12256 15206
rect 12280 15204 12336 15206
rect 12360 15204 12416 15206
rect 12440 15204 12496 15206
rect 12070 15000 12126 15056
rect 13082 16768 13138 16824
rect 12990 16632 13046 16688
rect 12254 14592 12310 14648
rect 12162 14492 12164 14512
rect 12164 14492 12216 14512
rect 12216 14492 12218 14512
rect 12162 14456 12218 14492
rect 12714 15000 12770 15056
rect 12346 14320 12402 14376
rect 12200 14170 12256 14172
rect 12280 14170 12336 14172
rect 12360 14170 12416 14172
rect 12440 14170 12496 14172
rect 12200 14118 12246 14170
rect 12246 14118 12256 14170
rect 12280 14118 12310 14170
rect 12310 14118 12322 14170
rect 12322 14118 12336 14170
rect 12360 14118 12374 14170
rect 12374 14118 12386 14170
rect 12386 14118 12416 14170
rect 12440 14118 12450 14170
rect 12450 14118 12496 14170
rect 12200 14116 12256 14118
rect 12280 14116 12336 14118
rect 12360 14116 12416 14118
rect 12440 14116 12496 14118
rect 12622 14492 12624 14512
rect 12624 14492 12676 14512
rect 12676 14492 12678 14512
rect 12622 14456 12678 14492
rect 12530 13912 12586 13968
rect 12714 13776 12770 13832
rect 12438 13640 12494 13696
rect 13082 16224 13138 16280
rect 13266 15952 13322 16008
rect 12200 13082 12256 13084
rect 12280 13082 12336 13084
rect 12360 13082 12416 13084
rect 12440 13082 12496 13084
rect 12200 13030 12246 13082
rect 12246 13030 12256 13082
rect 12280 13030 12310 13082
rect 12310 13030 12322 13082
rect 12322 13030 12336 13082
rect 12360 13030 12374 13082
rect 12374 13030 12386 13082
rect 12386 13030 12416 13082
rect 12440 13030 12450 13082
rect 12450 13030 12496 13082
rect 12200 13028 12256 13030
rect 12280 13028 12336 13030
rect 12360 13028 12416 13030
rect 12440 13028 12496 13030
rect 12346 12280 12402 12336
rect 12530 12280 12586 12336
rect 11334 7656 11390 7712
rect 11334 7248 11390 7304
rect 11334 6976 11390 7032
rect 11242 6568 11298 6624
rect 11518 6568 11574 6624
rect 11334 6160 11390 6216
rect 11058 4120 11114 4176
rect 11058 3848 11114 3904
rect 10966 3440 11022 3496
rect 10782 3032 10838 3088
rect 10326 2746 10382 2748
rect 10406 2746 10462 2748
rect 10486 2746 10542 2748
rect 10566 2746 10622 2748
rect 10326 2694 10372 2746
rect 10372 2694 10382 2746
rect 10406 2694 10436 2746
rect 10436 2694 10448 2746
rect 10448 2694 10462 2746
rect 10486 2694 10500 2746
rect 10500 2694 10512 2746
rect 10512 2694 10542 2746
rect 10566 2694 10576 2746
rect 10576 2694 10622 2746
rect 10326 2692 10382 2694
rect 10406 2692 10462 2694
rect 10486 2692 10542 2694
rect 10566 2692 10622 2694
rect 10782 2372 10838 2408
rect 10782 2352 10784 2372
rect 10784 2352 10836 2372
rect 10836 2352 10838 2372
rect 10690 1672 10746 1728
rect 11426 5344 11482 5400
rect 11518 4256 11574 4312
rect 11426 4120 11482 4176
rect 11334 3984 11390 4040
rect 11334 2796 11336 2816
rect 11336 2796 11388 2816
rect 11388 2796 11390 2816
rect 11334 2760 11390 2796
rect 11426 2624 11482 2680
rect 12200 11994 12256 11996
rect 12280 11994 12336 11996
rect 12360 11994 12416 11996
rect 12440 11994 12496 11996
rect 12200 11942 12246 11994
rect 12246 11942 12256 11994
rect 12280 11942 12310 11994
rect 12310 11942 12322 11994
rect 12322 11942 12336 11994
rect 12360 11942 12374 11994
rect 12374 11942 12386 11994
rect 12386 11942 12416 11994
rect 12440 11942 12450 11994
rect 12450 11942 12496 11994
rect 12200 11940 12256 11942
rect 12280 11940 12336 11942
rect 12360 11940 12416 11942
rect 12440 11940 12496 11942
rect 12200 10906 12256 10908
rect 12280 10906 12336 10908
rect 12360 10906 12416 10908
rect 12440 10906 12496 10908
rect 12200 10854 12246 10906
rect 12246 10854 12256 10906
rect 12280 10854 12310 10906
rect 12310 10854 12322 10906
rect 12322 10854 12336 10906
rect 12360 10854 12374 10906
rect 12374 10854 12386 10906
rect 12386 10854 12416 10906
rect 12440 10854 12450 10906
rect 12450 10854 12496 10906
rect 12200 10852 12256 10854
rect 12280 10852 12336 10854
rect 12360 10852 12416 10854
rect 12440 10852 12496 10854
rect 12070 10240 12126 10296
rect 11978 9424 12034 9480
rect 12200 9818 12256 9820
rect 12280 9818 12336 9820
rect 12360 9818 12416 9820
rect 12440 9818 12496 9820
rect 12200 9766 12246 9818
rect 12246 9766 12256 9818
rect 12280 9766 12310 9818
rect 12310 9766 12322 9818
rect 12322 9766 12336 9818
rect 12360 9766 12374 9818
rect 12374 9766 12386 9818
rect 12386 9766 12416 9818
rect 12440 9766 12450 9818
rect 12450 9766 12496 9818
rect 12200 9764 12256 9766
rect 12280 9764 12336 9766
rect 12360 9764 12416 9766
rect 12440 9764 12496 9766
rect 12070 9288 12126 9344
rect 13910 17040 13966 17096
rect 13266 13096 13322 13152
rect 13542 13640 13598 13696
rect 13542 13524 13598 13560
rect 13542 13504 13544 13524
rect 13544 13504 13596 13524
rect 13596 13504 13598 13524
rect 12806 9968 12862 10024
rect 12714 9832 12770 9888
rect 12990 10532 13046 10568
rect 12990 10512 12992 10532
rect 12992 10512 13044 10532
rect 13044 10512 13046 10532
rect 12806 9444 12862 9480
rect 12806 9424 12808 9444
rect 12808 9424 12860 9444
rect 12860 9424 12862 9444
rect 13358 12824 13414 12880
rect 13358 11736 13414 11792
rect 14074 16890 14130 16892
rect 14154 16890 14210 16892
rect 14234 16890 14290 16892
rect 14314 16890 14370 16892
rect 14074 16838 14120 16890
rect 14120 16838 14130 16890
rect 14154 16838 14184 16890
rect 14184 16838 14196 16890
rect 14196 16838 14210 16890
rect 14234 16838 14248 16890
rect 14248 16838 14260 16890
rect 14260 16838 14290 16890
rect 14314 16838 14324 16890
rect 14324 16838 14370 16890
rect 14074 16836 14130 16838
rect 14154 16836 14210 16838
rect 14234 16836 14290 16838
rect 14314 16836 14370 16838
rect 14002 15988 14004 16008
rect 14004 15988 14056 16008
rect 14056 15988 14058 16008
rect 14002 15952 14058 15988
rect 14074 15802 14130 15804
rect 14154 15802 14210 15804
rect 14234 15802 14290 15804
rect 14314 15802 14370 15804
rect 14074 15750 14120 15802
rect 14120 15750 14130 15802
rect 14154 15750 14184 15802
rect 14184 15750 14196 15802
rect 14196 15750 14210 15802
rect 14234 15750 14248 15802
rect 14248 15750 14260 15802
rect 14260 15750 14290 15802
rect 14314 15750 14324 15802
rect 14324 15750 14370 15802
rect 14074 15748 14130 15750
rect 14154 15748 14210 15750
rect 14234 15748 14290 15750
rect 14314 15748 14370 15750
rect 14462 15580 14464 15600
rect 14464 15580 14516 15600
rect 14516 15580 14518 15600
rect 14462 15544 14518 15580
rect 14074 14714 14130 14716
rect 14154 14714 14210 14716
rect 14234 14714 14290 14716
rect 14314 14714 14370 14716
rect 14074 14662 14120 14714
rect 14120 14662 14130 14714
rect 14154 14662 14184 14714
rect 14184 14662 14196 14714
rect 14196 14662 14210 14714
rect 14234 14662 14248 14714
rect 14248 14662 14260 14714
rect 14260 14662 14290 14714
rect 14314 14662 14324 14714
rect 14324 14662 14370 14714
rect 14074 14660 14130 14662
rect 14154 14660 14210 14662
rect 14234 14660 14290 14662
rect 14314 14660 14370 14662
rect 13818 13524 13874 13560
rect 13818 13504 13820 13524
rect 13820 13504 13872 13524
rect 13872 13504 13874 13524
rect 14074 13626 14130 13628
rect 14154 13626 14210 13628
rect 14234 13626 14290 13628
rect 14314 13626 14370 13628
rect 14074 13574 14120 13626
rect 14120 13574 14130 13626
rect 14154 13574 14184 13626
rect 14184 13574 14196 13626
rect 14196 13574 14210 13626
rect 14234 13574 14248 13626
rect 14248 13574 14260 13626
rect 14260 13574 14290 13626
rect 14314 13574 14324 13626
rect 14324 13574 14370 13626
rect 14074 13572 14130 13574
rect 14154 13572 14210 13574
rect 14234 13572 14290 13574
rect 14314 13572 14370 13574
rect 14646 15272 14702 15328
rect 14462 13368 14518 13424
rect 14278 13132 14280 13152
rect 14280 13132 14332 13152
rect 14332 13132 14334 13152
rect 14278 13096 14334 13132
rect 14074 12538 14130 12540
rect 14154 12538 14210 12540
rect 14234 12538 14290 12540
rect 14314 12538 14370 12540
rect 14074 12486 14120 12538
rect 14120 12486 14130 12538
rect 14154 12486 14184 12538
rect 14184 12486 14196 12538
rect 14196 12486 14210 12538
rect 14234 12486 14248 12538
rect 14248 12486 14260 12538
rect 14260 12486 14290 12538
rect 14314 12486 14324 12538
rect 14324 12486 14370 12538
rect 14074 12484 14130 12486
rect 14154 12484 14210 12486
rect 14234 12484 14290 12486
rect 14314 12484 14370 12486
rect 14646 13232 14702 13288
rect 15014 16088 15070 16144
rect 14074 11450 14130 11452
rect 14154 11450 14210 11452
rect 14234 11450 14290 11452
rect 14314 11450 14370 11452
rect 14074 11398 14120 11450
rect 14120 11398 14130 11450
rect 14154 11398 14184 11450
rect 14184 11398 14196 11450
rect 14196 11398 14210 11450
rect 14234 11398 14248 11450
rect 14248 11398 14260 11450
rect 14260 11398 14290 11450
rect 14314 11398 14324 11450
rect 14324 11398 14370 11450
rect 14074 11396 14130 11398
rect 14154 11396 14210 11398
rect 14234 11396 14290 11398
rect 14314 11396 14370 11398
rect 13266 10124 13322 10160
rect 13266 10104 13268 10124
rect 13268 10104 13320 10124
rect 13320 10104 13322 10124
rect 11978 8744 12034 8800
rect 12200 8730 12256 8732
rect 12280 8730 12336 8732
rect 12360 8730 12416 8732
rect 12440 8730 12496 8732
rect 12200 8678 12246 8730
rect 12246 8678 12256 8730
rect 12280 8678 12310 8730
rect 12310 8678 12322 8730
rect 12322 8678 12336 8730
rect 12360 8678 12374 8730
rect 12374 8678 12386 8730
rect 12386 8678 12416 8730
rect 12440 8678 12450 8730
rect 12450 8678 12496 8730
rect 12200 8676 12256 8678
rect 12280 8676 12336 8678
rect 12360 8676 12416 8678
rect 12440 8676 12496 8678
rect 11886 8492 11942 8528
rect 11886 8472 11888 8492
rect 11888 8472 11940 8492
rect 11940 8472 11942 8492
rect 12070 8472 12126 8528
rect 11794 6860 11850 6896
rect 11794 6840 11796 6860
rect 11796 6840 11848 6860
rect 11848 6840 11850 6860
rect 11886 6704 11942 6760
rect 12346 8356 12402 8392
rect 12346 8336 12348 8356
rect 12348 8336 12400 8356
rect 12400 8336 12402 8356
rect 12162 7948 12218 7984
rect 12162 7928 12164 7948
rect 12164 7928 12216 7948
rect 12216 7928 12218 7948
rect 12530 7792 12586 7848
rect 12200 7642 12256 7644
rect 12280 7642 12336 7644
rect 12360 7642 12416 7644
rect 12440 7642 12496 7644
rect 12200 7590 12246 7642
rect 12246 7590 12256 7642
rect 12280 7590 12310 7642
rect 12310 7590 12322 7642
rect 12322 7590 12336 7642
rect 12360 7590 12374 7642
rect 12374 7590 12386 7642
rect 12386 7590 12416 7642
rect 12440 7590 12450 7642
rect 12450 7590 12496 7642
rect 12200 7588 12256 7590
rect 12280 7588 12336 7590
rect 12360 7588 12416 7590
rect 12440 7588 12496 7590
rect 12346 7384 12402 7440
rect 12162 7248 12218 7304
rect 12162 7112 12218 7168
rect 12070 6976 12126 7032
rect 12200 6554 12256 6556
rect 12280 6554 12336 6556
rect 12360 6554 12416 6556
rect 12440 6554 12496 6556
rect 12200 6502 12246 6554
rect 12246 6502 12256 6554
rect 12280 6502 12310 6554
rect 12310 6502 12322 6554
rect 12322 6502 12336 6554
rect 12360 6502 12374 6554
rect 12374 6502 12386 6554
rect 12386 6502 12416 6554
rect 12440 6502 12450 6554
rect 12450 6502 12496 6554
rect 12200 6500 12256 6502
rect 12280 6500 12336 6502
rect 12360 6500 12416 6502
rect 12440 6500 12496 6502
rect 11886 6024 11942 6080
rect 11794 5616 11850 5672
rect 11978 5652 11980 5672
rect 11980 5652 12032 5672
rect 12032 5652 12034 5672
rect 11978 5616 12034 5652
rect 11978 4936 12034 4992
rect 12438 6160 12494 6216
rect 12898 7420 12900 7440
rect 12900 7420 12952 7440
rect 12952 7420 12954 7440
rect 12898 7384 12954 7420
rect 13450 9968 13506 10024
rect 13358 9832 13414 9888
rect 12714 6316 12770 6352
rect 12714 6296 12716 6316
rect 12716 6296 12768 6316
rect 12768 6296 12770 6316
rect 12622 6196 12624 6216
rect 12624 6196 12676 6216
rect 12676 6196 12678 6216
rect 12622 6160 12678 6196
rect 12898 5752 12954 5808
rect 12530 5616 12586 5672
rect 12200 5466 12256 5468
rect 12280 5466 12336 5468
rect 12360 5466 12416 5468
rect 12440 5466 12496 5468
rect 12200 5414 12246 5466
rect 12246 5414 12256 5466
rect 12280 5414 12310 5466
rect 12310 5414 12322 5466
rect 12322 5414 12336 5466
rect 12360 5414 12374 5466
rect 12374 5414 12386 5466
rect 12386 5414 12416 5466
rect 12440 5414 12450 5466
rect 12450 5414 12496 5466
rect 12200 5412 12256 5414
rect 12280 5412 12336 5414
rect 12360 5412 12416 5414
rect 12440 5412 12496 5414
rect 12162 4800 12218 4856
rect 11978 3984 12034 4040
rect 11794 3032 11850 3088
rect 11518 1400 11574 1456
rect 12346 5072 12402 5128
rect 12200 4378 12256 4380
rect 12280 4378 12336 4380
rect 12360 4378 12416 4380
rect 12440 4378 12496 4380
rect 12200 4326 12246 4378
rect 12246 4326 12256 4378
rect 12280 4326 12310 4378
rect 12310 4326 12322 4378
rect 12322 4326 12336 4378
rect 12360 4326 12374 4378
rect 12374 4326 12386 4378
rect 12386 4326 12416 4378
rect 12440 4326 12450 4378
rect 12450 4326 12496 4378
rect 12200 4324 12256 4326
rect 12280 4324 12336 4326
rect 12360 4324 12416 4326
rect 12440 4324 12496 4326
rect 12254 3984 12310 4040
rect 12162 3576 12218 3632
rect 12200 3290 12256 3292
rect 12280 3290 12336 3292
rect 12360 3290 12416 3292
rect 12440 3290 12496 3292
rect 12200 3238 12246 3290
rect 12246 3238 12256 3290
rect 12280 3238 12310 3290
rect 12310 3238 12322 3290
rect 12322 3238 12336 3290
rect 12360 3238 12374 3290
rect 12374 3238 12386 3290
rect 12386 3238 12416 3290
rect 12440 3238 12450 3290
rect 12450 3238 12496 3290
rect 12200 3236 12256 3238
rect 12280 3236 12336 3238
rect 12360 3236 12416 3238
rect 12440 3236 12496 3238
rect 12898 5228 12954 5264
rect 12898 5208 12900 5228
rect 12900 5208 12952 5228
rect 12952 5208 12954 5228
rect 12714 4256 12770 4312
rect 13174 6432 13230 6488
rect 12990 4936 13046 4992
rect 12990 4800 13046 4856
rect 14074 10362 14130 10364
rect 14154 10362 14210 10364
rect 14234 10362 14290 10364
rect 14314 10362 14370 10364
rect 14074 10310 14120 10362
rect 14120 10310 14130 10362
rect 14154 10310 14184 10362
rect 14184 10310 14196 10362
rect 14196 10310 14210 10362
rect 14234 10310 14248 10362
rect 14248 10310 14260 10362
rect 14260 10310 14290 10362
rect 14314 10310 14324 10362
rect 14324 10310 14370 10362
rect 14074 10308 14130 10310
rect 14154 10308 14210 10310
rect 14234 10308 14290 10310
rect 14314 10308 14370 10310
rect 13818 10240 13874 10296
rect 13542 9152 13598 9208
rect 13634 8880 13690 8936
rect 13450 7692 13452 7712
rect 13452 7692 13504 7712
rect 13504 7692 13506 7712
rect 13450 7656 13506 7692
rect 13634 6704 13690 6760
rect 13542 5752 13598 5808
rect 13450 5616 13506 5672
rect 13358 4936 13414 4992
rect 13358 4684 13414 4720
rect 13358 4664 13360 4684
rect 13360 4664 13412 4684
rect 13412 4664 13414 4684
rect 12898 4392 12954 4448
rect 13266 4392 13322 4448
rect 12254 3052 12310 3088
rect 12254 3032 12256 3052
rect 12256 3032 12308 3052
rect 12308 3032 12310 3052
rect 12200 2202 12256 2204
rect 12280 2202 12336 2204
rect 12360 2202 12416 2204
rect 12440 2202 12496 2204
rect 12200 2150 12246 2202
rect 12246 2150 12256 2202
rect 12280 2150 12310 2202
rect 12310 2150 12322 2202
rect 12322 2150 12336 2202
rect 12360 2150 12374 2202
rect 12374 2150 12386 2202
rect 12386 2150 12416 2202
rect 12440 2150 12450 2202
rect 12450 2150 12496 2202
rect 12200 2148 12256 2150
rect 12280 2148 12336 2150
rect 12360 2148 12416 2150
rect 12440 2148 12496 2150
rect 12806 3440 12862 3496
rect 12898 3168 12954 3224
rect 13358 3032 13414 3088
rect 13266 2488 13322 2544
rect 14646 11600 14702 11656
rect 15382 14864 15438 14920
rect 14462 9580 14518 9616
rect 14462 9560 14464 9580
rect 14464 9560 14516 9580
rect 14516 9560 14518 9580
rect 14002 9424 14058 9480
rect 14074 9274 14130 9276
rect 14154 9274 14210 9276
rect 14234 9274 14290 9276
rect 14314 9274 14370 9276
rect 14074 9222 14120 9274
rect 14120 9222 14130 9274
rect 14154 9222 14184 9274
rect 14184 9222 14196 9274
rect 14196 9222 14210 9274
rect 14234 9222 14248 9274
rect 14248 9222 14260 9274
rect 14260 9222 14290 9274
rect 14314 9222 14324 9274
rect 14324 9222 14370 9274
rect 14074 9220 14130 9222
rect 14154 9220 14210 9222
rect 14234 9220 14290 9222
rect 14314 9220 14370 9222
rect 14186 9016 14242 9072
rect 14370 9016 14426 9072
rect 14094 8780 14096 8800
rect 14096 8780 14148 8800
rect 14148 8780 14150 8800
rect 14094 8744 14150 8780
rect 14738 9968 14794 10024
rect 14554 9016 14610 9072
rect 14074 8186 14130 8188
rect 14154 8186 14210 8188
rect 14234 8186 14290 8188
rect 14314 8186 14370 8188
rect 14074 8134 14120 8186
rect 14120 8134 14130 8186
rect 14154 8134 14184 8186
rect 14184 8134 14196 8186
rect 14196 8134 14210 8186
rect 14234 8134 14248 8186
rect 14248 8134 14260 8186
rect 14260 8134 14290 8186
rect 14314 8134 14324 8186
rect 14324 8134 14370 8186
rect 14074 8132 14130 8134
rect 14154 8132 14210 8134
rect 14234 8132 14290 8134
rect 14314 8132 14370 8134
rect 13910 7948 13966 7984
rect 13910 7928 13912 7948
rect 13912 7928 13964 7948
rect 13964 7928 13966 7948
rect 13818 6740 13820 6760
rect 13820 6740 13872 6760
rect 13872 6740 13874 6760
rect 13818 6704 13874 6740
rect 13818 6296 13874 6352
rect 14646 7656 14702 7712
rect 14554 7520 14610 7576
rect 14370 7248 14426 7304
rect 14074 7098 14130 7100
rect 14154 7098 14210 7100
rect 14234 7098 14290 7100
rect 14314 7098 14370 7100
rect 14074 7046 14120 7098
rect 14120 7046 14130 7098
rect 14154 7046 14184 7098
rect 14184 7046 14196 7098
rect 14196 7046 14210 7098
rect 14234 7046 14248 7098
rect 14248 7046 14260 7098
rect 14260 7046 14290 7098
rect 14314 7046 14324 7098
rect 14324 7046 14370 7098
rect 14074 7044 14130 7046
rect 14154 7044 14210 7046
rect 14234 7044 14290 7046
rect 14314 7044 14370 7046
rect 13818 5888 13874 5944
rect 13634 3304 13690 3360
rect 13542 2624 13598 2680
rect 14094 6568 14150 6624
rect 14094 6452 14150 6488
rect 14094 6432 14096 6452
rect 14096 6432 14148 6452
rect 14148 6432 14150 6452
rect 14278 6160 14334 6216
rect 14074 6010 14130 6012
rect 14154 6010 14210 6012
rect 14234 6010 14290 6012
rect 14314 6010 14370 6012
rect 14074 5958 14120 6010
rect 14120 5958 14130 6010
rect 14154 5958 14184 6010
rect 14184 5958 14196 6010
rect 14196 5958 14210 6010
rect 14234 5958 14248 6010
rect 14248 5958 14260 6010
rect 14260 5958 14290 6010
rect 14314 5958 14324 6010
rect 14324 5958 14370 6010
rect 14074 5956 14130 5958
rect 14154 5956 14210 5958
rect 14234 5956 14290 5958
rect 14314 5956 14370 5958
rect 13910 5208 13966 5264
rect 14186 5752 14242 5808
rect 14094 5652 14096 5672
rect 14096 5652 14148 5672
rect 14148 5652 14150 5672
rect 14094 5616 14150 5652
rect 14094 5364 14150 5400
rect 14094 5344 14096 5364
rect 14096 5344 14148 5364
rect 14148 5344 14150 5364
rect 14370 5516 14372 5536
rect 14372 5516 14424 5536
rect 14424 5516 14426 5536
rect 14370 5480 14426 5516
rect 14074 4922 14130 4924
rect 14154 4922 14210 4924
rect 14234 4922 14290 4924
rect 14314 4922 14370 4924
rect 14074 4870 14120 4922
rect 14120 4870 14130 4922
rect 14154 4870 14184 4922
rect 14184 4870 14196 4922
rect 14196 4870 14210 4922
rect 14234 4870 14248 4922
rect 14248 4870 14260 4922
rect 14260 4870 14290 4922
rect 14314 4870 14324 4922
rect 14324 4870 14370 4922
rect 14074 4868 14130 4870
rect 14154 4868 14210 4870
rect 14234 4868 14290 4870
rect 14314 4868 14370 4870
rect 14002 3984 14058 4040
rect 14074 3834 14130 3836
rect 14154 3834 14210 3836
rect 14234 3834 14290 3836
rect 14314 3834 14370 3836
rect 14074 3782 14120 3834
rect 14120 3782 14130 3834
rect 14154 3782 14184 3834
rect 14184 3782 14196 3834
rect 14196 3782 14210 3834
rect 14234 3782 14248 3834
rect 14248 3782 14260 3834
rect 14260 3782 14290 3834
rect 14314 3782 14324 3834
rect 14324 3782 14370 3834
rect 14074 3780 14130 3782
rect 14154 3780 14210 3782
rect 14234 3780 14290 3782
rect 14314 3780 14370 3782
rect 14646 6704 14702 6760
rect 14646 6452 14702 6488
rect 14646 6432 14648 6452
rect 14648 6432 14700 6452
rect 14700 6432 14702 6452
rect 14646 6060 14648 6080
rect 14648 6060 14700 6080
rect 14700 6060 14702 6080
rect 14646 6024 14702 6060
rect 14646 4120 14702 4176
rect 14094 3576 14150 3632
rect 15106 9968 15162 10024
rect 15106 7656 15162 7712
rect 14922 5480 14978 5536
rect 14922 4256 14978 4312
rect 14462 3440 14518 3496
rect 14554 3304 14610 3360
rect 13910 2760 13966 2816
rect 13818 2216 13874 2272
rect 14074 2746 14130 2748
rect 14154 2746 14210 2748
rect 14234 2746 14290 2748
rect 14314 2746 14370 2748
rect 14074 2694 14120 2746
rect 14120 2694 14130 2746
rect 14154 2694 14184 2746
rect 14184 2694 14196 2746
rect 14196 2694 14210 2746
rect 14234 2694 14248 2746
rect 14248 2694 14260 2746
rect 14260 2694 14290 2746
rect 14314 2694 14324 2746
rect 14324 2694 14370 2746
rect 14074 2692 14130 2694
rect 14154 2692 14210 2694
rect 14234 2692 14290 2694
rect 14314 2692 14370 2694
rect 14370 2508 14426 2544
rect 14370 2488 14372 2508
rect 14372 2488 14424 2508
rect 14424 2488 14426 2508
rect 14646 1808 14702 1864
rect 15474 5364 15530 5400
rect 15474 5344 15476 5364
rect 15476 5344 15528 5364
rect 15528 5344 15530 5364
rect 16118 14320 16174 14376
rect 16118 8608 16174 8664
rect 16026 7248 16082 7304
rect 15934 6432 15990 6488
rect 15566 3304 15622 3360
rect 16210 7928 16266 7984
rect 16486 5752 16542 5808
rect 16854 12688 16910 12744
rect 16854 3576 16910 3632
rect 16670 3032 16726 3088
<< metal3 >>
rect 0 19002 800 19032
rect 1485 19002 1551 19005
rect 0 19000 1551 19002
rect 0 18944 1490 19000
rect 1546 18944 1551 19000
rect 0 18942 1551 18944
rect 0 18912 800 18942
rect 1485 18939 1551 18942
rect 0 18050 800 18080
rect 1853 18050 1919 18053
rect 0 18048 1919 18050
rect 0 17992 1858 18048
rect 1914 17992 1919 18048
rect 0 17990 1919 17992
rect 0 17960 800 17990
rect 1853 17987 1919 17990
rect 4694 17440 5010 17441
rect 4694 17376 4700 17440
rect 4764 17376 4780 17440
rect 4844 17376 4860 17440
rect 4924 17376 4940 17440
rect 5004 17376 5010 17440
rect 4694 17375 5010 17376
rect 8442 17440 8758 17441
rect 8442 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8758 17440
rect 8442 17375 8758 17376
rect 12190 17440 12506 17441
rect 12190 17376 12196 17440
rect 12260 17376 12276 17440
rect 12340 17376 12356 17440
rect 12420 17376 12436 17440
rect 12500 17376 12506 17440
rect 12190 17375 12506 17376
rect 5625 17234 5691 17237
rect 11462 17234 11468 17236
rect 5625 17232 11468 17234
rect 5625 17176 5630 17232
rect 5686 17176 11468 17232
rect 5625 17174 11468 17176
rect 5625 17171 5691 17174
rect 11462 17172 11468 17174
rect 11532 17172 11538 17236
rect 0 17008 800 17128
rect 2037 17098 2103 17101
rect 13905 17098 13971 17101
rect 2037 17096 13971 17098
rect 2037 17040 2042 17096
rect 2098 17040 13910 17096
rect 13966 17040 13971 17096
rect 2037 17038 13971 17040
rect 2037 17035 2103 17038
rect 13905 17035 13971 17038
rect 2820 16896 3136 16897
rect 2820 16832 2826 16896
rect 2890 16832 2906 16896
rect 2970 16832 2986 16896
rect 3050 16832 3066 16896
rect 3130 16832 3136 16896
rect 2820 16831 3136 16832
rect 6568 16896 6884 16897
rect 6568 16832 6574 16896
rect 6638 16832 6654 16896
rect 6718 16832 6734 16896
rect 6798 16832 6814 16896
rect 6878 16832 6884 16896
rect 6568 16831 6884 16832
rect 10316 16896 10632 16897
rect 10316 16832 10322 16896
rect 10386 16832 10402 16896
rect 10466 16832 10482 16896
rect 10546 16832 10562 16896
rect 10626 16832 10632 16896
rect 10316 16831 10632 16832
rect 14064 16896 14380 16897
rect 14064 16832 14070 16896
rect 14134 16832 14150 16896
rect 14214 16832 14230 16896
rect 14294 16832 14310 16896
rect 14374 16832 14380 16896
rect 14064 16831 14380 16832
rect 13077 16826 13143 16829
rect 13670 16826 13676 16828
rect 13077 16824 13676 16826
rect 13077 16768 13082 16824
rect 13138 16768 13676 16824
rect 13077 16766 13676 16768
rect 13077 16763 13143 16766
rect 13670 16764 13676 16766
rect 13740 16764 13746 16828
rect 9806 16628 9812 16692
rect 9876 16690 9882 16692
rect 10501 16690 10567 16693
rect 9876 16688 10567 16690
rect 9876 16632 10506 16688
rect 10562 16632 10567 16688
rect 9876 16630 10567 16632
rect 9876 16628 9882 16630
rect 10501 16627 10567 16630
rect 12985 16690 13051 16693
rect 13486 16690 13492 16692
rect 12985 16688 13492 16690
rect 12985 16632 12990 16688
rect 13046 16632 13492 16688
rect 12985 16630 13492 16632
rect 12985 16627 13051 16630
rect 13486 16628 13492 16630
rect 13556 16628 13562 16692
rect 16400 16600 17200 16720
rect 2129 16554 2195 16557
rect 7281 16554 7347 16557
rect 8385 16554 8451 16557
rect 2129 16552 8451 16554
rect 2129 16496 2134 16552
rect 2190 16496 7286 16552
rect 7342 16496 8390 16552
rect 8446 16496 8451 16552
rect 2129 16494 8451 16496
rect 2129 16491 2195 16494
rect 7281 16491 7347 16494
rect 8385 16491 8451 16494
rect 10777 16554 10843 16557
rect 12433 16554 12499 16557
rect 12750 16554 12756 16556
rect 10777 16552 12756 16554
rect 10777 16496 10782 16552
rect 10838 16496 12438 16552
rect 12494 16496 12756 16552
rect 10777 16494 12756 16496
rect 10777 16491 10843 16494
rect 12433 16491 12499 16494
rect 12750 16492 12756 16494
rect 12820 16492 12826 16556
rect 10041 16418 10107 16421
rect 11881 16418 11947 16421
rect 10041 16416 11947 16418
rect 10041 16360 10046 16416
rect 10102 16360 11886 16416
rect 11942 16360 11947 16416
rect 10041 16358 11947 16360
rect 10041 16355 10107 16358
rect 11881 16355 11947 16358
rect 4694 16352 5010 16353
rect 4694 16288 4700 16352
rect 4764 16288 4780 16352
rect 4844 16288 4860 16352
rect 4924 16288 4940 16352
rect 5004 16288 5010 16352
rect 4694 16287 5010 16288
rect 8442 16352 8758 16353
rect 8442 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8758 16352
rect 8442 16287 8758 16288
rect 12190 16352 12506 16353
rect 12190 16288 12196 16352
rect 12260 16288 12276 16352
rect 12340 16288 12356 16352
rect 12420 16288 12436 16352
rect 12500 16288 12506 16352
rect 12190 16287 12506 16288
rect 13077 16282 13143 16285
rect 14590 16282 14596 16284
rect 13077 16280 14596 16282
rect 13077 16224 13082 16280
rect 13138 16224 14596 16280
rect 13077 16222 14596 16224
rect 13077 16219 13143 16222
rect 14590 16220 14596 16222
rect 14660 16220 14666 16284
rect 0 16146 800 16176
rect 1485 16146 1551 16149
rect 0 16144 1551 16146
rect 0 16088 1490 16144
rect 1546 16088 1551 16144
rect 0 16086 1551 16088
rect 0 16056 800 16086
rect 1485 16083 1551 16086
rect 3049 16146 3115 16149
rect 15009 16146 15075 16149
rect 3049 16144 15075 16146
rect 3049 16088 3054 16144
rect 3110 16088 15014 16144
rect 15070 16088 15075 16144
rect 3049 16086 15075 16088
rect 3049 16083 3115 16086
rect 15009 16083 15075 16086
rect 5625 16010 5691 16013
rect 8569 16010 8635 16013
rect 5625 16008 8635 16010
rect 5625 15952 5630 16008
rect 5686 15952 8574 16008
rect 8630 15952 8635 16008
rect 5625 15950 8635 15952
rect 5625 15947 5691 15950
rect 8569 15947 8635 15950
rect 11973 16010 12039 16013
rect 13261 16012 13327 16013
rect 13261 16010 13308 16012
rect 11973 16008 13308 16010
rect 13372 16010 13378 16012
rect 11973 15952 11978 16008
rect 12034 15952 13266 16008
rect 11973 15950 13308 15952
rect 11973 15947 12039 15950
rect 13261 15948 13308 15950
rect 13372 15950 13454 16010
rect 13372 15948 13378 15950
rect 13854 15948 13860 16012
rect 13924 16010 13930 16012
rect 13997 16010 14063 16013
rect 13924 16008 14063 16010
rect 13924 15952 14002 16008
rect 14058 15952 14063 16008
rect 13924 15950 14063 15952
rect 13924 15948 13930 15950
rect 13261 15947 13327 15948
rect 13997 15947 14063 15950
rect 3877 15874 3943 15877
rect 6361 15874 6427 15877
rect 3877 15872 6427 15874
rect 3877 15816 3882 15872
rect 3938 15816 6366 15872
rect 6422 15816 6427 15872
rect 3877 15814 6427 15816
rect 3877 15811 3943 15814
rect 6361 15811 6427 15814
rect 2820 15808 3136 15809
rect 2820 15744 2826 15808
rect 2890 15744 2906 15808
rect 2970 15744 2986 15808
rect 3050 15744 3066 15808
rect 3130 15744 3136 15808
rect 2820 15743 3136 15744
rect 6568 15808 6884 15809
rect 6568 15744 6574 15808
rect 6638 15744 6654 15808
rect 6718 15744 6734 15808
rect 6798 15744 6814 15808
rect 6878 15744 6884 15808
rect 6568 15743 6884 15744
rect 10316 15808 10632 15809
rect 10316 15744 10322 15808
rect 10386 15744 10402 15808
rect 10466 15744 10482 15808
rect 10546 15744 10562 15808
rect 10626 15744 10632 15808
rect 10316 15743 10632 15744
rect 14064 15808 14380 15809
rect 14064 15744 14070 15808
rect 14134 15744 14150 15808
rect 14214 15744 14230 15808
rect 14294 15744 14310 15808
rect 14374 15744 14380 15808
rect 14064 15743 14380 15744
rect 2681 15602 2747 15605
rect 14457 15602 14523 15605
rect 2681 15600 14523 15602
rect 2681 15544 2686 15600
rect 2742 15544 14462 15600
rect 14518 15544 14523 15600
rect 2681 15542 14523 15544
rect 2681 15539 2747 15542
rect 14457 15539 14523 15542
rect 8158 15406 9506 15466
rect 1710 15268 1716 15332
rect 1780 15330 1786 15332
rect 2221 15330 2287 15333
rect 1780 15328 2287 15330
rect 1780 15272 2226 15328
rect 2282 15272 2287 15328
rect 1780 15270 2287 15272
rect 1780 15268 1786 15270
rect 2221 15267 2287 15270
rect 2405 15332 2471 15333
rect 2405 15328 2452 15332
rect 2516 15330 2522 15332
rect 2405 15272 2410 15328
rect 2405 15268 2452 15272
rect 2516 15270 2562 15330
rect 2516 15268 2522 15270
rect 6310 15268 6316 15332
rect 6380 15330 6386 15332
rect 6821 15330 6887 15333
rect 8158 15330 8218 15406
rect 6380 15328 8218 15330
rect 6380 15272 6826 15328
rect 6882 15272 8218 15328
rect 6380 15270 8218 15272
rect 6380 15268 6386 15270
rect 2405 15267 2471 15268
rect 6821 15267 6887 15270
rect 4694 15264 5010 15265
rect 0 15194 800 15224
rect 4694 15200 4700 15264
rect 4764 15200 4780 15264
rect 4844 15200 4860 15264
rect 4924 15200 4940 15264
rect 5004 15200 5010 15264
rect 4694 15199 5010 15200
rect 8442 15264 8758 15265
rect 8442 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8758 15264
rect 8442 15199 8758 15200
rect 1485 15194 1551 15197
rect 0 15192 1551 15194
rect 0 15136 1490 15192
rect 1546 15136 1551 15192
rect 0 15134 1551 15136
rect 9446 15194 9506 15406
rect 14641 15330 14707 15333
rect 15326 15330 15332 15332
rect 14641 15328 15332 15330
rect 14641 15272 14646 15328
rect 14702 15272 15332 15328
rect 14641 15270 15332 15272
rect 14641 15267 14707 15270
rect 15326 15268 15332 15270
rect 15396 15268 15402 15332
rect 12190 15264 12506 15265
rect 12190 15200 12196 15264
rect 12260 15200 12276 15264
rect 12340 15200 12356 15264
rect 12420 15200 12436 15264
rect 12500 15200 12506 15264
rect 12190 15199 12506 15200
rect 9765 15194 9831 15197
rect 9446 15192 9831 15194
rect 9446 15136 9770 15192
rect 9826 15136 9831 15192
rect 9446 15134 9831 15136
rect 0 15104 800 15134
rect 1485 15131 1551 15134
rect 9765 15131 9831 15134
rect 2405 15058 2471 15061
rect 10225 15058 10291 15061
rect 2405 15056 10291 15058
rect 2405 15000 2410 15056
rect 2466 15000 10230 15056
rect 10286 15000 10291 15056
rect 2405 14998 10291 15000
rect 2405 14995 2471 14998
rect 10225 14995 10291 14998
rect 12065 15058 12131 15061
rect 12709 15058 12775 15061
rect 12065 15056 12775 15058
rect 12065 15000 12070 15056
rect 12126 15000 12714 15056
rect 12770 15000 12775 15056
rect 12065 14998 12775 15000
rect 12065 14995 12131 14998
rect 12709 14995 12775 14998
rect 9581 14922 9647 14925
rect 12014 14922 12020 14924
rect 9581 14920 12020 14922
rect 9581 14864 9586 14920
rect 9642 14864 12020 14920
rect 9581 14862 12020 14864
rect 9581 14859 9647 14862
rect 12014 14860 12020 14862
rect 12084 14860 12090 14924
rect 15377 14922 15443 14925
rect 12206 14920 15443 14922
rect 12206 14864 15382 14920
rect 15438 14864 15443 14920
rect 12206 14862 15443 14864
rect 11697 14786 11763 14789
rect 12206 14786 12266 14862
rect 15377 14859 15443 14862
rect 11697 14784 12266 14786
rect 11697 14728 11702 14784
rect 11758 14728 12266 14784
rect 11697 14726 12266 14728
rect 11697 14723 11763 14726
rect 2820 14720 3136 14721
rect 2820 14656 2826 14720
rect 2890 14656 2906 14720
rect 2970 14656 2986 14720
rect 3050 14656 3066 14720
rect 3130 14656 3136 14720
rect 2820 14655 3136 14656
rect 6568 14720 6884 14721
rect 6568 14656 6574 14720
rect 6638 14656 6654 14720
rect 6718 14656 6734 14720
rect 6798 14656 6814 14720
rect 6878 14656 6884 14720
rect 6568 14655 6884 14656
rect 10316 14720 10632 14721
rect 10316 14656 10322 14720
rect 10386 14656 10402 14720
rect 10466 14656 10482 14720
rect 10546 14656 10562 14720
rect 10626 14656 10632 14720
rect 10316 14655 10632 14656
rect 14064 14720 14380 14721
rect 14064 14656 14070 14720
rect 14134 14656 14150 14720
rect 14214 14656 14230 14720
rect 14294 14656 14310 14720
rect 14374 14656 14380 14720
rect 14064 14655 14380 14656
rect 10869 14650 10935 14653
rect 12249 14650 12315 14653
rect 10869 14648 12315 14650
rect 10869 14592 10874 14648
rect 10930 14592 12254 14648
rect 12310 14592 12315 14648
rect 10869 14590 12315 14592
rect 10869 14587 10935 14590
rect 12249 14587 12315 14590
rect 1945 14514 2011 14517
rect 11789 14514 11855 14517
rect 1945 14512 11855 14514
rect 1945 14456 1950 14512
rect 2006 14456 11794 14512
rect 11850 14456 11855 14512
rect 1945 14454 11855 14456
rect 1945 14451 2011 14454
rect 11789 14451 11855 14454
rect 12157 14514 12223 14517
rect 12617 14514 12683 14517
rect 12157 14512 12683 14514
rect 12157 14456 12162 14512
rect 12218 14456 12622 14512
rect 12678 14456 12683 14512
rect 12157 14454 12683 14456
rect 12157 14451 12223 14454
rect 12617 14451 12683 14454
rect 10961 14378 11027 14381
rect 12341 14378 12407 14381
rect 16113 14378 16179 14381
rect 10961 14376 16179 14378
rect 10961 14320 10966 14376
rect 11022 14320 12346 14376
rect 12402 14320 16118 14376
rect 16174 14320 16179 14376
rect 10961 14318 16179 14320
rect 10961 14315 11027 14318
rect 12341 14315 12407 14318
rect 16113 14315 16179 14318
rect 0 14242 800 14272
rect 1485 14242 1551 14245
rect 0 14240 1551 14242
rect 0 14184 1490 14240
rect 1546 14184 1551 14240
rect 0 14182 1551 14184
rect 0 14152 800 14182
rect 1485 14179 1551 14182
rect 2865 14242 2931 14245
rect 4061 14244 4127 14245
rect 4061 14242 4108 14244
rect 2865 14240 4108 14242
rect 2865 14184 2870 14240
rect 2926 14184 4066 14240
rect 2865 14182 4108 14184
rect 2865 14179 2931 14182
rect 4061 14180 4108 14182
rect 4172 14180 4178 14244
rect 7414 14180 7420 14244
rect 7484 14242 7490 14244
rect 7649 14242 7715 14245
rect 7484 14240 7715 14242
rect 7484 14184 7654 14240
rect 7710 14184 7715 14240
rect 7484 14182 7715 14184
rect 7484 14180 7490 14182
rect 4061 14179 4127 14180
rect 7649 14179 7715 14182
rect 10777 14242 10843 14245
rect 10961 14242 11027 14245
rect 10777 14240 11027 14242
rect 10777 14184 10782 14240
rect 10838 14184 10966 14240
rect 11022 14184 11027 14240
rect 10777 14182 11027 14184
rect 10777 14179 10843 14182
rect 10961 14179 11027 14182
rect 4694 14176 5010 14177
rect 4694 14112 4700 14176
rect 4764 14112 4780 14176
rect 4844 14112 4860 14176
rect 4924 14112 4940 14176
rect 5004 14112 5010 14176
rect 4694 14111 5010 14112
rect 8442 14176 8758 14177
rect 8442 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8758 14176
rect 8442 14111 8758 14112
rect 12190 14176 12506 14177
rect 12190 14112 12196 14176
rect 12260 14112 12276 14176
rect 12340 14112 12356 14176
rect 12420 14112 12436 14176
rect 12500 14112 12506 14176
rect 12190 14111 12506 14112
rect 2405 13970 2471 13973
rect 12525 13970 12591 13973
rect 2405 13968 12591 13970
rect 2405 13912 2410 13968
rect 2466 13912 12530 13968
rect 12586 13912 12591 13968
rect 2405 13910 12591 13912
rect 2405 13907 2471 13910
rect 12525 13907 12591 13910
rect 6637 13834 6703 13837
rect 9254 13834 9260 13836
rect 6637 13832 9260 13834
rect 6637 13776 6642 13832
rect 6698 13776 9260 13832
rect 6637 13774 9260 13776
rect 6637 13771 6703 13774
rect 9254 13772 9260 13774
rect 9324 13772 9330 13836
rect 9489 13834 9555 13837
rect 12566 13834 12572 13836
rect 9489 13832 12572 13834
rect 9489 13776 9494 13832
rect 9550 13776 12572 13832
rect 9489 13774 12572 13776
rect 9489 13771 9555 13774
rect 12566 13772 12572 13774
rect 12636 13834 12642 13836
rect 12709 13834 12775 13837
rect 12636 13832 12775 13834
rect 12636 13776 12714 13832
rect 12770 13776 12775 13832
rect 12636 13774 12775 13776
rect 12636 13772 12642 13774
rect 12709 13771 12775 13774
rect 9305 13698 9371 13701
rect 9489 13698 9555 13701
rect 9305 13696 9555 13698
rect 9305 13640 9310 13696
rect 9366 13640 9494 13696
rect 9550 13640 9555 13696
rect 9305 13638 9555 13640
rect 9305 13635 9371 13638
rect 9489 13635 9555 13638
rect 10133 13698 10199 13701
rect 11421 13698 11487 13701
rect 12433 13698 12499 13701
rect 13537 13698 13603 13701
rect 10133 13696 10242 13698
rect 10133 13640 10138 13696
rect 10194 13640 10242 13696
rect 10133 13635 10242 13640
rect 11421 13696 12499 13698
rect 11421 13640 11426 13696
rect 11482 13640 12438 13696
rect 12494 13640 12499 13696
rect 11421 13638 12499 13640
rect 11421 13635 11487 13638
rect 12433 13635 12499 13638
rect 13356 13696 13603 13698
rect 13356 13640 13542 13696
rect 13598 13640 13603 13696
rect 13356 13638 13603 13640
rect 2820 13632 3136 13633
rect 2820 13568 2826 13632
rect 2890 13568 2906 13632
rect 2970 13568 2986 13632
rect 3050 13568 3066 13632
rect 3130 13568 3136 13632
rect 2820 13567 3136 13568
rect 6568 13632 6884 13633
rect 6568 13568 6574 13632
rect 6638 13568 6654 13632
rect 6718 13568 6734 13632
rect 6798 13568 6814 13632
rect 6878 13568 6884 13632
rect 6568 13567 6884 13568
rect 9673 13426 9739 13429
rect 10182 13426 10242 13635
rect 10316 13632 10632 13633
rect 10316 13568 10322 13632
rect 10386 13568 10402 13632
rect 10466 13568 10482 13632
rect 10546 13568 10562 13632
rect 10626 13568 10632 13632
rect 10316 13567 10632 13568
rect 12014 13500 12020 13564
rect 12084 13562 12090 13564
rect 13356 13562 13416 13638
rect 13537 13635 13603 13638
rect 14064 13632 14380 13633
rect 14064 13568 14070 13632
rect 14134 13568 14150 13632
rect 14214 13568 14230 13632
rect 14294 13568 14310 13632
rect 14374 13568 14380 13632
rect 14064 13567 14380 13568
rect 13537 13564 13603 13565
rect 12084 13502 13416 13562
rect 12084 13500 12090 13502
rect 13486 13500 13492 13564
rect 13556 13562 13603 13564
rect 13813 13564 13879 13565
rect 13813 13562 13860 13564
rect 13556 13560 13648 13562
rect 13598 13504 13648 13560
rect 13556 13502 13648 13504
rect 13768 13560 13860 13562
rect 13768 13504 13818 13560
rect 13768 13502 13860 13504
rect 13556 13500 13603 13502
rect 13537 13499 13603 13500
rect 13813 13500 13860 13502
rect 13924 13500 13930 13564
rect 13813 13499 13879 13500
rect 14457 13426 14523 13429
rect 9673 13424 14523 13426
rect 9673 13368 9678 13424
rect 9734 13368 14462 13424
rect 14518 13368 14523 13424
rect 9673 13366 14523 13368
rect 9673 13363 9739 13366
rect 14457 13363 14523 13366
rect 0 13290 800 13320
rect 1485 13290 1551 13293
rect 0 13288 1551 13290
rect 0 13232 1490 13288
rect 1546 13232 1551 13288
rect 0 13230 1551 13232
rect 0 13200 800 13230
rect 1485 13227 1551 13230
rect 1761 13290 1827 13293
rect 11053 13290 11119 13293
rect 14641 13290 14707 13293
rect 1761 13288 11119 13290
rect 1761 13232 1766 13288
rect 1822 13232 11058 13288
rect 11114 13232 11119 13288
rect 1761 13230 11119 13232
rect 1761 13227 1827 13230
rect 11053 13227 11119 13230
rect 12068 13288 14707 13290
rect 12068 13232 14646 13288
rect 14702 13232 14707 13288
rect 12068 13230 14707 13232
rect 9949 13154 10015 13157
rect 12068 13154 12128 13230
rect 14641 13227 14707 13230
rect 9949 13152 12128 13154
rect 9949 13096 9954 13152
rect 10010 13096 12128 13152
rect 9949 13094 12128 13096
rect 13261 13154 13327 13157
rect 13486 13154 13492 13156
rect 13261 13152 13492 13154
rect 13261 13096 13266 13152
rect 13322 13096 13492 13152
rect 13261 13094 13492 13096
rect 9949 13091 10015 13094
rect 13261 13091 13327 13094
rect 13486 13092 13492 13094
rect 13556 13092 13562 13156
rect 13670 13092 13676 13156
rect 13740 13154 13746 13156
rect 14273 13154 14339 13157
rect 13740 13152 14339 13154
rect 13740 13096 14278 13152
rect 14334 13096 14339 13152
rect 13740 13094 14339 13096
rect 13740 13092 13746 13094
rect 14273 13091 14339 13094
rect 4694 13088 5010 13089
rect 4694 13024 4700 13088
rect 4764 13024 4780 13088
rect 4844 13024 4860 13088
rect 4924 13024 4940 13088
rect 5004 13024 5010 13088
rect 4694 13023 5010 13024
rect 8442 13088 8758 13089
rect 8442 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8758 13088
rect 8442 13023 8758 13024
rect 12190 13088 12506 13089
rect 12190 13024 12196 13088
rect 12260 13024 12276 13088
rect 12340 13024 12356 13088
rect 12420 13024 12436 13088
rect 12500 13024 12506 13088
rect 12190 13023 12506 13024
rect 7649 12882 7715 12885
rect 13353 12882 13419 12885
rect 7649 12880 13419 12882
rect 7649 12824 7654 12880
rect 7710 12824 13358 12880
rect 13414 12824 13419 12880
rect 7649 12822 13419 12824
rect 7649 12819 7715 12822
rect 13353 12819 13419 12822
rect 5257 12746 5323 12749
rect 8886 12746 8892 12748
rect 5257 12744 8892 12746
rect 5257 12688 5262 12744
rect 5318 12688 8892 12744
rect 5257 12686 8892 12688
rect 5257 12683 5323 12686
rect 8886 12684 8892 12686
rect 8956 12684 8962 12748
rect 10225 12746 10291 12749
rect 16849 12746 16915 12749
rect 10225 12744 16915 12746
rect 10225 12688 10230 12744
rect 10286 12688 16854 12744
rect 16910 12688 16915 12744
rect 10225 12686 16915 12688
rect 10225 12683 10291 12686
rect 16849 12683 16915 12686
rect 4245 12610 4311 12613
rect 6126 12610 6132 12612
rect 4245 12608 6132 12610
rect 4245 12552 4250 12608
rect 4306 12552 6132 12608
rect 4245 12550 6132 12552
rect 4245 12547 4311 12550
rect 6126 12548 6132 12550
rect 6196 12548 6202 12612
rect 6361 12610 6427 12613
rect 6318 12608 6427 12610
rect 6318 12552 6366 12608
rect 6422 12552 6427 12608
rect 6318 12547 6427 12552
rect 2820 12544 3136 12545
rect 2820 12480 2826 12544
rect 2890 12480 2906 12544
rect 2970 12480 2986 12544
rect 3050 12480 3066 12544
rect 3130 12480 3136 12544
rect 2820 12479 3136 12480
rect 5625 12474 5691 12477
rect 6318 12474 6378 12547
rect 6568 12544 6884 12545
rect 6568 12480 6574 12544
rect 6638 12480 6654 12544
rect 6718 12480 6734 12544
rect 6798 12480 6814 12544
rect 6878 12480 6884 12544
rect 6568 12479 6884 12480
rect 10316 12544 10632 12545
rect 10316 12480 10322 12544
rect 10386 12480 10402 12544
rect 10466 12480 10482 12544
rect 10546 12480 10562 12544
rect 10626 12480 10632 12544
rect 10316 12479 10632 12480
rect 14064 12544 14380 12545
rect 14064 12480 14070 12544
rect 14134 12480 14150 12544
rect 14214 12480 14230 12544
rect 14294 12480 14310 12544
rect 14374 12480 14380 12544
rect 14064 12479 14380 12480
rect 9857 12474 9923 12477
rect 5625 12472 6378 12474
rect 5625 12416 5630 12472
rect 5686 12416 6378 12472
rect 5625 12414 6378 12416
rect 9446 12472 9923 12474
rect 9446 12416 9862 12472
rect 9918 12416 9923 12472
rect 9446 12414 9923 12416
rect 5625 12411 5691 12414
rect 0 12338 800 12368
rect 1485 12338 1551 12341
rect 0 12336 1551 12338
rect 0 12280 1490 12336
rect 1546 12280 1551 12336
rect 0 12278 1551 12280
rect 0 12248 800 12278
rect 1485 12275 1551 12278
rect 7557 12338 7623 12341
rect 9446 12340 9506 12414
rect 9857 12411 9923 12414
rect 9438 12338 9444 12340
rect 7557 12336 9444 12338
rect 7557 12280 7562 12336
rect 7618 12280 9444 12336
rect 7557 12278 9444 12280
rect 7557 12275 7623 12278
rect 9438 12276 9444 12278
rect 9508 12276 9514 12340
rect 10910 12276 10916 12340
rect 10980 12338 10986 12340
rect 12341 12338 12407 12341
rect 10980 12336 12407 12338
rect 10980 12280 12346 12336
rect 12402 12280 12407 12336
rect 10980 12278 12407 12280
rect 10980 12276 10986 12278
rect 12341 12275 12407 12278
rect 12525 12338 12591 12341
rect 12750 12338 12756 12340
rect 12525 12336 12756 12338
rect 12525 12280 12530 12336
rect 12586 12280 12756 12336
rect 12525 12278 12756 12280
rect 12525 12275 12591 12278
rect 12750 12276 12756 12278
rect 12820 12276 12826 12340
rect 9673 12202 9739 12205
rect 9806 12202 9812 12204
rect 9673 12200 9812 12202
rect 9673 12144 9678 12200
rect 9734 12144 9812 12200
rect 9673 12142 9812 12144
rect 9673 12139 9739 12142
rect 9806 12140 9812 12142
rect 9876 12140 9882 12204
rect 4694 12000 5010 12001
rect 4694 11936 4700 12000
rect 4764 11936 4780 12000
rect 4844 11936 4860 12000
rect 4924 11936 4940 12000
rect 5004 11936 5010 12000
rect 4694 11935 5010 11936
rect 8442 12000 8758 12001
rect 8442 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8758 12000
rect 8442 11935 8758 11936
rect 12190 12000 12506 12001
rect 12190 11936 12196 12000
rect 12260 11936 12276 12000
rect 12340 11936 12356 12000
rect 12420 11936 12436 12000
rect 12500 11936 12506 12000
rect 12190 11935 12506 11936
rect 10174 11868 10180 11932
rect 10244 11930 10250 11932
rect 10317 11930 10383 11933
rect 10244 11928 10383 11930
rect 10244 11872 10322 11928
rect 10378 11872 10383 11928
rect 10244 11870 10383 11872
rect 10244 11868 10250 11870
rect 10317 11867 10383 11870
rect 10685 11930 10751 11933
rect 10869 11930 10935 11933
rect 11513 11932 11579 11933
rect 10685 11928 10935 11930
rect 10685 11872 10690 11928
rect 10746 11872 10874 11928
rect 10930 11872 10935 11928
rect 10685 11870 10935 11872
rect 10685 11867 10751 11870
rect 10869 11867 10935 11870
rect 11462 11868 11468 11932
rect 11532 11930 11579 11932
rect 11532 11928 11624 11930
rect 11574 11872 11624 11928
rect 11532 11870 11624 11872
rect 11532 11868 11579 11870
rect 11513 11867 11579 11868
rect 4153 11794 4219 11797
rect 11697 11794 11763 11797
rect 13353 11794 13419 11797
rect 4153 11792 13419 11794
rect 4153 11736 4158 11792
rect 4214 11736 11702 11792
rect 11758 11736 13358 11792
rect 13414 11736 13419 11792
rect 4153 11734 13419 11736
rect 4153 11731 4219 11734
rect 11697 11731 11763 11734
rect 13353 11731 13419 11734
rect 7741 11658 7807 11661
rect 14641 11658 14707 11661
rect 7741 11656 14707 11658
rect 7741 11600 7746 11656
rect 7802 11600 14646 11656
rect 14702 11600 14707 11656
rect 7741 11598 14707 11600
rect 7741 11595 7807 11598
rect 14641 11595 14707 11598
rect 2820 11456 3136 11457
rect 0 11386 800 11416
rect 2820 11392 2826 11456
rect 2890 11392 2906 11456
rect 2970 11392 2986 11456
rect 3050 11392 3066 11456
rect 3130 11392 3136 11456
rect 2820 11391 3136 11392
rect 6568 11456 6884 11457
rect 6568 11392 6574 11456
rect 6638 11392 6654 11456
rect 6718 11392 6734 11456
rect 6798 11392 6814 11456
rect 6878 11392 6884 11456
rect 6568 11391 6884 11392
rect 10316 11456 10632 11457
rect 10316 11392 10322 11456
rect 10386 11392 10402 11456
rect 10466 11392 10482 11456
rect 10546 11392 10562 11456
rect 10626 11392 10632 11456
rect 10316 11391 10632 11392
rect 14064 11456 14380 11457
rect 14064 11392 14070 11456
rect 14134 11392 14150 11456
rect 14214 11392 14230 11456
rect 14294 11392 14310 11456
rect 14374 11392 14380 11456
rect 14064 11391 14380 11392
rect 1485 11386 1551 11389
rect 0 11384 1551 11386
rect 0 11328 1490 11384
rect 1546 11328 1551 11384
rect 0 11326 1551 11328
rect 0 11296 800 11326
rect 1485 11323 1551 11326
rect 4705 11114 4771 11117
rect 9673 11114 9739 11117
rect 4705 11112 9739 11114
rect 4705 11056 4710 11112
rect 4766 11056 9678 11112
rect 9734 11056 9739 11112
rect 4705 11054 9739 11056
rect 4705 11051 4771 11054
rect 9673 11051 9739 11054
rect 4694 10912 5010 10913
rect 4694 10848 4700 10912
rect 4764 10848 4780 10912
rect 4844 10848 4860 10912
rect 4924 10848 4940 10912
rect 5004 10848 5010 10912
rect 4694 10847 5010 10848
rect 8442 10912 8758 10913
rect 8442 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8758 10912
rect 8442 10847 8758 10848
rect 12190 10912 12506 10913
rect 12190 10848 12196 10912
rect 12260 10848 12276 10912
rect 12340 10848 12356 10912
rect 12420 10848 12436 10912
rect 12500 10848 12506 10912
rect 12190 10847 12506 10848
rect 3233 10570 3299 10573
rect 12985 10570 13051 10573
rect 3233 10568 13051 10570
rect 3233 10512 3238 10568
rect 3294 10512 12990 10568
rect 13046 10512 13051 10568
rect 3233 10510 13051 10512
rect 3233 10507 3299 10510
rect 12985 10507 13051 10510
rect 0 10434 800 10464
rect 1485 10434 1551 10437
rect 0 10432 1551 10434
rect 0 10376 1490 10432
rect 1546 10376 1551 10432
rect 0 10374 1551 10376
rect 0 10344 800 10374
rect 1485 10371 1551 10374
rect 2820 10368 3136 10369
rect 2820 10304 2826 10368
rect 2890 10304 2906 10368
rect 2970 10304 2986 10368
rect 3050 10304 3066 10368
rect 3130 10304 3136 10368
rect 2820 10303 3136 10304
rect 6568 10368 6884 10369
rect 6568 10304 6574 10368
rect 6638 10304 6654 10368
rect 6718 10304 6734 10368
rect 6798 10304 6814 10368
rect 6878 10304 6884 10368
rect 6568 10303 6884 10304
rect 10316 10368 10632 10369
rect 10316 10304 10322 10368
rect 10386 10304 10402 10368
rect 10466 10304 10482 10368
rect 10546 10304 10562 10368
rect 10626 10304 10632 10368
rect 10316 10303 10632 10304
rect 14064 10368 14380 10369
rect 14064 10304 14070 10368
rect 14134 10304 14150 10368
rect 14214 10304 14230 10368
rect 14294 10304 14310 10368
rect 14374 10304 14380 10368
rect 14064 10303 14380 10304
rect 12065 10298 12131 10301
rect 13813 10300 13879 10301
rect 13813 10298 13860 10300
rect 12065 10296 13860 10298
rect 12065 10240 12070 10296
rect 12126 10240 13818 10296
rect 12065 10238 13860 10240
rect 12065 10235 12131 10238
rect 13813 10236 13860 10238
rect 13924 10236 13930 10300
rect 13813 10235 13879 10236
rect 13118 10100 13124 10164
rect 13188 10162 13194 10164
rect 13261 10162 13327 10165
rect 13188 10160 13327 10162
rect 13188 10104 13266 10160
rect 13322 10104 13327 10160
rect 13188 10102 13327 10104
rect 13188 10100 13194 10102
rect 13261 10099 13327 10102
rect 11237 10026 11303 10029
rect 12801 10026 12867 10029
rect 13445 10028 13511 10029
rect 13445 10026 13492 10028
rect 11237 10024 12867 10026
rect 11237 9968 11242 10024
rect 11298 9968 12806 10024
rect 12862 9968 12867 10024
rect 11237 9966 12867 9968
rect 13400 10024 13492 10026
rect 13400 9968 13450 10024
rect 13400 9966 13492 9968
rect 11237 9963 11303 9966
rect 12801 9963 12867 9966
rect 13445 9964 13492 9966
rect 13556 9964 13562 10028
rect 14590 9964 14596 10028
rect 14660 10026 14666 10028
rect 14733 10026 14799 10029
rect 14660 10024 14799 10026
rect 14660 9968 14738 10024
rect 14794 9968 14799 10024
rect 14660 9966 14799 9968
rect 14660 9964 14666 9966
rect 13445 9963 13511 9964
rect 14733 9963 14799 9966
rect 15101 10026 15167 10029
rect 16400 10026 17200 10056
rect 15101 10024 17200 10026
rect 15101 9968 15106 10024
rect 15162 9968 17200 10024
rect 15101 9966 17200 9968
rect 15101 9963 15167 9966
rect 16400 9936 17200 9966
rect 9489 9890 9555 9893
rect 11094 9890 11100 9892
rect 9489 9888 11100 9890
rect 9489 9832 9494 9888
rect 9550 9832 11100 9888
rect 9489 9830 11100 9832
rect 9489 9827 9555 9830
rect 11094 9828 11100 9830
rect 11164 9828 11170 9892
rect 12709 9890 12775 9893
rect 13353 9890 13419 9893
rect 12709 9888 13419 9890
rect 12709 9832 12714 9888
rect 12770 9832 13358 9888
rect 13414 9832 13419 9888
rect 12709 9830 13419 9832
rect 12709 9827 12775 9830
rect 13353 9827 13419 9830
rect 4694 9824 5010 9825
rect 4694 9760 4700 9824
rect 4764 9760 4780 9824
rect 4844 9760 4860 9824
rect 4924 9760 4940 9824
rect 5004 9760 5010 9824
rect 4694 9759 5010 9760
rect 8442 9824 8758 9825
rect 8442 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8758 9824
rect 8442 9759 8758 9760
rect 12190 9824 12506 9825
rect 12190 9760 12196 9824
rect 12260 9760 12276 9824
rect 12340 9760 12356 9824
rect 12420 9760 12436 9824
rect 12500 9760 12506 9824
rect 12190 9759 12506 9760
rect 9630 9630 10058 9690
rect 4102 9556 4108 9620
rect 4172 9618 4178 9620
rect 9630 9618 9690 9630
rect 4172 9558 9690 9618
rect 9998 9618 10058 9630
rect 13486 9618 13492 9620
rect 9998 9558 13492 9618
rect 4172 9556 4178 9558
rect 13486 9556 13492 9558
rect 13556 9618 13562 9620
rect 14457 9618 14523 9621
rect 13556 9616 14523 9618
rect 13556 9560 14462 9616
rect 14518 9560 14523 9616
rect 13556 9558 14523 9560
rect 13556 9556 13562 9558
rect 14457 9555 14523 9558
rect 0 9482 800 9512
rect 1485 9482 1551 9485
rect 0 9480 1551 9482
rect 0 9424 1490 9480
rect 1546 9424 1551 9480
rect 0 9422 1551 9424
rect 0 9392 800 9422
rect 1485 9419 1551 9422
rect 4429 9482 4495 9485
rect 11973 9482 12039 9485
rect 12801 9482 12867 9485
rect 4429 9480 9322 9482
rect 4429 9424 4434 9480
rect 4490 9424 9322 9480
rect 4429 9422 9322 9424
rect 4429 9419 4495 9422
rect 2820 9280 3136 9281
rect 2820 9216 2826 9280
rect 2890 9216 2906 9280
rect 2970 9216 2986 9280
rect 3050 9216 3066 9280
rect 3130 9216 3136 9280
rect 2820 9215 3136 9216
rect 6568 9280 6884 9281
rect 6568 9216 6574 9280
rect 6638 9216 6654 9280
rect 6718 9216 6734 9280
rect 6798 9216 6814 9280
rect 6878 9216 6884 9280
rect 6568 9215 6884 9216
rect 7966 9148 7972 9212
rect 8036 9210 8042 9212
rect 8293 9210 8359 9213
rect 8036 9208 8359 9210
rect 8036 9152 8298 9208
rect 8354 9152 8359 9208
rect 8036 9150 8359 9152
rect 8036 9148 8042 9150
rect 8293 9147 8359 9150
rect 5390 9012 5396 9076
rect 5460 9074 5466 9076
rect 8886 9074 8892 9076
rect 5460 9014 8892 9074
rect 5460 9012 5466 9014
rect 8886 9012 8892 9014
rect 8956 9074 8962 9076
rect 9121 9074 9187 9077
rect 8956 9072 9187 9074
rect 8956 9016 9126 9072
rect 9182 9016 9187 9072
rect 8956 9014 9187 9016
rect 9262 9074 9322 9422
rect 11973 9480 12867 9482
rect 11973 9424 11978 9480
rect 12034 9424 12806 9480
rect 12862 9424 12867 9480
rect 11973 9422 12867 9424
rect 11973 9419 12039 9422
rect 12801 9419 12867 9422
rect 13670 9420 13676 9484
rect 13740 9482 13746 9484
rect 13997 9482 14063 9485
rect 13740 9480 14063 9482
rect 13740 9424 14002 9480
rect 14058 9424 14063 9480
rect 13740 9422 14063 9424
rect 13740 9420 13746 9422
rect 13997 9419 14063 9422
rect 11278 9284 11284 9348
rect 11348 9346 11354 9348
rect 12065 9346 12131 9349
rect 11348 9344 12131 9346
rect 11348 9288 12070 9344
rect 12126 9288 12131 9344
rect 11348 9286 12131 9288
rect 11348 9284 11354 9286
rect 12065 9283 12131 9286
rect 10316 9280 10632 9281
rect 10316 9216 10322 9280
rect 10386 9216 10402 9280
rect 10466 9216 10482 9280
rect 10546 9216 10562 9280
rect 10626 9216 10632 9280
rect 10316 9215 10632 9216
rect 14064 9280 14380 9281
rect 14064 9216 14070 9280
rect 14134 9216 14150 9280
rect 14214 9216 14230 9280
rect 14294 9216 14310 9280
rect 14374 9216 14380 9280
rect 14064 9215 14380 9216
rect 11462 9148 11468 9212
rect 11532 9210 11538 9212
rect 12014 9210 12020 9212
rect 11532 9150 12020 9210
rect 11532 9148 11538 9150
rect 12014 9148 12020 9150
rect 12084 9210 12090 9212
rect 13537 9210 13603 9213
rect 12084 9208 13603 9210
rect 12084 9152 13542 9208
rect 13598 9152 13603 9208
rect 12084 9150 13603 9152
rect 12084 9148 12090 9150
rect 13537 9147 13603 9150
rect 14181 9074 14247 9077
rect 9262 9072 14247 9074
rect 9262 9016 14186 9072
rect 14242 9016 14247 9072
rect 9262 9014 14247 9016
rect 8956 9012 8962 9014
rect 9121 9011 9187 9014
rect 14181 9011 14247 9014
rect 14365 9074 14431 9077
rect 14549 9074 14615 9077
rect 14365 9072 14615 9074
rect 14365 9016 14370 9072
rect 14426 9016 14554 9072
rect 14610 9016 14615 9072
rect 14365 9014 14615 9016
rect 14365 9011 14431 9014
rect 14549 9011 14615 9014
rect 1853 8938 1919 8941
rect 13629 8938 13695 8941
rect 1853 8936 13695 8938
rect 1853 8880 1858 8936
rect 1914 8880 13634 8936
rect 13690 8880 13695 8936
rect 1853 8878 13695 8880
rect 1853 8875 1919 8878
rect 13629 8875 13695 8878
rect 8150 8740 8156 8804
rect 8220 8802 8226 8804
rect 8293 8802 8359 8805
rect 8220 8800 8359 8802
rect 8220 8744 8298 8800
rect 8354 8744 8359 8800
rect 8220 8742 8359 8744
rect 8220 8740 8226 8742
rect 8293 8739 8359 8742
rect 9765 8802 9831 8805
rect 11973 8802 12039 8805
rect 9765 8800 12039 8802
rect 9765 8744 9770 8800
rect 9826 8744 11978 8800
rect 12034 8744 12039 8800
rect 9765 8742 12039 8744
rect 9765 8739 9831 8742
rect 11973 8739 12039 8742
rect 13670 8740 13676 8804
rect 13740 8802 13746 8804
rect 14089 8802 14155 8805
rect 13740 8800 14155 8802
rect 13740 8744 14094 8800
rect 14150 8744 14155 8800
rect 13740 8742 14155 8744
rect 13740 8740 13746 8742
rect 14089 8739 14155 8742
rect 4694 8736 5010 8737
rect 4694 8672 4700 8736
rect 4764 8672 4780 8736
rect 4844 8672 4860 8736
rect 4924 8672 4940 8736
rect 5004 8672 5010 8736
rect 4694 8671 5010 8672
rect 8442 8736 8758 8737
rect 8442 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8758 8736
rect 8442 8671 8758 8672
rect 12190 8736 12506 8737
rect 12190 8672 12196 8736
rect 12260 8672 12276 8736
rect 12340 8672 12356 8736
rect 12420 8672 12436 8736
rect 12500 8672 12506 8736
rect 12190 8671 12506 8672
rect 8845 8666 8911 8669
rect 10593 8666 10659 8669
rect 16113 8666 16179 8669
rect 8845 8664 10659 8666
rect 8845 8608 8850 8664
rect 8906 8608 10598 8664
rect 10654 8608 10659 8664
rect 8845 8606 10659 8608
rect 8845 8603 8911 8606
rect 10593 8603 10659 8606
rect 13494 8664 16179 8666
rect 13494 8608 16118 8664
rect 16174 8608 16179 8664
rect 13494 8606 16179 8608
rect 0 8530 800 8560
rect 1485 8530 1551 8533
rect 0 8528 1551 8530
rect 0 8472 1490 8528
rect 1546 8472 1551 8528
rect 0 8470 1551 8472
rect 0 8440 800 8470
rect 1485 8467 1551 8470
rect 6729 8530 6795 8533
rect 9581 8530 9647 8533
rect 6729 8528 9647 8530
rect 6729 8472 6734 8528
rect 6790 8472 9586 8528
rect 9642 8472 9647 8528
rect 6729 8470 9647 8472
rect 6729 8467 6795 8470
rect 9581 8467 9647 8470
rect 9806 8468 9812 8532
rect 9876 8530 9882 8532
rect 9949 8530 10015 8533
rect 11881 8532 11947 8533
rect 9876 8528 10015 8530
rect 9876 8472 9954 8528
rect 10010 8472 10015 8528
rect 9876 8470 10015 8472
rect 9876 8468 9882 8470
rect 9949 8467 10015 8470
rect 11830 8468 11836 8532
rect 11900 8530 11947 8532
rect 12065 8530 12131 8533
rect 12566 8530 12572 8532
rect 11900 8528 11992 8530
rect 11942 8472 11992 8528
rect 11900 8470 11992 8472
rect 12065 8528 12572 8530
rect 12065 8472 12070 8528
rect 12126 8472 12572 8528
rect 12065 8470 12572 8472
rect 11900 8468 11947 8470
rect 11881 8467 11947 8468
rect 12065 8467 12131 8470
rect 12566 8468 12572 8470
rect 12636 8530 12642 8532
rect 13494 8530 13554 8606
rect 16113 8603 16179 8606
rect 12636 8470 13554 8530
rect 12636 8468 12642 8470
rect 1945 8394 2011 8397
rect 12341 8394 12407 8397
rect 1945 8392 12407 8394
rect 1945 8336 1950 8392
rect 2006 8336 12346 8392
rect 12402 8336 12407 8392
rect 1945 8334 12407 8336
rect 1945 8331 2011 8334
rect 12341 8331 12407 8334
rect 2820 8192 3136 8193
rect 2820 8128 2826 8192
rect 2890 8128 2906 8192
rect 2970 8128 2986 8192
rect 3050 8128 3066 8192
rect 3130 8128 3136 8192
rect 2820 8127 3136 8128
rect 6568 8192 6884 8193
rect 6568 8128 6574 8192
rect 6638 8128 6654 8192
rect 6718 8128 6734 8192
rect 6798 8128 6814 8192
rect 6878 8128 6884 8192
rect 6568 8127 6884 8128
rect 10316 8192 10632 8193
rect 10316 8128 10322 8192
rect 10386 8128 10402 8192
rect 10466 8128 10482 8192
rect 10546 8128 10562 8192
rect 10626 8128 10632 8192
rect 10316 8127 10632 8128
rect 14064 8192 14380 8193
rect 14064 8128 14070 8192
rect 14134 8128 14150 8192
rect 14214 8128 14230 8192
rect 14294 8128 14310 8192
rect 14374 8128 14380 8192
rect 14064 8127 14380 8128
rect 9622 8060 9628 8124
rect 9692 8122 9698 8124
rect 9765 8122 9831 8125
rect 9692 8120 9831 8122
rect 9692 8064 9770 8120
rect 9826 8064 9831 8120
rect 9692 8062 9831 8064
rect 9692 8060 9698 8062
rect 9765 8059 9831 8062
rect 7005 7986 7071 7989
rect 10726 7986 10732 7988
rect 7005 7984 10732 7986
rect 7005 7928 7010 7984
rect 7066 7928 10732 7984
rect 7005 7926 10732 7928
rect 7005 7923 7071 7926
rect 10726 7924 10732 7926
rect 10796 7986 10802 7988
rect 12157 7986 12223 7989
rect 13905 7988 13971 7989
rect 13854 7986 13860 7988
rect 10796 7984 12223 7986
rect 10796 7928 12162 7984
rect 12218 7928 12223 7984
rect 10796 7926 12223 7928
rect 13778 7926 13860 7986
rect 13924 7986 13971 7988
rect 16205 7986 16271 7989
rect 13924 7984 16271 7986
rect 13966 7928 16210 7984
rect 16266 7928 16271 7984
rect 10796 7924 10802 7926
rect 12157 7923 12223 7926
rect 13854 7924 13860 7926
rect 13924 7926 16271 7928
rect 13924 7924 13971 7926
rect 13905 7923 13971 7924
rect 16205 7923 16271 7926
rect 5165 7850 5231 7853
rect 11053 7850 11119 7853
rect 5165 7848 11119 7850
rect 5165 7792 5170 7848
rect 5226 7792 11058 7848
rect 11114 7792 11119 7848
rect 5165 7790 11119 7792
rect 5165 7787 5231 7790
rect 11053 7787 11119 7790
rect 12525 7850 12591 7853
rect 12525 7848 12634 7850
rect 12525 7792 12530 7848
rect 12586 7792 12634 7848
rect 12525 7787 12634 7792
rect 9765 7714 9831 7717
rect 11329 7714 11395 7717
rect 12574 7716 12634 7787
rect 9765 7712 11395 7714
rect 9765 7656 9770 7712
rect 9826 7656 11334 7712
rect 11390 7656 11395 7712
rect 9765 7654 11395 7656
rect 9765 7651 9831 7654
rect 11329 7651 11395 7654
rect 12566 7652 12572 7716
rect 12636 7714 12642 7716
rect 13445 7714 13511 7717
rect 12636 7712 13511 7714
rect 12636 7656 13450 7712
rect 13506 7656 13511 7712
rect 12636 7654 13511 7656
rect 12636 7652 12642 7654
rect 13445 7651 13511 7654
rect 14641 7714 14707 7717
rect 15101 7714 15167 7717
rect 14641 7712 15167 7714
rect 14641 7656 14646 7712
rect 14702 7656 15106 7712
rect 15162 7656 15167 7712
rect 14641 7654 15167 7656
rect 14641 7651 14707 7654
rect 15101 7651 15167 7654
rect 4694 7648 5010 7649
rect 0 7578 800 7608
rect 4694 7584 4700 7648
rect 4764 7584 4780 7648
rect 4844 7584 4860 7648
rect 4924 7584 4940 7648
rect 5004 7584 5010 7648
rect 4694 7583 5010 7584
rect 8442 7648 8758 7649
rect 8442 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8758 7648
rect 8442 7583 8758 7584
rect 12190 7648 12506 7649
rect 12190 7584 12196 7648
rect 12260 7584 12276 7648
rect 12340 7584 12356 7648
rect 12420 7584 12436 7648
rect 12500 7584 12506 7648
rect 12190 7583 12506 7584
rect 1485 7578 1551 7581
rect 0 7576 1551 7578
rect 0 7520 1490 7576
rect 1546 7520 1551 7576
rect 0 7518 1551 7520
rect 0 7488 800 7518
rect 1485 7515 1551 7518
rect 8845 7580 8911 7581
rect 8845 7576 8892 7580
rect 8956 7578 8962 7580
rect 14549 7578 14615 7581
rect 8845 7520 8850 7576
rect 8845 7516 8892 7520
rect 8956 7518 9002 7578
rect 12574 7576 14615 7578
rect 12574 7520 14554 7576
rect 14610 7520 14615 7576
rect 12574 7518 14615 7520
rect 8956 7516 8962 7518
rect 8845 7515 8911 7516
rect 5942 7380 5948 7444
rect 6012 7442 6018 7444
rect 12341 7442 12407 7445
rect 6012 7440 12407 7442
rect 6012 7384 12346 7440
rect 12402 7384 12407 7440
rect 6012 7382 12407 7384
rect 6012 7380 6018 7382
rect 12341 7379 12407 7382
rect 3877 7306 3943 7309
rect 10174 7306 10180 7308
rect 3877 7304 10180 7306
rect 3877 7248 3882 7304
rect 3938 7248 10180 7304
rect 3877 7246 10180 7248
rect 3877 7243 3943 7246
rect 10174 7244 10180 7246
rect 10244 7244 10250 7308
rect 11329 7306 11395 7309
rect 12157 7306 12223 7309
rect 11329 7304 12223 7306
rect 11329 7248 11334 7304
rect 11390 7248 12162 7304
rect 12218 7248 12223 7304
rect 11329 7246 12223 7248
rect 11329 7243 11395 7246
rect 12157 7243 12223 7246
rect 7833 7170 7899 7173
rect 7008 7168 7899 7170
rect 7008 7112 7838 7168
rect 7894 7112 7899 7168
rect 7008 7110 7899 7112
rect 2820 7104 3136 7105
rect 2820 7040 2826 7104
rect 2890 7040 2906 7104
rect 2970 7040 2986 7104
rect 3050 7040 3066 7104
rect 3130 7040 3136 7104
rect 2820 7039 3136 7040
rect 6568 7104 6884 7105
rect 6568 7040 6574 7104
rect 6638 7040 6654 7104
rect 6718 7040 6734 7104
rect 6798 7040 6814 7104
rect 6878 7040 6884 7104
rect 6568 7039 6884 7040
rect 6126 6836 6132 6900
rect 6196 6898 6202 6900
rect 6361 6898 6427 6901
rect 6637 6898 6703 6901
rect 6196 6896 6703 6898
rect 6196 6840 6366 6896
rect 6422 6840 6642 6896
rect 6698 6840 6703 6896
rect 6196 6838 6703 6840
rect 6196 6836 6202 6838
rect 6361 6835 6427 6838
rect 6637 6835 6703 6838
rect 2221 6762 2287 6765
rect 7008 6762 7068 7110
rect 7833 7107 7899 7110
rect 8293 7170 8359 7173
rect 10133 7170 10199 7173
rect 8293 7168 10199 7170
rect 8293 7112 8298 7168
rect 8354 7112 10138 7168
rect 10194 7112 10199 7168
rect 8293 7110 10199 7112
rect 8293 7107 8359 7110
rect 10133 7107 10199 7110
rect 12157 7170 12223 7173
rect 12574 7170 12634 7518
rect 14549 7515 14615 7518
rect 12893 7444 12959 7445
rect 12893 7442 12940 7444
rect 12848 7440 12940 7442
rect 12848 7384 12898 7440
rect 12848 7382 12940 7384
rect 12893 7380 12940 7382
rect 13004 7380 13010 7444
rect 12893 7379 12959 7380
rect 14365 7306 14431 7309
rect 16021 7306 16087 7309
rect 14365 7304 16087 7306
rect 14365 7248 14370 7304
rect 14426 7248 16026 7304
rect 16082 7248 16087 7304
rect 14365 7246 16087 7248
rect 14365 7243 14431 7246
rect 16021 7243 16087 7246
rect 12157 7168 12634 7170
rect 12157 7112 12162 7168
rect 12218 7112 12634 7168
rect 12157 7110 12634 7112
rect 12157 7107 12223 7110
rect 10316 7104 10632 7105
rect 10316 7040 10322 7104
rect 10386 7040 10402 7104
rect 10466 7040 10482 7104
rect 10546 7040 10562 7104
rect 10626 7040 10632 7104
rect 10316 7039 10632 7040
rect 14064 7104 14380 7105
rect 14064 7040 14070 7104
rect 14134 7040 14150 7104
rect 14214 7040 14230 7104
rect 14294 7040 14310 7104
rect 14374 7040 14380 7104
rect 14064 7039 14380 7040
rect 7925 7034 7991 7037
rect 8385 7034 8451 7037
rect 7925 7032 8451 7034
rect 7925 6976 7930 7032
rect 7986 6976 8390 7032
rect 8446 6976 8451 7032
rect 7925 6974 8451 6976
rect 7925 6971 7991 6974
rect 8385 6971 8451 6974
rect 8937 7034 9003 7037
rect 9397 7034 9463 7037
rect 9857 7036 9923 7037
rect 9852 7034 9858 7036
rect 8937 7032 9463 7034
rect 8937 6976 8942 7032
rect 8998 6976 9402 7032
rect 9458 6976 9463 7032
rect 8937 6974 9463 6976
rect 9766 6974 9858 7034
rect 8937 6971 9003 6974
rect 9397 6971 9463 6974
rect 9852 6972 9858 6974
rect 9922 6972 9928 7036
rect 11329 7034 11395 7037
rect 12065 7036 12131 7037
rect 11646 7034 11652 7036
rect 11329 7032 11652 7034
rect 11329 6976 11334 7032
rect 11390 6976 11652 7032
rect 11329 6974 11652 6976
rect 9857 6971 9923 6972
rect 11329 6971 11395 6974
rect 11646 6972 11652 6974
rect 11716 6972 11722 7036
rect 12014 7034 12020 7036
rect 11974 6974 12020 7034
rect 12084 7032 12131 7036
rect 12126 6976 12131 7032
rect 12014 6972 12020 6974
rect 12084 6972 12131 6976
rect 12065 6971 12131 6972
rect 7373 6898 7439 6901
rect 11789 6898 11855 6901
rect 7373 6896 11855 6898
rect 7373 6840 7378 6896
rect 7434 6840 11794 6896
rect 11850 6840 11855 6896
rect 7373 6838 11855 6840
rect 7373 6835 7439 6838
rect 11789 6835 11855 6838
rect 2221 6760 7068 6762
rect 2221 6704 2226 6760
rect 2282 6704 7068 6760
rect 2221 6702 7068 6704
rect 7465 6762 7531 6765
rect 7598 6762 7604 6764
rect 7465 6760 7604 6762
rect 7465 6704 7470 6760
rect 7526 6704 7604 6760
rect 7465 6702 7604 6704
rect 2221 6699 2287 6702
rect 7465 6699 7531 6702
rect 7598 6700 7604 6702
rect 7668 6700 7674 6764
rect 7782 6700 7788 6764
rect 7852 6762 7858 6764
rect 9990 6762 9996 6764
rect 7852 6702 9996 6762
rect 7852 6700 7858 6702
rect 9990 6700 9996 6702
rect 10060 6700 10066 6764
rect 10133 6762 10199 6765
rect 11881 6762 11947 6765
rect 10133 6760 11947 6762
rect 10133 6704 10138 6760
rect 10194 6704 11886 6760
rect 11942 6704 11947 6760
rect 10133 6702 11947 6704
rect 10133 6699 10199 6702
rect 11881 6699 11947 6702
rect 13629 6762 13695 6765
rect 13813 6762 13879 6765
rect 14641 6762 14707 6765
rect 13629 6760 13738 6762
rect 13629 6704 13634 6760
rect 13690 6704 13738 6760
rect 13629 6699 13738 6704
rect 13813 6760 14707 6762
rect 13813 6704 13818 6760
rect 13874 6704 14646 6760
rect 14702 6704 14707 6760
rect 13813 6702 14707 6704
rect 13813 6699 13879 6702
rect 14641 6699 14707 6702
rect 0 6626 800 6656
rect 1485 6626 1551 6629
rect 0 6624 1551 6626
rect 0 6568 1490 6624
rect 1546 6568 1551 6624
rect 0 6566 1551 6568
rect 0 6536 800 6566
rect 1485 6563 1551 6566
rect 7230 6564 7236 6628
rect 7300 6626 7306 6628
rect 7741 6626 7807 6629
rect 7300 6624 7807 6626
rect 7300 6568 7746 6624
rect 7802 6568 7807 6624
rect 7300 6566 7807 6568
rect 7300 6564 7306 6566
rect 7741 6563 7807 6566
rect 9254 6564 9260 6628
rect 9324 6626 9330 6628
rect 9489 6626 9555 6629
rect 11237 6628 11303 6629
rect 11237 6626 11284 6628
rect 9324 6624 9555 6626
rect 9324 6568 9494 6624
rect 9550 6568 9555 6624
rect 9324 6566 9555 6568
rect 9324 6564 9330 6566
rect 9489 6563 9555 6566
rect 9630 6566 10656 6626
rect 11192 6624 11284 6626
rect 11348 6626 11354 6628
rect 11513 6626 11579 6629
rect 11348 6624 11579 6626
rect 11192 6568 11242 6624
rect 11348 6568 11518 6624
rect 11574 6568 11579 6624
rect 11192 6566 11284 6568
rect 4694 6560 5010 6561
rect 4694 6496 4700 6560
rect 4764 6496 4780 6560
rect 4844 6496 4860 6560
rect 4924 6496 4940 6560
rect 5004 6496 5010 6560
rect 4694 6495 5010 6496
rect 8442 6560 8758 6561
rect 8442 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8758 6560
rect 8442 6495 8758 6496
rect 3734 6428 3740 6492
rect 3804 6490 3810 6492
rect 4061 6490 4127 6493
rect 3804 6488 4127 6490
rect 3804 6432 4066 6488
rect 4122 6432 4127 6488
rect 3804 6430 4127 6432
rect 3804 6428 3810 6430
rect 4061 6427 4127 6430
rect 5165 6490 5231 6493
rect 7097 6490 7163 6493
rect 9630 6490 9690 6566
rect 5165 6488 7163 6490
rect 5165 6432 5170 6488
rect 5226 6432 7102 6488
rect 7158 6432 7163 6488
rect 5165 6430 7163 6432
rect 5165 6427 5231 6430
rect 7097 6427 7163 6430
rect 8894 6430 9690 6490
rect 3877 6354 3943 6357
rect 8894 6354 8954 6430
rect 3877 6352 8954 6354
rect 3877 6296 3882 6352
rect 3938 6296 8954 6352
rect 3877 6294 8954 6296
rect 10041 6354 10107 6357
rect 10225 6354 10291 6357
rect 10041 6352 10291 6354
rect 10041 6296 10046 6352
rect 10102 6296 10230 6352
rect 10286 6296 10291 6352
rect 10041 6294 10291 6296
rect 3877 6291 3943 6294
rect 10041 6291 10107 6294
rect 10225 6291 10291 6294
rect 4470 6156 4476 6220
rect 4540 6218 4546 6220
rect 8937 6218 9003 6221
rect 9121 6218 9187 6221
rect 4540 6158 8632 6218
rect 4540 6156 4546 6158
rect 7598 6020 7604 6084
rect 7668 6082 7674 6084
rect 8385 6082 8451 6085
rect 7668 6080 8451 6082
rect 7668 6024 8390 6080
rect 8446 6024 8451 6080
rect 7668 6022 8451 6024
rect 8572 6082 8632 6158
rect 8937 6216 9187 6218
rect 8937 6160 8942 6216
rect 8998 6160 9126 6216
rect 9182 6160 9187 6216
rect 8937 6158 9187 6160
rect 10596 6218 10656 6566
rect 11237 6564 11284 6566
rect 11348 6566 11579 6568
rect 11348 6564 11354 6566
rect 11237 6563 11303 6564
rect 11513 6563 11579 6566
rect 12190 6560 12506 6561
rect 12190 6496 12196 6560
rect 12260 6496 12276 6560
rect 12340 6496 12356 6560
rect 12420 6496 12436 6560
rect 12500 6496 12506 6560
rect 12190 6495 12506 6496
rect 13169 6492 13235 6493
rect 13118 6490 13124 6492
rect 13078 6430 13124 6490
rect 13188 6488 13235 6492
rect 13230 6432 13235 6488
rect 13118 6428 13124 6430
rect 13188 6428 13235 6432
rect 13169 6427 13235 6428
rect 11278 6292 11284 6356
rect 11348 6354 11354 6356
rect 12709 6354 12775 6357
rect 11348 6352 12775 6354
rect 11348 6296 12714 6352
rect 12770 6296 12775 6352
rect 11348 6294 12775 6296
rect 13678 6354 13738 6699
rect 14089 6626 14155 6629
rect 14089 6624 14704 6626
rect 14089 6568 14094 6624
rect 14150 6568 14704 6624
rect 14089 6566 14704 6568
rect 14089 6563 14155 6566
rect 14644 6493 14704 6566
rect 13854 6428 13860 6492
rect 13924 6490 13930 6492
rect 14089 6490 14155 6493
rect 13924 6488 14155 6490
rect 13924 6432 14094 6488
rect 14150 6432 14155 6488
rect 13924 6430 14155 6432
rect 13924 6428 13930 6430
rect 14089 6427 14155 6430
rect 14641 6490 14707 6493
rect 15929 6490 15995 6493
rect 14641 6488 15995 6490
rect 14641 6432 14646 6488
rect 14702 6432 15934 6488
rect 15990 6432 15995 6488
rect 14641 6430 15995 6432
rect 14641 6427 14707 6430
rect 15929 6427 15995 6430
rect 13813 6354 13879 6357
rect 13678 6352 13879 6354
rect 13678 6296 13818 6352
rect 13874 6296 13879 6352
rect 13678 6294 13879 6296
rect 11348 6292 11354 6294
rect 12709 6291 12775 6294
rect 13813 6291 13879 6294
rect 11329 6218 11395 6221
rect 12433 6218 12499 6221
rect 12617 6220 12683 6221
rect 10596 6158 10794 6218
rect 8937 6155 9003 6158
rect 9121 6155 9187 6158
rect 9254 6082 9260 6084
rect 8572 6022 9260 6082
rect 7668 6020 7674 6022
rect 8385 6019 8451 6022
rect 9254 6020 9260 6022
rect 9324 6020 9330 6084
rect 2820 6016 3136 6017
rect 2820 5952 2826 6016
rect 2890 5952 2906 6016
rect 2970 5952 2986 6016
rect 3050 5952 3066 6016
rect 3130 5952 3136 6016
rect 2820 5951 3136 5952
rect 6568 6016 6884 6017
rect 6568 5952 6574 6016
rect 6638 5952 6654 6016
rect 6718 5952 6734 6016
rect 6798 5952 6814 6016
rect 6878 5952 6884 6016
rect 6568 5951 6884 5952
rect 10316 6016 10632 6017
rect 10316 5952 10322 6016
rect 10386 5952 10402 6016
rect 10466 5952 10482 6016
rect 10546 5952 10562 6016
rect 10626 5952 10632 6016
rect 10316 5951 10632 5952
rect 3366 5884 3372 5948
rect 3436 5946 3442 5948
rect 5901 5946 5967 5949
rect 3436 5944 5967 5946
rect 3436 5888 5906 5944
rect 5962 5888 5967 5944
rect 3436 5886 5967 5888
rect 3436 5884 3442 5886
rect 2221 5810 2287 5813
rect 3374 5810 3434 5884
rect 5901 5883 5967 5886
rect 7097 5946 7163 5949
rect 9305 5946 9371 5949
rect 10041 5946 10107 5949
rect 7097 5944 9371 5946
rect 7097 5888 7102 5944
rect 7158 5888 9310 5944
rect 9366 5888 9371 5944
rect 7097 5886 9371 5888
rect 7097 5883 7163 5886
rect 9305 5883 9371 5886
rect 9446 5944 10107 5946
rect 9446 5888 10046 5944
rect 10102 5888 10107 5944
rect 9446 5886 10107 5888
rect 9446 5813 9506 5886
rect 10041 5883 10107 5886
rect 2221 5808 3434 5810
rect 2221 5752 2226 5808
rect 2282 5752 3434 5808
rect 2221 5750 3434 5752
rect 4337 5810 4403 5813
rect 8293 5810 8359 5813
rect 4337 5808 8359 5810
rect 4337 5752 4342 5808
rect 4398 5752 8298 5808
rect 8354 5752 8359 5808
rect 4337 5750 8359 5752
rect 2221 5747 2287 5750
rect 4337 5747 4403 5750
rect 8293 5747 8359 5750
rect 8480 5750 9092 5810
rect 0 5674 800 5704
rect 1485 5674 1551 5677
rect 0 5672 1551 5674
rect 0 5616 1490 5672
rect 1546 5616 1551 5672
rect 0 5614 1551 5616
rect 0 5584 800 5614
rect 1485 5611 1551 5614
rect 4981 5674 5047 5677
rect 5206 5674 5212 5676
rect 4981 5672 5212 5674
rect 4981 5616 4986 5672
rect 5042 5616 5212 5672
rect 4981 5614 5212 5616
rect 4981 5611 5047 5614
rect 5206 5612 5212 5614
rect 5276 5612 5282 5676
rect 5533 5674 5599 5677
rect 5533 5672 8310 5674
rect 5533 5616 5538 5672
rect 5594 5640 8310 5672
rect 8480 5640 8540 5750
rect 5594 5616 8540 5640
rect 5533 5614 8540 5616
rect 9032 5674 9092 5750
rect 9397 5808 9506 5813
rect 9397 5752 9402 5808
rect 9458 5752 9506 5808
rect 9397 5750 9506 5752
rect 9397 5747 9463 5750
rect 9622 5748 9628 5812
rect 9692 5810 9698 5812
rect 9765 5810 9831 5813
rect 9692 5808 9831 5810
rect 9692 5752 9770 5808
rect 9826 5752 9831 5808
rect 9692 5750 9831 5752
rect 9692 5748 9698 5750
rect 9765 5747 9831 5750
rect 10593 5810 10659 5813
rect 10734 5810 10794 6158
rect 11329 6216 12499 6218
rect 11329 6160 11334 6216
rect 11390 6160 12438 6216
rect 12494 6160 12499 6216
rect 11329 6158 12499 6160
rect 11329 6155 11395 6158
rect 12433 6155 12499 6158
rect 12566 6156 12572 6220
rect 12636 6218 12683 6220
rect 14273 6218 14339 6221
rect 12636 6216 12728 6218
rect 12678 6160 12728 6216
rect 12636 6158 12728 6160
rect 13862 6216 14339 6218
rect 13862 6160 14278 6216
rect 14334 6160 14339 6216
rect 13862 6158 14339 6160
rect 12636 6156 12683 6158
rect 12617 6155 12683 6156
rect 11881 6082 11947 6085
rect 13862 6082 13922 6158
rect 14273 6155 14339 6158
rect 11881 6080 13922 6082
rect 11881 6024 11886 6080
rect 11942 6024 13922 6080
rect 11881 6022 13922 6024
rect 14641 6082 14707 6085
rect 14774 6082 14780 6084
rect 14641 6080 14780 6082
rect 14641 6024 14646 6080
rect 14702 6024 14780 6080
rect 14641 6022 14780 6024
rect 11881 6019 11947 6022
rect 14641 6019 14707 6022
rect 14774 6020 14780 6022
rect 14844 6020 14850 6084
rect 14064 6016 14380 6017
rect 14064 5952 14070 6016
rect 14134 5952 14150 6016
rect 14214 5952 14230 6016
rect 14294 5952 14310 6016
rect 14374 5952 14380 6016
rect 14064 5951 14380 5952
rect 10961 5946 11027 5949
rect 11094 5946 11100 5948
rect 10961 5944 11100 5946
rect 10961 5888 10966 5944
rect 11022 5888 11100 5944
rect 10961 5886 11100 5888
rect 10961 5883 11027 5886
rect 11094 5884 11100 5886
rect 11164 5884 11170 5948
rect 13813 5946 13879 5949
rect 11516 5944 13879 5946
rect 11516 5888 13818 5944
rect 13874 5888 13879 5944
rect 11516 5886 13879 5888
rect 10593 5808 10794 5810
rect 10593 5752 10598 5808
rect 10654 5752 10794 5808
rect 10593 5750 10794 5752
rect 10593 5747 10659 5750
rect 11094 5748 11100 5812
rect 11164 5810 11170 5812
rect 11516 5810 11576 5886
rect 13813 5883 13879 5886
rect 12893 5810 12959 5813
rect 13537 5810 13603 5813
rect 11164 5750 11576 5810
rect 11654 5808 13603 5810
rect 11654 5752 12898 5808
rect 12954 5752 13542 5808
rect 13598 5752 13603 5808
rect 11654 5750 13603 5752
rect 11164 5748 11170 5750
rect 10685 5674 10751 5677
rect 9032 5672 10751 5674
rect 9032 5616 10690 5672
rect 10746 5616 10751 5672
rect 9032 5614 10751 5616
rect 5533 5611 5599 5614
rect 8250 5580 8540 5614
rect 10685 5611 10751 5614
rect 10961 5674 11027 5677
rect 11654 5674 11714 5750
rect 12893 5747 12959 5750
rect 13537 5747 13603 5750
rect 14181 5810 14247 5813
rect 16481 5810 16547 5813
rect 14181 5808 16547 5810
rect 14181 5752 14186 5808
rect 14242 5752 16486 5808
rect 16542 5752 16547 5808
rect 14181 5750 16547 5752
rect 14181 5747 14247 5750
rect 16481 5747 16547 5750
rect 10961 5672 11714 5674
rect 10961 5616 10966 5672
rect 11022 5616 11714 5672
rect 10961 5614 11714 5616
rect 11789 5672 11855 5677
rect 11789 5616 11794 5672
rect 11850 5616 11855 5672
rect 10961 5611 11027 5614
rect 11789 5611 11855 5616
rect 11973 5674 12039 5677
rect 12525 5674 12591 5677
rect 11973 5672 12591 5674
rect 11973 5616 11978 5672
rect 12034 5616 12530 5672
rect 12586 5616 12591 5672
rect 11973 5614 12591 5616
rect 11973 5611 12039 5614
rect 12525 5611 12591 5614
rect 13118 5612 13124 5676
rect 13188 5674 13194 5676
rect 13445 5674 13511 5677
rect 14089 5674 14155 5677
rect 13188 5672 14155 5674
rect 13188 5616 13450 5672
rect 13506 5616 14094 5672
rect 14150 5616 14155 5672
rect 13188 5614 14155 5616
rect 13188 5612 13194 5614
rect 13445 5611 13511 5614
rect 14089 5611 14155 5614
rect 5257 5538 5323 5541
rect 6126 5538 6132 5540
rect 5257 5536 6132 5538
rect 5257 5480 5262 5536
rect 5318 5480 6132 5536
rect 5257 5478 6132 5480
rect 5257 5475 5323 5478
rect 6126 5476 6132 5478
rect 6196 5476 6202 5540
rect 6913 5538 6979 5541
rect 7046 5538 7052 5540
rect 6913 5536 7052 5538
rect 6913 5480 6918 5536
rect 6974 5480 7052 5536
rect 6913 5478 7052 5480
rect 6913 5475 6979 5478
rect 7046 5476 7052 5478
rect 7116 5476 7122 5540
rect 8845 5536 8911 5541
rect 8845 5480 8850 5536
rect 8906 5480 8911 5536
rect 8845 5475 8911 5480
rect 9254 5476 9260 5540
rect 9324 5538 9330 5540
rect 9581 5538 9647 5541
rect 9324 5536 9647 5538
rect 9324 5480 9586 5536
rect 9642 5480 9647 5536
rect 9324 5478 9647 5480
rect 9324 5476 9330 5478
rect 9581 5475 9647 5478
rect 9765 5538 9831 5541
rect 11792 5538 11852 5611
rect 9765 5536 11852 5538
rect 9765 5480 9770 5536
rect 9826 5480 11852 5536
rect 9765 5478 11852 5480
rect 14365 5538 14431 5541
rect 14590 5538 14596 5540
rect 14365 5536 14596 5538
rect 14365 5480 14370 5536
rect 14426 5480 14596 5536
rect 14365 5478 14596 5480
rect 9765 5475 9831 5478
rect 14365 5475 14431 5478
rect 14590 5476 14596 5478
rect 14660 5538 14666 5540
rect 14917 5538 14983 5541
rect 14660 5536 14983 5538
rect 14660 5480 14922 5536
rect 14978 5480 14983 5536
rect 14660 5478 14983 5480
rect 14660 5476 14666 5478
rect 14917 5475 14983 5478
rect 4694 5472 5010 5473
rect 4694 5408 4700 5472
rect 4764 5408 4780 5472
rect 4844 5408 4860 5472
rect 4924 5408 4940 5472
rect 5004 5408 5010 5472
rect 4694 5407 5010 5408
rect 8442 5472 8758 5473
rect 8442 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8758 5472
rect 8442 5407 8758 5408
rect 5901 5402 5967 5405
rect 7782 5402 7788 5404
rect 5214 5400 7788 5402
rect 5214 5344 5906 5400
rect 5962 5344 7788 5400
rect 5214 5342 7788 5344
rect 3693 5266 3759 5269
rect 5214 5266 5274 5342
rect 5901 5339 5967 5342
rect 7782 5340 7788 5342
rect 7852 5340 7858 5404
rect 8848 5402 8908 5475
rect 12190 5472 12506 5473
rect 12190 5408 12196 5472
rect 12260 5408 12276 5472
rect 12340 5408 12356 5472
rect 12420 5408 12436 5472
rect 12500 5408 12506 5472
rect 12190 5407 12506 5408
rect 9397 5402 9463 5405
rect 8848 5400 9463 5402
rect 8848 5344 9402 5400
rect 9458 5344 9463 5400
rect 8848 5342 9463 5344
rect 9397 5339 9463 5342
rect 9581 5404 9647 5405
rect 9581 5400 9628 5404
rect 9692 5402 9698 5404
rect 10409 5402 10475 5405
rect 11421 5402 11487 5405
rect 9581 5344 9586 5400
rect 9581 5340 9628 5344
rect 9692 5342 9738 5402
rect 10409 5400 11487 5402
rect 10409 5344 10414 5400
rect 10470 5344 11426 5400
rect 11482 5344 11487 5400
rect 10409 5342 11487 5344
rect 9692 5340 9698 5342
rect 9581 5339 9647 5340
rect 10409 5339 10475 5342
rect 11421 5339 11487 5342
rect 12566 5340 12572 5404
rect 12636 5402 12642 5404
rect 13854 5402 13860 5404
rect 12636 5342 13860 5402
rect 12636 5340 12642 5342
rect 13854 5340 13860 5342
rect 13924 5402 13930 5404
rect 14089 5402 14155 5405
rect 13924 5400 14155 5402
rect 13924 5344 14094 5400
rect 14150 5344 14155 5400
rect 13924 5342 14155 5344
rect 13924 5340 13930 5342
rect 14089 5339 14155 5342
rect 15326 5340 15332 5404
rect 15396 5402 15402 5404
rect 15469 5402 15535 5405
rect 15396 5400 15535 5402
rect 15396 5344 15474 5400
rect 15530 5344 15535 5400
rect 15396 5342 15535 5344
rect 15396 5340 15402 5342
rect 15469 5339 15535 5342
rect 5441 5268 5507 5269
rect 5390 5266 5396 5268
rect 3693 5264 5274 5266
rect 3693 5208 3698 5264
rect 3754 5208 5274 5264
rect 3693 5206 5274 5208
rect 5350 5206 5396 5266
rect 5460 5264 5507 5268
rect 5502 5208 5507 5264
rect 3693 5203 3759 5206
rect 5390 5204 5396 5206
rect 5460 5204 5507 5208
rect 5441 5203 5507 5204
rect 6085 5266 6151 5269
rect 8477 5266 8543 5269
rect 9581 5266 9647 5269
rect 9806 5266 9812 5268
rect 6085 5264 8402 5266
rect 6085 5208 6090 5264
rect 6146 5208 8402 5264
rect 6085 5206 8402 5208
rect 6085 5203 6151 5206
rect 2221 5130 2287 5133
rect 8201 5130 8267 5133
rect 2221 5128 8267 5130
rect 2221 5072 2226 5128
rect 2282 5072 8206 5128
rect 8262 5072 8267 5128
rect 2221 5070 8267 5072
rect 8342 5130 8402 5206
rect 8477 5264 9506 5266
rect 8477 5208 8482 5264
rect 8538 5208 9506 5264
rect 8477 5206 9506 5208
rect 8477 5203 8543 5206
rect 9029 5130 9095 5133
rect 8342 5128 9095 5130
rect 8342 5072 9034 5128
rect 9090 5072 9095 5128
rect 8342 5070 9095 5072
rect 2221 5067 2287 5070
rect 8201 5067 8267 5070
rect 9029 5067 9095 5070
rect 9213 5128 9279 5133
rect 9213 5072 9218 5128
rect 9274 5072 9279 5128
rect 9213 5067 9279 5072
rect 9446 5130 9506 5206
rect 9581 5264 9812 5266
rect 9581 5208 9586 5264
rect 9642 5208 9812 5264
rect 9581 5206 9812 5208
rect 9581 5203 9647 5206
rect 9806 5204 9812 5206
rect 9876 5204 9882 5268
rect 10174 5204 10180 5268
rect 10244 5266 10250 5268
rect 10685 5266 10751 5269
rect 12893 5266 12959 5269
rect 13905 5268 13971 5269
rect 10244 5264 12959 5266
rect 10244 5208 10690 5264
rect 10746 5208 12898 5264
rect 12954 5208 12959 5264
rect 10244 5206 12959 5208
rect 10244 5204 10250 5206
rect 10685 5203 10751 5206
rect 12893 5203 12959 5206
rect 13854 5204 13860 5268
rect 13924 5266 13971 5268
rect 13924 5264 14016 5266
rect 13966 5208 14016 5264
rect 13924 5206 14016 5208
rect 13924 5204 13971 5206
rect 13905 5203 13971 5204
rect 12341 5130 12407 5133
rect 9446 5128 12407 5130
rect 9446 5072 12346 5128
rect 12402 5072 12407 5128
rect 9446 5070 12407 5072
rect 12341 5067 12407 5070
rect 4889 4994 4955 4997
rect 6085 4994 6151 4997
rect 4889 4992 6151 4994
rect 4889 4936 4894 4992
rect 4950 4936 6090 4992
rect 6146 4936 6151 4992
rect 4889 4934 6151 4936
rect 4889 4931 4955 4934
rect 6085 4931 6151 4934
rect 7189 4994 7255 4997
rect 8569 4994 8635 4997
rect 7189 4992 8635 4994
rect 7189 4936 7194 4992
rect 7250 4936 8574 4992
rect 8630 4936 8635 4992
rect 7189 4934 8635 4936
rect 7189 4931 7255 4934
rect 8569 4931 8635 4934
rect 2820 4928 3136 4929
rect 2820 4864 2826 4928
rect 2890 4864 2906 4928
rect 2970 4864 2986 4928
rect 3050 4864 3066 4928
rect 3130 4864 3136 4928
rect 2820 4863 3136 4864
rect 6568 4928 6884 4929
rect 6568 4864 6574 4928
rect 6638 4864 6654 4928
rect 6718 4864 6734 4928
rect 6798 4864 6814 4928
rect 6878 4864 6884 4928
rect 6568 4863 6884 4864
rect 2405 4860 2471 4861
rect 3693 4860 3759 4861
rect 2405 4858 2452 4860
rect 2360 4856 2452 4858
rect 2360 4800 2410 4856
rect 2360 4798 2452 4800
rect 2405 4796 2452 4798
rect 2516 4796 2522 4860
rect 3693 4856 3740 4860
rect 3804 4858 3810 4860
rect 3693 4800 3698 4856
rect 3693 4796 3740 4800
rect 3804 4798 3850 4858
rect 3804 4796 3810 4798
rect 3918 4796 3924 4860
rect 3988 4858 3994 4860
rect 4061 4858 4127 4861
rect 3988 4856 4127 4858
rect 3988 4800 4066 4856
rect 4122 4800 4127 4856
rect 3988 4798 4127 4800
rect 3988 4796 3994 4798
rect 2405 4795 2471 4796
rect 3693 4795 3759 4796
rect 4061 4795 4127 4798
rect 4429 4858 4495 4861
rect 6310 4858 6316 4860
rect 4429 4856 6316 4858
rect 4429 4800 4434 4856
rect 4490 4800 6316 4856
rect 4429 4798 6316 4800
rect 4429 4795 4495 4798
rect 6310 4796 6316 4798
rect 6380 4796 6386 4860
rect 0 4722 800 4752
rect 9216 4725 9276 5067
rect 11973 4994 12039 4997
rect 12985 4994 13051 4997
rect 11973 4992 13051 4994
rect 11973 4936 11978 4992
rect 12034 4936 12990 4992
rect 13046 4936 13051 4992
rect 11973 4934 13051 4936
rect 11973 4931 12039 4934
rect 12985 4931 13051 4934
rect 13353 4994 13419 4997
rect 13353 4992 13554 4994
rect 13353 4936 13358 4992
rect 13414 4936 13554 4992
rect 13353 4934 13554 4936
rect 13353 4931 13419 4934
rect 10316 4928 10632 4929
rect 10316 4864 10322 4928
rect 10386 4864 10402 4928
rect 10466 4864 10482 4928
rect 10546 4864 10562 4928
rect 10626 4864 10632 4928
rect 10316 4863 10632 4864
rect 9489 4858 9555 4861
rect 9622 4858 9628 4860
rect 9489 4856 9628 4858
rect 9489 4800 9494 4856
rect 9550 4800 9628 4856
rect 9489 4798 9628 4800
rect 9489 4795 9555 4798
rect 9622 4796 9628 4798
rect 9692 4796 9698 4860
rect 9765 4858 9831 4861
rect 9990 4858 9996 4860
rect 9765 4856 9996 4858
rect 9765 4800 9770 4856
rect 9826 4800 9996 4856
rect 9765 4798 9996 4800
rect 9765 4795 9831 4798
rect 9990 4796 9996 4798
rect 10060 4796 10066 4860
rect 12157 4858 12223 4861
rect 12985 4860 13051 4861
rect 12566 4858 12572 4860
rect 12157 4856 12572 4858
rect 12157 4800 12162 4856
rect 12218 4800 12572 4856
rect 12157 4798 12572 4800
rect 12157 4795 12223 4798
rect 12566 4796 12572 4798
rect 12636 4796 12642 4860
rect 12934 4796 12940 4860
rect 13004 4858 13051 4860
rect 13004 4856 13096 4858
rect 13046 4800 13096 4856
rect 13004 4798 13096 4800
rect 13004 4796 13051 4798
rect 12985 4795 13051 4796
rect 1485 4722 1551 4725
rect 0 4720 1551 4722
rect 0 4664 1490 4720
rect 1546 4664 1551 4720
rect 0 4662 1551 4664
rect 0 4632 800 4662
rect 1485 4659 1551 4662
rect 2313 4722 2379 4725
rect 8753 4722 8819 4725
rect 2313 4720 8819 4722
rect 2313 4664 2318 4720
rect 2374 4664 8758 4720
rect 8814 4664 8819 4720
rect 2313 4662 8819 4664
rect 2313 4659 2379 4662
rect 8753 4659 8819 4662
rect 9213 4720 9279 4725
rect 9213 4664 9218 4720
rect 9274 4664 9279 4720
rect 9213 4659 9279 4664
rect 9857 4722 9923 4725
rect 13353 4722 13419 4725
rect 9857 4720 13419 4722
rect 9857 4664 9862 4720
rect 9918 4664 13358 4720
rect 13414 4664 13419 4720
rect 9857 4662 13419 4664
rect 9857 4659 9923 4662
rect 13353 4659 13419 4662
rect 3785 4586 3851 4589
rect 4286 4586 4292 4588
rect 3785 4584 4292 4586
rect 3785 4528 3790 4584
rect 3846 4528 4292 4584
rect 3785 4526 4292 4528
rect 3785 4523 3851 4526
rect 4286 4524 4292 4526
rect 4356 4524 4362 4588
rect 4981 4586 5047 4589
rect 7281 4586 7347 4589
rect 9397 4586 9463 4589
rect 10593 4586 10659 4589
rect 13494 4586 13554 4934
rect 14064 4928 14380 4929
rect 14064 4864 14070 4928
rect 14134 4864 14150 4928
rect 14214 4864 14230 4928
rect 14294 4864 14310 4928
rect 14374 4864 14380 4928
rect 14064 4863 14380 4864
rect 4981 4584 8954 4586
rect 4981 4528 4986 4584
rect 5042 4528 7286 4584
rect 7342 4528 8954 4584
rect 4981 4526 8954 4528
rect 4981 4523 5047 4526
rect 7281 4523 7347 4526
rect 3325 4450 3391 4453
rect 4470 4450 4476 4452
rect 3325 4448 4476 4450
rect 3325 4392 3330 4448
rect 3386 4392 4476 4448
rect 3325 4390 4476 4392
rect 3325 4387 3391 4390
rect 4470 4388 4476 4390
rect 4540 4388 4546 4452
rect 6453 4450 6519 4453
rect 5444 4448 6519 4450
rect 5444 4392 6458 4448
rect 6514 4392 6519 4448
rect 5444 4390 6519 4392
rect 8894 4450 8954 4526
rect 9397 4584 10659 4586
rect 9397 4528 9402 4584
rect 9458 4528 10598 4584
rect 10654 4528 10659 4584
rect 9397 4526 10659 4528
rect 9397 4523 9463 4526
rect 10593 4523 10659 4526
rect 10780 4526 13554 4586
rect 10780 4450 10840 4526
rect 11278 4450 11284 4452
rect 8894 4390 10840 4450
rect 11056 4390 11284 4450
rect 4694 4384 5010 4385
rect 4694 4320 4700 4384
rect 4764 4320 4780 4384
rect 4844 4320 4860 4384
rect 4924 4320 4940 4384
rect 5004 4320 5010 4384
rect 4694 4319 5010 4320
rect 5444 4317 5504 4390
rect 6453 4387 6519 4390
rect 8442 4384 8758 4385
rect 8442 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8758 4384
rect 8442 4319 8758 4320
rect 3233 4314 3299 4317
rect 4061 4314 4127 4317
rect 3233 4312 4127 4314
rect 3233 4256 3238 4312
rect 3294 4256 4066 4312
rect 4122 4256 4127 4312
rect 3233 4254 4127 4256
rect 3233 4251 3299 4254
rect 4061 4251 4127 4254
rect 5441 4312 5507 4317
rect 7189 4314 7255 4317
rect 5441 4256 5446 4312
rect 5502 4256 5507 4312
rect 5441 4251 5507 4256
rect 5996 4312 7255 4314
rect 5996 4256 7194 4312
rect 7250 4256 7255 4312
rect 5996 4254 7255 4256
rect 2865 4178 2931 4181
rect 4153 4178 4219 4181
rect 2865 4176 4219 4178
rect 2865 4120 2870 4176
rect 2926 4120 4158 4176
rect 4214 4120 4219 4176
rect 2865 4118 4219 4120
rect 2865 4115 2931 4118
rect 4153 4115 4219 4118
rect 4613 4178 4679 4181
rect 5996 4178 6056 4254
rect 7189 4251 7255 4254
rect 7557 4314 7623 4317
rect 8937 4314 9003 4317
rect 9305 4314 9371 4317
rect 7557 4312 7988 4314
rect 7557 4256 7562 4312
rect 7618 4256 7988 4312
rect 7557 4254 7988 4256
rect 7557 4251 7623 4254
rect 6637 4178 6703 4181
rect 7465 4178 7531 4181
rect 7928 4178 7988 4254
rect 8937 4312 9371 4314
rect 8937 4256 8942 4312
rect 8998 4256 9310 4312
rect 9366 4256 9371 4312
rect 8937 4254 9371 4256
rect 8937 4251 9003 4254
rect 9305 4251 9371 4254
rect 9622 4252 9628 4316
rect 9692 4314 9698 4316
rect 9765 4314 9831 4317
rect 9692 4312 9831 4314
rect 9692 4256 9770 4312
rect 9826 4256 9831 4312
rect 9692 4254 9831 4256
rect 9692 4252 9698 4254
rect 9765 4251 9831 4254
rect 10317 4314 10383 4317
rect 10726 4314 10732 4316
rect 10317 4312 10732 4314
rect 10317 4256 10322 4312
rect 10378 4256 10732 4312
rect 10317 4254 10732 4256
rect 10317 4251 10383 4254
rect 10726 4252 10732 4254
rect 10796 4252 10802 4316
rect 11056 4181 11116 4390
rect 11278 4388 11284 4390
rect 11348 4388 11354 4452
rect 12566 4388 12572 4452
rect 12636 4450 12642 4452
rect 12893 4450 12959 4453
rect 12636 4448 12959 4450
rect 12636 4392 12898 4448
rect 12954 4392 12959 4448
rect 12636 4390 12959 4392
rect 12636 4388 12642 4390
rect 12893 4387 12959 4390
rect 13261 4450 13327 4453
rect 13670 4450 13676 4452
rect 13261 4448 13676 4450
rect 13261 4392 13266 4448
rect 13322 4392 13676 4448
rect 13261 4390 13676 4392
rect 13261 4387 13327 4390
rect 13670 4388 13676 4390
rect 13740 4388 13746 4452
rect 12190 4384 12506 4385
rect 12190 4320 12196 4384
rect 12260 4320 12276 4384
rect 12340 4320 12356 4384
rect 12420 4320 12436 4384
rect 12500 4320 12506 4384
rect 12190 4319 12506 4320
rect 11278 4252 11284 4316
rect 11348 4314 11354 4316
rect 11513 4314 11579 4317
rect 11348 4312 11579 4314
rect 11348 4256 11518 4312
rect 11574 4256 11579 4312
rect 11348 4254 11579 4256
rect 11348 4252 11354 4254
rect 11513 4251 11579 4254
rect 12709 4314 12775 4317
rect 14917 4314 14983 4317
rect 12709 4312 14983 4314
rect 12709 4256 12714 4312
rect 12770 4256 14922 4312
rect 14978 4256 14983 4312
rect 12709 4254 14983 4256
rect 12709 4251 12775 4254
rect 14917 4251 14983 4254
rect 8477 4178 8543 4181
rect 4613 4176 6056 4178
rect 4613 4120 4618 4176
rect 4674 4120 6056 4176
rect 4613 4118 6056 4120
rect 6134 4176 6703 4178
rect 6134 4120 6642 4176
rect 6698 4120 6703 4176
rect 6134 4118 6703 4120
rect 4613 4115 4679 4118
rect 1761 4044 1827 4045
rect 1710 4042 1716 4044
rect 1670 3982 1716 4042
rect 1780 4040 1827 4044
rect 1822 3984 1827 4040
rect 1710 3980 1716 3982
rect 1780 3980 1827 3984
rect 1761 3979 1827 3980
rect 3417 4042 3483 4045
rect 6134 4042 6194 4118
rect 6637 4115 6703 4118
rect 6870 4176 7850 4178
rect 6870 4120 7470 4176
rect 7526 4120 7850 4176
rect 6870 4118 7850 4120
rect 7928 4176 8543 4178
rect 7928 4120 8482 4176
rect 8538 4120 8543 4176
rect 7928 4118 8543 4120
rect 3417 4040 6194 4042
rect 3417 3984 3422 4040
rect 3478 3984 6194 4040
rect 3417 3982 6194 3984
rect 6545 4042 6611 4045
rect 6870 4042 6930 4118
rect 7465 4115 7531 4118
rect 7465 4044 7531 4045
rect 7414 4042 7420 4044
rect 6545 4040 6930 4042
rect 6545 3984 6550 4040
rect 6606 3984 6930 4040
rect 6545 3982 6930 3984
rect 7374 3982 7420 4042
rect 7484 4040 7531 4044
rect 7526 3984 7531 4040
rect 3417 3979 3483 3982
rect 6545 3979 6611 3982
rect 7414 3980 7420 3982
rect 7484 3980 7531 3984
rect 7790 4042 7850 4118
rect 8477 4115 8543 4118
rect 8661 4178 8727 4181
rect 11053 4178 11119 4181
rect 8661 4176 11119 4178
rect 8661 4120 8666 4176
rect 8722 4120 11058 4176
rect 11114 4120 11119 4176
rect 8661 4118 11119 4120
rect 8661 4115 8727 4118
rect 11053 4115 11119 4118
rect 11421 4178 11487 4181
rect 14641 4178 14707 4181
rect 11421 4176 14707 4178
rect 11421 4120 11426 4176
rect 11482 4120 14646 4176
rect 14702 4120 14707 4176
rect 11421 4118 14707 4120
rect 11421 4115 11487 4118
rect 14641 4115 14707 4118
rect 11329 4042 11395 4045
rect 7790 4040 11395 4042
rect 7790 3984 11334 4040
rect 11390 3984 11395 4040
rect 7790 3982 11395 3984
rect 7465 3979 7531 3980
rect 11329 3979 11395 3982
rect 11462 3980 11468 4044
rect 11532 4042 11538 4044
rect 11973 4042 12039 4045
rect 11532 4040 12039 4042
rect 11532 3984 11978 4040
rect 12034 3984 12039 4040
rect 11532 3982 12039 3984
rect 11532 3980 11538 3982
rect 11973 3979 12039 3982
rect 12249 4042 12315 4045
rect 13997 4042 14063 4045
rect 12249 4040 14063 4042
rect 12249 3984 12254 4040
rect 12310 3984 14002 4040
rect 14058 3984 14063 4040
rect 12249 3982 14063 3984
rect 12249 3979 12315 3982
rect 13997 3979 14063 3982
rect 6269 3906 6335 3909
rect 8017 3908 8083 3909
rect 3742 3904 6335 3906
rect 3742 3848 6274 3904
rect 6330 3848 6335 3904
rect 3742 3846 6335 3848
rect 2820 3840 3136 3841
rect 0 3770 800 3800
rect 2820 3776 2826 3840
rect 2890 3776 2906 3840
rect 2970 3776 2986 3840
rect 3050 3776 3066 3840
rect 3130 3776 3136 3840
rect 2820 3775 3136 3776
rect 1485 3770 1551 3773
rect 0 3768 1551 3770
rect 0 3712 1490 3768
rect 1546 3712 1551 3768
rect 0 3710 1551 3712
rect 0 3680 800 3710
rect 1485 3707 1551 3710
rect 2865 3634 2931 3637
rect 3366 3634 3372 3636
rect 2865 3632 3372 3634
rect 2865 3576 2870 3632
rect 2926 3576 3372 3632
rect 2865 3574 3372 3576
rect 2865 3571 2931 3574
rect 3366 3572 3372 3574
rect 3436 3572 3442 3636
rect 1945 3498 2011 3501
rect 3742 3498 3802 3846
rect 6269 3843 6335 3846
rect 7966 3844 7972 3908
rect 8036 3906 8083 3908
rect 8201 3906 8267 3909
rect 9121 3906 9187 3909
rect 8036 3904 8128 3906
rect 8078 3848 8128 3904
rect 8036 3846 8128 3848
rect 8201 3904 9187 3906
rect 8201 3848 8206 3904
rect 8262 3848 9126 3904
rect 9182 3848 9187 3904
rect 8201 3846 9187 3848
rect 8036 3844 8083 3846
rect 8017 3843 8083 3844
rect 8201 3843 8267 3846
rect 9121 3843 9187 3846
rect 10777 3906 10843 3909
rect 10910 3906 10916 3908
rect 10777 3904 10916 3906
rect 10777 3848 10782 3904
rect 10838 3848 10916 3904
rect 10777 3846 10916 3848
rect 10777 3843 10843 3846
rect 10910 3844 10916 3846
rect 10980 3844 10986 3908
rect 11053 3906 11119 3909
rect 11053 3904 13968 3906
rect 11053 3848 11058 3904
rect 11114 3848 13968 3904
rect 11053 3846 13968 3848
rect 11053 3843 11119 3846
rect 6568 3840 6884 3841
rect 6568 3776 6574 3840
rect 6638 3776 6654 3840
rect 6718 3776 6734 3840
rect 6798 3776 6814 3840
rect 6878 3776 6884 3840
rect 6568 3775 6884 3776
rect 10316 3840 10632 3841
rect 10316 3776 10322 3840
rect 10386 3776 10402 3840
rect 10466 3776 10482 3840
rect 10546 3776 10562 3840
rect 10626 3776 10632 3840
rect 10316 3775 10632 3776
rect 3969 3770 4035 3773
rect 6361 3770 6427 3773
rect 7373 3772 7439 3773
rect 7373 3770 7420 3772
rect 3969 3768 6427 3770
rect 3969 3712 3974 3768
rect 4030 3712 6366 3768
rect 6422 3712 6427 3768
rect 3969 3710 6427 3712
rect 7328 3768 7420 3770
rect 7328 3712 7378 3768
rect 7328 3710 7420 3712
rect 3969 3707 4035 3710
rect 6361 3707 6427 3710
rect 7373 3708 7420 3710
rect 7484 3708 7490 3772
rect 7649 3770 7715 3773
rect 10041 3770 10107 3773
rect 7649 3768 10107 3770
rect 7649 3712 7654 3768
rect 7710 3712 10046 3768
rect 10102 3712 10107 3768
rect 7649 3710 10107 3712
rect 7373 3707 7439 3708
rect 7649 3707 7715 3710
rect 10041 3707 10107 3710
rect 10777 3770 10843 3773
rect 12750 3770 12756 3772
rect 10777 3768 12756 3770
rect 10777 3712 10782 3768
rect 10838 3712 12756 3768
rect 10777 3710 12756 3712
rect 10777 3707 10843 3710
rect 12750 3708 12756 3710
rect 12820 3708 12826 3772
rect 6126 3572 6132 3636
rect 6196 3634 6202 3636
rect 6269 3634 6335 3637
rect 6637 3634 6703 3637
rect 6196 3632 6703 3634
rect 6196 3576 6274 3632
rect 6330 3576 6642 3632
rect 6698 3576 6703 3632
rect 6196 3574 6703 3576
rect 6196 3572 6202 3574
rect 6269 3571 6335 3574
rect 6637 3571 6703 3574
rect 6821 3634 6887 3637
rect 8150 3634 8156 3636
rect 6821 3632 8156 3634
rect 6821 3576 6826 3632
rect 6882 3576 8156 3632
rect 6821 3574 8156 3576
rect 6821 3571 6887 3574
rect 8150 3572 8156 3574
rect 8220 3572 8226 3636
rect 9213 3634 9279 3637
rect 9438 3634 9444 3636
rect 8296 3632 9444 3634
rect 8296 3576 9218 3632
rect 9274 3576 9444 3632
rect 8296 3574 9444 3576
rect 1945 3496 3802 3498
rect 1945 3440 1950 3496
rect 2006 3440 3802 3496
rect 1945 3438 3802 3440
rect 5809 3498 5875 3501
rect 7097 3498 7163 3501
rect 5809 3496 7163 3498
rect 5809 3440 5814 3496
rect 5870 3440 7102 3496
rect 7158 3440 7163 3496
rect 5809 3438 7163 3440
rect 1945 3435 2011 3438
rect 5809 3435 5875 3438
rect 7097 3435 7163 3438
rect 7281 3498 7347 3501
rect 7833 3498 7899 3501
rect 7281 3496 7899 3498
rect 7281 3440 7286 3496
rect 7342 3440 7838 3496
rect 7894 3440 7899 3496
rect 7281 3438 7899 3440
rect 7281 3435 7347 3438
rect 7833 3435 7899 3438
rect 5441 3362 5507 3365
rect 8109 3362 8175 3365
rect 5441 3360 8175 3362
rect 5441 3304 5446 3360
rect 5502 3304 8114 3360
rect 8170 3304 8175 3360
rect 5441 3302 8175 3304
rect 5441 3299 5507 3302
rect 8109 3299 8175 3302
rect 4694 3296 5010 3297
rect 4694 3232 4700 3296
rect 4764 3232 4780 3296
rect 4844 3232 4860 3296
rect 4924 3232 4940 3296
rect 5004 3232 5010 3296
rect 4694 3231 5010 3232
rect 5441 3226 5507 3229
rect 8296 3226 8356 3574
rect 9213 3571 9279 3574
rect 9438 3572 9444 3574
rect 9508 3572 9514 3636
rect 10409 3634 10475 3637
rect 11278 3634 11284 3636
rect 10409 3632 11284 3634
rect 10409 3576 10414 3632
rect 10470 3576 11284 3632
rect 10409 3574 11284 3576
rect 10409 3571 10475 3574
rect 11278 3572 11284 3574
rect 11348 3572 11354 3636
rect 12157 3634 12223 3637
rect 13908 3634 13968 3846
rect 14064 3840 14380 3841
rect 14064 3776 14070 3840
rect 14134 3776 14150 3840
rect 14214 3776 14230 3840
rect 14294 3776 14310 3840
rect 14374 3776 14380 3840
rect 14064 3775 14380 3776
rect 14089 3634 14155 3637
rect 16849 3634 16915 3637
rect 12157 3632 13002 3634
rect 12157 3576 12162 3632
rect 12218 3576 13002 3632
rect 12157 3574 13002 3576
rect 13908 3632 14155 3634
rect 13908 3576 14094 3632
rect 14150 3576 14155 3632
rect 13908 3574 14155 3576
rect 12157 3571 12223 3574
rect 8477 3498 8543 3501
rect 10961 3498 11027 3501
rect 8477 3496 11027 3498
rect 8477 3440 8482 3496
rect 8538 3440 10966 3496
rect 11022 3440 11027 3496
rect 8477 3438 11027 3440
rect 8477 3435 8543 3438
rect 10961 3435 11027 3438
rect 11646 3436 11652 3500
rect 11716 3498 11722 3500
rect 12801 3498 12867 3501
rect 11716 3496 12867 3498
rect 11716 3440 12806 3496
rect 12862 3440 12867 3496
rect 11716 3438 12867 3440
rect 12942 3498 13002 3574
rect 14089 3571 14155 3574
rect 14230 3632 16915 3634
rect 14230 3576 16854 3632
rect 16910 3576 16915 3632
rect 14230 3574 16915 3576
rect 14230 3498 14290 3574
rect 16849 3571 16915 3574
rect 12942 3438 14290 3498
rect 14457 3498 14523 3501
rect 14590 3498 14596 3500
rect 14457 3496 14596 3498
rect 14457 3440 14462 3496
rect 14518 3440 14596 3496
rect 14457 3438 14596 3440
rect 11716 3436 11722 3438
rect 12801 3435 12867 3438
rect 14457 3435 14523 3438
rect 14590 3436 14596 3438
rect 14660 3436 14666 3500
rect 12934 3300 12940 3364
rect 13004 3362 13010 3364
rect 13629 3362 13695 3365
rect 13004 3360 13695 3362
rect 13004 3304 13634 3360
rect 13690 3304 13695 3360
rect 13004 3302 13695 3304
rect 13004 3300 13010 3302
rect 13629 3299 13695 3302
rect 14549 3362 14615 3365
rect 14774 3362 14780 3364
rect 14549 3360 14780 3362
rect 14549 3304 14554 3360
rect 14610 3304 14780 3360
rect 14549 3302 14780 3304
rect 14549 3299 14615 3302
rect 14774 3300 14780 3302
rect 14844 3300 14850 3364
rect 15561 3362 15627 3365
rect 16400 3362 17200 3392
rect 15561 3360 17200 3362
rect 15561 3304 15566 3360
rect 15622 3304 17200 3360
rect 15561 3302 17200 3304
rect 15561 3299 15627 3302
rect 8442 3296 8758 3297
rect 8442 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8758 3296
rect 8442 3231 8758 3232
rect 12190 3296 12506 3297
rect 12190 3232 12196 3296
rect 12260 3232 12276 3296
rect 12340 3232 12356 3296
rect 12420 3232 12436 3296
rect 12500 3232 12506 3296
rect 16400 3272 17200 3302
rect 12190 3231 12506 3232
rect 5441 3224 8356 3226
rect 5441 3168 5446 3224
rect 5502 3168 8356 3224
rect 5441 3166 8356 3168
rect 5441 3163 5507 3166
rect 12750 3164 12756 3228
rect 12820 3226 12826 3228
rect 12893 3226 12959 3229
rect 12820 3224 15578 3226
rect 12820 3168 12898 3224
rect 12954 3168 15578 3224
rect 12820 3166 15578 3168
rect 12820 3164 12826 3166
rect 12893 3163 12959 3166
rect 6177 3090 6243 3093
rect 7281 3092 7347 3093
rect 6177 3088 7068 3090
rect 6177 3032 6182 3088
rect 6238 3032 7068 3088
rect 6177 3030 7068 3032
rect 6177 3027 6243 3030
rect 2313 2954 2379 2957
rect 6821 2954 6887 2957
rect 2313 2952 6887 2954
rect 2313 2896 2318 2952
rect 2374 2896 6826 2952
rect 6882 2896 6887 2952
rect 2313 2894 6887 2896
rect 2313 2891 2379 2894
rect 6821 2891 6887 2894
rect 0 2818 800 2848
rect 1485 2818 1551 2821
rect 0 2816 1551 2818
rect 0 2760 1490 2816
rect 1546 2760 1551 2816
rect 0 2758 1551 2760
rect 0 2728 800 2758
rect 1485 2755 1551 2758
rect 4337 2818 4403 2821
rect 5574 2818 5580 2820
rect 4337 2816 5580 2818
rect 4337 2760 4342 2816
rect 4398 2760 5580 2816
rect 4337 2758 5580 2760
rect 4337 2755 4403 2758
rect 5574 2756 5580 2758
rect 5644 2756 5650 2820
rect 7008 2818 7068 3030
rect 7230 3028 7236 3092
rect 7300 3090 7347 3092
rect 8109 3090 8175 3093
rect 9806 3090 9812 3092
rect 7300 3088 7392 3090
rect 7342 3032 7392 3088
rect 7300 3030 7392 3032
rect 8109 3088 9812 3090
rect 8109 3032 8114 3088
rect 8170 3032 9812 3088
rect 8109 3030 9812 3032
rect 7300 3028 7347 3030
rect 7281 3027 7347 3028
rect 8109 3027 8175 3030
rect 9806 3028 9812 3030
rect 9876 3090 9882 3092
rect 10501 3090 10567 3093
rect 9876 3088 10567 3090
rect 9876 3032 10506 3088
rect 10562 3032 10567 3088
rect 9876 3030 10567 3032
rect 9876 3028 9882 3030
rect 10501 3027 10567 3030
rect 10777 3090 10843 3093
rect 11789 3092 11855 3093
rect 11094 3090 11100 3092
rect 10777 3088 11100 3090
rect 10777 3032 10782 3088
rect 10838 3032 11100 3088
rect 10777 3030 11100 3032
rect 10777 3027 10843 3030
rect 11094 3028 11100 3030
rect 11164 3028 11170 3092
rect 11789 3088 11836 3092
rect 11900 3090 11906 3092
rect 11789 3032 11794 3088
rect 11789 3028 11836 3032
rect 11900 3030 11946 3090
rect 11900 3028 11906 3030
rect 12014 3028 12020 3092
rect 12084 3090 12090 3092
rect 12249 3090 12315 3093
rect 12084 3088 12315 3090
rect 12084 3032 12254 3088
rect 12310 3032 12315 3088
rect 12084 3030 12315 3032
rect 12084 3028 12090 3030
rect 11789 3027 11855 3028
rect 12249 3027 12315 3030
rect 13118 3028 13124 3092
rect 13188 3090 13194 3092
rect 13353 3090 13419 3093
rect 15326 3090 15332 3092
rect 13188 3088 13419 3090
rect 13188 3032 13358 3088
rect 13414 3032 13419 3088
rect 13188 3030 13419 3032
rect 13188 3028 13194 3030
rect 13353 3027 13419 3030
rect 13678 3030 15332 3090
rect 9397 2954 9463 2957
rect 13678 2954 13738 3030
rect 15326 3028 15332 3030
rect 15396 3028 15402 3092
rect 15518 3090 15578 3166
rect 16665 3090 16731 3093
rect 15518 3088 16731 3090
rect 15518 3032 16670 3088
rect 16726 3032 16731 3088
rect 15518 3030 16731 3032
rect 16665 3027 16731 3030
rect 9397 2952 13738 2954
rect 9397 2896 9402 2952
rect 9458 2896 13738 2952
rect 9397 2894 13738 2896
rect 9397 2891 9463 2894
rect 11329 2818 11395 2821
rect 13905 2820 13971 2821
rect 12566 2818 12572 2820
rect 7008 2758 10242 2818
rect 2820 2752 3136 2753
rect 2820 2688 2826 2752
rect 2890 2688 2906 2752
rect 2970 2688 2986 2752
rect 3050 2688 3066 2752
rect 3130 2688 3136 2752
rect 2820 2687 3136 2688
rect 6568 2752 6884 2753
rect 6568 2688 6574 2752
rect 6638 2688 6654 2752
rect 6718 2688 6734 2752
rect 6798 2688 6814 2752
rect 6878 2688 6884 2752
rect 6568 2687 6884 2688
rect 5809 2682 5875 2685
rect 5942 2682 5948 2684
rect 5809 2680 5948 2682
rect 5809 2624 5814 2680
rect 5870 2624 5948 2680
rect 5809 2622 5948 2624
rect 5809 2619 5875 2622
rect 5942 2620 5948 2622
rect 6012 2620 6018 2684
rect 7046 2620 7052 2684
rect 7116 2682 7122 2684
rect 7189 2682 7255 2685
rect 7116 2680 7255 2682
rect 7116 2624 7194 2680
rect 7250 2624 7255 2680
rect 7116 2622 7255 2624
rect 7116 2620 7122 2622
rect 7189 2619 7255 2622
rect 7373 2684 7439 2685
rect 7373 2680 7420 2684
rect 7484 2682 7490 2684
rect 7373 2624 7378 2680
rect 7373 2620 7420 2624
rect 7484 2622 7530 2682
rect 7484 2620 7490 2622
rect 7373 2619 7439 2620
rect 4889 2546 4955 2549
rect 5206 2546 5212 2548
rect 4889 2544 5212 2546
rect 4889 2488 4894 2544
rect 4950 2488 5212 2544
rect 4889 2486 5212 2488
rect 4889 2483 4955 2486
rect 5206 2484 5212 2486
rect 5276 2546 5282 2548
rect 5533 2546 5599 2549
rect 5276 2544 5599 2546
rect 5276 2488 5538 2544
rect 5594 2488 5599 2544
rect 5276 2486 5599 2488
rect 5276 2484 5282 2486
rect 5533 2483 5599 2486
rect 5942 2484 5948 2548
rect 6012 2546 6018 2548
rect 7465 2546 7531 2549
rect 6012 2544 7531 2546
rect 6012 2488 7470 2544
rect 7526 2488 7531 2544
rect 6012 2486 7531 2488
rect 6012 2484 6018 2486
rect 7465 2483 7531 2486
rect 8293 2546 8359 2549
rect 8845 2548 8911 2549
rect 8845 2546 8892 2548
rect 8293 2544 8892 2546
rect 8293 2488 8298 2544
rect 8354 2488 8850 2544
rect 8293 2486 8892 2488
rect 8293 2483 8359 2486
rect 8845 2484 8892 2486
rect 8956 2484 8962 2548
rect 10182 2546 10242 2758
rect 11329 2816 12572 2818
rect 11329 2760 11334 2816
rect 11390 2760 12572 2816
rect 11329 2758 12572 2760
rect 11329 2755 11395 2758
rect 12566 2756 12572 2758
rect 12636 2756 12642 2820
rect 13854 2818 13860 2820
rect 13814 2758 13860 2818
rect 13924 2816 13971 2820
rect 13966 2760 13971 2816
rect 13854 2756 13860 2758
rect 13924 2756 13971 2760
rect 13905 2755 13971 2756
rect 10316 2752 10632 2753
rect 10316 2688 10322 2752
rect 10386 2688 10402 2752
rect 10466 2688 10482 2752
rect 10546 2688 10562 2752
rect 10626 2688 10632 2752
rect 10316 2687 10632 2688
rect 14064 2752 14380 2753
rect 14064 2688 14070 2752
rect 14134 2688 14150 2752
rect 14214 2688 14230 2752
rect 14294 2688 14310 2752
rect 14374 2688 14380 2752
rect 14064 2687 14380 2688
rect 11421 2682 11487 2685
rect 13537 2682 13603 2685
rect 11421 2680 13603 2682
rect 11421 2624 11426 2680
rect 11482 2624 13542 2680
rect 13598 2624 13603 2680
rect 11421 2622 13603 2624
rect 11421 2619 11487 2622
rect 13537 2619 13603 2622
rect 13261 2546 13327 2549
rect 10182 2544 13327 2546
rect 10182 2488 13266 2544
rect 13322 2488 13327 2544
rect 10182 2486 13327 2488
rect 8845 2483 8911 2484
rect 13261 2483 13327 2486
rect 13486 2484 13492 2548
rect 13556 2546 13562 2548
rect 14365 2546 14431 2549
rect 13556 2544 14431 2546
rect 13556 2488 14370 2544
rect 14426 2488 14431 2544
rect 13556 2486 14431 2488
rect 13556 2484 13562 2486
rect 14365 2483 14431 2486
rect 4286 2348 4292 2412
rect 4356 2410 4362 2412
rect 7005 2410 7071 2413
rect 10777 2410 10843 2413
rect 14590 2410 14596 2412
rect 4356 2350 6930 2410
rect 4356 2348 4362 2350
rect 6870 2274 6930 2350
rect 7005 2408 10843 2410
rect 7005 2352 7010 2408
rect 7066 2352 10782 2408
rect 10838 2352 10843 2408
rect 7005 2350 10843 2352
rect 7005 2347 7071 2350
rect 10777 2347 10843 2350
rect 12068 2350 14596 2410
rect 7465 2274 7531 2277
rect 6870 2272 7531 2274
rect 6870 2216 7470 2272
rect 7526 2216 7531 2272
rect 6870 2214 7531 2216
rect 7465 2211 7531 2214
rect 9121 2274 9187 2277
rect 12068 2274 12128 2350
rect 14590 2348 14596 2350
rect 14660 2348 14666 2412
rect 9121 2272 12128 2274
rect 9121 2216 9126 2272
rect 9182 2216 12128 2272
rect 9121 2214 12128 2216
rect 9121 2211 9187 2214
rect 13670 2212 13676 2276
rect 13740 2274 13746 2276
rect 13813 2274 13879 2277
rect 13740 2272 13879 2274
rect 13740 2216 13818 2272
rect 13874 2216 13879 2272
rect 13740 2214 13879 2216
rect 13740 2212 13746 2214
rect 13813 2211 13879 2214
rect 4694 2208 5010 2209
rect 4694 2144 4700 2208
rect 4764 2144 4780 2208
rect 4844 2144 4860 2208
rect 4924 2144 4940 2208
rect 5004 2144 5010 2208
rect 4694 2143 5010 2144
rect 8442 2208 8758 2209
rect 8442 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8758 2208
rect 8442 2143 8758 2144
rect 12190 2208 12506 2209
rect 12190 2144 12196 2208
rect 12260 2144 12276 2208
rect 12340 2144 12356 2208
rect 12420 2144 12436 2208
rect 12500 2144 12506 2208
rect 12190 2143 12506 2144
rect 7741 2138 7807 2141
rect 8109 2138 8175 2141
rect 6180 2136 8175 2138
rect 6180 2080 7746 2136
rect 7802 2080 8114 2136
rect 8170 2080 8175 2136
rect 6180 2078 8175 2080
rect 2405 2002 2471 2005
rect 2405 2000 2790 2002
rect 2405 1944 2410 2000
rect 2466 1944 2790 2000
rect 2405 1942 2790 1944
rect 2405 1939 2471 1942
rect 0 1866 800 1896
rect 1853 1866 1919 1869
rect 0 1864 1919 1866
rect 0 1808 1858 1864
rect 1914 1808 1919 1864
rect 0 1806 1919 1808
rect 0 1776 800 1806
rect 1853 1803 1919 1806
rect 2730 1458 2790 1942
rect 3918 1940 3924 2004
rect 3988 2002 3994 2004
rect 6180 2002 6240 2078
rect 7741 2075 7807 2078
rect 8109 2075 8175 2078
rect 3988 1942 6240 2002
rect 6361 2002 6427 2005
rect 9254 2002 9260 2004
rect 6361 2000 9260 2002
rect 6361 1944 6366 2000
rect 6422 1944 9260 2000
rect 6361 1942 9260 1944
rect 3988 1940 3994 1942
rect 6361 1939 6427 1942
rect 9254 1940 9260 1942
rect 9324 1940 9330 2004
rect 3601 1866 3667 1869
rect 6085 1866 6151 1869
rect 9857 1866 9923 1869
rect 14641 1866 14707 1869
rect 3601 1864 9923 1866
rect 3601 1808 3606 1864
rect 3662 1808 6090 1864
rect 6146 1808 9862 1864
rect 9918 1808 9923 1864
rect 3601 1806 9923 1808
rect 3601 1803 3667 1806
rect 6085 1803 6151 1806
rect 9857 1803 9923 1806
rect 12390 1864 14707 1866
rect 12390 1808 14646 1864
rect 14702 1808 14707 1864
rect 12390 1806 14707 1808
rect 3877 1730 3943 1733
rect 10685 1730 10751 1733
rect 3877 1728 10751 1730
rect 3877 1672 3882 1728
rect 3938 1672 10690 1728
rect 10746 1672 10751 1728
rect 3877 1670 10751 1672
rect 3877 1667 3943 1670
rect 10685 1667 10751 1670
rect 5349 1594 5415 1597
rect 12390 1594 12450 1806
rect 14641 1803 14707 1806
rect 5349 1592 12450 1594
rect 5349 1536 5354 1592
rect 5410 1536 12450 1592
rect 5349 1534 12450 1536
rect 5349 1531 5415 1534
rect 11513 1458 11579 1461
rect 2730 1456 11579 1458
rect 2730 1400 11518 1456
rect 11574 1400 11579 1456
rect 2730 1398 11579 1400
rect 11513 1395 11579 1398
rect 0 914 800 944
rect 1393 914 1459 917
rect 0 912 1459 914
rect 0 856 1398 912
rect 1454 856 1459 912
rect 0 854 1459 856
rect 0 824 800 854
rect 1393 851 1459 854
<< via3 >>
rect 4700 17436 4764 17440
rect 4700 17380 4704 17436
rect 4704 17380 4760 17436
rect 4760 17380 4764 17436
rect 4700 17376 4764 17380
rect 4780 17436 4844 17440
rect 4780 17380 4784 17436
rect 4784 17380 4840 17436
rect 4840 17380 4844 17436
rect 4780 17376 4844 17380
rect 4860 17436 4924 17440
rect 4860 17380 4864 17436
rect 4864 17380 4920 17436
rect 4920 17380 4924 17436
rect 4860 17376 4924 17380
rect 4940 17436 5004 17440
rect 4940 17380 4944 17436
rect 4944 17380 5000 17436
rect 5000 17380 5004 17436
rect 4940 17376 5004 17380
rect 8448 17436 8512 17440
rect 8448 17380 8452 17436
rect 8452 17380 8508 17436
rect 8508 17380 8512 17436
rect 8448 17376 8512 17380
rect 8528 17436 8592 17440
rect 8528 17380 8532 17436
rect 8532 17380 8588 17436
rect 8588 17380 8592 17436
rect 8528 17376 8592 17380
rect 8608 17436 8672 17440
rect 8608 17380 8612 17436
rect 8612 17380 8668 17436
rect 8668 17380 8672 17436
rect 8608 17376 8672 17380
rect 8688 17436 8752 17440
rect 8688 17380 8692 17436
rect 8692 17380 8748 17436
rect 8748 17380 8752 17436
rect 8688 17376 8752 17380
rect 12196 17436 12260 17440
rect 12196 17380 12200 17436
rect 12200 17380 12256 17436
rect 12256 17380 12260 17436
rect 12196 17376 12260 17380
rect 12276 17436 12340 17440
rect 12276 17380 12280 17436
rect 12280 17380 12336 17436
rect 12336 17380 12340 17436
rect 12276 17376 12340 17380
rect 12356 17436 12420 17440
rect 12356 17380 12360 17436
rect 12360 17380 12416 17436
rect 12416 17380 12420 17436
rect 12356 17376 12420 17380
rect 12436 17436 12500 17440
rect 12436 17380 12440 17436
rect 12440 17380 12496 17436
rect 12496 17380 12500 17436
rect 12436 17376 12500 17380
rect 11468 17172 11532 17236
rect 2826 16892 2890 16896
rect 2826 16836 2830 16892
rect 2830 16836 2886 16892
rect 2886 16836 2890 16892
rect 2826 16832 2890 16836
rect 2906 16892 2970 16896
rect 2906 16836 2910 16892
rect 2910 16836 2966 16892
rect 2966 16836 2970 16892
rect 2906 16832 2970 16836
rect 2986 16892 3050 16896
rect 2986 16836 2990 16892
rect 2990 16836 3046 16892
rect 3046 16836 3050 16892
rect 2986 16832 3050 16836
rect 3066 16892 3130 16896
rect 3066 16836 3070 16892
rect 3070 16836 3126 16892
rect 3126 16836 3130 16892
rect 3066 16832 3130 16836
rect 6574 16892 6638 16896
rect 6574 16836 6578 16892
rect 6578 16836 6634 16892
rect 6634 16836 6638 16892
rect 6574 16832 6638 16836
rect 6654 16892 6718 16896
rect 6654 16836 6658 16892
rect 6658 16836 6714 16892
rect 6714 16836 6718 16892
rect 6654 16832 6718 16836
rect 6734 16892 6798 16896
rect 6734 16836 6738 16892
rect 6738 16836 6794 16892
rect 6794 16836 6798 16892
rect 6734 16832 6798 16836
rect 6814 16892 6878 16896
rect 6814 16836 6818 16892
rect 6818 16836 6874 16892
rect 6874 16836 6878 16892
rect 6814 16832 6878 16836
rect 10322 16892 10386 16896
rect 10322 16836 10326 16892
rect 10326 16836 10382 16892
rect 10382 16836 10386 16892
rect 10322 16832 10386 16836
rect 10402 16892 10466 16896
rect 10402 16836 10406 16892
rect 10406 16836 10462 16892
rect 10462 16836 10466 16892
rect 10402 16832 10466 16836
rect 10482 16892 10546 16896
rect 10482 16836 10486 16892
rect 10486 16836 10542 16892
rect 10542 16836 10546 16892
rect 10482 16832 10546 16836
rect 10562 16892 10626 16896
rect 10562 16836 10566 16892
rect 10566 16836 10622 16892
rect 10622 16836 10626 16892
rect 10562 16832 10626 16836
rect 14070 16892 14134 16896
rect 14070 16836 14074 16892
rect 14074 16836 14130 16892
rect 14130 16836 14134 16892
rect 14070 16832 14134 16836
rect 14150 16892 14214 16896
rect 14150 16836 14154 16892
rect 14154 16836 14210 16892
rect 14210 16836 14214 16892
rect 14150 16832 14214 16836
rect 14230 16892 14294 16896
rect 14230 16836 14234 16892
rect 14234 16836 14290 16892
rect 14290 16836 14294 16892
rect 14230 16832 14294 16836
rect 14310 16892 14374 16896
rect 14310 16836 14314 16892
rect 14314 16836 14370 16892
rect 14370 16836 14374 16892
rect 14310 16832 14374 16836
rect 13676 16764 13740 16828
rect 9812 16628 9876 16692
rect 13492 16628 13556 16692
rect 12756 16492 12820 16556
rect 4700 16348 4764 16352
rect 4700 16292 4704 16348
rect 4704 16292 4760 16348
rect 4760 16292 4764 16348
rect 4700 16288 4764 16292
rect 4780 16348 4844 16352
rect 4780 16292 4784 16348
rect 4784 16292 4840 16348
rect 4840 16292 4844 16348
rect 4780 16288 4844 16292
rect 4860 16348 4924 16352
rect 4860 16292 4864 16348
rect 4864 16292 4920 16348
rect 4920 16292 4924 16348
rect 4860 16288 4924 16292
rect 4940 16348 5004 16352
rect 4940 16292 4944 16348
rect 4944 16292 5000 16348
rect 5000 16292 5004 16348
rect 4940 16288 5004 16292
rect 8448 16348 8512 16352
rect 8448 16292 8452 16348
rect 8452 16292 8508 16348
rect 8508 16292 8512 16348
rect 8448 16288 8512 16292
rect 8528 16348 8592 16352
rect 8528 16292 8532 16348
rect 8532 16292 8588 16348
rect 8588 16292 8592 16348
rect 8528 16288 8592 16292
rect 8608 16348 8672 16352
rect 8608 16292 8612 16348
rect 8612 16292 8668 16348
rect 8668 16292 8672 16348
rect 8608 16288 8672 16292
rect 8688 16348 8752 16352
rect 8688 16292 8692 16348
rect 8692 16292 8748 16348
rect 8748 16292 8752 16348
rect 8688 16288 8752 16292
rect 12196 16348 12260 16352
rect 12196 16292 12200 16348
rect 12200 16292 12256 16348
rect 12256 16292 12260 16348
rect 12196 16288 12260 16292
rect 12276 16348 12340 16352
rect 12276 16292 12280 16348
rect 12280 16292 12336 16348
rect 12336 16292 12340 16348
rect 12276 16288 12340 16292
rect 12356 16348 12420 16352
rect 12356 16292 12360 16348
rect 12360 16292 12416 16348
rect 12416 16292 12420 16348
rect 12356 16288 12420 16292
rect 12436 16348 12500 16352
rect 12436 16292 12440 16348
rect 12440 16292 12496 16348
rect 12496 16292 12500 16348
rect 12436 16288 12500 16292
rect 14596 16220 14660 16284
rect 13308 16008 13372 16012
rect 13308 15952 13322 16008
rect 13322 15952 13372 16008
rect 13308 15948 13372 15952
rect 13860 15948 13924 16012
rect 2826 15804 2890 15808
rect 2826 15748 2830 15804
rect 2830 15748 2886 15804
rect 2886 15748 2890 15804
rect 2826 15744 2890 15748
rect 2906 15804 2970 15808
rect 2906 15748 2910 15804
rect 2910 15748 2966 15804
rect 2966 15748 2970 15804
rect 2906 15744 2970 15748
rect 2986 15804 3050 15808
rect 2986 15748 2990 15804
rect 2990 15748 3046 15804
rect 3046 15748 3050 15804
rect 2986 15744 3050 15748
rect 3066 15804 3130 15808
rect 3066 15748 3070 15804
rect 3070 15748 3126 15804
rect 3126 15748 3130 15804
rect 3066 15744 3130 15748
rect 6574 15804 6638 15808
rect 6574 15748 6578 15804
rect 6578 15748 6634 15804
rect 6634 15748 6638 15804
rect 6574 15744 6638 15748
rect 6654 15804 6718 15808
rect 6654 15748 6658 15804
rect 6658 15748 6714 15804
rect 6714 15748 6718 15804
rect 6654 15744 6718 15748
rect 6734 15804 6798 15808
rect 6734 15748 6738 15804
rect 6738 15748 6794 15804
rect 6794 15748 6798 15804
rect 6734 15744 6798 15748
rect 6814 15804 6878 15808
rect 6814 15748 6818 15804
rect 6818 15748 6874 15804
rect 6874 15748 6878 15804
rect 6814 15744 6878 15748
rect 10322 15804 10386 15808
rect 10322 15748 10326 15804
rect 10326 15748 10382 15804
rect 10382 15748 10386 15804
rect 10322 15744 10386 15748
rect 10402 15804 10466 15808
rect 10402 15748 10406 15804
rect 10406 15748 10462 15804
rect 10462 15748 10466 15804
rect 10402 15744 10466 15748
rect 10482 15804 10546 15808
rect 10482 15748 10486 15804
rect 10486 15748 10542 15804
rect 10542 15748 10546 15804
rect 10482 15744 10546 15748
rect 10562 15804 10626 15808
rect 10562 15748 10566 15804
rect 10566 15748 10622 15804
rect 10622 15748 10626 15804
rect 10562 15744 10626 15748
rect 14070 15804 14134 15808
rect 14070 15748 14074 15804
rect 14074 15748 14130 15804
rect 14130 15748 14134 15804
rect 14070 15744 14134 15748
rect 14150 15804 14214 15808
rect 14150 15748 14154 15804
rect 14154 15748 14210 15804
rect 14210 15748 14214 15804
rect 14150 15744 14214 15748
rect 14230 15804 14294 15808
rect 14230 15748 14234 15804
rect 14234 15748 14290 15804
rect 14290 15748 14294 15804
rect 14230 15744 14294 15748
rect 14310 15804 14374 15808
rect 14310 15748 14314 15804
rect 14314 15748 14370 15804
rect 14370 15748 14374 15804
rect 14310 15744 14374 15748
rect 1716 15268 1780 15332
rect 2452 15328 2516 15332
rect 2452 15272 2466 15328
rect 2466 15272 2516 15328
rect 2452 15268 2516 15272
rect 6316 15268 6380 15332
rect 4700 15260 4764 15264
rect 4700 15204 4704 15260
rect 4704 15204 4760 15260
rect 4760 15204 4764 15260
rect 4700 15200 4764 15204
rect 4780 15260 4844 15264
rect 4780 15204 4784 15260
rect 4784 15204 4840 15260
rect 4840 15204 4844 15260
rect 4780 15200 4844 15204
rect 4860 15260 4924 15264
rect 4860 15204 4864 15260
rect 4864 15204 4920 15260
rect 4920 15204 4924 15260
rect 4860 15200 4924 15204
rect 4940 15260 5004 15264
rect 4940 15204 4944 15260
rect 4944 15204 5000 15260
rect 5000 15204 5004 15260
rect 4940 15200 5004 15204
rect 8448 15260 8512 15264
rect 8448 15204 8452 15260
rect 8452 15204 8508 15260
rect 8508 15204 8512 15260
rect 8448 15200 8512 15204
rect 8528 15260 8592 15264
rect 8528 15204 8532 15260
rect 8532 15204 8588 15260
rect 8588 15204 8592 15260
rect 8528 15200 8592 15204
rect 8608 15260 8672 15264
rect 8608 15204 8612 15260
rect 8612 15204 8668 15260
rect 8668 15204 8672 15260
rect 8608 15200 8672 15204
rect 8688 15260 8752 15264
rect 8688 15204 8692 15260
rect 8692 15204 8748 15260
rect 8748 15204 8752 15260
rect 8688 15200 8752 15204
rect 15332 15268 15396 15332
rect 12196 15260 12260 15264
rect 12196 15204 12200 15260
rect 12200 15204 12256 15260
rect 12256 15204 12260 15260
rect 12196 15200 12260 15204
rect 12276 15260 12340 15264
rect 12276 15204 12280 15260
rect 12280 15204 12336 15260
rect 12336 15204 12340 15260
rect 12276 15200 12340 15204
rect 12356 15260 12420 15264
rect 12356 15204 12360 15260
rect 12360 15204 12416 15260
rect 12416 15204 12420 15260
rect 12356 15200 12420 15204
rect 12436 15260 12500 15264
rect 12436 15204 12440 15260
rect 12440 15204 12496 15260
rect 12496 15204 12500 15260
rect 12436 15200 12500 15204
rect 12020 14860 12084 14924
rect 2826 14716 2890 14720
rect 2826 14660 2830 14716
rect 2830 14660 2886 14716
rect 2886 14660 2890 14716
rect 2826 14656 2890 14660
rect 2906 14716 2970 14720
rect 2906 14660 2910 14716
rect 2910 14660 2966 14716
rect 2966 14660 2970 14716
rect 2906 14656 2970 14660
rect 2986 14716 3050 14720
rect 2986 14660 2990 14716
rect 2990 14660 3046 14716
rect 3046 14660 3050 14716
rect 2986 14656 3050 14660
rect 3066 14716 3130 14720
rect 3066 14660 3070 14716
rect 3070 14660 3126 14716
rect 3126 14660 3130 14716
rect 3066 14656 3130 14660
rect 6574 14716 6638 14720
rect 6574 14660 6578 14716
rect 6578 14660 6634 14716
rect 6634 14660 6638 14716
rect 6574 14656 6638 14660
rect 6654 14716 6718 14720
rect 6654 14660 6658 14716
rect 6658 14660 6714 14716
rect 6714 14660 6718 14716
rect 6654 14656 6718 14660
rect 6734 14716 6798 14720
rect 6734 14660 6738 14716
rect 6738 14660 6794 14716
rect 6794 14660 6798 14716
rect 6734 14656 6798 14660
rect 6814 14716 6878 14720
rect 6814 14660 6818 14716
rect 6818 14660 6874 14716
rect 6874 14660 6878 14716
rect 6814 14656 6878 14660
rect 10322 14716 10386 14720
rect 10322 14660 10326 14716
rect 10326 14660 10382 14716
rect 10382 14660 10386 14716
rect 10322 14656 10386 14660
rect 10402 14716 10466 14720
rect 10402 14660 10406 14716
rect 10406 14660 10462 14716
rect 10462 14660 10466 14716
rect 10402 14656 10466 14660
rect 10482 14716 10546 14720
rect 10482 14660 10486 14716
rect 10486 14660 10542 14716
rect 10542 14660 10546 14716
rect 10482 14656 10546 14660
rect 10562 14716 10626 14720
rect 10562 14660 10566 14716
rect 10566 14660 10622 14716
rect 10622 14660 10626 14716
rect 10562 14656 10626 14660
rect 14070 14716 14134 14720
rect 14070 14660 14074 14716
rect 14074 14660 14130 14716
rect 14130 14660 14134 14716
rect 14070 14656 14134 14660
rect 14150 14716 14214 14720
rect 14150 14660 14154 14716
rect 14154 14660 14210 14716
rect 14210 14660 14214 14716
rect 14150 14656 14214 14660
rect 14230 14716 14294 14720
rect 14230 14660 14234 14716
rect 14234 14660 14290 14716
rect 14290 14660 14294 14716
rect 14230 14656 14294 14660
rect 14310 14716 14374 14720
rect 14310 14660 14314 14716
rect 14314 14660 14370 14716
rect 14370 14660 14374 14716
rect 14310 14656 14374 14660
rect 4108 14240 4172 14244
rect 4108 14184 4122 14240
rect 4122 14184 4172 14240
rect 4108 14180 4172 14184
rect 7420 14180 7484 14244
rect 4700 14172 4764 14176
rect 4700 14116 4704 14172
rect 4704 14116 4760 14172
rect 4760 14116 4764 14172
rect 4700 14112 4764 14116
rect 4780 14172 4844 14176
rect 4780 14116 4784 14172
rect 4784 14116 4840 14172
rect 4840 14116 4844 14172
rect 4780 14112 4844 14116
rect 4860 14172 4924 14176
rect 4860 14116 4864 14172
rect 4864 14116 4920 14172
rect 4920 14116 4924 14172
rect 4860 14112 4924 14116
rect 4940 14172 5004 14176
rect 4940 14116 4944 14172
rect 4944 14116 5000 14172
rect 5000 14116 5004 14172
rect 4940 14112 5004 14116
rect 8448 14172 8512 14176
rect 8448 14116 8452 14172
rect 8452 14116 8508 14172
rect 8508 14116 8512 14172
rect 8448 14112 8512 14116
rect 8528 14172 8592 14176
rect 8528 14116 8532 14172
rect 8532 14116 8588 14172
rect 8588 14116 8592 14172
rect 8528 14112 8592 14116
rect 8608 14172 8672 14176
rect 8608 14116 8612 14172
rect 8612 14116 8668 14172
rect 8668 14116 8672 14172
rect 8608 14112 8672 14116
rect 8688 14172 8752 14176
rect 8688 14116 8692 14172
rect 8692 14116 8748 14172
rect 8748 14116 8752 14172
rect 8688 14112 8752 14116
rect 12196 14172 12260 14176
rect 12196 14116 12200 14172
rect 12200 14116 12256 14172
rect 12256 14116 12260 14172
rect 12196 14112 12260 14116
rect 12276 14172 12340 14176
rect 12276 14116 12280 14172
rect 12280 14116 12336 14172
rect 12336 14116 12340 14172
rect 12276 14112 12340 14116
rect 12356 14172 12420 14176
rect 12356 14116 12360 14172
rect 12360 14116 12416 14172
rect 12416 14116 12420 14172
rect 12356 14112 12420 14116
rect 12436 14172 12500 14176
rect 12436 14116 12440 14172
rect 12440 14116 12496 14172
rect 12496 14116 12500 14172
rect 12436 14112 12500 14116
rect 9260 13772 9324 13836
rect 12572 13772 12636 13836
rect 2826 13628 2890 13632
rect 2826 13572 2830 13628
rect 2830 13572 2886 13628
rect 2886 13572 2890 13628
rect 2826 13568 2890 13572
rect 2906 13628 2970 13632
rect 2906 13572 2910 13628
rect 2910 13572 2966 13628
rect 2966 13572 2970 13628
rect 2906 13568 2970 13572
rect 2986 13628 3050 13632
rect 2986 13572 2990 13628
rect 2990 13572 3046 13628
rect 3046 13572 3050 13628
rect 2986 13568 3050 13572
rect 3066 13628 3130 13632
rect 3066 13572 3070 13628
rect 3070 13572 3126 13628
rect 3126 13572 3130 13628
rect 3066 13568 3130 13572
rect 6574 13628 6638 13632
rect 6574 13572 6578 13628
rect 6578 13572 6634 13628
rect 6634 13572 6638 13628
rect 6574 13568 6638 13572
rect 6654 13628 6718 13632
rect 6654 13572 6658 13628
rect 6658 13572 6714 13628
rect 6714 13572 6718 13628
rect 6654 13568 6718 13572
rect 6734 13628 6798 13632
rect 6734 13572 6738 13628
rect 6738 13572 6794 13628
rect 6794 13572 6798 13628
rect 6734 13568 6798 13572
rect 6814 13628 6878 13632
rect 6814 13572 6818 13628
rect 6818 13572 6874 13628
rect 6874 13572 6878 13628
rect 6814 13568 6878 13572
rect 10322 13628 10386 13632
rect 10322 13572 10326 13628
rect 10326 13572 10382 13628
rect 10382 13572 10386 13628
rect 10322 13568 10386 13572
rect 10402 13628 10466 13632
rect 10402 13572 10406 13628
rect 10406 13572 10462 13628
rect 10462 13572 10466 13628
rect 10402 13568 10466 13572
rect 10482 13628 10546 13632
rect 10482 13572 10486 13628
rect 10486 13572 10542 13628
rect 10542 13572 10546 13628
rect 10482 13568 10546 13572
rect 10562 13628 10626 13632
rect 10562 13572 10566 13628
rect 10566 13572 10622 13628
rect 10622 13572 10626 13628
rect 10562 13568 10626 13572
rect 12020 13500 12084 13564
rect 14070 13628 14134 13632
rect 14070 13572 14074 13628
rect 14074 13572 14130 13628
rect 14130 13572 14134 13628
rect 14070 13568 14134 13572
rect 14150 13628 14214 13632
rect 14150 13572 14154 13628
rect 14154 13572 14210 13628
rect 14210 13572 14214 13628
rect 14150 13568 14214 13572
rect 14230 13628 14294 13632
rect 14230 13572 14234 13628
rect 14234 13572 14290 13628
rect 14290 13572 14294 13628
rect 14230 13568 14294 13572
rect 14310 13628 14374 13632
rect 14310 13572 14314 13628
rect 14314 13572 14370 13628
rect 14370 13572 14374 13628
rect 14310 13568 14374 13572
rect 13492 13560 13556 13564
rect 13492 13504 13542 13560
rect 13542 13504 13556 13560
rect 13492 13500 13556 13504
rect 13860 13560 13924 13564
rect 13860 13504 13874 13560
rect 13874 13504 13924 13560
rect 13860 13500 13924 13504
rect 13492 13092 13556 13156
rect 13676 13092 13740 13156
rect 4700 13084 4764 13088
rect 4700 13028 4704 13084
rect 4704 13028 4760 13084
rect 4760 13028 4764 13084
rect 4700 13024 4764 13028
rect 4780 13084 4844 13088
rect 4780 13028 4784 13084
rect 4784 13028 4840 13084
rect 4840 13028 4844 13084
rect 4780 13024 4844 13028
rect 4860 13084 4924 13088
rect 4860 13028 4864 13084
rect 4864 13028 4920 13084
rect 4920 13028 4924 13084
rect 4860 13024 4924 13028
rect 4940 13084 5004 13088
rect 4940 13028 4944 13084
rect 4944 13028 5000 13084
rect 5000 13028 5004 13084
rect 4940 13024 5004 13028
rect 8448 13084 8512 13088
rect 8448 13028 8452 13084
rect 8452 13028 8508 13084
rect 8508 13028 8512 13084
rect 8448 13024 8512 13028
rect 8528 13084 8592 13088
rect 8528 13028 8532 13084
rect 8532 13028 8588 13084
rect 8588 13028 8592 13084
rect 8528 13024 8592 13028
rect 8608 13084 8672 13088
rect 8608 13028 8612 13084
rect 8612 13028 8668 13084
rect 8668 13028 8672 13084
rect 8608 13024 8672 13028
rect 8688 13084 8752 13088
rect 8688 13028 8692 13084
rect 8692 13028 8748 13084
rect 8748 13028 8752 13084
rect 8688 13024 8752 13028
rect 12196 13084 12260 13088
rect 12196 13028 12200 13084
rect 12200 13028 12256 13084
rect 12256 13028 12260 13084
rect 12196 13024 12260 13028
rect 12276 13084 12340 13088
rect 12276 13028 12280 13084
rect 12280 13028 12336 13084
rect 12336 13028 12340 13084
rect 12276 13024 12340 13028
rect 12356 13084 12420 13088
rect 12356 13028 12360 13084
rect 12360 13028 12416 13084
rect 12416 13028 12420 13084
rect 12356 13024 12420 13028
rect 12436 13084 12500 13088
rect 12436 13028 12440 13084
rect 12440 13028 12496 13084
rect 12496 13028 12500 13084
rect 12436 13024 12500 13028
rect 8892 12684 8956 12748
rect 6132 12548 6196 12612
rect 2826 12540 2890 12544
rect 2826 12484 2830 12540
rect 2830 12484 2886 12540
rect 2886 12484 2890 12540
rect 2826 12480 2890 12484
rect 2906 12540 2970 12544
rect 2906 12484 2910 12540
rect 2910 12484 2966 12540
rect 2966 12484 2970 12540
rect 2906 12480 2970 12484
rect 2986 12540 3050 12544
rect 2986 12484 2990 12540
rect 2990 12484 3046 12540
rect 3046 12484 3050 12540
rect 2986 12480 3050 12484
rect 3066 12540 3130 12544
rect 3066 12484 3070 12540
rect 3070 12484 3126 12540
rect 3126 12484 3130 12540
rect 3066 12480 3130 12484
rect 6574 12540 6638 12544
rect 6574 12484 6578 12540
rect 6578 12484 6634 12540
rect 6634 12484 6638 12540
rect 6574 12480 6638 12484
rect 6654 12540 6718 12544
rect 6654 12484 6658 12540
rect 6658 12484 6714 12540
rect 6714 12484 6718 12540
rect 6654 12480 6718 12484
rect 6734 12540 6798 12544
rect 6734 12484 6738 12540
rect 6738 12484 6794 12540
rect 6794 12484 6798 12540
rect 6734 12480 6798 12484
rect 6814 12540 6878 12544
rect 6814 12484 6818 12540
rect 6818 12484 6874 12540
rect 6874 12484 6878 12540
rect 6814 12480 6878 12484
rect 10322 12540 10386 12544
rect 10322 12484 10326 12540
rect 10326 12484 10382 12540
rect 10382 12484 10386 12540
rect 10322 12480 10386 12484
rect 10402 12540 10466 12544
rect 10402 12484 10406 12540
rect 10406 12484 10462 12540
rect 10462 12484 10466 12540
rect 10402 12480 10466 12484
rect 10482 12540 10546 12544
rect 10482 12484 10486 12540
rect 10486 12484 10542 12540
rect 10542 12484 10546 12540
rect 10482 12480 10546 12484
rect 10562 12540 10626 12544
rect 10562 12484 10566 12540
rect 10566 12484 10622 12540
rect 10622 12484 10626 12540
rect 10562 12480 10626 12484
rect 14070 12540 14134 12544
rect 14070 12484 14074 12540
rect 14074 12484 14130 12540
rect 14130 12484 14134 12540
rect 14070 12480 14134 12484
rect 14150 12540 14214 12544
rect 14150 12484 14154 12540
rect 14154 12484 14210 12540
rect 14210 12484 14214 12540
rect 14150 12480 14214 12484
rect 14230 12540 14294 12544
rect 14230 12484 14234 12540
rect 14234 12484 14290 12540
rect 14290 12484 14294 12540
rect 14230 12480 14294 12484
rect 14310 12540 14374 12544
rect 14310 12484 14314 12540
rect 14314 12484 14370 12540
rect 14370 12484 14374 12540
rect 14310 12480 14374 12484
rect 9444 12276 9508 12340
rect 10916 12276 10980 12340
rect 12756 12276 12820 12340
rect 9812 12140 9876 12204
rect 4700 11996 4764 12000
rect 4700 11940 4704 11996
rect 4704 11940 4760 11996
rect 4760 11940 4764 11996
rect 4700 11936 4764 11940
rect 4780 11996 4844 12000
rect 4780 11940 4784 11996
rect 4784 11940 4840 11996
rect 4840 11940 4844 11996
rect 4780 11936 4844 11940
rect 4860 11996 4924 12000
rect 4860 11940 4864 11996
rect 4864 11940 4920 11996
rect 4920 11940 4924 11996
rect 4860 11936 4924 11940
rect 4940 11996 5004 12000
rect 4940 11940 4944 11996
rect 4944 11940 5000 11996
rect 5000 11940 5004 11996
rect 4940 11936 5004 11940
rect 8448 11996 8512 12000
rect 8448 11940 8452 11996
rect 8452 11940 8508 11996
rect 8508 11940 8512 11996
rect 8448 11936 8512 11940
rect 8528 11996 8592 12000
rect 8528 11940 8532 11996
rect 8532 11940 8588 11996
rect 8588 11940 8592 11996
rect 8528 11936 8592 11940
rect 8608 11996 8672 12000
rect 8608 11940 8612 11996
rect 8612 11940 8668 11996
rect 8668 11940 8672 11996
rect 8608 11936 8672 11940
rect 8688 11996 8752 12000
rect 8688 11940 8692 11996
rect 8692 11940 8748 11996
rect 8748 11940 8752 11996
rect 8688 11936 8752 11940
rect 12196 11996 12260 12000
rect 12196 11940 12200 11996
rect 12200 11940 12256 11996
rect 12256 11940 12260 11996
rect 12196 11936 12260 11940
rect 12276 11996 12340 12000
rect 12276 11940 12280 11996
rect 12280 11940 12336 11996
rect 12336 11940 12340 11996
rect 12276 11936 12340 11940
rect 12356 11996 12420 12000
rect 12356 11940 12360 11996
rect 12360 11940 12416 11996
rect 12416 11940 12420 11996
rect 12356 11936 12420 11940
rect 12436 11996 12500 12000
rect 12436 11940 12440 11996
rect 12440 11940 12496 11996
rect 12496 11940 12500 11996
rect 12436 11936 12500 11940
rect 10180 11868 10244 11932
rect 11468 11928 11532 11932
rect 11468 11872 11518 11928
rect 11518 11872 11532 11928
rect 11468 11868 11532 11872
rect 2826 11452 2890 11456
rect 2826 11396 2830 11452
rect 2830 11396 2886 11452
rect 2886 11396 2890 11452
rect 2826 11392 2890 11396
rect 2906 11452 2970 11456
rect 2906 11396 2910 11452
rect 2910 11396 2966 11452
rect 2966 11396 2970 11452
rect 2906 11392 2970 11396
rect 2986 11452 3050 11456
rect 2986 11396 2990 11452
rect 2990 11396 3046 11452
rect 3046 11396 3050 11452
rect 2986 11392 3050 11396
rect 3066 11452 3130 11456
rect 3066 11396 3070 11452
rect 3070 11396 3126 11452
rect 3126 11396 3130 11452
rect 3066 11392 3130 11396
rect 6574 11452 6638 11456
rect 6574 11396 6578 11452
rect 6578 11396 6634 11452
rect 6634 11396 6638 11452
rect 6574 11392 6638 11396
rect 6654 11452 6718 11456
rect 6654 11396 6658 11452
rect 6658 11396 6714 11452
rect 6714 11396 6718 11452
rect 6654 11392 6718 11396
rect 6734 11452 6798 11456
rect 6734 11396 6738 11452
rect 6738 11396 6794 11452
rect 6794 11396 6798 11452
rect 6734 11392 6798 11396
rect 6814 11452 6878 11456
rect 6814 11396 6818 11452
rect 6818 11396 6874 11452
rect 6874 11396 6878 11452
rect 6814 11392 6878 11396
rect 10322 11452 10386 11456
rect 10322 11396 10326 11452
rect 10326 11396 10382 11452
rect 10382 11396 10386 11452
rect 10322 11392 10386 11396
rect 10402 11452 10466 11456
rect 10402 11396 10406 11452
rect 10406 11396 10462 11452
rect 10462 11396 10466 11452
rect 10402 11392 10466 11396
rect 10482 11452 10546 11456
rect 10482 11396 10486 11452
rect 10486 11396 10542 11452
rect 10542 11396 10546 11452
rect 10482 11392 10546 11396
rect 10562 11452 10626 11456
rect 10562 11396 10566 11452
rect 10566 11396 10622 11452
rect 10622 11396 10626 11452
rect 10562 11392 10626 11396
rect 14070 11452 14134 11456
rect 14070 11396 14074 11452
rect 14074 11396 14130 11452
rect 14130 11396 14134 11452
rect 14070 11392 14134 11396
rect 14150 11452 14214 11456
rect 14150 11396 14154 11452
rect 14154 11396 14210 11452
rect 14210 11396 14214 11452
rect 14150 11392 14214 11396
rect 14230 11452 14294 11456
rect 14230 11396 14234 11452
rect 14234 11396 14290 11452
rect 14290 11396 14294 11452
rect 14230 11392 14294 11396
rect 14310 11452 14374 11456
rect 14310 11396 14314 11452
rect 14314 11396 14370 11452
rect 14370 11396 14374 11452
rect 14310 11392 14374 11396
rect 4700 10908 4764 10912
rect 4700 10852 4704 10908
rect 4704 10852 4760 10908
rect 4760 10852 4764 10908
rect 4700 10848 4764 10852
rect 4780 10908 4844 10912
rect 4780 10852 4784 10908
rect 4784 10852 4840 10908
rect 4840 10852 4844 10908
rect 4780 10848 4844 10852
rect 4860 10908 4924 10912
rect 4860 10852 4864 10908
rect 4864 10852 4920 10908
rect 4920 10852 4924 10908
rect 4860 10848 4924 10852
rect 4940 10908 5004 10912
rect 4940 10852 4944 10908
rect 4944 10852 5000 10908
rect 5000 10852 5004 10908
rect 4940 10848 5004 10852
rect 8448 10908 8512 10912
rect 8448 10852 8452 10908
rect 8452 10852 8508 10908
rect 8508 10852 8512 10908
rect 8448 10848 8512 10852
rect 8528 10908 8592 10912
rect 8528 10852 8532 10908
rect 8532 10852 8588 10908
rect 8588 10852 8592 10908
rect 8528 10848 8592 10852
rect 8608 10908 8672 10912
rect 8608 10852 8612 10908
rect 8612 10852 8668 10908
rect 8668 10852 8672 10908
rect 8608 10848 8672 10852
rect 8688 10908 8752 10912
rect 8688 10852 8692 10908
rect 8692 10852 8748 10908
rect 8748 10852 8752 10908
rect 8688 10848 8752 10852
rect 12196 10908 12260 10912
rect 12196 10852 12200 10908
rect 12200 10852 12256 10908
rect 12256 10852 12260 10908
rect 12196 10848 12260 10852
rect 12276 10908 12340 10912
rect 12276 10852 12280 10908
rect 12280 10852 12336 10908
rect 12336 10852 12340 10908
rect 12276 10848 12340 10852
rect 12356 10908 12420 10912
rect 12356 10852 12360 10908
rect 12360 10852 12416 10908
rect 12416 10852 12420 10908
rect 12356 10848 12420 10852
rect 12436 10908 12500 10912
rect 12436 10852 12440 10908
rect 12440 10852 12496 10908
rect 12496 10852 12500 10908
rect 12436 10848 12500 10852
rect 2826 10364 2890 10368
rect 2826 10308 2830 10364
rect 2830 10308 2886 10364
rect 2886 10308 2890 10364
rect 2826 10304 2890 10308
rect 2906 10364 2970 10368
rect 2906 10308 2910 10364
rect 2910 10308 2966 10364
rect 2966 10308 2970 10364
rect 2906 10304 2970 10308
rect 2986 10364 3050 10368
rect 2986 10308 2990 10364
rect 2990 10308 3046 10364
rect 3046 10308 3050 10364
rect 2986 10304 3050 10308
rect 3066 10364 3130 10368
rect 3066 10308 3070 10364
rect 3070 10308 3126 10364
rect 3126 10308 3130 10364
rect 3066 10304 3130 10308
rect 6574 10364 6638 10368
rect 6574 10308 6578 10364
rect 6578 10308 6634 10364
rect 6634 10308 6638 10364
rect 6574 10304 6638 10308
rect 6654 10364 6718 10368
rect 6654 10308 6658 10364
rect 6658 10308 6714 10364
rect 6714 10308 6718 10364
rect 6654 10304 6718 10308
rect 6734 10364 6798 10368
rect 6734 10308 6738 10364
rect 6738 10308 6794 10364
rect 6794 10308 6798 10364
rect 6734 10304 6798 10308
rect 6814 10364 6878 10368
rect 6814 10308 6818 10364
rect 6818 10308 6874 10364
rect 6874 10308 6878 10364
rect 6814 10304 6878 10308
rect 10322 10364 10386 10368
rect 10322 10308 10326 10364
rect 10326 10308 10382 10364
rect 10382 10308 10386 10364
rect 10322 10304 10386 10308
rect 10402 10364 10466 10368
rect 10402 10308 10406 10364
rect 10406 10308 10462 10364
rect 10462 10308 10466 10364
rect 10402 10304 10466 10308
rect 10482 10364 10546 10368
rect 10482 10308 10486 10364
rect 10486 10308 10542 10364
rect 10542 10308 10546 10364
rect 10482 10304 10546 10308
rect 10562 10364 10626 10368
rect 10562 10308 10566 10364
rect 10566 10308 10622 10364
rect 10622 10308 10626 10364
rect 10562 10304 10626 10308
rect 14070 10364 14134 10368
rect 14070 10308 14074 10364
rect 14074 10308 14130 10364
rect 14130 10308 14134 10364
rect 14070 10304 14134 10308
rect 14150 10364 14214 10368
rect 14150 10308 14154 10364
rect 14154 10308 14210 10364
rect 14210 10308 14214 10364
rect 14150 10304 14214 10308
rect 14230 10364 14294 10368
rect 14230 10308 14234 10364
rect 14234 10308 14290 10364
rect 14290 10308 14294 10364
rect 14230 10304 14294 10308
rect 14310 10364 14374 10368
rect 14310 10308 14314 10364
rect 14314 10308 14370 10364
rect 14370 10308 14374 10364
rect 14310 10304 14374 10308
rect 13860 10296 13924 10300
rect 13860 10240 13874 10296
rect 13874 10240 13924 10296
rect 13860 10236 13924 10240
rect 13124 10100 13188 10164
rect 13492 10024 13556 10028
rect 13492 9968 13506 10024
rect 13506 9968 13556 10024
rect 13492 9964 13556 9968
rect 14596 9964 14660 10028
rect 11100 9828 11164 9892
rect 4700 9820 4764 9824
rect 4700 9764 4704 9820
rect 4704 9764 4760 9820
rect 4760 9764 4764 9820
rect 4700 9760 4764 9764
rect 4780 9820 4844 9824
rect 4780 9764 4784 9820
rect 4784 9764 4840 9820
rect 4840 9764 4844 9820
rect 4780 9760 4844 9764
rect 4860 9820 4924 9824
rect 4860 9764 4864 9820
rect 4864 9764 4920 9820
rect 4920 9764 4924 9820
rect 4860 9760 4924 9764
rect 4940 9820 5004 9824
rect 4940 9764 4944 9820
rect 4944 9764 5000 9820
rect 5000 9764 5004 9820
rect 4940 9760 5004 9764
rect 8448 9820 8512 9824
rect 8448 9764 8452 9820
rect 8452 9764 8508 9820
rect 8508 9764 8512 9820
rect 8448 9760 8512 9764
rect 8528 9820 8592 9824
rect 8528 9764 8532 9820
rect 8532 9764 8588 9820
rect 8588 9764 8592 9820
rect 8528 9760 8592 9764
rect 8608 9820 8672 9824
rect 8608 9764 8612 9820
rect 8612 9764 8668 9820
rect 8668 9764 8672 9820
rect 8608 9760 8672 9764
rect 8688 9820 8752 9824
rect 8688 9764 8692 9820
rect 8692 9764 8748 9820
rect 8748 9764 8752 9820
rect 8688 9760 8752 9764
rect 12196 9820 12260 9824
rect 12196 9764 12200 9820
rect 12200 9764 12256 9820
rect 12256 9764 12260 9820
rect 12196 9760 12260 9764
rect 12276 9820 12340 9824
rect 12276 9764 12280 9820
rect 12280 9764 12336 9820
rect 12336 9764 12340 9820
rect 12276 9760 12340 9764
rect 12356 9820 12420 9824
rect 12356 9764 12360 9820
rect 12360 9764 12416 9820
rect 12416 9764 12420 9820
rect 12356 9760 12420 9764
rect 12436 9820 12500 9824
rect 12436 9764 12440 9820
rect 12440 9764 12496 9820
rect 12496 9764 12500 9820
rect 12436 9760 12500 9764
rect 4108 9556 4172 9620
rect 13492 9556 13556 9620
rect 2826 9276 2890 9280
rect 2826 9220 2830 9276
rect 2830 9220 2886 9276
rect 2886 9220 2890 9276
rect 2826 9216 2890 9220
rect 2906 9276 2970 9280
rect 2906 9220 2910 9276
rect 2910 9220 2966 9276
rect 2966 9220 2970 9276
rect 2906 9216 2970 9220
rect 2986 9276 3050 9280
rect 2986 9220 2990 9276
rect 2990 9220 3046 9276
rect 3046 9220 3050 9276
rect 2986 9216 3050 9220
rect 3066 9276 3130 9280
rect 3066 9220 3070 9276
rect 3070 9220 3126 9276
rect 3126 9220 3130 9276
rect 3066 9216 3130 9220
rect 6574 9276 6638 9280
rect 6574 9220 6578 9276
rect 6578 9220 6634 9276
rect 6634 9220 6638 9276
rect 6574 9216 6638 9220
rect 6654 9276 6718 9280
rect 6654 9220 6658 9276
rect 6658 9220 6714 9276
rect 6714 9220 6718 9276
rect 6654 9216 6718 9220
rect 6734 9276 6798 9280
rect 6734 9220 6738 9276
rect 6738 9220 6794 9276
rect 6794 9220 6798 9276
rect 6734 9216 6798 9220
rect 6814 9276 6878 9280
rect 6814 9220 6818 9276
rect 6818 9220 6874 9276
rect 6874 9220 6878 9276
rect 6814 9216 6878 9220
rect 7972 9148 8036 9212
rect 5396 9012 5460 9076
rect 8892 9012 8956 9076
rect 13676 9420 13740 9484
rect 11284 9284 11348 9348
rect 10322 9276 10386 9280
rect 10322 9220 10326 9276
rect 10326 9220 10382 9276
rect 10382 9220 10386 9276
rect 10322 9216 10386 9220
rect 10402 9276 10466 9280
rect 10402 9220 10406 9276
rect 10406 9220 10462 9276
rect 10462 9220 10466 9276
rect 10402 9216 10466 9220
rect 10482 9276 10546 9280
rect 10482 9220 10486 9276
rect 10486 9220 10542 9276
rect 10542 9220 10546 9276
rect 10482 9216 10546 9220
rect 10562 9276 10626 9280
rect 10562 9220 10566 9276
rect 10566 9220 10622 9276
rect 10622 9220 10626 9276
rect 10562 9216 10626 9220
rect 14070 9276 14134 9280
rect 14070 9220 14074 9276
rect 14074 9220 14130 9276
rect 14130 9220 14134 9276
rect 14070 9216 14134 9220
rect 14150 9276 14214 9280
rect 14150 9220 14154 9276
rect 14154 9220 14210 9276
rect 14210 9220 14214 9276
rect 14150 9216 14214 9220
rect 14230 9276 14294 9280
rect 14230 9220 14234 9276
rect 14234 9220 14290 9276
rect 14290 9220 14294 9276
rect 14230 9216 14294 9220
rect 14310 9276 14374 9280
rect 14310 9220 14314 9276
rect 14314 9220 14370 9276
rect 14370 9220 14374 9276
rect 14310 9216 14374 9220
rect 11468 9148 11532 9212
rect 12020 9148 12084 9212
rect 8156 8740 8220 8804
rect 13676 8740 13740 8804
rect 4700 8732 4764 8736
rect 4700 8676 4704 8732
rect 4704 8676 4760 8732
rect 4760 8676 4764 8732
rect 4700 8672 4764 8676
rect 4780 8732 4844 8736
rect 4780 8676 4784 8732
rect 4784 8676 4840 8732
rect 4840 8676 4844 8732
rect 4780 8672 4844 8676
rect 4860 8732 4924 8736
rect 4860 8676 4864 8732
rect 4864 8676 4920 8732
rect 4920 8676 4924 8732
rect 4860 8672 4924 8676
rect 4940 8732 5004 8736
rect 4940 8676 4944 8732
rect 4944 8676 5000 8732
rect 5000 8676 5004 8732
rect 4940 8672 5004 8676
rect 8448 8732 8512 8736
rect 8448 8676 8452 8732
rect 8452 8676 8508 8732
rect 8508 8676 8512 8732
rect 8448 8672 8512 8676
rect 8528 8732 8592 8736
rect 8528 8676 8532 8732
rect 8532 8676 8588 8732
rect 8588 8676 8592 8732
rect 8528 8672 8592 8676
rect 8608 8732 8672 8736
rect 8608 8676 8612 8732
rect 8612 8676 8668 8732
rect 8668 8676 8672 8732
rect 8608 8672 8672 8676
rect 8688 8732 8752 8736
rect 8688 8676 8692 8732
rect 8692 8676 8748 8732
rect 8748 8676 8752 8732
rect 8688 8672 8752 8676
rect 12196 8732 12260 8736
rect 12196 8676 12200 8732
rect 12200 8676 12256 8732
rect 12256 8676 12260 8732
rect 12196 8672 12260 8676
rect 12276 8732 12340 8736
rect 12276 8676 12280 8732
rect 12280 8676 12336 8732
rect 12336 8676 12340 8732
rect 12276 8672 12340 8676
rect 12356 8732 12420 8736
rect 12356 8676 12360 8732
rect 12360 8676 12416 8732
rect 12416 8676 12420 8732
rect 12356 8672 12420 8676
rect 12436 8732 12500 8736
rect 12436 8676 12440 8732
rect 12440 8676 12496 8732
rect 12496 8676 12500 8732
rect 12436 8672 12500 8676
rect 9812 8468 9876 8532
rect 11836 8528 11900 8532
rect 11836 8472 11886 8528
rect 11886 8472 11900 8528
rect 11836 8468 11900 8472
rect 12572 8468 12636 8532
rect 2826 8188 2890 8192
rect 2826 8132 2830 8188
rect 2830 8132 2886 8188
rect 2886 8132 2890 8188
rect 2826 8128 2890 8132
rect 2906 8188 2970 8192
rect 2906 8132 2910 8188
rect 2910 8132 2966 8188
rect 2966 8132 2970 8188
rect 2906 8128 2970 8132
rect 2986 8188 3050 8192
rect 2986 8132 2990 8188
rect 2990 8132 3046 8188
rect 3046 8132 3050 8188
rect 2986 8128 3050 8132
rect 3066 8188 3130 8192
rect 3066 8132 3070 8188
rect 3070 8132 3126 8188
rect 3126 8132 3130 8188
rect 3066 8128 3130 8132
rect 6574 8188 6638 8192
rect 6574 8132 6578 8188
rect 6578 8132 6634 8188
rect 6634 8132 6638 8188
rect 6574 8128 6638 8132
rect 6654 8188 6718 8192
rect 6654 8132 6658 8188
rect 6658 8132 6714 8188
rect 6714 8132 6718 8188
rect 6654 8128 6718 8132
rect 6734 8188 6798 8192
rect 6734 8132 6738 8188
rect 6738 8132 6794 8188
rect 6794 8132 6798 8188
rect 6734 8128 6798 8132
rect 6814 8188 6878 8192
rect 6814 8132 6818 8188
rect 6818 8132 6874 8188
rect 6874 8132 6878 8188
rect 6814 8128 6878 8132
rect 10322 8188 10386 8192
rect 10322 8132 10326 8188
rect 10326 8132 10382 8188
rect 10382 8132 10386 8188
rect 10322 8128 10386 8132
rect 10402 8188 10466 8192
rect 10402 8132 10406 8188
rect 10406 8132 10462 8188
rect 10462 8132 10466 8188
rect 10402 8128 10466 8132
rect 10482 8188 10546 8192
rect 10482 8132 10486 8188
rect 10486 8132 10542 8188
rect 10542 8132 10546 8188
rect 10482 8128 10546 8132
rect 10562 8188 10626 8192
rect 10562 8132 10566 8188
rect 10566 8132 10622 8188
rect 10622 8132 10626 8188
rect 10562 8128 10626 8132
rect 14070 8188 14134 8192
rect 14070 8132 14074 8188
rect 14074 8132 14130 8188
rect 14130 8132 14134 8188
rect 14070 8128 14134 8132
rect 14150 8188 14214 8192
rect 14150 8132 14154 8188
rect 14154 8132 14210 8188
rect 14210 8132 14214 8188
rect 14150 8128 14214 8132
rect 14230 8188 14294 8192
rect 14230 8132 14234 8188
rect 14234 8132 14290 8188
rect 14290 8132 14294 8188
rect 14230 8128 14294 8132
rect 14310 8188 14374 8192
rect 14310 8132 14314 8188
rect 14314 8132 14370 8188
rect 14370 8132 14374 8188
rect 14310 8128 14374 8132
rect 9628 8060 9692 8124
rect 10732 7924 10796 7988
rect 13860 7984 13924 7988
rect 13860 7928 13910 7984
rect 13910 7928 13924 7984
rect 13860 7924 13924 7928
rect 12572 7652 12636 7716
rect 4700 7644 4764 7648
rect 4700 7588 4704 7644
rect 4704 7588 4760 7644
rect 4760 7588 4764 7644
rect 4700 7584 4764 7588
rect 4780 7644 4844 7648
rect 4780 7588 4784 7644
rect 4784 7588 4840 7644
rect 4840 7588 4844 7644
rect 4780 7584 4844 7588
rect 4860 7644 4924 7648
rect 4860 7588 4864 7644
rect 4864 7588 4920 7644
rect 4920 7588 4924 7644
rect 4860 7584 4924 7588
rect 4940 7644 5004 7648
rect 4940 7588 4944 7644
rect 4944 7588 5000 7644
rect 5000 7588 5004 7644
rect 4940 7584 5004 7588
rect 8448 7644 8512 7648
rect 8448 7588 8452 7644
rect 8452 7588 8508 7644
rect 8508 7588 8512 7644
rect 8448 7584 8512 7588
rect 8528 7644 8592 7648
rect 8528 7588 8532 7644
rect 8532 7588 8588 7644
rect 8588 7588 8592 7644
rect 8528 7584 8592 7588
rect 8608 7644 8672 7648
rect 8608 7588 8612 7644
rect 8612 7588 8668 7644
rect 8668 7588 8672 7644
rect 8608 7584 8672 7588
rect 8688 7644 8752 7648
rect 8688 7588 8692 7644
rect 8692 7588 8748 7644
rect 8748 7588 8752 7644
rect 8688 7584 8752 7588
rect 12196 7644 12260 7648
rect 12196 7588 12200 7644
rect 12200 7588 12256 7644
rect 12256 7588 12260 7644
rect 12196 7584 12260 7588
rect 12276 7644 12340 7648
rect 12276 7588 12280 7644
rect 12280 7588 12336 7644
rect 12336 7588 12340 7644
rect 12276 7584 12340 7588
rect 12356 7644 12420 7648
rect 12356 7588 12360 7644
rect 12360 7588 12416 7644
rect 12416 7588 12420 7644
rect 12356 7584 12420 7588
rect 12436 7644 12500 7648
rect 12436 7588 12440 7644
rect 12440 7588 12496 7644
rect 12496 7588 12500 7644
rect 12436 7584 12500 7588
rect 8892 7576 8956 7580
rect 8892 7520 8906 7576
rect 8906 7520 8956 7576
rect 8892 7516 8956 7520
rect 5948 7380 6012 7444
rect 10180 7244 10244 7308
rect 2826 7100 2890 7104
rect 2826 7044 2830 7100
rect 2830 7044 2886 7100
rect 2886 7044 2890 7100
rect 2826 7040 2890 7044
rect 2906 7100 2970 7104
rect 2906 7044 2910 7100
rect 2910 7044 2966 7100
rect 2966 7044 2970 7100
rect 2906 7040 2970 7044
rect 2986 7100 3050 7104
rect 2986 7044 2990 7100
rect 2990 7044 3046 7100
rect 3046 7044 3050 7100
rect 2986 7040 3050 7044
rect 3066 7100 3130 7104
rect 3066 7044 3070 7100
rect 3070 7044 3126 7100
rect 3126 7044 3130 7100
rect 3066 7040 3130 7044
rect 6574 7100 6638 7104
rect 6574 7044 6578 7100
rect 6578 7044 6634 7100
rect 6634 7044 6638 7100
rect 6574 7040 6638 7044
rect 6654 7100 6718 7104
rect 6654 7044 6658 7100
rect 6658 7044 6714 7100
rect 6714 7044 6718 7100
rect 6654 7040 6718 7044
rect 6734 7100 6798 7104
rect 6734 7044 6738 7100
rect 6738 7044 6794 7100
rect 6794 7044 6798 7100
rect 6734 7040 6798 7044
rect 6814 7100 6878 7104
rect 6814 7044 6818 7100
rect 6818 7044 6874 7100
rect 6874 7044 6878 7100
rect 6814 7040 6878 7044
rect 6132 6836 6196 6900
rect 12940 7440 13004 7444
rect 12940 7384 12954 7440
rect 12954 7384 13004 7440
rect 12940 7380 13004 7384
rect 10322 7100 10386 7104
rect 10322 7044 10326 7100
rect 10326 7044 10382 7100
rect 10382 7044 10386 7100
rect 10322 7040 10386 7044
rect 10402 7100 10466 7104
rect 10402 7044 10406 7100
rect 10406 7044 10462 7100
rect 10462 7044 10466 7100
rect 10402 7040 10466 7044
rect 10482 7100 10546 7104
rect 10482 7044 10486 7100
rect 10486 7044 10542 7100
rect 10542 7044 10546 7100
rect 10482 7040 10546 7044
rect 10562 7100 10626 7104
rect 10562 7044 10566 7100
rect 10566 7044 10622 7100
rect 10622 7044 10626 7100
rect 10562 7040 10626 7044
rect 14070 7100 14134 7104
rect 14070 7044 14074 7100
rect 14074 7044 14130 7100
rect 14130 7044 14134 7100
rect 14070 7040 14134 7044
rect 14150 7100 14214 7104
rect 14150 7044 14154 7100
rect 14154 7044 14210 7100
rect 14210 7044 14214 7100
rect 14150 7040 14214 7044
rect 14230 7100 14294 7104
rect 14230 7044 14234 7100
rect 14234 7044 14290 7100
rect 14290 7044 14294 7100
rect 14230 7040 14294 7044
rect 14310 7100 14374 7104
rect 14310 7044 14314 7100
rect 14314 7044 14370 7100
rect 14370 7044 14374 7100
rect 14310 7040 14374 7044
rect 9858 7032 9922 7036
rect 9858 6976 9862 7032
rect 9862 6976 9918 7032
rect 9918 6976 9922 7032
rect 9858 6972 9922 6976
rect 11652 6972 11716 7036
rect 12020 7032 12084 7036
rect 12020 6976 12070 7032
rect 12070 6976 12084 7032
rect 12020 6972 12084 6976
rect 7604 6700 7668 6764
rect 7788 6700 7852 6764
rect 9996 6700 10060 6764
rect 7236 6564 7300 6628
rect 9260 6564 9324 6628
rect 11284 6624 11348 6628
rect 11284 6568 11298 6624
rect 11298 6568 11348 6624
rect 4700 6556 4764 6560
rect 4700 6500 4704 6556
rect 4704 6500 4760 6556
rect 4760 6500 4764 6556
rect 4700 6496 4764 6500
rect 4780 6556 4844 6560
rect 4780 6500 4784 6556
rect 4784 6500 4840 6556
rect 4840 6500 4844 6556
rect 4780 6496 4844 6500
rect 4860 6556 4924 6560
rect 4860 6500 4864 6556
rect 4864 6500 4920 6556
rect 4920 6500 4924 6556
rect 4860 6496 4924 6500
rect 4940 6556 5004 6560
rect 4940 6500 4944 6556
rect 4944 6500 5000 6556
rect 5000 6500 5004 6556
rect 4940 6496 5004 6500
rect 8448 6556 8512 6560
rect 8448 6500 8452 6556
rect 8452 6500 8508 6556
rect 8508 6500 8512 6556
rect 8448 6496 8512 6500
rect 8528 6556 8592 6560
rect 8528 6500 8532 6556
rect 8532 6500 8588 6556
rect 8588 6500 8592 6556
rect 8528 6496 8592 6500
rect 8608 6556 8672 6560
rect 8608 6500 8612 6556
rect 8612 6500 8668 6556
rect 8668 6500 8672 6556
rect 8608 6496 8672 6500
rect 8688 6556 8752 6560
rect 8688 6500 8692 6556
rect 8692 6500 8748 6556
rect 8748 6500 8752 6556
rect 8688 6496 8752 6500
rect 3740 6428 3804 6492
rect 4476 6156 4540 6220
rect 7604 6020 7668 6084
rect 11284 6564 11348 6568
rect 12196 6556 12260 6560
rect 12196 6500 12200 6556
rect 12200 6500 12256 6556
rect 12256 6500 12260 6556
rect 12196 6496 12260 6500
rect 12276 6556 12340 6560
rect 12276 6500 12280 6556
rect 12280 6500 12336 6556
rect 12336 6500 12340 6556
rect 12276 6496 12340 6500
rect 12356 6556 12420 6560
rect 12356 6500 12360 6556
rect 12360 6500 12416 6556
rect 12416 6500 12420 6556
rect 12356 6496 12420 6500
rect 12436 6556 12500 6560
rect 12436 6500 12440 6556
rect 12440 6500 12496 6556
rect 12496 6500 12500 6556
rect 12436 6496 12500 6500
rect 13124 6488 13188 6492
rect 13124 6432 13174 6488
rect 13174 6432 13188 6488
rect 13124 6428 13188 6432
rect 11284 6292 11348 6356
rect 13860 6428 13924 6492
rect 9260 6020 9324 6084
rect 2826 6012 2890 6016
rect 2826 5956 2830 6012
rect 2830 5956 2886 6012
rect 2886 5956 2890 6012
rect 2826 5952 2890 5956
rect 2906 6012 2970 6016
rect 2906 5956 2910 6012
rect 2910 5956 2966 6012
rect 2966 5956 2970 6012
rect 2906 5952 2970 5956
rect 2986 6012 3050 6016
rect 2986 5956 2990 6012
rect 2990 5956 3046 6012
rect 3046 5956 3050 6012
rect 2986 5952 3050 5956
rect 3066 6012 3130 6016
rect 3066 5956 3070 6012
rect 3070 5956 3126 6012
rect 3126 5956 3130 6012
rect 3066 5952 3130 5956
rect 6574 6012 6638 6016
rect 6574 5956 6578 6012
rect 6578 5956 6634 6012
rect 6634 5956 6638 6012
rect 6574 5952 6638 5956
rect 6654 6012 6718 6016
rect 6654 5956 6658 6012
rect 6658 5956 6714 6012
rect 6714 5956 6718 6012
rect 6654 5952 6718 5956
rect 6734 6012 6798 6016
rect 6734 5956 6738 6012
rect 6738 5956 6794 6012
rect 6794 5956 6798 6012
rect 6734 5952 6798 5956
rect 6814 6012 6878 6016
rect 6814 5956 6818 6012
rect 6818 5956 6874 6012
rect 6874 5956 6878 6012
rect 6814 5952 6878 5956
rect 10322 6012 10386 6016
rect 10322 5956 10326 6012
rect 10326 5956 10382 6012
rect 10382 5956 10386 6012
rect 10322 5952 10386 5956
rect 10402 6012 10466 6016
rect 10402 5956 10406 6012
rect 10406 5956 10462 6012
rect 10462 5956 10466 6012
rect 10402 5952 10466 5956
rect 10482 6012 10546 6016
rect 10482 5956 10486 6012
rect 10486 5956 10542 6012
rect 10542 5956 10546 6012
rect 10482 5952 10546 5956
rect 10562 6012 10626 6016
rect 10562 5956 10566 6012
rect 10566 5956 10622 6012
rect 10622 5956 10626 6012
rect 10562 5952 10626 5956
rect 3372 5884 3436 5948
rect 5212 5612 5276 5676
rect 9628 5748 9692 5812
rect 12572 6216 12636 6220
rect 12572 6160 12622 6216
rect 12622 6160 12636 6216
rect 12572 6156 12636 6160
rect 14780 6020 14844 6084
rect 14070 6012 14134 6016
rect 14070 5956 14074 6012
rect 14074 5956 14130 6012
rect 14130 5956 14134 6012
rect 14070 5952 14134 5956
rect 14150 6012 14214 6016
rect 14150 5956 14154 6012
rect 14154 5956 14210 6012
rect 14210 5956 14214 6012
rect 14150 5952 14214 5956
rect 14230 6012 14294 6016
rect 14230 5956 14234 6012
rect 14234 5956 14290 6012
rect 14290 5956 14294 6012
rect 14230 5952 14294 5956
rect 14310 6012 14374 6016
rect 14310 5956 14314 6012
rect 14314 5956 14370 6012
rect 14370 5956 14374 6012
rect 14310 5952 14374 5956
rect 11100 5884 11164 5948
rect 11100 5748 11164 5812
rect 13124 5612 13188 5676
rect 6132 5476 6196 5540
rect 7052 5476 7116 5540
rect 9260 5476 9324 5540
rect 14596 5476 14660 5540
rect 4700 5468 4764 5472
rect 4700 5412 4704 5468
rect 4704 5412 4760 5468
rect 4760 5412 4764 5468
rect 4700 5408 4764 5412
rect 4780 5468 4844 5472
rect 4780 5412 4784 5468
rect 4784 5412 4840 5468
rect 4840 5412 4844 5468
rect 4780 5408 4844 5412
rect 4860 5468 4924 5472
rect 4860 5412 4864 5468
rect 4864 5412 4920 5468
rect 4920 5412 4924 5468
rect 4860 5408 4924 5412
rect 4940 5468 5004 5472
rect 4940 5412 4944 5468
rect 4944 5412 5000 5468
rect 5000 5412 5004 5468
rect 4940 5408 5004 5412
rect 8448 5468 8512 5472
rect 8448 5412 8452 5468
rect 8452 5412 8508 5468
rect 8508 5412 8512 5468
rect 8448 5408 8512 5412
rect 8528 5468 8592 5472
rect 8528 5412 8532 5468
rect 8532 5412 8588 5468
rect 8588 5412 8592 5468
rect 8528 5408 8592 5412
rect 8608 5468 8672 5472
rect 8608 5412 8612 5468
rect 8612 5412 8668 5468
rect 8668 5412 8672 5468
rect 8608 5408 8672 5412
rect 8688 5468 8752 5472
rect 8688 5412 8692 5468
rect 8692 5412 8748 5468
rect 8748 5412 8752 5468
rect 8688 5408 8752 5412
rect 7788 5340 7852 5404
rect 12196 5468 12260 5472
rect 12196 5412 12200 5468
rect 12200 5412 12256 5468
rect 12256 5412 12260 5468
rect 12196 5408 12260 5412
rect 12276 5468 12340 5472
rect 12276 5412 12280 5468
rect 12280 5412 12336 5468
rect 12336 5412 12340 5468
rect 12276 5408 12340 5412
rect 12356 5468 12420 5472
rect 12356 5412 12360 5468
rect 12360 5412 12416 5468
rect 12416 5412 12420 5468
rect 12356 5408 12420 5412
rect 12436 5468 12500 5472
rect 12436 5412 12440 5468
rect 12440 5412 12496 5468
rect 12496 5412 12500 5468
rect 12436 5408 12500 5412
rect 9628 5400 9692 5404
rect 9628 5344 9642 5400
rect 9642 5344 9692 5400
rect 9628 5340 9692 5344
rect 12572 5340 12636 5404
rect 13860 5340 13924 5404
rect 15332 5340 15396 5404
rect 5396 5264 5460 5268
rect 5396 5208 5446 5264
rect 5446 5208 5460 5264
rect 5396 5204 5460 5208
rect 9812 5204 9876 5268
rect 10180 5204 10244 5268
rect 13860 5264 13924 5268
rect 13860 5208 13910 5264
rect 13910 5208 13924 5264
rect 13860 5204 13924 5208
rect 2826 4924 2890 4928
rect 2826 4868 2830 4924
rect 2830 4868 2886 4924
rect 2886 4868 2890 4924
rect 2826 4864 2890 4868
rect 2906 4924 2970 4928
rect 2906 4868 2910 4924
rect 2910 4868 2966 4924
rect 2966 4868 2970 4924
rect 2906 4864 2970 4868
rect 2986 4924 3050 4928
rect 2986 4868 2990 4924
rect 2990 4868 3046 4924
rect 3046 4868 3050 4924
rect 2986 4864 3050 4868
rect 3066 4924 3130 4928
rect 3066 4868 3070 4924
rect 3070 4868 3126 4924
rect 3126 4868 3130 4924
rect 3066 4864 3130 4868
rect 6574 4924 6638 4928
rect 6574 4868 6578 4924
rect 6578 4868 6634 4924
rect 6634 4868 6638 4924
rect 6574 4864 6638 4868
rect 6654 4924 6718 4928
rect 6654 4868 6658 4924
rect 6658 4868 6714 4924
rect 6714 4868 6718 4924
rect 6654 4864 6718 4868
rect 6734 4924 6798 4928
rect 6734 4868 6738 4924
rect 6738 4868 6794 4924
rect 6794 4868 6798 4924
rect 6734 4864 6798 4868
rect 6814 4924 6878 4928
rect 6814 4868 6818 4924
rect 6818 4868 6874 4924
rect 6874 4868 6878 4924
rect 6814 4864 6878 4868
rect 2452 4856 2516 4860
rect 2452 4800 2466 4856
rect 2466 4800 2516 4856
rect 2452 4796 2516 4800
rect 3740 4856 3804 4860
rect 3740 4800 3754 4856
rect 3754 4800 3804 4856
rect 3740 4796 3804 4800
rect 3924 4796 3988 4860
rect 6316 4796 6380 4860
rect 10322 4924 10386 4928
rect 10322 4868 10326 4924
rect 10326 4868 10382 4924
rect 10382 4868 10386 4924
rect 10322 4864 10386 4868
rect 10402 4924 10466 4928
rect 10402 4868 10406 4924
rect 10406 4868 10462 4924
rect 10462 4868 10466 4924
rect 10402 4864 10466 4868
rect 10482 4924 10546 4928
rect 10482 4868 10486 4924
rect 10486 4868 10542 4924
rect 10542 4868 10546 4924
rect 10482 4864 10546 4868
rect 10562 4924 10626 4928
rect 10562 4868 10566 4924
rect 10566 4868 10622 4924
rect 10622 4868 10626 4924
rect 10562 4864 10626 4868
rect 9628 4796 9692 4860
rect 9996 4796 10060 4860
rect 12572 4796 12636 4860
rect 12940 4856 13004 4860
rect 12940 4800 12990 4856
rect 12990 4800 13004 4856
rect 12940 4796 13004 4800
rect 4292 4524 4356 4588
rect 14070 4924 14134 4928
rect 14070 4868 14074 4924
rect 14074 4868 14130 4924
rect 14130 4868 14134 4924
rect 14070 4864 14134 4868
rect 14150 4924 14214 4928
rect 14150 4868 14154 4924
rect 14154 4868 14210 4924
rect 14210 4868 14214 4924
rect 14150 4864 14214 4868
rect 14230 4924 14294 4928
rect 14230 4868 14234 4924
rect 14234 4868 14290 4924
rect 14290 4868 14294 4924
rect 14230 4864 14294 4868
rect 14310 4924 14374 4928
rect 14310 4868 14314 4924
rect 14314 4868 14370 4924
rect 14370 4868 14374 4924
rect 14310 4864 14374 4868
rect 4476 4388 4540 4452
rect 4700 4380 4764 4384
rect 4700 4324 4704 4380
rect 4704 4324 4760 4380
rect 4760 4324 4764 4380
rect 4700 4320 4764 4324
rect 4780 4380 4844 4384
rect 4780 4324 4784 4380
rect 4784 4324 4840 4380
rect 4840 4324 4844 4380
rect 4780 4320 4844 4324
rect 4860 4380 4924 4384
rect 4860 4324 4864 4380
rect 4864 4324 4920 4380
rect 4920 4324 4924 4380
rect 4860 4320 4924 4324
rect 4940 4380 5004 4384
rect 4940 4324 4944 4380
rect 4944 4324 5000 4380
rect 5000 4324 5004 4380
rect 4940 4320 5004 4324
rect 8448 4380 8512 4384
rect 8448 4324 8452 4380
rect 8452 4324 8508 4380
rect 8508 4324 8512 4380
rect 8448 4320 8512 4324
rect 8528 4380 8592 4384
rect 8528 4324 8532 4380
rect 8532 4324 8588 4380
rect 8588 4324 8592 4380
rect 8528 4320 8592 4324
rect 8608 4380 8672 4384
rect 8608 4324 8612 4380
rect 8612 4324 8668 4380
rect 8668 4324 8672 4380
rect 8608 4320 8672 4324
rect 8688 4380 8752 4384
rect 8688 4324 8692 4380
rect 8692 4324 8748 4380
rect 8748 4324 8752 4380
rect 8688 4320 8752 4324
rect 9628 4252 9692 4316
rect 10732 4252 10796 4316
rect 11284 4388 11348 4452
rect 12572 4388 12636 4452
rect 13676 4388 13740 4452
rect 12196 4380 12260 4384
rect 12196 4324 12200 4380
rect 12200 4324 12256 4380
rect 12256 4324 12260 4380
rect 12196 4320 12260 4324
rect 12276 4380 12340 4384
rect 12276 4324 12280 4380
rect 12280 4324 12336 4380
rect 12336 4324 12340 4380
rect 12276 4320 12340 4324
rect 12356 4380 12420 4384
rect 12356 4324 12360 4380
rect 12360 4324 12416 4380
rect 12416 4324 12420 4380
rect 12356 4320 12420 4324
rect 12436 4380 12500 4384
rect 12436 4324 12440 4380
rect 12440 4324 12496 4380
rect 12496 4324 12500 4380
rect 12436 4320 12500 4324
rect 11284 4252 11348 4316
rect 1716 4040 1780 4044
rect 1716 3984 1766 4040
rect 1766 3984 1780 4040
rect 1716 3980 1780 3984
rect 7420 4040 7484 4044
rect 7420 3984 7470 4040
rect 7470 3984 7484 4040
rect 7420 3980 7484 3984
rect 11468 3980 11532 4044
rect 2826 3836 2890 3840
rect 2826 3780 2830 3836
rect 2830 3780 2886 3836
rect 2886 3780 2890 3836
rect 2826 3776 2890 3780
rect 2906 3836 2970 3840
rect 2906 3780 2910 3836
rect 2910 3780 2966 3836
rect 2966 3780 2970 3836
rect 2906 3776 2970 3780
rect 2986 3836 3050 3840
rect 2986 3780 2990 3836
rect 2990 3780 3046 3836
rect 3046 3780 3050 3836
rect 2986 3776 3050 3780
rect 3066 3836 3130 3840
rect 3066 3780 3070 3836
rect 3070 3780 3126 3836
rect 3126 3780 3130 3836
rect 3066 3776 3130 3780
rect 3372 3572 3436 3636
rect 7972 3904 8036 3908
rect 7972 3848 8022 3904
rect 8022 3848 8036 3904
rect 7972 3844 8036 3848
rect 10916 3844 10980 3908
rect 6574 3836 6638 3840
rect 6574 3780 6578 3836
rect 6578 3780 6634 3836
rect 6634 3780 6638 3836
rect 6574 3776 6638 3780
rect 6654 3836 6718 3840
rect 6654 3780 6658 3836
rect 6658 3780 6714 3836
rect 6714 3780 6718 3836
rect 6654 3776 6718 3780
rect 6734 3836 6798 3840
rect 6734 3780 6738 3836
rect 6738 3780 6794 3836
rect 6794 3780 6798 3836
rect 6734 3776 6798 3780
rect 6814 3836 6878 3840
rect 6814 3780 6818 3836
rect 6818 3780 6874 3836
rect 6874 3780 6878 3836
rect 6814 3776 6878 3780
rect 10322 3836 10386 3840
rect 10322 3780 10326 3836
rect 10326 3780 10382 3836
rect 10382 3780 10386 3836
rect 10322 3776 10386 3780
rect 10402 3836 10466 3840
rect 10402 3780 10406 3836
rect 10406 3780 10462 3836
rect 10462 3780 10466 3836
rect 10402 3776 10466 3780
rect 10482 3836 10546 3840
rect 10482 3780 10486 3836
rect 10486 3780 10542 3836
rect 10542 3780 10546 3836
rect 10482 3776 10546 3780
rect 10562 3836 10626 3840
rect 10562 3780 10566 3836
rect 10566 3780 10622 3836
rect 10622 3780 10626 3836
rect 10562 3776 10626 3780
rect 7420 3768 7484 3772
rect 7420 3712 7434 3768
rect 7434 3712 7484 3768
rect 7420 3708 7484 3712
rect 12756 3708 12820 3772
rect 6132 3572 6196 3636
rect 8156 3572 8220 3636
rect 4700 3292 4764 3296
rect 4700 3236 4704 3292
rect 4704 3236 4760 3292
rect 4760 3236 4764 3292
rect 4700 3232 4764 3236
rect 4780 3292 4844 3296
rect 4780 3236 4784 3292
rect 4784 3236 4840 3292
rect 4840 3236 4844 3292
rect 4780 3232 4844 3236
rect 4860 3292 4924 3296
rect 4860 3236 4864 3292
rect 4864 3236 4920 3292
rect 4920 3236 4924 3292
rect 4860 3232 4924 3236
rect 4940 3292 5004 3296
rect 4940 3236 4944 3292
rect 4944 3236 5000 3292
rect 5000 3236 5004 3292
rect 4940 3232 5004 3236
rect 9444 3572 9508 3636
rect 11284 3572 11348 3636
rect 14070 3836 14134 3840
rect 14070 3780 14074 3836
rect 14074 3780 14130 3836
rect 14130 3780 14134 3836
rect 14070 3776 14134 3780
rect 14150 3836 14214 3840
rect 14150 3780 14154 3836
rect 14154 3780 14210 3836
rect 14210 3780 14214 3836
rect 14150 3776 14214 3780
rect 14230 3836 14294 3840
rect 14230 3780 14234 3836
rect 14234 3780 14290 3836
rect 14290 3780 14294 3836
rect 14230 3776 14294 3780
rect 14310 3836 14374 3840
rect 14310 3780 14314 3836
rect 14314 3780 14370 3836
rect 14370 3780 14374 3836
rect 14310 3776 14374 3780
rect 11652 3436 11716 3500
rect 14596 3436 14660 3500
rect 12940 3300 13004 3364
rect 14780 3300 14844 3364
rect 8448 3292 8512 3296
rect 8448 3236 8452 3292
rect 8452 3236 8508 3292
rect 8508 3236 8512 3292
rect 8448 3232 8512 3236
rect 8528 3292 8592 3296
rect 8528 3236 8532 3292
rect 8532 3236 8588 3292
rect 8588 3236 8592 3292
rect 8528 3232 8592 3236
rect 8608 3292 8672 3296
rect 8608 3236 8612 3292
rect 8612 3236 8668 3292
rect 8668 3236 8672 3292
rect 8608 3232 8672 3236
rect 8688 3292 8752 3296
rect 8688 3236 8692 3292
rect 8692 3236 8748 3292
rect 8748 3236 8752 3292
rect 8688 3232 8752 3236
rect 12196 3292 12260 3296
rect 12196 3236 12200 3292
rect 12200 3236 12256 3292
rect 12256 3236 12260 3292
rect 12196 3232 12260 3236
rect 12276 3292 12340 3296
rect 12276 3236 12280 3292
rect 12280 3236 12336 3292
rect 12336 3236 12340 3292
rect 12276 3232 12340 3236
rect 12356 3292 12420 3296
rect 12356 3236 12360 3292
rect 12360 3236 12416 3292
rect 12416 3236 12420 3292
rect 12356 3232 12420 3236
rect 12436 3292 12500 3296
rect 12436 3236 12440 3292
rect 12440 3236 12496 3292
rect 12496 3236 12500 3292
rect 12436 3232 12500 3236
rect 12756 3164 12820 3228
rect 5580 2756 5644 2820
rect 7236 3088 7300 3092
rect 7236 3032 7286 3088
rect 7286 3032 7300 3088
rect 7236 3028 7300 3032
rect 9812 3028 9876 3092
rect 11100 3028 11164 3092
rect 11836 3088 11900 3092
rect 11836 3032 11850 3088
rect 11850 3032 11900 3088
rect 11836 3028 11900 3032
rect 12020 3028 12084 3092
rect 13124 3028 13188 3092
rect 15332 3028 15396 3092
rect 2826 2748 2890 2752
rect 2826 2692 2830 2748
rect 2830 2692 2886 2748
rect 2886 2692 2890 2748
rect 2826 2688 2890 2692
rect 2906 2748 2970 2752
rect 2906 2692 2910 2748
rect 2910 2692 2966 2748
rect 2966 2692 2970 2748
rect 2906 2688 2970 2692
rect 2986 2748 3050 2752
rect 2986 2692 2990 2748
rect 2990 2692 3046 2748
rect 3046 2692 3050 2748
rect 2986 2688 3050 2692
rect 3066 2748 3130 2752
rect 3066 2692 3070 2748
rect 3070 2692 3126 2748
rect 3126 2692 3130 2748
rect 3066 2688 3130 2692
rect 6574 2748 6638 2752
rect 6574 2692 6578 2748
rect 6578 2692 6634 2748
rect 6634 2692 6638 2748
rect 6574 2688 6638 2692
rect 6654 2748 6718 2752
rect 6654 2692 6658 2748
rect 6658 2692 6714 2748
rect 6714 2692 6718 2748
rect 6654 2688 6718 2692
rect 6734 2748 6798 2752
rect 6734 2692 6738 2748
rect 6738 2692 6794 2748
rect 6794 2692 6798 2748
rect 6734 2688 6798 2692
rect 6814 2748 6878 2752
rect 6814 2692 6818 2748
rect 6818 2692 6874 2748
rect 6874 2692 6878 2748
rect 6814 2688 6878 2692
rect 5948 2620 6012 2684
rect 7052 2620 7116 2684
rect 7420 2680 7484 2684
rect 7420 2624 7434 2680
rect 7434 2624 7484 2680
rect 7420 2620 7484 2624
rect 5212 2484 5276 2548
rect 5948 2484 6012 2548
rect 8892 2544 8956 2548
rect 8892 2488 8906 2544
rect 8906 2488 8956 2544
rect 8892 2484 8956 2488
rect 12572 2756 12636 2820
rect 13860 2816 13924 2820
rect 13860 2760 13910 2816
rect 13910 2760 13924 2816
rect 13860 2756 13924 2760
rect 10322 2748 10386 2752
rect 10322 2692 10326 2748
rect 10326 2692 10382 2748
rect 10382 2692 10386 2748
rect 10322 2688 10386 2692
rect 10402 2748 10466 2752
rect 10402 2692 10406 2748
rect 10406 2692 10462 2748
rect 10462 2692 10466 2748
rect 10402 2688 10466 2692
rect 10482 2748 10546 2752
rect 10482 2692 10486 2748
rect 10486 2692 10542 2748
rect 10542 2692 10546 2748
rect 10482 2688 10546 2692
rect 10562 2748 10626 2752
rect 10562 2692 10566 2748
rect 10566 2692 10622 2748
rect 10622 2692 10626 2748
rect 10562 2688 10626 2692
rect 14070 2748 14134 2752
rect 14070 2692 14074 2748
rect 14074 2692 14130 2748
rect 14130 2692 14134 2748
rect 14070 2688 14134 2692
rect 14150 2748 14214 2752
rect 14150 2692 14154 2748
rect 14154 2692 14210 2748
rect 14210 2692 14214 2748
rect 14150 2688 14214 2692
rect 14230 2748 14294 2752
rect 14230 2692 14234 2748
rect 14234 2692 14290 2748
rect 14290 2692 14294 2748
rect 14230 2688 14294 2692
rect 14310 2748 14374 2752
rect 14310 2692 14314 2748
rect 14314 2692 14370 2748
rect 14370 2692 14374 2748
rect 14310 2688 14374 2692
rect 13492 2484 13556 2548
rect 4292 2348 4356 2412
rect 14596 2348 14660 2412
rect 13676 2212 13740 2276
rect 4700 2204 4764 2208
rect 4700 2148 4704 2204
rect 4704 2148 4760 2204
rect 4760 2148 4764 2204
rect 4700 2144 4764 2148
rect 4780 2204 4844 2208
rect 4780 2148 4784 2204
rect 4784 2148 4840 2204
rect 4840 2148 4844 2204
rect 4780 2144 4844 2148
rect 4860 2204 4924 2208
rect 4860 2148 4864 2204
rect 4864 2148 4920 2204
rect 4920 2148 4924 2204
rect 4860 2144 4924 2148
rect 4940 2204 5004 2208
rect 4940 2148 4944 2204
rect 4944 2148 5000 2204
rect 5000 2148 5004 2204
rect 4940 2144 5004 2148
rect 8448 2204 8512 2208
rect 8448 2148 8452 2204
rect 8452 2148 8508 2204
rect 8508 2148 8512 2204
rect 8448 2144 8512 2148
rect 8528 2204 8592 2208
rect 8528 2148 8532 2204
rect 8532 2148 8588 2204
rect 8588 2148 8592 2204
rect 8528 2144 8592 2148
rect 8608 2204 8672 2208
rect 8608 2148 8612 2204
rect 8612 2148 8668 2204
rect 8668 2148 8672 2204
rect 8608 2144 8672 2148
rect 8688 2204 8752 2208
rect 8688 2148 8692 2204
rect 8692 2148 8748 2204
rect 8748 2148 8752 2204
rect 8688 2144 8752 2148
rect 12196 2204 12260 2208
rect 12196 2148 12200 2204
rect 12200 2148 12256 2204
rect 12256 2148 12260 2204
rect 12196 2144 12260 2148
rect 12276 2204 12340 2208
rect 12276 2148 12280 2204
rect 12280 2148 12336 2204
rect 12336 2148 12340 2204
rect 12276 2144 12340 2148
rect 12356 2204 12420 2208
rect 12356 2148 12360 2204
rect 12360 2148 12416 2204
rect 12416 2148 12420 2204
rect 12356 2144 12420 2148
rect 12436 2204 12500 2208
rect 12436 2148 12440 2204
rect 12440 2148 12496 2204
rect 12496 2148 12500 2204
rect 12436 2144 12500 2148
rect 3924 1940 3988 2004
rect 9260 1940 9324 2004
<< metal4 >>
rect 2818 16896 3138 17456
rect 2818 16832 2826 16896
rect 2890 16832 2906 16896
rect 2970 16832 2986 16896
rect 3050 16832 3066 16896
rect 3130 16832 3138 16896
rect 2818 15808 3138 16832
rect 2818 15744 2826 15808
rect 2890 15744 2906 15808
rect 2970 15744 2986 15808
rect 3050 15744 3066 15808
rect 3130 15744 3138 15808
rect 1715 15332 1781 15333
rect 1715 15268 1716 15332
rect 1780 15268 1781 15332
rect 1715 15267 1781 15268
rect 2451 15332 2517 15333
rect 2451 15268 2452 15332
rect 2516 15268 2517 15332
rect 2451 15267 2517 15268
rect 1718 4045 1778 15267
rect 2454 4861 2514 15267
rect 2818 14720 3138 15744
rect 2818 14656 2826 14720
rect 2890 14656 2906 14720
rect 2970 14656 2986 14720
rect 3050 14656 3066 14720
rect 3130 14656 3138 14720
rect 2818 13632 3138 14656
rect 4692 17440 5012 17456
rect 4692 17376 4700 17440
rect 4764 17376 4780 17440
rect 4844 17376 4860 17440
rect 4924 17376 4940 17440
rect 5004 17376 5012 17440
rect 4692 16352 5012 17376
rect 4692 16288 4700 16352
rect 4764 16288 4780 16352
rect 4844 16288 4860 16352
rect 4924 16288 4940 16352
rect 5004 16288 5012 16352
rect 4692 15264 5012 16288
rect 6566 16896 6886 17456
rect 6566 16832 6574 16896
rect 6638 16832 6654 16896
rect 6718 16832 6734 16896
rect 6798 16832 6814 16896
rect 6878 16832 6886 16896
rect 6566 15808 6886 16832
rect 6566 15744 6574 15808
rect 6638 15744 6654 15808
rect 6718 15744 6734 15808
rect 6798 15744 6814 15808
rect 6878 15744 6886 15808
rect 6315 15332 6381 15333
rect 6315 15268 6316 15332
rect 6380 15268 6381 15332
rect 6315 15267 6381 15268
rect 4692 15200 4700 15264
rect 4764 15200 4780 15264
rect 4844 15200 4860 15264
rect 4924 15200 4940 15264
rect 5004 15200 5012 15264
rect 4107 14244 4173 14245
rect 4107 14180 4108 14244
rect 4172 14180 4173 14244
rect 4107 14179 4173 14180
rect 2818 13568 2826 13632
rect 2890 13568 2906 13632
rect 2970 13568 2986 13632
rect 3050 13568 3066 13632
rect 3130 13568 3138 13632
rect 2818 12544 3138 13568
rect 2818 12480 2826 12544
rect 2890 12480 2906 12544
rect 2970 12480 2986 12544
rect 3050 12480 3066 12544
rect 3130 12480 3138 12544
rect 2818 11456 3138 12480
rect 2818 11392 2826 11456
rect 2890 11392 2906 11456
rect 2970 11392 2986 11456
rect 3050 11392 3066 11456
rect 3130 11392 3138 11456
rect 2818 10368 3138 11392
rect 2818 10304 2826 10368
rect 2890 10304 2906 10368
rect 2970 10304 2986 10368
rect 3050 10304 3066 10368
rect 3130 10304 3138 10368
rect 2818 9280 3138 10304
rect 4110 9621 4170 14179
rect 4692 14176 5012 15200
rect 4692 14112 4700 14176
rect 4764 14112 4780 14176
rect 4844 14112 4860 14176
rect 4924 14112 4940 14176
rect 5004 14112 5012 14176
rect 4692 13088 5012 14112
rect 4692 13024 4700 13088
rect 4764 13024 4780 13088
rect 4844 13024 4860 13088
rect 4924 13024 4940 13088
rect 5004 13024 5012 13088
rect 4692 12000 5012 13024
rect 6131 12612 6197 12613
rect 6131 12548 6132 12612
rect 6196 12548 6197 12612
rect 6131 12547 6197 12548
rect 4692 11936 4700 12000
rect 4764 11936 4780 12000
rect 4844 11936 4860 12000
rect 4924 11936 4940 12000
rect 5004 11936 5012 12000
rect 4692 10912 5012 11936
rect 4692 10848 4700 10912
rect 4764 10848 4780 10912
rect 4844 10848 4860 10912
rect 4924 10848 4940 10912
rect 5004 10848 5012 10912
rect 4692 9824 5012 10848
rect 4692 9760 4700 9824
rect 4764 9760 4780 9824
rect 4844 9760 4860 9824
rect 4924 9760 4940 9824
rect 5004 9760 5012 9824
rect 4107 9620 4173 9621
rect 4107 9556 4108 9620
rect 4172 9556 4173 9620
rect 4107 9555 4173 9556
rect 2818 9216 2826 9280
rect 2890 9216 2906 9280
rect 2970 9216 2986 9280
rect 3050 9216 3066 9280
rect 3130 9216 3138 9280
rect 2818 8192 3138 9216
rect 2818 8128 2826 8192
rect 2890 8128 2906 8192
rect 2970 8128 2986 8192
rect 3050 8128 3066 8192
rect 3130 8128 3138 8192
rect 2818 7104 3138 8128
rect 2818 7040 2826 7104
rect 2890 7040 2906 7104
rect 2970 7040 2986 7104
rect 3050 7040 3066 7104
rect 3130 7040 3138 7104
rect 2818 6016 3138 7040
rect 4692 8736 5012 9760
rect 5395 9076 5461 9077
rect 5395 9012 5396 9076
rect 5460 9012 5461 9076
rect 5395 9011 5461 9012
rect 4692 8672 4700 8736
rect 4764 8672 4780 8736
rect 4844 8672 4860 8736
rect 4924 8672 4940 8736
rect 5004 8672 5012 8736
rect 4692 7648 5012 8672
rect 4692 7584 4700 7648
rect 4764 7584 4780 7648
rect 4844 7584 4860 7648
rect 4924 7584 4940 7648
rect 5004 7584 5012 7648
rect 4692 6560 5012 7584
rect 4692 6496 4700 6560
rect 4764 6496 4780 6560
rect 4844 6496 4860 6560
rect 4924 6496 4940 6560
rect 5004 6496 5012 6560
rect 3739 6492 3805 6493
rect 3739 6428 3740 6492
rect 3804 6428 3805 6492
rect 3739 6427 3805 6428
rect 2818 5952 2826 6016
rect 2890 5952 2906 6016
rect 2970 5952 2986 6016
rect 3050 5952 3066 6016
rect 3130 5952 3138 6016
rect 2818 4928 3138 5952
rect 3371 5948 3437 5949
rect 3371 5884 3372 5948
rect 3436 5884 3437 5948
rect 3371 5883 3437 5884
rect 2818 4864 2826 4928
rect 2890 4864 2906 4928
rect 2970 4864 2986 4928
rect 3050 4864 3066 4928
rect 3130 4864 3138 4928
rect 2451 4860 2517 4861
rect 2451 4796 2452 4860
rect 2516 4796 2517 4860
rect 2451 4795 2517 4796
rect 1715 4044 1781 4045
rect 1715 3980 1716 4044
rect 1780 3980 1781 4044
rect 1715 3979 1781 3980
rect 2818 3840 3138 4864
rect 2818 3776 2826 3840
rect 2890 3776 2906 3840
rect 2970 3776 2986 3840
rect 3050 3776 3066 3840
rect 3130 3776 3138 3840
rect 2818 2752 3138 3776
rect 3374 3637 3434 5883
rect 3742 4861 3802 6427
rect 4475 6220 4541 6221
rect 4475 6156 4476 6220
rect 4540 6156 4541 6220
rect 4475 6155 4541 6156
rect 3739 4860 3805 4861
rect 3739 4796 3740 4860
rect 3804 4796 3805 4860
rect 3739 4795 3805 4796
rect 3923 4860 3989 4861
rect 3923 4796 3924 4860
rect 3988 4796 3989 4860
rect 3923 4795 3989 4796
rect 3371 3636 3437 3637
rect 3371 3572 3372 3636
rect 3436 3572 3437 3636
rect 3371 3571 3437 3572
rect 2818 2688 2826 2752
rect 2890 2688 2906 2752
rect 2970 2688 2986 2752
rect 3050 2688 3066 2752
rect 3130 2688 3138 2752
rect 2818 2128 3138 2688
rect 3926 2005 3986 4795
rect 4291 4588 4357 4589
rect 4291 4524 4292 4588
rect 4356 4524 4357 4588
rect 4291 4523 4357 4524
rect 4294 2413 4354 4523
rect 4478 4453 4538 6155
rect 4692 5472 5012 6496
rect 5211 5676 5277 5677
rect 5211 5612 5212 5676
rect 5276 5612 5277 5676
rect 5211 5611 5277 5612
rect 4692 5408 4700 5472
rect 4764 5408 4780 5472
rect 4844 5408 4860 5472
rect 4924 5408 4940 5472
rect 5004 5408 5012 5472
rect 4475 4452 4541 4453
rect 4475 4388 4476 4452
rect 4540 4388 4541 4452
rect 4475 4387 4541 4388
rect 4692 4384 5012 5408
rect 4692 4320 4700 4384
rect 4764 4320 4780 4384
rect 4844 4320 4860 4384
rect 4924 4320 4940 4384
rect 5004 4320 5012 4384
rect 4692 3296 5012 4320
rect 4692 3232 4700 3296
rect 4764 3232 4780 3296
rect 4844 3232 4860 3296
rect 4924 3232 4940 3296
rect 5004 3232 5012 3296
rect 4291 2412 4357 2413
rect 4291 2348 4292 2412
rect 4356 2348 4357 2412
rect 4291 2347 4357 2348
rect 4692 2208 5012 3232
rect 5214 2549 5274 5611
rect 5398 5269 5458 9011
rect 5947 7444 6013 7445
rect 5947 7380 5948 7444
rect 6012 7380 6013 7444
rect 5947 7379 6013 7380
rect 5395 5268 5461 5269
rect 5395 5204 5396 5268
rect 5460 5204 5461 5268
rect 5395 5203 5461 5204
rect 5579 2820 5645 2821
rect 5579 2756 5580 2820
rect 5644 2756 5645 2820
rect 5579 2755 5645 2756
rect 5211 2548 5277 2549
rect 5211 2484 5212 2548
rect 5276 2484 5277 2548
rect 5211 2483 5277 2484
rect 5582 2410 5642 2755
rect 5950 2685 6010 7379
rect 6134 6901 6194 12547
rect 6131 6900 6197 6901
rect 6131 6836 6132 6900
rect 6196 6836 6197 6900
rect 6131 6835 6197 6836
rect 6131 5540 6197 5541
rect 6131 5476 6132 5540
rect 6196 5476 6197 5540
rect 6131 5475 6197 5476
rect 6134 3637 6194 5475
rect 6318 4861 6378 15267
rect 6566 14720 6886 15744
rect 6566 14656 6574 14720
rect 6638 14656 6654 14720
rect 6718 14656 6734 14720
rect 6798 14656 6814 14720
rect 6878 14656 6886 14720
rect 6566 13632 6886 14656
rect 8440 17440 8760 17456
rect 8440 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8760 17440
rect 8440 16352 8760 17376
rect 10314 16896 10634 17456
rect 12188 17440 12508 17456
rect 12188 17376 12196 17440
rect 12260 17376 12276 17440
rect 12340 17376 12356 17440
rect 12420 17376 12436 17440
rect 12500 17376 12508 17440
rect 11467 17236 11533 17237
rect 11467 17172 11468 17236
rect 11532 17172 11533 17236
rect 11467 17171 11533 17172
rect 10314 16832 10322 16896
rect 10386 16832 10402 16896
rect 10466 16832 10482 16896
rect 10546 16832 10562 16896
rect 10626 16832 10634 16896
rect 9811 16692 9877 16693
rect 9811 16628 9812 16692
rect 9876 16628 9877 16692
rect 9811 16627 9877 16628
rect 8440 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8760 16352
rect 8440 15264 8760 16288
rect 8440 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8760 15264
rect 7419 14244 7485 14245
rect 7419 14180 7420 14244
rect 7484 14180 7485 14244
rect 7419 14179 7485 14180
rect 6566 13568 6574 13632
rect 6638 13568 6654 13632
rect 6718 13568 6734 13632
rect 6798 13568 6814 13632
rect 6878 13568 6886 13632
rect 6566 12544 6886 13568
rect 6566 12480 6574 12544
rect 6638 12480 6654 12544
rect 6718 12480 6734 12544
rect 6798 12480 6814 12544
rect 6878 12480 6886 12544
rect 6566 11456 6886 12480
rect 6566 11392 6574 11456
rect 6638 11392 6654 11456
rect 6718 11392 6734 11456
rect 6798 11392 6814 11456
rect 6878 11392 6886 11456
rect 6566 10368 6886 11392
rect 6566 10304 6574 10368
rect 6638 10304 6654 10368
rect 6718 10304 6734 10368
rect 6798 10304 6814 10368
rect 6878 10304 6886 10368
rect 6566 9280 6886 10304
rect 6566 9216 6574 9280
rect 6638 9216 6654 9280
rect 6718 9216 6734 9280
rect 6798 9216 6814 9280
rect 6878 9216 6886 9280
rect 6566 8192 6886 9216
rect 6566 8128 6574 8192
rect 6638 8128 6654 8192
rect 6718 8128 6734 8192
rect 6798 8128 6814 8192
rect 6878 8128 6886 8192
rect 6566 7104 6886 8128
rect 6566 7040 6574 7104
rect 6638 7040 6654 7104
rect 6718 7040 6734 7104
rect 6798 7040 6814 7104
rect 6878 7040 6886 7104
rect 6566 6016 6886 7040
rect 7235 6628 7301 6629
rect 7235 6564 7236 6628
rect 7300 6564 7301 6628
rect 7235 6563 7301 6564
rect 6566 5952 6574 6016
rect 6638 5952 6654 6016
rect 6718 5952 6734 6016
rect 6798 5952 6814 6016
rect 6878 5952 6886 6016
rect 6566 4928 6886 5952
rect 7051 5540 7117 5541
rect 7051 5476 7052 5540
rect 7116 5476 7117 5540
rect 7051 5475 7117 5476
rect 6566 4864 6574 4928
rect 6638 4864 6654 4928
rect 6718 4864 6734 4928
rect 6798 4864 6814 4928
rect 6878 4864 6886 4928
rect 6315 4860 6381 4861
rect 6315 4796 6316 4860
rect 6380 4796 6381 4860
rect 6315 4795 6381 4796
rect 6566 3840 6886 4864
rect 6566 3776 6574 3840
rect 6638 3776 6654 3840
rect 6718 3776 6734 3840
rect 6798 3776 6814 3840
rect 6878 3776 6886 3840
rect 6131 3636 6197 3637
rect 6131 3572 6132 3636
rect 6196 3572 6197 3636
rect 6131 3571 6197 3572
rect 6566 2752 6886 3776
rect 6566 2688 6574 2752
rect 6638 2688 6654 2752
rect 6718 2688 6734 2752
rect 6798 2688 6814 2752
rect 6878 2688 6886 2752
rect 5947 2684 6013 2685
rect 5947 2620 5948 2684
rect 6012 2620 6013 2684
rect 5947 2619 6013 2620
rect 5947 2548 6013 2549
rect 5947 2484 5948 2548
rect 6012 2484 6013 2548
rect 5947 2483 6013 2484
rect 5950 2410 6010 2483
rect 5582 2350 6010 2410
rect 4692 2144 4700 2208
rect 4764 2144 4780 2208
rect 4844 2144 4860 2208
rect 4924 2144 4940 2208
rect 5004 2144 5012 2208
rect 4692 2128 5012 2144
rect 6566 2128 6886 2688
rect 7054 2685 7114 5475
rect 7238 3093 7298 6563
rect 7422 4045 7482 14179
rect 8440 14176 8760 15200
rect 9814 15210 9874 16627
rect 10314 15808 10634 16832
rect 10314 15744 10322 15808
rect 10386 15744 10402 15808
rect 10466 15744 10482 15808
rect 10546 15744 10562 15808
rect 10626 15744 10634 15808
rect 9814 15150 10058 15210
rect 8440 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8760 14176
rect 8440 13088 8760 14112
rect 9259 13836 9325 13837
rect 9259 13772 9260 13836
rect 9324 13772 9325 13836
rect 9259 13771 9325 13772
rect 8440 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8760 13088
rect 8440 12000 8760 13024
rect 8891 12748 8957 12749
rect 8891 12684 8892 12748
rect 8956 12684 8957 12748
rect 8891 12683 8957 12684
rect 8440 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8760 12000
rect 8440 10912 8760 11936
rect 8440 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8760 10912
rect 8440 9824 8760 10848
rect 8440 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8760 9824
rect 7971 9212 8037 9213
rect 7971 9148 7972 9212
rect 8036 9148 8037 9212
rect 7971 9147 8037 9148
rect 7603 6764 7669 6765
rect 7603 6700 7604 6764
rect 7668 6700 7669 6764
rect 7603 6699 7669 6700
rect 7787 6764 7853 6765
rect 7787 6700 7788 6764
rect 7852 6700 7853 6764
rect 7787 6699 7853 6700
rect 7606 6085 7666 6699
rect 7603 6084 7669 6085
rect 7603 6020 7604 6084
rect 7668 6020 7669 6084
rect 7603 6019 7669 6020
rect 7790 5405 7850 6699
rect 7787 5404 7853 5405
rect 7787 5340 7788 5404
rect 7852 5340 7853 5404
rect 7787 5339 7853 5340
rect 7419 4044 7485 4045
rect 7419 3980 7420 4044
rect 7484 3980 7485 4044
rect 7419 3979 7485 3980
rect 7974 3909 8034 9147
rect 8155 8804 8221 8805
rect 8155 8740 8156 8804
rect 8220 8740 8221 8804
rect 8155 8739 8221 8740
rect 7971 3908 8037 3909
rect 7971 3844 7972 3908
rect 8036 3844 8037 3908
rect 7971 3843 8037 3844
rect 7419 3772 7485 3773
rect 7419 3708 7420 3772
rect 7484 3708 7485 3772
rect 7419 3707 7485 3708
rect 7235 3092 7301 3093
rect 7235 3028 7236 3092
rect 7300 3028 7301 3092
rect 7235 3027 7301 3028
rect 7422 2685 7482 3707
rect 8158 3637 8218 8739
rect 8440 8736 8760 9760
rect 8894 9077 8954 12683
rect 8891 9076 8957 9077
rect 8891 9012 8892 9076
rect 8956 9012 8957 9076
rect 8891 9011 8957 9012
rect 8440 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8760 8736
rect 8440 7648 8760 8672
rect 8440 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8760 7648
rect 8440 6560 8760 7584
rect 8891 7580 8957 7581
rect 8891 7516 8892 7580
rect 8956 7516 8957 7580
rect 8891 7515 8957 7516
rect 8440 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8760 6560
rect 8440 5472 8760 6496
rect 8440 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8760 5472
rect 8440 4384 8760 5408
rect 8440 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8760 4384
rect 8155 3636 8221 3637
rect 8155 3572 8156 3636
rect 8220 3572 8221 3636
rect 8155 3571 8221 3572
rect 8440 3296 8760 4320
rect 8440 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8760 3296
rect 7051 2684 7117 2685
rect 7051 2620 7052 2684
rect 7116 2620 7117 2684
rect 7051 2619 7117 2620
rect 7419 2684 7485 2685
rect 7419 2620 7420 2684
rect 7484 2620 7485 2684
rect 7419 2619 7485 2620
rect 8440 2208 8760 3232
rect 8894 2549 8954 7515
rect 9262 6629 9322 13771
rect 9443 12340 9509 12341
rect 9443 12276 9444 12340
rect 9508 12276 9509 12340
rect 9443 12275 9509 12276
rect 9259 6628 9325 6629
rect 9259 6564 9260 6628
rect 9324 6564 9325 6628
rect 9259 6563 9325 6564
rect 9262 6085 9322 6563
rect 9259 6084 9325 6085
rect 9259 6020 9260 6084
rect 9324 6020 9325 6084
rect 9259 6019 9325 6020
rect 9259 5540 9325 5541
rect 9259 5476 9260 5540
rect 9324 5476 9325 5540
rect 9259 5475 9325 5476
rect 8891 2548 8957 2549
rect 8891 2484 8892 2548
rect 8956 2484 8957 2548
rect 8891 2483 8957 2484
rect 8440 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8760 2208
rect 8440 2128 8760 2144
rect 9262 2005 9322 5475
rect 9446 3637 9506 12275
rect 9811 12204 9877 12205
rect 9811 12140 9812 12204
rect 9876 12140 9877 12204
rect 9811 12139 9877 12140
rect 9814 8533 9874 12139
rect 9811 8532 9877 8533
rect 9811 8468 9812 8532
rect 9876 8468 9877 8532
rect 9811 8467 9877 8468
rect 9627 8124 9693 8125
rect 9627 8060 9628 8124
rect 9692 8060 9693 8124
rect 9627 8059 9693 8060
rect 9630 5813 9690 8059
rect 9857 7036 9923 7037
rect 9857 7034 9858 7036
rect 9814 6972 9858 7034
rect 9922 6972 9923 7036
rect 9814 6971 9923 6972
rect 9627 5812 9693 5813
rect 9627 5748 9628 5812
rect 9692 5748 9693 5812
rect 9627 5747 9693 5748
rect 9627 5404 9693 5405
rect 9627 5340 9628 5404
rect 9692 5340 9693 5404
rect 9627 5339 9693 5340
rect 9630 5130 9690 5339
rect 9814 5269 9874 6971
rect 9998 6765 10058 15150
rect 10314 14720 10634 15744
rect 10314 14656 10322 14720
rect 10386 14656 10402 14720
rect 10466 14656 10482 14720
rect 10546 14656 10562 14720
rect 10626 14656 10634 14720
rect 10314 13632 10634 14656
rect 10314 13568 10322 13632
rect 10386 13568 10402 13632
rect 10466 13568 10482 13632
rect 10546 13568 10562 13632
rect 10626 13568 10634 13632
rect 10314 12544 10634 13568
rect 10314 12480 10322 12544
rect 10386 12480 10402 12544
rect 10466 12480 10482 12544
rect 10546 12480 10562 12544
rect 10626 12480 10634 12544
rect 10179 11932 10245 11933
rect 10179 11868 10180 11932
rect 10244 11868 10245 11932
rect 10179 11867 10245 11868
rect 10182 7309 10242 11867
rect 10314 11456 10634 12480
rect 10915 12340 10981 12341
rect 10915 12276 10916 12340
rect 10980 12276 10981 12340
rect 10915 12275 10981 12276
rect 10314 11392 10322 11456
rect 10386 11392 10402 11456
rect 10466 11392 10482 11456
rect 10546 11392 10562 11456
rect 10626 11392 10634 11456
rect 10314 10368 10634 11392
rect 10314 10304 10322 10368
rect 10386 10304 10402 10368
rect 10466 10304 10482 10368
rect 10546 10304 10562 10368
rect 10626 10304 10634 10368
rect 10314 9280 10634 10304
rect 10314 9216 10322 9280
rect 10386 9216 10402 9280
rect 10466 9216 10482 9280
rect 10546 9216 10562 9280
rect 10626 9216 10634 9280
rect 10314 8192 10634 9216
rect 10314 8128 10322 8192
rect 10386 8128 10402 8192
rect 10466 8128 10482 8192
rect 10546 8128 10562 8192
rect 10626 8128 10634 8192
rect 10179 7308 10245 7309
rect 10179 7244 10180 7308
rect 10244 7244 10245 7308
rect 10179 7243 10245 7244
rect 9995 6764 10061 6765
rect 9995 6700 9996 6764
rect 10060 6700 10061 6764
rect 9995 6699 10061 6700
rect 9811 5268 9877 5269
rect 9811 5204 9812 5268
rect 9876 5204 9877 5268
rect 9811 5203 9877 5204
rect 9630 5070 9874 5130
rect 9627 4860 9693 4861
rect 9627 4796 9628 4860
rect 9692 4796 9693 4860
rect 9627 4795 9693 4796
rect 9630 4317 9690 4795
rect 9627 4316 9693 4317
rect 9627 4252 9628 4316
rect 9692 4252 9693 4316
rect 9627 4251 9693 4252
rect 9443 3636 9509 3637
rect 9443 3572 9444 3636
rect 9508 3572 9509 3636
rect 9443 3571 9509 3572
rect 9814 3093 9874 5070
rect 9998 4861 10058 6699
rect 10182 5269 10242 7243
rect 10314 7104 10634 8128
rect 10731 7988 10797 7989
rect 10731 7924 10732 7988
rect 10796 7924 10797 7988
rect 10731 7923 10797 7924
rect 10314 7040 10322 7104
rect 10386 7040 10402 7104
rect 10466 7040 10482 7104
rect 10546 7040 10562 7104
rect 10626 7040 10634 7104
rect 10314 6016 10634 7040
rect 10314 5952 10322 6016
rect 10386 5952 10402 6016
rect 10466 5952 10482 6016
rect 10546 5952 10562 6016
rect 10626 5952 10634 6016
rect 10179 5268 10245 5269
rect 10179 5204 10180 5268
rect 10244 5204 10245 5268
rect 10179 5203 10245 5204
rect 10314 4928 10634 5952
rect 10314 4864 10322 4928
rect 10386 4864 10402 4928
rect 10466 4864 10482 4928
rect 10546 4864 10562 4928
rect 10626 4864 10634 4928
rect 9995 4860 10061 4861
rect 9995 4796 9996 4860
rect 10060 4796 10061 4860
rect 9995 4795 10061 4796
rect 10314 3840 10634 4864
rect 10734 4317 10794 7923
rect 10731 4316 10797 4317
rect 10731 4252 10732 4316
rect 10796 4252 10797 4316
rect 10731 4251 10797 4252
rect 10918 3909 10978 12275
rect 11470 11933 11530 17171
rect 12188 16352 12508 17376
rect 14062 16896 14382 17456
rect 14062 16832 14070 16896
rect 14134 16832 14150 16896
rect 14214 16832 14230 16896
rect 14294 16832 14310 16896
rect 14374 16832 14382 16896
rect 13675 16828 13741 16829
rect 13675 16764 13676 16828
rect 13740 16764 13741 16828
rect 13675 16763 13741 16764
rect 13491 16692 13557 16693
rect 13491 16628 13492 16692
rect 13556 16628 13557 16692
rect 13491 16627 13557 16628
rect 12755 16556 12821 16557
rect 12755 16492 12756 16556
rect 12820 16492 12821 16556
rect 12755 16491 12821 16492
rect 12188 16288 12196 16352
rect 12260 16288 12276 16352
rect 12340 16288 12356 16352
rect 12420 16288 12436 16352
rect 12500 16288 12508 16352
rect 12188 15264 12508 16288
rect 12188 15200 12196 15264
rect 12260 15200 12276 15264
rect 12340 15200 12356 15264
rect 12420 15200 12436 15264
rect 12500 15200 12508 15264
rect 12019 14924 12085 14925
rect 12019 14860 12020 14924
rect 12084 14860 12085 14924
rect 12019 14859 12085 14860
rect 12022 13565 12082 14859
rect 12188 14176 12508 15200
rect 12188 14112 12196 14176
rect 12260 14112 12276 14176
rect 12340 14112 12356 14176
rect 12420 14112 12436 14176
rect 12500 14112 12508 14176
rect 12019 13564 12085 13565
rect 12019 13500 12020 13564
rect 12084 13500 12085 13564
rect 12019 13499 12085 13500
rect 11467 11932 11533 11933
rect 11467 11868 11468 11932
rect 11532 11868 11533 11932
rect 11467 11867 11533 11868
rect 11099 9892 11165 9893
rect 11099 9828 11100 9892
rect 11164 9828 11165 9892
rect 11099 9827 11165 9828
rect 11102 5949 11162 9827
rect 11283 9348 11349 9349
rect 11283 9284 11284 9348
rect 11348 9284 11349 9348
rect 11283 9283 11349 9284
rect 11286 6629 11346 9283
rect 12022 9213 12082 13499
rect 12188 13088 12508 14112
rect 12571 13836 12637 13837
rect 12571 13772 12572 13836
rect 12636 13772 12637 13836
rect 12571 13771 12637 13772
rect 12188 13024 12196 13088
rect 12260 13024 12276 13088
rect 12340 13024 12356 13088
rect 12420 13024 12436 13088
rect 12500 13024 12508 13088
rect 12188 12000 12508 13024
rect 12188 11936 12196 12000
rect 12260 11936 12276 12000
rect 12340 11936 12356 12000
rect 12420 11936 12436 12000
rect 12500 11936 12508 12000
rect 12188 10912 12508 11936
rect 12188 10848 12196 10912
rect 12260 10848 12276 10912
rect 12340 10848 12356 10912
rect 12420 10848 12436 10912
rect 12500 10848 12508 10912
rect 12188 9824 12508 10848
rect 12188 9760 12196 9824
rect 12260 9760 12276 9824
rect 12340 9760 12356 9824
rect 12420 9760 12436 9824
rect 12500 9760 12508 9824
rect 11467 9212 11533 9213
rect 11467 9148 11468 9212
rect 11532 9148 11533 9212
rect 11467 9147 11533 9148
rect 12019 9212 12085 9213
rect 12019 9148 12020 9212
rect 12084 9148 12085 9212
rect 12019 9147 12085 9148
rect 11283 6628 11349 6629
rect 11283 6564 11284 6628
rect 11348 6564 11349 6628
rect 11283 6563 11349 6564
rect 11283 6356 11349 6357
rect 11283 6292 11284 6356
rect 11348 6292 11349 6356
rect 11283 6291 11349 6292
rect 11099 5948 11165 5949
rect 11099 5884 11100 5948
rect 11164 5884 11165 5948
rect 11099 5883 11165 5884
rect 11099 5812 11165 5813
rect 11099 5748 11100 5812
rect 11164 5748 11165 5812
rect 11099 5747 11165 5748
rect 10915 3908 10981 3909
rect 10915 3844 10916 3908
rect 10980 3844 10981 3908
rect 10915 3843 10981 3844
rect 10314 3776 10322 3840
rect 10386 3776 10402 3840
rect 10466 3776 10482 3840
rect 10546 3776 10562 3840
rect 10626 3776 10634 3840
rect 9811 3092 9877 3093
rect 9811 3028 9812 3092
rect 9876 3028 9877 3092
rect 9811 3027 9877 3028
rect 10314 2752 10634 3776
rect 11102 3093 11162 5747
rect 11286 4453 11346 6291
rect 11283 4452 11349 4453
rect 11283 4388 11284 4452
rect 11348 4388 11349 4452
rect 11283 4387 11349 4388
rect 11283 4316 11349 4317
rect 11283 4252 11284 4316
rect 11348 4252 11349 4316
rect 11283 4251 11349 4252
rect 11286 3637 11346 4251
rect 11470 4045 11530 9147
rect 12188 8736 12508 9760
rect 12188 8672 12196 8736
rect 12260 8672 12276 8736
rect 12340 8672 12356 8736
rect 12420 8672 12436 8736
rect 12500 8672 12508 8736
rect 11835 8532 11901 8533
rect 11835 8468 11836 8532
rect 11900 8468 11901 8532
rect 11835 8467 11901 8468
rect 11651 7036 11717 7037
rect 11651 6972 11652 7036
rect 11716 6972 11717 7036
rect 11651 6971 11717 6972
rect 11467 4044 11533 4045
rect 11467 3980 11468 4044
rect 11532 3980 11533 4044
rect 11467 3979 11533 3980
rect 11283 3636 11349 3637
rect 11283 3572 11284 3636
rect 11348 3572 11349 3636
rect 11283 3571 11349 3572
rect 11654 3501 11714 6971
rect 11651 3500 11717 3501
rect 11651 3436 11652 3500
rect 11716 3436 11717 3500
rect 11651 3435 11717 3436
rect 11838 3093 11898 8467
rect 12188 7648 12508 8672
rect 12574 8533 12634 13771
rect 12758 12341 12818 16491
rect 13307 16012 13373 16013
rect 13307 15948 13308 16012
rect 13372 15948 13373 16012
rect 13307 15947 13373 15948
rect 13310 12450 13370 15947
rect 13494 13565 13554 16627
rect 13491 13564 13557 13565
rect 13491 13500 13492 13564
rect 13556 13500 13557 13564
rect 13491 13499 13557 13500
rect 13678 13157 13738 16763
rect 13859 16012 13925 16013
rect 13859 15948 13860 16012
rect 13924 15948 13925 16012
rect 13859 15947 13925 15948
rect 13862 13565 13922 15947
rect 14062 15808 14382 16832
rect 14595 16284 14661 16285
rect 14595 16220 14596 16284
rect 14660 16220 14661 16284
rect 14595 16219 14661 16220
rect 14062 15744 14070 15808
rect 14134 15744 14150 15808
rect 14214 15744 14230 15808
rect 14294 15744 14310 15808
rect 14374 15744 14382 15808
rect 14062 14720 14382 15744
rect 14062 14656 14070 14720
rect 14134 14656 14150 14720
rect 14214 14656 14230 14720
rect 14294 14656 14310 14720
rect 14374 14656 14382 14720
rect 14062 13632 14382 14656
rect 14062 13568 14070 13632
rect 14134 13568 14150 13632
rect 14214 13568 14230 13632
rect 14294 13568 14310 13632
rect 14374 13568 14382 13632
rect 13859 13564 13925 13565
rect 13859 13500 13860 13564
rect 13924 13500 13925 13564
rect 13859 13499 13925 13500
rect 13491 13156 13557 13157
rect 13491 13092 13492 13156
rect 13556 13092 13557 13156
rect 13491 13091 13557 13092
rect 13675 13156 13741 13157
rect 13675 13092 13676 13156
rect 13740 13092 13741 13156
rect 13675 13091 13741 13092
rect 13126 12390 13370 12450
rect 12755 12340 12821 12341
rect 12755 12276 12756 12340
rect 12820 12276 12821 12340
rect 12755 12275 12821 12276
rect 13126 10165 13186 12390
rect 13123 10164 13189 10165
rect 13123 10100 13124 10164
rect 13188 10100 13189 10164
rect 13123 10099 13189 10100
rect 12571 8532 12637 8533
rect 12571 8468 12572 8532
rect 12636 8468 12637 8532
rect 12571 8467 12637 8468
rect 12571 7716 12637 7717
rect 12571 7652 12572 7716
rect 12636 7652 12637 7716
rect 12571 7651 12637 7652
rect 12188 7584 12196 7648
rect 12260 7584 12276 7648
rect 12340 7584 12356 7648
rect 12420 7584 12436 7648
rect 12500 7584 12508 7648
rect 12019 7036 12085 7037
rect 12019 6972 12020 7036
rect 12084 6972 12085 7036
rect 12019 6971 12085 6972
rect 12022 3093 12082 6971
rect 12188 6560 12508 7584
rect 12188 6496 12196 6560
rect 12260 6496 12276 6560
rect 12340 6496 12356 6560
rect 12420 6496 12436 6560
rect 12500 6496 12508 6560
rect 12188 5472 12508 6496
rect 12574 6221 12634 7651
rect 12939 7444 13005 7445
rect 12939 7380 12940 7444
rect 13004 7380 13005 7444
rect 12939 7379 13005 7380
rect 12571 6220 12637 6221
rect 12571 6156 12572 6220
rect 12636 6156 12637 6220
rect 12571 6155 12637 6156
rect 12188 5408 12196 5472
rect 12260 5408 12276 5472
rect 12340 5408 12356 5472
rect 12420 5408 12436 5472
rect 12500 5408 12508 5472
rect 12188 4384 12508 5408
rect 12571 5404 12637 5405
rect 12571 5340 12572 5404
rect 12636 5340 12637 5404
rect 12571 5339 12637 5340
rect 12574 4861 12634 5339
rect 12942 4861 13002 7379
rect 13126 6493 13186 10099
rect 13494 10029 13554 13091
rect 13862 10301 13922 13499
rect 14062 12544 14382 13568
rect 14062 12480 14070 12544
rect 14134 12480 14150 12544
rect 14214 12480 14230 12544
rect 14294 12480 14310 12544
rect 14374 12480 14382 12544
rect 14062 11456 14382 12480
rect 14062 11392 14070 11456
rect 14134 11392 14150 11456
rect 14214 11392 14230 11456
rect 14294 11392 14310 11456
rect 14374 11392 14382 11456
rect 14062 10368 14382 11392
rect 14062 10304 14070 10368
rect 14134 10304 14150 10368
rect 14214 10304 14230 10368
rect 14294 10304 14310 10368
rect 14374 10304 14382 10368
rect 13859 10300 13925 10301
rect 13859 10236 13860 10300
rect 13924 10236 13925 10300
rect 13859 10235 13925 10236
rect 13491 10028 13557 10029
rect 13491 9964 13492 10028
rect 13556 9964 13557 10028
rect 13491 9963 13557 9964
rect 13494 9890 13554 9963
rect 13310 9830 13554 9890
rect 13123 6492 13189 6493
rect 13123 6428 13124 6492
rect 13188 6428 13189 6492
rect 13123 6427 13189 6428
rect 13123 5676 13189 5677
rect 13123 5612 13124 5676
rect 13188 5612 13189 5676
rect 13123 5611 13189 5612
rect 12571 4860 12637 4861
rect 12571 4796 12572 4860
rect 12636 4796 12637 4860
rect 12571 4795 12637 4796
rect 12939 4860 13005 4861
rect 12939 4796 12940 4860
rect 13004 4796 13005 4860
rect 12939 4795 13005 4796
rect 12571 4452 12637 4453
rect 12571 4388 12572 4452
rect 12636 4388 12637 4452
rect 12571 4387 12637 4388
rect 12188 4320 12196 4384
rect 12260 4320 12276 4384
rect 12340 4320 12356 4384
rect 12420 4320 12436 4384
rect 12500 4320 12508 4384
rect 12188 3296 12508 4320
rect 12188 3232 12196 3296
rect 12260 3232 12276 3296
rect 12340 3232 12356 3296
rect 12420 3232 12436 3296
rect 12500 3232 12508 3296
rect 11099 3092 11165 3093
rect 11099 3028 11100 3092
rect 11164 3028 11165 3092
rect 11099 3027 11165 3028
rect 11835 3092 11901 3093
rect 11835 3028 11836 3092
rect 11900 3028 11901 3092
rect 11835 3027 11901 3028
rect 12019 3092 12085 3093
rect 12019 3028 12020 3092
rect 12084 3028 12085 3092
rect 12019 3027 12085 3028
rect 10314 2688 10322 2752
rect 10386 2688 10402 2752
rect 10466 2688 10482 2752
rect 10546 2688 10562 2752
rect 10626 2688 10634 2752
rect 10314 2128 10634 2688
rect 12188 2208 12508 3232
rect 12574 2821 12634 4387
rect 12755 3772 12821 3773
rect 12755 3708 12756 3772
rect 12820 3708 12821 3772
rect 12755 3707 12821 3708
rect 12758 3229 12818 3707
rect 12942 3365 13002 4795
rect 12939 3364 13005 3365
rect 12939 3300 12940 3364
rect 13004 3300 13005 3364
rect 12939 3299 13005 3300
rect 12755 3228 12821 3229
rect 12755 3164 12756 3228
rect 12820 3164 12821 3228
rect 12755 3163 12821 3164
rect 13126 3093 13186 5611
rect 13123 3092 13189 3093
rect 13123 3028 13124 3092
rect 13188 3028 13189 3092
rect 13123 3027 13189 3028
rect 12571 2820 12637 2821
rect 12571 2756 12572 2820
rect 12636 2756 12637 2820
rect 12571 2755 12637 2756
rect 13310 2790 13370 9830
rect 13491 9620 13557 9621
rect 13491 9556 13492 9620
rect 13556 9556 13557 9620
rect 13491 9555 13557 9556
rect 13494 2954 13554 9555
rect 13675 9484 13741 9485
rect 13675 9420 13676 9484
rect 13740 9420 13741 9484
rect 13675 9419 13741 9420
rect 13678 8805 13738 9419
rect 14062 9280 14382 10304
rect 14598 10029 14658 16219
rect 15331 15332 15397 15333
rect 15331 15268 15332 15332
rect 15396 15268 15397 15332
rect 15331 15267 15397 15268
rect 14595 10028 14661 10029
rect 14595 9964 14596 10028
rect 14660 9964 14661 10028
rect 14595 9963 14661 9964
rect 14062 9216 14070 9280
rect 14134 9216 14150 9280
rect 14214 9216 14230 9280
rect 14294 9216 14310 9280
rect 14374 9216 14382 9280
rect 13675 8804 13741 8805
rect 13675 8740 13676 8804
rect 13740 8740 13741 8804
rect 13675 8739 13741 8740
rect 13678 4453 13738 8739
rect 14062 8192 14382 9216
rect 14062 8128 14070 8192
rect 14134 8128 14150 8192
rect 14214 8128 14230 8192
rect 14294 8128 14310 8192
rect 14374 8128 14382 8192
rect 13859 7988 13925 7989
rect 13859 7924 13860 7988
rect 13924 7924 13925 7988
rect 13859 7923 13925 7924
rect 13862 6493 13922 7923
rect 14062 7104 14382 8128
rect 14062 7040 14070 7104
rect 14134 7040 14150 7104
rect 14214 7040 14230 7104
rect 14294 7040 14310 7104
rect 14374 7040 14382 7104
rect 13859 6492 13925 6493
rect 13859 6428 13860 6492
rect 13924 6428 13925 6492
rect 13859 6427 13925 6428
rect 13862 5405 13922 6427
rect 14062 6016 14382 7040
rect 14779 6084 14845 6085
rect 14779 6020 14780 6084
rect 14844 6020 14845 6084
rect 14779 6019 14845 6020
rect 14062 5952 14070 6016
rect 14134 5952 14150 6016
rect 14214 5952 14230 6016
rect 14294 5952 14310 6016
rect 14374 5952 14382 6016
rect 13859 5404 13925 5405
rect 13859 5340 13860 5404
rect 13924 5340 13925 5404
rect 13859 5339 13925 5340
rect 13859 5268 13925 5269
rect 13859 5204 13860 5268
rect 13924 5204 13925 5268
rect 13859 5203 13925 5204
rect 13675 4452 13741 4453
rect 13675 4388 13676 4452
rect 13740 4388 13741 4452
rect 13675 4387 13741 4388
rect 13494 2894 13738 2954
rect 13310 2730 13554 2790
rect 13494 2549 13554 2730
rect 13491 2548 13557 2549
rect 13491 2484 13492 2548
rect 13556 2484 13557 2548
rect 13491 2483 13557 2484
rect 13678 2277 13738 2894
rect 13862 2821 13922 5203
rect 14062 4928 14382 5952
rect 14595 5540 14661 5541
rect 14595 5476 14596 5540
rect 14660 5476 14661 5540
rect 14595 5475 14661 5476
rect 14062 4864 14070 4928
rect 14134 4864 14150 4928
rect 14214 4864 14230 4928
rect 14294 4864 14310 4928
rect 14374 4864 14382 4928
rect 14062 3840 14382 4864
rect 14062 3776 14070 3840
rect 14134 3776 14150 3840
rect 14214 3776 14230 3840
rect 14294 3776 14310 3840
rect 14374 3776 14382 3840
rect 13859 2820 13925 2821
rect 13859 2756 13860 2820
rect 13924 2756 13925 2820
rect 13859 2755 13925 2756
rect 14062 2752 14382 3776
rect 14598 3501 14658 5475
rect 14595 3500 14661 3501
rect 14595 3436 14596 3500
rect 14660 3436 14661 3500
rect 14595 3435 14661 3436
rect 14062 2688 14070 2752
rect 14134 2688 14150 2752
rect 14214 2688 14230 2752
rect 14294 2688 14310 2752
rect 14374 2688 14382 2752
rect 13675 2276 13741 2277
rect 13675 2212 13676 2276
rect 13740 2212 13741 2276
rect 13675 2211 13741 2212
rect 12188 2144 12196 2208
rect 12260 2144 12276 2208
rect 12340 2144 12356 2208
rect 12420 2144 12436 2208
rect 12500 2144 12508 2208
rect 12188 2128 12508 2144
rect 14062 2128 14382 2688
rect 14598 2413 14658 3435
rect 14782 3365 14842 6019
rect 15334 5405 15394 15267
rect 15331 5404 15397 5405
rect 15331 5340 15332 5404
rect 15396 5340 15397 5404
rect 15331 5339 15397 5340
rect 14779 3364 14845 3365
rect 14779 3300 14780 3364
rect 14844 3300 14845 3364
rect 14779 3299 14845 3300
rect 15334 3093 15394 5339
rect 15331 3092 15397 3093
rect 15331 3028 15332 3092
rect 15396 3028 15397 3092
rect 15331 3027 15397 3028
rect 14595 2412 14661 2413
rect 14595 2348 14596 2412
rect 14660 2348 14661 2412
rect 14595 2347 14661 2348
rect 3923 2004 3989 2005
rect 3923 1940 3924 2004
rect 3988 1940 3989 2004
rect 3923 1939 3989 1940
rect 9259 2004 9325 2005
rect 9259 1940 9260 2004
rect 9324 1940 9325 2004
rect 9259 1939 9325 1940
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_E_FTB01_A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14352 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_N_FTB01_A
timestamp 1649977179
transform 1 0 2760 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_W_FTB01_A
timestamp 1649977179
transform 1 0 4140 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1649977179
transform 1 0 3956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1649977179
transform -1 0 2668 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1649977179
transform -1 0 2300 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1649977179
transform -1 0 5796 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1649977179
transform -1 0 6532 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1649977179
transform -1 0 4692 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1649977179
transform -1 0 5060 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1649977179
transform -1 0 6256 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1649977179
transform 1 0 9292 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1649977179
transform 1 0 12512 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1649977179
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1649977179
transform -1 0 2208 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1649977179
transform -1 0 3036 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1649977179
transform 1 0 3956 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1649977179
transform 1 0 4508 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1649977179
transform -1 0 5888 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1649977179
transform 1 0 5704 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1649977179
transform -1 0 7176 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1649977179
transform -1 0 7176 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1649977179
transform 1 0 7820 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 1564 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform 1 0 8096 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 14260 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 10488 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 10672 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 10856 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 11960 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 14628 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 12144 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 12512 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 11408 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 11408 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 3680 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 3312 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 4876 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 4784 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 2668 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 5520 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 9936 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 5428 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform 1 0 10212 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 15732 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 14628 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 13800 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 15732 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 15548 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 14444 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 13708 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 15732 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 15732 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 13892 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 13616 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 15732 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 14444 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 13892 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 13524 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 10488 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 11408 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 13156 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 13340 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 15548 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 14260 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 2760 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 6900 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 8280 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 4600 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 2392 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 5244 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5428 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 4324 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 3036 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 4416 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 3864 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 4784 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform -1 0 6256 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 5612 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1649977179
transform 1 0 7912 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9200 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5612 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 5428 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 8924 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7176 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 4048 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 4232 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 9384 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9108 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 3864 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 4600 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 8648 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 4232 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 2668 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 4416 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 6348 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 9016 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9292 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 4324 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 4416 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 2944 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9200 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 7360 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 4048 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 6900 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 4140 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 3128 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5336 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9384 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 4232 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 3680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 10580 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9200 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6900 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 8280 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 8832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 7176 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 9108 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7084 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 7176 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 7176 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 6900 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 9568 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 9568 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 6532 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 11040 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 4968 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 4600 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 11040 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 10304 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 2668 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 6532 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 10488 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 14904 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 13708 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__S
timestamp 1649977179
transform -1 0 15732 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 11960 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 12696 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 12328 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 13616 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 13432 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__S
timestamp 1649977179
transform 1 0 11592 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_0__S
timestamp 1649977179
transform 1 0 12144 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_1__S
timestamp 1649977179
transform -1 0 9108 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 5888 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 4876 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 1564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 2944 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__S
timestamp 1649977179
transform -1 0 12696 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 10856 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__S
timestamp 1649977179
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 9200 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 12788 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 7176 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 5244 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 13708 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 15732 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 13984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 14352 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 14260 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 14352 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 14536 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 3128 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 3772 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 12420 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 13432 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 13340 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 3036 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 12420 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 12052 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 13892 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 12328 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 14352 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 13708 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 11684 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 10488 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 15180 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 9108 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 9108 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 10764 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 14260 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 13616 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 12604 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l4_in_0__S
timestamp 1649977179
transform 1 0 12328 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output50_A
timestamp 1649977179
transform 1 0 12144 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform 1 0 3312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_N_FTB01_A
timestamp 1649977179
transform 1 0 1748 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_S_FTB01_A
timestamp 1649977179
transform 1 0 11776 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater128_A
timestamp 1649977179
transform -1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_70
timestamp 1649977179
transform 1 0 7544 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_158
timestamp 1649977179
transform 1 0 15640 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_71
timestamp 1649977179
transform 1 0 7636 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_90
timestamp 1649977179
transform 1 0 9384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_19
timestamp 1649977179
transform 1 0 2852 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_87
timestamp 1649977179
transform 1 0 9108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1649977179
transform 1 0 1748 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_26
timestamp 1649977179
transform 1 0 3496 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_36
timestamp 1649977179
transform 1 0 4416 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_10
timestamp 1649977179
transform 1 0 2024 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_24
timestamp 1649977179
transform 1 0 3312 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_113
timestamp 1649977179
transform 1 0 11500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_14 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2392 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_33 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4140 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_37
timestamp 1649977179
transform 1 0 4508 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_40 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4784 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_53
timestamp 1649977179
transform 1 0 5980 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_158
timestamp 1649977179
transform 1 0 15640 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7
timestamp 1649977179
transform 1 0 1748 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_17 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2668 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_35
timestamp 1649977179
transform 1 0 4324 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_38 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4600 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_50
timestamp 1649977179
transform 1 0 5704 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_56
timestamp 1649977179
transform 1 0 6256 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_96
timestamp 1649977179
transform 1 0 9936 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_99
timestamp 1649977179
transform 1 0 10212 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_108
timestamp 1649977179
transform 1 0 11040 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_136
timestamp 1649977179
transform 1 0 13616 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_10
timestamp 1649977179
transform 1 0 2024 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_18
timestamp 1649977179
transform 1 0 2760 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_65
timestamp 1649977179
transform 1 0 7084 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_122
timestamp 1649977179
transform 1 0 12328 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_36
timestamp 1649977179
transform 1 0 4416 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_72
timestamp 1649977179
transform 1 0 7728 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1649977179
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_106
timestamp 1649977179
transform 1 0 10856 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_145
timestamp 1649977179
transform 1 0 14444 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_13
timestamp 1649977179
transform 1 0 2300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_48
timestamp 1649977179
transform 1 0 5520 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_74
timestamp 1649977179
transform 1 0 7912 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_104
timestamp 1649977179
transform 1 0 10672 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_151
timestamp 1649977179
transform 1 0 14996 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_10
timestamp 1649977179
transform 1 0 2024 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_49
timestamp 1649977179
transform 1 0 5612 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_61
timestamp 1649977179
transform 1 0 6716 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_106
timestamp 1649977179
transform 1 0 10856 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_114
timestamp 1649977179
transform 1 0 11592 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_143
timestamp 1649977179
transform 1 0 14260 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_146
timestamp 1649977179
transform 1 0 14536 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_10
timestamp 1649977179
transform 1 0 2024 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_53
timestamp 1649977179
transform 1 0 5980 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_73
timestamp 1649977179
transform 1 0 7820 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_86
timestamp 1649977179
transform 1 0 9016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_145
timestamp 1649977179
transform 1 0 14444 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_158
timestamp 1649977179
transform 1 0 15640 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_7
timestamp 1649977179
transform 1 0 1748 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_19
timestamp 1649977179
transform 1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_37
timestamp 1649977179
transform 1 0 4508 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_45
timestamp 1649977179
transform 1 0 5244 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_64
timestamp 1649977179
transform 1 0 6992 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_23
timestamp 1649977179
transform 1 0 3220 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_46
timestamp 1649977179
transform 1 0 5336 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1649977179
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_82
timestamp 1649977179
transform 1 0 8648 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1649977179
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_138
timestamp 1649977179
transform 1 0 13800 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_158
timestamp 1649977179
transform 1 0 15640 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_7
timestamp 1649977179
transform 1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_38
timestamp 1649977179
transform 1 0 4600 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_46
timestamp 1649977179
transform 1 0 5336 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_67
timestamp 1649977179
transform 1 0 7268 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_105
timestamp 1649977179
transform 1 0 10764 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_121
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_146
timestamp 1649977179
transform 1 0 14536 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_158
timestamp 1649977179
transform 1 0 15640 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_7
timestamp 1649977179
transform 1 0 1748 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_50
timestamp 1649977179
transform 1 0 5704 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_76
timestamp 1649977179
transform 1 0 8096 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_88
timestamp 1649977179
transform 1 0 9200 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1649977179
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_31
timestamp 1649977179
transform 1 0 3956 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_57
timestamp 1649977179
transform 1 0 6348 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_10
timestamp 1649977179
transform 1 0 2024 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_16
timestamp 1649977179
transform 1 0 2576 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1649977179
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_83
timestamp 1649977179
transform 1 0 8740 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_86
timestamp 1649977179
transform 1 0 9016 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_107
timestamp 1649977179
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_117
timestamp 1649977179
transform 1 0 11868 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 1649977179
transform 1 0 12236 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_153
timestamp 1649977179
transform 1 0 15180 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_9
timestamp 1649977179
transform 1 0 1932 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 1649977179
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_67
timestamp 1649977179
transform 1 0 7268 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_102
timestamp 1649977179
transform 1 0 10488 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_20
timestamp 1649977179
transform 1 0 2944 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_40
timestamp 1649977179
transform 1 0 4784 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_46
timestamp 1649977179
transform 1 0 5336 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_59
timestamp 1649977179
transform 1 0 6532 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_87
timestamp 1649977179
transform 1 0 9108 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_106
timestamp 1649977179
transform 1 0 10856 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_147
timestamp 1649977179
transform 1 0 14628 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_35
timestamp 1649977179
transform 1 0 4324 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_75
timestamp 1649977179
transform 1 0 8004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_148
timestamp 1649977179
transform 1 0 14720 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_41
timestamp 1649977179
transform 1 0 4876 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_47
timestamp 1649977179
transform 1 0 5428 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1649977179
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_139
timestamp 1649977179
transform 1 0 13892 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_46
timestamp 1649977179
transform 1 0 5336 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_63
timestamp 1649977179
transform 1 0 6900 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_158
timestamp 1649977179
transform 1 0 15640 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_46
timestamp 1649977179
transform 1 0 5336 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_102
timestamp 1649977179
transform 1 0 10488 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 16008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 16008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 16008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 16008 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 16008 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 16008 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 16008 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 16008 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 16008 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 16008 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 16008 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 16008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 16008 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 16008 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 16008 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 16008 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 16008 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 16008 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 16008 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 16008 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 16008 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 16008 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 16008 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 16008 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 16008 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 16008 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 16008 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 16008 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  Test_en_E_FTB01 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 14812 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Test_en_N_FTB01
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Test_en_W_FTB01
timestamp 1649977179
transform 1 0 2576 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _32_
timestamp 1649977179
transform 1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _33_
timestamp 1649977179
transform 1 0 3220 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _34_
timestamp 1649977179
transform 1 0 2944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1649977179
transform 1 0 2392 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _36_
timestamp 1649977179
transform 1 0 2944 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _37_
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp 1649977179
transform 1 0 2668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp 1649977179
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1649977179
transform 1 0 6256 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _43_
timestamp 1649977179
transform 1 0 14260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _44_
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _45_
timestamp 1649977179
transform 1 0 7176 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _46_
timestamp 1649977179
transform 1 0 8280 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _47_
timestamp 1649977179
transform 1 0 15456 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1649977179
transform 1 0 9752 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1649977179
transform 1 0 14352 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1649977179
transform 1 0 3312 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1649977179
transform -1 0 2392 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1649977179
transform -1 0 3312 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1649977179
transform -1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1649977179
transform -1 0 3864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1649977179
transform -1 0 3680 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1649977179
transform -1 0 4140 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1649977179
transform -1 0 4416 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 1649977179
transform 1 0 5428 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1649977179
transform 1 0 7176 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 1649977179
transform 1 0 7544 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1649977179
transform 1 0 7636 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1649977179
transform 1 0 8004 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1649977179
transform 1 0 8464 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1649977179
transform 1 0 9108 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1649977179
transform 1 0 15272 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1649977179
transform 1 0 13432 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1649977179
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_2_N_FTB01
timestamp 1649977179
transform -1 0 2484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_2_S_FTB01
timestamp 1649977179
transform -1 0 14260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_3_N_FTB01
timestamp 1649977179
transform 1 0 14996 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_3_S_FTB01
timestamp 1649977179
transform 1 0 15364 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 8832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1649977179
transform -1 0 11224 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10488 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1649977179
transform 1 0 12420 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1649977179
transform -1 0 12420 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1649977179
transform 1 0 12420 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1649977179
transform 1 0 12420 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 1649977179
transform 1 0 13340 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1649977179
transform -1 0 7728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform -1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1649977179
transform 1 0 7728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1649977179
transform 1 0 8464 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1649977179
transform -1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1649977179
transform -1 0 8832 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1649977179
transform 1 0 9384 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1649977179
transform 1 0 9568 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1649977179
transform -1 0 9568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform -1 0 10488 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1649977179
transform 1 0 13616 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform 1 0 15272 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1649977179
transform 1 0 14536 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1649977179
transform 1 0 14720 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform -1 0 15732 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input30
timestamp 1649977179
transform -1 0 13616 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1649977179
transform -1 0 12512 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1649977179
transform -1 0 11408 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1649977179
transform -1 0 15732 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform -1 0 13984 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform 1 0 12328 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform -1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input37
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1649977179
transform -1 0 13708 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1649977179
transform -1 0 13340 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1649977179
transform -1 0 13432 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input41
timestamp 1649977179
transform 1 0 14076 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1649977179
transform -1 0 13432 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1649977179
transform -1 0 14352 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1649977179
transform 1 0 15456 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1649977179
transform -1 0 14536 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2208 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2944 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 7084 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 10212 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8004 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 6348 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 5336 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 6532 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 5428 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10580 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 2208 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 3680 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 3220 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 2116 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 5336 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 5796 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10856 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5336 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 5796 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 10580 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8832 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 4048 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 2208 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 11040 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10764 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4048 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4784 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 10580 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 5888 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 2852 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 6532 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 9200 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10948 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 7820 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 5980 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 6072 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 4600 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 5428 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 7728 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10856 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 9108 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4232 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 8832 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 5796 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 2760 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 5520 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 7360 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11040 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 2668 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 3864 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 12052 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10856 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7084 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 7912 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 9016 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10764 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 8832 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 10764 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7268 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7360 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 8832 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 7084 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8004 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9384 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8004 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 7544 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 9936 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 10580 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_0.mux_l2_in_3__138 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11224 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 7452 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1649977179
transform 1 0 6808 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5152 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4508 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 3772 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_2_
timestamp 1649977179
transform -1 0 8556 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_1.mux_l2_in_3__139
timestamp 1649977179
transform 1 0 9384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_3_
timestamp 1649977179
transform -1 0 8556 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_0_
timestamp 1649977179
transform -1 0 4324 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l4_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 2668 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2668 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_2_
timestamp 1649977179
transform 1 0 6716 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_2.mux_l2_in_3__146
timestamp 1649977179
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_3_
timestamp 1649977179
transform 1 0 7636 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2668 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_1_
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l4_in_0_
timestamp 1649977179
transform -1 0 2392 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2392 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12328 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_1_
timestamp 1649977179
transform -1 0 15364 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_2_
timestamp 1649977179
transform -1 0 14904 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14904 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14260 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_2_
timestamp 1649977179
transform 1 0 13616 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_3_
timestamp 1649977179
transform 1 0 11776 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_3.mux_l2_in_3__147
timestamp 1649977179
transform 1 0 14260 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 12328 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_1_
timestamp 1649977179
transform -1 0 10580 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l4_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5152 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 4324 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 5796 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 4876 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5428 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_2_
timestamp 1649977179
transform 1 0 11408 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_4.mux_l2_in_3__148
timestamp 1649977179
transform 1 0 10764 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 10028 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 5428 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_1_
timestamp 1649977179
transform 1 0 9108 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l4_in_0_
timestamp 1649977179
transform 1 0 5428 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 4600 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10304 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10580 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_1_
timestamp 1649977179
transform -1 0 10580 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_2_
timestamp 1649977179
transform 1 0 13156 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_5.mux_l2_in_3__133
timestamp 1649977179
transform 1 0 13524 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 12696 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_0_
timestamp 1649977179
transform -1 0 11408 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_1_
timestamp 1649977179
transform 1 0 12328 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l4_in_0_
timestamp 1649977179
transform 1 0 10580 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6900 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6624 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_1_
timestamp 1649977179
transform -1 0 5612 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_2_
timestamp 1649977179
transform 1 0 12052 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_6.mux_l2_in_3__134
timestamp 1649977179
transform 1 0 13524 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_3_
timestamp 1649977179
transform 1 0 12696 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6164 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_1_
timestamp 1649977179
transform 1 0 10672 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l4_in_0_
timestamp 1649977179
transform 1 0 5060 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1748 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14628 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 14536 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_2_
timestamp 1649977179
transform -1 0 15364 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_0_
timestamp 1649977179
transform 1 0 13524 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14628 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_2_
timestamp 1649977179
transform 1 0 12880 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_7.mux_l2_in_3__135
timestamp 1649977179
transform 1 0 15088 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14720 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_0_
timestamp 1649977179
transform 1 0 12788 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_1_
timestamp 1649977179
transform 1 0 12512 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12328 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1748 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 11040 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_1_
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_2_
timestamp 1649977179
transform 1 0 11868 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_1_
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_2_
timestamp 1649977179
transform -1 0 13708 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_8.mux_l2_in_3__136
timestamp 1649977179
transform 1 0 14628 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14168 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_0_
timestamp 1649977179
transform 1 0 10948 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_1_
timestamp 1649977179
transform 1 0 13616 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l4_in_0_
timestamp 1649977179
transform -1 0 2300 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1748 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2300 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_1_
timestamp 1649977179
transform 1 0 2944 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_2_
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_9.mux_l2_in_3__137
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_3_
timestamp 1649977179
transform 1 0 13432 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 1564 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_1_
timestamp 1649977179
transform 1 0 11960 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l4_in_0_
timestamp 1649977179
transform -1 0 2208 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1748 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l1_in_0_
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_0_
timestamp 1649977179
transform -1 0 2208 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_1_
timestamp 1649977179
transform 1 0 2208 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_2_
timestamp 1649977179
transform 1 0 11592 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_10.mux_l2_in_3__140
timestamp 1649977179
transform 1 0 12328 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_3_
timestamp 1649977179
transform 1 0 11224 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_0_
timestamp 1649977179
transform -1 0 2208 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_1_
timestamp 1649977179
transform 1 0 11040 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l4_in_0_
timestamp 1649977179
transform -1 0 2208 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1748 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_0_
timestamp 1649977179
transform -1 0 15548 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_1_
timestamp 1649977179
transform -1 0 15732 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_2_
timestamp 1649977179
transform -1 0 13340 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14904 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_1_
timestamp 1649977179
transform -1 0 15364 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_2_
timestamp 1649977179
transform -1 0 13984 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_11.mux_l2_in_3__141
timestamp 1649977179
transform -1 0 15364 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12972 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1472 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_0_
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_1_
timestamp 1649977179
transform -1 0 13156 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_2_
timestamp 1649977179
transform 1 0 11868 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_0_
timestamp 1649977179
transform 1 0 13156 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_1_
timestamp 1649977179
transform -1 0 12328 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_2_
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_3_
timestamp 1649977179
transform 1 0 12328 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_12.mux_l2_in_3__142
timestamp 1649977179
transform 1 0 13156 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_1_
timestamp 1649977179
transform 1 0 10948 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l4_in_0_
timestamp 1649977179
transform 1 0 10580 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2208 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14812 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_1_
timestamp 1649977179
transform -1 0 11500 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_2_
timestamp 1649977179
transform 1 0 14168 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_13.mux_l2_in_3__143
timestamp 1649977179
transform 1 0 14996 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_3_
timestamp 1649977179
transform -1 0 10488 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_0_
timestamp 1649977179
transform 1 0 13800 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_1_
timestamp 1649977179
transform -1 0 11408 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12512 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2208 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10396 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7912 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_1_
timestamp 1649977179
transform 1 0 9384 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_2_
timestamp 1649977179
transform 1 0 12696 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_14.mux_l2_in_3__144
timestamp 1649977179
transform -1 0 12972 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_3_
timestamp 1649977179
transform 1 0 12788 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6808 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_1_
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l4_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1748 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14812 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_1_
timestamp 1649977179
transform 1 0 13984 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_2_
timestamp 1649977179
transform -1 0 13616 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_0_
timestamp 1649977179
transform 1 0 13340 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_1_
timestamp 1649977179
transform 1 0 13156 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_2_
timestamp 1649977179
transform 1 0 14628 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_15.mux_l2_in_3__145
timestamp 1649977179
transform 1 0 14444 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_3_
timestamp 1649977179
transform -1 0 12328 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_0_
timestamp 1649977179
transform 1 0 12604 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_1_
timestamp 1649977179
transform 1 0 12328 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l4_in_0_
timestamp 1649977179
transform 1 0 11776 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1748 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output47 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15364 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1649977179
transform -1 0 2208 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1649977179
transform -1 0 2116 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1649977179
transform 1 0 15364 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1649977179
transform -1 0 2116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1649977179
transform -1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1649977179
transform -1 0 5244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1649977179
transform -1 0 3680 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1649977179
transform -1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1649977179
transform -1 0 4508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1649977179
transform -1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1649977179
transform -1 0 6716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1649977179
transform -1 0 6256 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1649977179
transform -1 0 6992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1649977179
transform -1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1649977179
transform -1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1649977179
transform -1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform -1 0 2208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform -1 0 3036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform -1 0 3588 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform -1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform -1 0 3404 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform -1 0 2944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform -1 0 3772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform -1 0 2576 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform -1 0 5244 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform -1 0 6992 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform -1 0 6992 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform -1 0 7360 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform -1 0 7728 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform -1 0 8096 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform -1 0 8464 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform -1 0 8832 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform -1 0 9292 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform -1 0 9660 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform -1 0 2944 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform 1 0 2944 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform 1 0 3312 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform 1 0 3772 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform 1 0 4416 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform 1 0 4140 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform 1 0 4968 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform 1 0 4508 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform -1 0 6256 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform 1 0 2392 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform 1 0 14996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform -1 0 3128 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform 1 0 15364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform -1 0 2116 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform -1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform -1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform -1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform -1 0 1748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform -1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1649977179
transform -1 0 1748 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1649977179
transform -1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1649977179
transform -1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1649977179
transform -1 0 1748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1649977179
transform -1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1649977179
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1649977179
transform -1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1649977179
transform -1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output111
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output112
timestamp 1649977179
transform -1 0 11868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1649977179
transform -1 0 2392 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1649977179
transform 1 0 15364 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1649977179
transform -1 0 1840 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1649977179
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2024 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_N_FTB01 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1472 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_S_FTB01
timestamp 1649977179
transform 1 0 15088 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_2_N_FTB01
timestamp 1649977179
transform 1 0 14444 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_2_S_FTB01
timestamp 1649977179
transform -1 0 9752 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_3_N_FTB01
timestamp 1649977179
transform 1 0 14168 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_3_S_FTB01
timestamp 1649977179
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater117
timestamp 1649977179
transform 1 0 14812 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater118
timestamp 1649977179
transform 1 0 15272 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater119
timestamp 1649977179
transform 1 0 5244 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater120
timestamp 1649977179
transform 1 0 12788 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater121
timestamp 1649977179
transform 1 0 14812 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater122
timestamp 1649977179
transform 1 0 15456 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater123
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater124
timestamp 1649977179
transform -1 0 8096 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater125
timestamp 1649977179
transform 1 0 8004 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater126
timestamp 1649977179
transform 1 0 11224 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater127
timestamp 1649977179
transform -1 0 14812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater128
timestamp 1649977179
transform -1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater129
timestamp 1649977179
transform 1 0 7544 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater130
timestamp 1649977179
transform 1 0 6532 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater131
timestamp 1649977179
transform -1 0 14812 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater132
timestamp 1649977179
transform -1 0 6808 0 1 3264
box -38 -48 314 592
<< labels >>
flabel metal3 s 16400 16600 17200 16720 0 FreeSans 480 0 0 0 Test_en_E_in
port 0 nsew signal input
flabel metal3 s 16400 9936 17200 10056 0 FreeSans 480 0 0 0 Test_en_E_out
port 1 nsew signal tristate
flabel metal2 s 2134 19200 2190 20000 0 FreeSans 224 90 0 0 Test_en_N_out
port 2 nsew signal tristate
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 Test_en_S_in
port 3 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 Test_en_W_in
port 4 nsew signal input
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 Test_en_W_out
port 5 nsew signal tristate
flabel metal4 s 4692 2128 5012 17456 0 FreeSans 1920 90 0 0 VGND
port 6 nsew ground bidirectional
flabel metal4 s 8440 2128 8760 17456 0 FreeSans 1920 90 0 0 VGND
port 6 nsew ground bidirectional
flabel metal4 s 12188 2128 12508 17456 0 FreeSans 1920 90 0 0 VGND
port 6 nsew ground bidirectional
flabel metal4 s 2818 2128 3138 17456 0 FreeSans 1920 90 0 0 VPWR
port 7 nsew power bidirectional
flabel metal4 s 6566 2128 6886 17456 0 FreeSans 1920 90 0 0 VPWR
port 7 nsew power bidirectional
flabel metal4 s 10314 2128 10634 17456 0 FreeSans 1920 90 0 0 VPWR
port 7 nsew power bidirectional
flabel metal4 s 14062 2128 14382 17456 0 FreeSans 1920 90 0 0 VPWR
port 7 nsew power bidirectional
flabel metal3 s 0 824 800 944 0 FreeSans 480 0 0 0 ccff_head
port 8 nsew signal input
flabel metal3 s 16400 3272 17200 3392 0 FreeSans 480 0 0 0 ccff_tail
port 9 nsew signal tristate
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 10 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 11 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 12 nsew signal input
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 13 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 14 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 15 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 16 nsew signal input
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 17 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 18 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 19 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 20 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 21 nsew signal input
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 22 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 23 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 24 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 25 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 26 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 27 nsew signal input
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 28 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 29 nsew signal input
flabel metal2 s 1766 0 1822 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 30 nsew signal tristate
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 31 nsew signal tristate
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 32 nsew signal tristate
flabel metal2 s 5078 0 5134 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 33 nsew signal tristate
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 34 nsew signal tristate
flabel metal2 s 5630 0 5686 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 35 nsew signal tristate
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 36 nsew signal tristate
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 37 nsew signal tristate
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 38 nsew signal tristate
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 39 nsew signal tristate
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 40 nsew signal tristate
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 41 nsew signal tristate
flabel metal2 s 2318 0 2374 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 42 nsew signal tristate
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 43 nsew signal tristate
flabel metal2 s 2870 0 2926 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 44 nsew signal tristate
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 45 nsew signal tristate
flabel metal2 s 3422 0 3478 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 46 nsew signal tristate
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 47 nsew signal tristate
flabel metal2 s 3974 0 4030 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 48 nsew signal tristate
flabel metal2 s 4250 0 4306 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 49 nsew signal tristate
flabel metal2 s 9862 19200 9918 20000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 50 nsew signal input
flabel metal2 s 13542 19200 13598 20000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 51 nsew signal input
flabel metal2 s 13910 19200 13966 20000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 52 nsew signal input
flabel metal2 s 14278 19200 14334 20000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 53 nsew signal input
flabel metal2 s 14646 19200 14702 20000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 54 nsew signal input
flabel metal2 s 15014 19200 15070 20000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 55 nsew signal input
flabel metal2 s 15382 19200 15438 20000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 56 nsew signal input
flabel metal2 s 15750 19200 15806 20000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 57 nsew signal input
flabel metal2 s 16118 19200 16174 20000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 58 nsew signal input
flabel metal2 s 16486 19200 16542 20000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 59 nsew signal input
flabel metal2 s 16854 19200 16910 20000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 60 nsew signal input
flabel metal2 s 10230 19200 10286 20000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 61 nsew signal input
flabel metal2 s 10598 19200 10654 20000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 62 nsew signal input
flabel metal2 s 10966 19200 11022 20000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 63 nsew signal input
flabel metal2 s 11334 19200 11390 20000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 64 nsew signal input
flabel metal2 s 11702 19200 11758 20000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 65 nsew signal input
flabel metal2 s 12070 19200 12126 20000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 66 nsew signal input
flabel metal2 s 12438 19200 12494 20000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 67 nsew signal input
flabel metal2 s 12806 19200 12862 20000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 68 nsew signal input
flabel metal2 s 13174 19200 13230 20000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 69 nsew signal input
flabel metal2 s 2502 19200 2558 20000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 70 nsew signal tristate
flabel metal2 s 6182 19200 6238 20000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 71 nsew signal tristate
flabel metal2 s 6550 19200 6606 20000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 72 nsew signal tristate
flabel metal2 s 6918 19200 6974 20000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 73 nsew signal tristate
flabel metal2 s 7286 19200 7342 20000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 74 nsew signal tristate
flabel metal2 s 7654 19200 7710 20000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 75 nsew signal tristate
flabel metal2 s 8022 19200 8078 20000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 76 nsew signal tristate
flabel metal2 s 8390 19200 8446 20000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 77 nsew signal tristate
flabel metal2 s 8758 19200 8814 20000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 78 nsew signal tristate
flabel metal2 s 9126 19200 9182 20000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 79 nsew signal tristate
flabel metal2 s 9494 19200 9550 20000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 80 nsew signal tristate
flabel metal2 s 2870 19200 2926 20000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 81 nsew signal tristate
flabel metal2 s 3238 19200 3294 20000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 82 nsew signal tristate
flabel metal2 s 3606 19200 3662 20000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 83 nsew signal tristate
flabel metal2 s 3974 19200 4030 20000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 84 nsew signal tristate
flabel metal2 s 4342 19200 4398 20000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 85 nsew signal tristate
flabel metal2 s 4710 19200 4766 20000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 86 nsew signal tristate
flabel metal2 s 5078 19200 5134 20000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 87 nsew signal tristate
flabel metal2 s 5446 19200 5502 20000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 88 nsew signal tristate
flabel metal2 s 5814 19200 5870 20000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 89 nsew signal tristate
flabel metal2 s 294 19200 350 20000 0 FreeSans 224 90 0 0 clk_2_N_out
port 90 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 clk_2_S_in
port 91 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 clk_2_S_out
port 92 nsew signal tristate
flabel metal2 s 662 19200 718 20000 0 FreeSans 224 90 0 0 clk_3_N_out
port 93 nsew signal tristate
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 clk_3_S_in
port 94 nsew signal input
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 clk_3_S_out
port 95 nsew signal tristate
flabel metal3 s 0 1776 800 1896 0 FreeSans 480 0 0 0 left_grid_pin_16_
port 96 nsew signal tristate
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 left_grid_pin_17_
port 97 nsew signal tristate
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 left_grid_pin_18_
port 98 nsew signal tristate
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 left_grid_pin_19_
port 99 nsew signal tristate
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 left_grid_pin_20_
port 100 nsew signal tristate
flabel metal3 s 0 6536 800 6656 0 FreeSans 480 0 0 0 left_grid_pin_21_
port 101 nsew signal tristate
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 left_grid_pin_22_
port 102 nsew signal tristate
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 left_grid_pin_23_
port 103 nsew signal tristate
flabel metal3 s 0 9392 800 9512 0 FreeSans 480 0 0 0 left_grid_pin_24_
port 104 nsew signal tristate
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 left_grid_pin_25_
port 105 nsew signal tristate
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 left_grid_pin_26_
port 106 nsew signal tristate
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 left_grid_pin_27_
port 107 nsew signal tristate
flabel metal3 s 0 13200 800 13320 0 FreeSans 480 0 0 0 left_grid_pin_28_
port 108 nsew signal tristate
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 left_grid_pin_29_
port 109 nsew signal tristate
flabel metal3 s 0 15104 800 15224 0 FreeSans 480 0 0 0 left_grid_pin_30_
port 110 nsew signal tristate
flabel metal3 s 0 16056 800 16176 0 FreeSans 480 0 0 0 left_grid_pin_31_
port 111 nsew signal tristate
flabel metal2 s 1030 19200 1086 20000 0 FreeSans 224 90 0 0 prog_clk_0_N_out
port 112 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 prog_clk_0_S_out
port 113 nsew signal tristate
flabel metal3 s 0 18912 800 19032 0 FreeSans 480 0 0 0 prog_clk_0_W_in
port 114 nsew signal input
flabel metal2 s 1398 19200 1454 20000 0 FreeSans 224 90 0 0 prog_clk_2_N_out
port 115 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 prog_clk_2_S_in
port 116 nsew signal input
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 prog_clk_2_S_out
port 117 nsew signal tristate
flabel metal2 s 1766 19200 1822 20000 0 FreeSans 224 90 0 0 prog_clk_3_N_out
port 118 nsew signal tristate
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 prog_clk_3_S_in
port 119 nsew signal input
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 prog_clk_3_S_out
port 120 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 17200 20000
<< end >>
