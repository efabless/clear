magic
tech sky130A
magscale 1 2
timestamp 1656241705
<< viali >>
rect 3433 14569 3467 14603
rect 5733 14569 5767 14603
rect 6653 14569 6687 14603
rect 7021 14569 7055 14603
rect 7389 14569 7423 14603
rect 8677 14569 8711 14603
rect 9321 14569 9355 14603
rect 9965 14569 9999 14603
rect 10609 14569 10643 14603
rect 11805 14569 11839 14603
rect 12541 14569 12575 14603
rect 13185 14569 13219 14603
rect 10241 14501 10275 14535
rect 14289 14501 14323 14535
rect 3157 14433 3191 14467
rect 4629 14433 4663 14467
rect 6009 14433 6043 14467
rect 15117 14433 15151 14467
rect 16773 14433 16807 14467
rect 1961 14365 1995 14399
rect 2237 14365 2271 14399
rect 2881 14365 2915 14399
rect 3617 14365 3651 14399
rect 4353 14365 4387 14399
rect 4721 14365 4755 14399
rect 4997 14365 5031 14399
rect 5917 14365 5951 14399
rect 6561 14365 6595 14399
rect 6837 14365 6871 14399
rect 7481 14365 7515 14399
rect 9137 14365 9171 14399
rect 9597 14365 9631 14399
rect 10057 14365 10091 14399
rect 10885 14365 10919 14399
rect 11713 14365 11747 14399
rect 11989 14365 12023 14399
rect 12265 14365 12299 14399
rect 12817 14365 12851 14399
rect 13277 14365 13311 14399
rect 14105 14365 14139 14399
rect 14381 14365 14415 14399
rect 15301 14365 15335 14399
rect 15577 14365 15611 14399
rect 16221 14365 16255 14399
rect 16497 14365 16531 14399
rect 17049 14365 17083 14399
rect 17693 14365 17727 14399
rect 17969 14365 18003 14399
rect 6377 14229 6411 14263
rect 7665 14229 7699 14263
rect 8953 14229 8987 14263
rect 9413 14229 9447 14263
rect 10701 14229 10735 14263
rect 11529 14229 11563 14263
rect 12173 14229 12207 14263
rect 12633 14229 12667 14263
rect 13461 14229 13495 14263
rect 15393 14229 15427 14263
rect 4353 14025 4387 14059
rect 4721 14025 4755 14059
rect 4997 14025 5031 14059
rect 8125 14025 8159 14059
rect 8677 14025 8711 14059
rect 11069 14025 11103 14059
rect 12541 14025 12575 14059
rect 13277 14025 13311 14059
rect 14013 14025 14047 14059
rect 14933 14025 14967 14059
rect 10241 13957 10275 13991
rect 11621 13957 11655 13991
rect 1961 13889 1995 13923
rect 2237 13889 2271 13923
rect 2881 13889 2915 13923
rect 4077 13889 4111 13923
rect 4537 13889 4571 13923
rect 5181 13889 5215 13923
rect 5549 13889 5583 13923
rect 5825 13889 5859 13923
rect 6009 13889 6043 13923
rect 6377 13889 6411 13923
rect 6837 13889 6871 13923
rect 7021 13889 7055 13923
rect 7481 13889 7515 13923
rect 8033 13889 8067 13923
rect 8309 13889 8343 13923
rect 10057 13889 10091 13923
rect 11253 13889 11287 13923
rect 12725 13889 12759 13923
rect 13461 13889 13495 13923
rect 13837 13889 13871 13923
rect 15117 13889 15151 13923
rect 15945 13889 15979 13923
rect 16221 13889 16255 13923
rect 16497 13889 16531 13923
rect 17969 13889 18003 13923
rect 3157 13821 3191 13855
rect 3801 13821 3835 13855
rect 8493 13821 8527 13855
rect 16773 13821 16807 13855
rect 17049 13821 17083 13855
rect 17693 13821 17727 13855
rect 5365 13753 5399 13787
rect 6193 13753 6227 13787
rect 6561 13753 6595 13787
rect 7849 13753 7883 13787
rect 16037 13753 16071 13787
rect 5641 13685 5675 13719
rect 6653 13685 6687 13719
rect 7297 13685 7331 13719
rect 7665 13685 7699 13719
rect 9873 13685 9907 13719
rect 13645 13685 13679 13719
rect 16313 13685 16347 13719
rect 3341 13481 3375 13515
rect 4905 13481 4939 13515
rect 16681 13481 16715 13515
rect 3893 13413 3927 13447
rect 16313 13413 16347 13447
rect 1961 13345 1995 13379
rect 5733 13345 5767 13379
rect 6469 13345 6503 13379
rect 6561 13345 6595 13379
rect 7481 13345 7515 13379
rect 9781 13345 9815 13379
rect 11621 13345 11655 13379
rect 12449 13345 12483 13379
rect 16865 13345 16899 13379
rect 2237 13277 2271 13311
rect 2881 13277 2915 13311
rect 3157 13277 3191 13311
rect 3525 13277 3559 13311
rect 4077 13277 4111 13311
rect 4445 13277 4479 13311
rect 4813 13277 4847 13311
rect 7297 13277 7331 13311
rect 12173 13277 12207 13311
rect 16497 13277 16531 13311
rect 17693 13277 17727 13311
rect 17969 13277 18003 13311
rect 5549 13209 5583 13243
rect 9597 13209 9631 13243
rect 10057 13209 10091 13243
rect 17141 13209 17175 13243
rect 17509 13209 17543 13243
rect 4261 13141 4295 13175
rect 4629 13141 4663 13175
rect 5181 13141 5215 13175
rect 5641 13141 5675 13175
rect 6009 13141 6043 13175
rect 6377 13141 6411 13175
rect 6837 13141 6871 13175
rect 7205 13141 7239 13175
rect 9229 13141 9263 13175
rect 9689 13141 9723 13175
rect 10977 13141 11011 13175
rect 11345 13141 11379 13175
rect 11437 13141 11471 13175
rect 11805 13141 11839 13175
rect 12265 13141 12299 13175
rect 12633 13141 12667 13175
rect 13829 13141 13863 13175
rect 17049 13141 17083 13175
rect 17417 13141 17451 13175
rect 3893 12937 3927 12971
rect 4721 12937 4755 12971
rect 5181 12937 5215 12971
rect 6653 12937 6687 12971
rect 9229 12937 9263 12971
rect 9597 12937 9631 12971
rect 11621 12937 11655 12971
rect 11989 12937 12023 12971
rect 13553 12937 13587 12971
rect 13921 12937 13955 12971
rect 16865 12937 16899 12971
rect 5641 12869 5675 12903
rect 9965 12869 9999 12903
rect 10425 12869 10459 12903
rect 16957 12869 16991 12903
rect 17325 12869 17359 12903
rect 17601 12869 17635 12903
rect 3157 12801 3191 12835
rect 3433 12801 3467 12835
rect 4537 12801 4571 12835
rect 9137 12801 9171 12835
rect 10057 12801 10091 12835
rect 12081 12801 12115 12835
rect 13461 12801 13495 12835
rect 14289 12801 14323 12835
rect 14381 12801 14415 12835
rect 1961 12733 1995 12767
rect 2237 12733 2271 12767
rect 2881 12733 2915 12767
rect 3985 12733 4019 12767
rect 4077 12733 4111 12767
rect 5273 12733 5307 12767
rect 5365 12733 5399 12767
rect 9321 12733 9355 12767
rect 10241 12733 10275 12767
rect 12265 12733 12299 12767
rect 13645 12733 13679 12767
rect 14473 12733 14507 12767
rect 17233 12733 17267 12767
rect 17693 12733 17727 12767
rect 17969 12733 18003 12767
rect 6837 12665 6871 12699
rect 8677 12665 8711 12699
rect 12725 12665 12759 12699
rect 3249 12597 3283 12631
rect 3525 12597 3559 12631
rect 4353 12597 4387 12631
rect 4813 12597 4847 12631
rect 5825 12597 5859 12631
rect 8769 12597 8803 12631
rect 13093 12597 13127 12631
rect 14841 12597 14875 12631
rect 4077 12393 4111 12427
rect 9689 12393 9723 12427
rect 12817 12393 12851 12427
rect 14105 12393 14139 12427
rect 10885 12325 10919 12359
rect 13829 12325 13863 12359
rect 16589 12325 16623 12359
rect 17601 12325 17635 12359
rect 1961 12257 1995 12291
rect 3065 12257 3099 12291
rect 4997 12257 5031 12291
rect 6653 12257 6687 12291
rect 7481 12257 7515 12291
rect 8309 12257 8343 12291
rect 10241 12257 10275 12291
rect 11437 12257 11471 12291
rect 12449 12257 12483 12291
rect 12633 12257 12667 12291
rect 13369 12257 13403 12291
rect 14565 12257 14599 12291
rect 14657 12257 14691 12291
rect 16957 12257 16991 12291
rect 2237 12189 2271 12223
rect 5273 12189 5307 12223
rect 7297 12189 7331 12223
rect 11253 12189 11287 12223
rect 17417 12189 17451 12223
rect 17693 12189 17727 12223
rect 17969 12189 18003 12223
rect 2421 12121 2455 12155
rect 2697 12121 2731 12155
rect 3157 12121 3191 12155
rect 3249 12121 3283 12155
rect 3801 12121 3835 12155
rect 4261 12121 4295 12155
rect 4813 12121 4847 12155
rect 6469 12121 6503 12155
rect 8217 12121 8251 12155
rect 9505 12121 9539 12155
rect 10149 12121 10183 12155
rect 12357 12121 12391 12155
rect 15025 12121 15059 12155
rect 17141 12121 17175 12155
rect 2513 12053 2547 12087
rect 3617 12053 3651 12087
rect 4445 12053 4479 12087
rect 4905 12053 4939 12087
rect 6101 12053 6135 12087
rect 6561 12053 6595 12087
rect 6929 12053 6963 12087
rect 7389 12053 7423 12087
rect 7757 12053 7791 12087
rect 8125 12053 8159 12087
rect 8585 12053 8619 12087
rect 10057 12053 10091 12087
rect 10517 12053 10551 12087
rect 11345 12053 11379 12087
rect 11989 12053 12023 12087
rect 13185 12053 13219 12087
rect 13277 12053 13311 12087
rect 14473 12053 14507 12087
rect 15301 12053 15335 12087
rect 16405 12053 16439 12087
rect 17325 12053 17359 12087
rect 3341 11849 3375 11883
rect 3433 11849 3467 11883
rect 4353 11849 4387 11883
rect 5457 11849 5491 11883
rect 5917 11849 5951 11883
rect 8309 11849 8343 11883
rect 9137 11849 9171 11883
rect 9965 11849 9999 11883
rect 10425 11849 10459 11883
rect 13093 11849 13127 11883
rect 15025 11849 15059 11883
rect 16405 11849 16439 11883
rect 4445 11781 4479 11815
rect 6469 11781 6503 11815
rect 7113 11781 7147 11815
rect 12633 11781 12667 11815
rect 15945 11781 15979 11815
rect 17233 11781 17267 11815
rect 1961 11713 1995 11747
rect 2513 11713 2547 11747
rect 2789 11713 2823 11747
rect 5825 11713 5859 11747
rect 7021 11713 7055 11747
rect 9229 11713 9263 11747
rect 12725 11713 12759 11747
rect 13277 11713 13311 11747
rect 15117 11713 15151 11747
rect 17141 11713 17175 11747
rect 2237 11645 2271 11679
rect 3617 11645 3651 11679
rect 4537 11645 4571 11679
rect 6101 11645 6135 11679
rect 7205 11645 7239 11679
rect 7757 11645 7791 11679
rect 8125 11645 8159 11679
rect 8217 11645 8251 11679
rect 9413 11645 9447 11679
rect 10057 11645 10091 11679
rect 10241 11645 10275 11679
rect 12541 11645 12575 11679
rect 14933 11645 14967 11679
rect 16037 11645 16071 11679
rect 16129 11645 16163 11679
rect 17417 11645 17451 11679
rect 17693 11645 17727 11679
rect 17969 11645 18003 11679
rect 3801 11577 3835 11611
rect 6653 11577 6687 11611
rect 8769 11577 8803 11611
rect 2329 11509 2363 11543
rect 2605 11509 2639 11543
rect 2973 11509 3007 11543
rect 3985 11509 4019 11543
rect 7573 11509 7607 11543
rect 8677 11509 8711 11543
rect 9597 11509 9631 11543
rect 14565 11509 14599 11543
rect 15485 11509 15519 11543
rect 15577 11509 15611 11543
rect 16773 11509 16807 11543
rect 4537 11305 4571 11339
rect 7757 11305 7791 11339
rect 8953 11305 8987 11339
rect 14105 11305 14139 11339
rect 16037 11305 16071 11339
rect 2329 11237 2363 11271
rect 3341 11237 3375 11271
rect 16129 11237 16163 11271
rect 1961 11169 1995 11203
rect 2789 11169 2823 11203
rect 2881 11169 2915 11203
rect 8217 11169 8251 11203
rect 8309 11169 8343 11203
rect 9505 11169 9539 11203
rect 9781 11169 9815 11203
rect 14565 11169 14599 11203
rect 14749 11169 14783 11203
rect 15393 11169 15427 11203
rect 15485 11169 15519 11203
rect 16681 11169 16715 11203
rect 2237 11101 2271 11135
rect 2513 11101 2547 11135
rect 2973 11101 3007 11135
rect 3525 11101 3559 11135
rect 5650 11101 5684 11135
rect 5917 11101 5951 11135
rect 8585 11101 8619 11135
rect 9321 11101 9355 11135
rect 9413 11101 9447 11135
rect 11713 11101 11747 11135
rect 15301 11101 15335 11135
rect 16497 11101 16531 11135
rect 17049 11101 17083 11135
rect 17141 11101 17175 11135
rect 17417 11101 17451 11135
rect 17693 11101 17727 11135
rect 17969 11101 18003 11135
rect 3801 11033 3835 11067
rect 7665 11033 7699 11067
rect 11958 11033 11992 11067
rect 14473 11033 14507 11067
rect 16589 11033 16623 11067
rect 8125 10965 8159 10999
rect 13093 10965 13127 10999
rect 14933 10965 14967 10999
rect 17325 10965 17359 10999
rect 17601 10965 17635 10999
rect 2881 10761 2915 10795
rect 4353 10761 4387 10795
rect 8217 10761 8251 10795
rect 11529 10761 11563 10795
rect 14381 10761 14415 10795
rect 14657 10761 14691 10795
rect 15117 10761 15151 10795
rect 16681 10761 16715 10795
rect 17049 10761 17083 10795
rect 17509 10761 17543 10795
rect 5926 10693 5960 10727
rect 9422 10693 9456 10727
rect 13268 10693 13302 10727
rect 2789 10625 2823 10659
rect 3617 10625 3651 10659
rect 6193 10625 6227 10659
rect 6837 10625 6871 10659
rect 7093 10625 7127 10659
rect 10140 10625 10174 10659
rect 12642 10625 12676 10659
rect 14473 10625 14507 10659
rect 15025 10625 15059 10659
rect 1961 10557 1995 10591
rect 2237 10557 2271 10591
rect 2973 10557 3007 10591
rect 3709 10557 3743 10591
rect 3801 10557 3835 10591
rect 9689 10557 9723 10591
rect 9873 10557 9907 10591
rect 12909 10557 12943 10591
rect 13001 10557 13035 10591
rect 15209 10557 15243 10591
rect 17141 10557 17175 10591
rect 17233 10557 17267 10591
rect 17693 10557 17727 10591
rect 17969 10557 18003 10591
rect 8309 10489 8343 10523
rect 16497 10489 16531 10523
rect 2421 10421 2455 10455
rect 3249 10421 3283 10455
rect 4169 10421 4203 10455
rect 4813 10421 4847 10455
rect 11253 10421 11287 10455
rect 1593 10217 1627 10251
rect 3801 10217 3835 10251
rect 11437 10217 11471 10251
rect 16589 10217 16623 10251
rect 17417 10217 17451 10251
rect 18337 10217 18371 10251
rect 6561 10149 6595 10183
rect 9045 10149 9079 10183
rect 2513 10081 2547 10115
rect 2605 10081 2639 10115
rect 3157 10081 3191 10115
rect 16405 10081 16439 10115
rect 17049 10081 17083 10115
rect 17233 10081 17267 10115
rect 1501 10013 1535 10047
rect 1961 10013 1995 10047
rect 3249 10013 3283 10047
rect 3525 10013 3559 10047
rect 4537 10013 4571 10047
rect 7941 10013 7975 10047
rect 10158 10013 10192 10047
rect 10425 10013 10459 10047
rect 12817 10013 12851 10047
rect 16957 10013 16991 10047
rect 17785 10013 17819 10047
rect 17877 10013 17911 10047
rect 3985 9945 4019 9979
rect 4804 9945 4838 9979
rect 7674 9945 7708 9979
rect 12572 9945 12606 9979
rect 18429 9945 18463 9979
rect 1777 9877 1811 9911
rect 2053 9877 2087 9911
rect 2421 9877 2455 9911
rect 3433 9877 3467 9911
rect 5917 9877 5951 9911
rect 17601 9877 17635 9911
rect 18061 9877 18095 9911
rect 2053 9673 2087 9707
rect 3433 9673 3467 9707
rect 17417 9673 17451 9707
rect 3525 9605 3559 9639
rect 5580 9605 5614 9639
rect 13032 9605 13066 9639
rect 17141 9605 17175 9639
rect 18245 9605 18279 9639
rect 1501 9537 1535 9571
rect 1961 9537 1995 9571
rect 2605 9537 2639 9571
rect 7297 9537 7331 9571
rect 8401 9537 8435 9571
rect 8841 9537 8875 9571
rect 17601 9537 17635 9571
rect 17877 9537 17911 9571
rect 18429 9537 18463 9571
rect 2697 9469 2731 9503
rect 2881 9469 2915 9503
rect 3065 9469 3099 9503
rect 5825 9469 5859 9503
rect 7665 9469 7699 9503
rect 8585 9469 8619 9503
rect 13277 9469 13311 9503
rect 16957 9469 16991 9503
rect 1685 9401 1719 9435
rect 4445 9401 4479 9435
rect 17233 9401 17267 9435
rect 1777 9333 1811 9367
rect 2237 9333 2271 9367
rect 9965 9333 9999 9367
rect 11897 9333 11931 9367
rect 17785 9333 17819 9367
rect 18061 9333 18095 9367
rect 2513 9129 2547 9163
rect 3433 9129 3467 9163
rect 6837 9129 6871 9163
rect 8769 9129 8803 9163
rect 10149 9129 10183 9163
rect 11989 9129 12023 9163
rect 15301 9129 15335 9163
rect 17325 9129 17359 9163
rect 18337 9129 18371 9163
rect 17693 9061 17727 9095
rect 3157 8993 3191 9027
rect 14565 8993 14599 9027
rect 16037 8993 16071 9027
rect 17049 8993 17083 9027
rect 1685 8925 1719 8959
rect 2053 8925 2087 8959
rect 2145 8925 2179 8959
rect 2881 8925 2915 8959
rect 5365 8925 5399 8959
rect 5457 8925 5491 8959
rect 7389 8925 7423 8959
rect 11262 8925 11296 8959
rect 11529 8925 11563 8959
rect 13369 8925 13403 8959
rect 14749 8925 14783 8959
rect 15853 8925 15887 8959
rect 17509 8925 17543 8959
rect 17877 8925 17911 8959
rect 18245 8925 18279 8959
rect 18521 8925 18555 8959
rect 3525 8857 3559 8891
rect 5098 8857 5132 8891
rect 5724 8857 5758 8891
rect 7634 8857 7668 8891
rect 13124 8857 13158 8891
rect 15945 8857 15979 8891
rect 17233 8857 17267 8891
rect 1501 8789 1535 8823
rect 1869 8789 1903 8823
rect 2329 8789 2363 8823
rect 2973 8789 3007 8823
rect 3985 8789 4019 8823
rect 14289 8789 14323 8823
rect 14657 8789 14691 8823
rect 15117 8789 15151 8823
rect 15485 8789 15519 8823
rect 18061 8789 18095 8823
rect 2329 8585 2363 8619
rect 12909 8585 12943 8619
rect 14381 8585 14415 8619
rect 15761 8585 15795 8619
rect 17601 8585 17635 8619
rect 1869 8517 1903 8551
rect 2789 8517 2823 8551
rect 4988 8517 5022 8551
rect 9312 8517 9346 8551
rect 11774 8517 11808 8551
rect 13268 8517 13302 8551
rect 2697 8449 2731 8483
rect 3525 8449 3559 8483
rect 7490 8449 7524 8483
rect 7757 8449 7791 8483
rect 9045 8449 9079 8483
rect 13001 8449 13035 8483
rect 15853 8449 15887 8483
rect 17417 8449 17451 8483
rect 17785 8449 17819 8483
rect 17877 8449 17911 8483
rect 18245 8449 18279 8483
rect 1961 8381 1995 8415
rect 2145 8381 2179 8415
rect 2881 8381 2915 8415
rect 3617 8381 3651 8415
rect 3801 8381 3835 8415
rect 4721 8381 4755 8415
rect 11069 8381 11103 8415
rect 11529 8381 11563 8415
rect 16037 8381 16071 8415
rect 1501 8313 1535 8347
rect 6377 8313 6411 8347
rect 10425 8313 10459 8347
rect 18061 8313 18095 8347
rect 18429 8313 18463 8347
rect 3157 8245 3191 8279
rect 4077 8245 4111 8279
rect 6101 8245 6135 8279
rect 10517 8245 10551 8279
rect 15393 8245 15427 8279
rect 1501 8041 1535 8075
rect 2145 8041 2179 8075
rect 3249 8041 3283 8075
rect 11897 8041 11931 8075
rect 16957 8041 16991 8075
rect 17233 7973 17267 8007
rect 2789 7905 2823 7939
rect 3065 7905 3099 7939
rect 8953 7905 8987 7939
rect 12081 7905 12115 7939
rect 15025 7905 15059 7939
rect 15117 7905 15151 7939
rect 1685 7837 1719 7871
rect 2053 7837 2087 7871
rect 2605 7837 2639 7871
rect 4537 7837 4571 7871
rect 6193 7837 6227 7871
rect 6929 7837 6963 7871
rect 10517 7837 10551 7871
rect 10784 7837 10818 7871
rect 15209 7837 15243 7871
rect 17049 7837 17083 7871
rect 17509 7837 17543 7871
rect 18245 7837 18279 7871
rect 4782 7769 4816 7803
rect 6837 7769 6871 7803
rect 7174 7769 7208 7803
rect 9220 7769 9254 7803
rect 12348 7769 12382 7803
rect 1869 7701 1903 7735
rect 2513 7701 2547 7735
rect 5917 7701 5951 7735
rect 8309 7701 8343 7735
rect 10333 7701 10367 7735
rect 13461 7701 13495 7735
rect 15577 7701 15611 7735
rect 17601 7701 17635 7735
rect 18429 7701 18463 7735
rect 1777 7497 1811 7531
rect 2145 7497 2179 7531
rect 2513 7497 2547 7531
rect 2973 7497 3007 7531
rect 9137 7497 9171 7531
rect 14105 7497 14139 7531
rect 14565 7497 14599 7531
rect 14933 7497 14967 7531
rect 15393 7497 15427 7531
rect 16405 7497 16439 7531
rect 17049 7497 17083 7531
rect 18061 7497 18095 7531
rect 7880 7429 7914 7463
rect 10364 7429 10398 7463
rect 2605 7361 2639 7395
rect 4189 7361 4223 7395
rect 5661 7361 5695 7395
rect 5917 7361 5951 7395
rect 8125 7361 8159 7395
rect 10609 7361 10643 7395
rect 12348 7361 12382 7395
rect 14473 7361 14507 7395
rect 15301 7361 15335 7395
rect 17141 7361 17175 7395
rect 17601 7361 17635 7395
rect 17877 7361 17911 7395
rect 18245 7361 18279 7395
rect 1501 7293 1535 7327
rect 1685 7293 1719 7327
rect 2421 7293 2455 7327
rect 4445 7293 4479 7327
rect 8493 7293 8527 7327
rect 11253 7293 11287 7327
rect 12081 7293 12115 7327
rect 14657 7293 14691 7327
rect 15577 7293 15611 7327
rect 17233 7293 17267 7327
rect 3065 7225 3099 7259
rect 9229 7225 9263 7259
rect 16681 7225 16715 7259
rect 4537 7157 4571 7191
rect 6745 7157 6779 7191
rect 10701 7157 10735 7191
rect 13461 7157 13495 7191
rect 17785 7157 17819 7191
rect 18429 7157 18463 7191
rect 1501 6953 1535 6987
rect 1961 6953 1995 6987
rect 3525 6953 3559 6987
rect 5825 6953 5859 6987
rect 15393 6953 15427 6987
rect 17693 6953 17727 6987
rect 4169 6885 4203 6919
rect 2605 6817 2639 6851
rect 2973 6817 3007 6851
rect 4445 6817 4479 6851
rect 6009 6817 6043 6851
rect 12357 6817 12391 6851
rect 14841 6817 14875 6851
rect 14933 6817 14967 6851
rect 16221 6817 16255 6851
rect 16313 6817 16347 6851
rect 17141 6817 17175 6851
rect 1685 6749 1719 6783
rect 3801 6749 3835 6783
rect 4353 6749 4387 6783
rect 8493 6749 8527 6783
rect 9321 6749 9355 6783
rect 13829 6749 13863 6783
rect 17049 6749 17083 6783
rect 17877 6749 17911 6783
rect 18245 6749 18279 6783
rect 2421 6681 2455 6715
rect 4690 6681 4724 6715
rect 8237 6681 8271 6715
rect 9588 6681 9622 6715
rect 12090 6681 12124 6715
rect 13562 6681 13596 6715
rect 16129 6681 16163 6715
rect 16957 6681 16991 6715
rect 17417 6681 17451 6715
rect 1869 6613 1903 6647
rect 2329 6613 2363 6647
rect 3065 6613 3099 6647
rect 3157 6613 3191 6647
rect 3985 6613 4019 6647
rect 7113 6613 7147 6647
rect 10701 6613 10735 6647
rect 10977 6613 11011 6647
rect 12449 6613 12483 6647
rect 14473 6613 14507 6647
rect 15025 6613 15059 6647
rect 15761 6613 15795 6647
rect 16589 6613 16623 6647
rect 18061 6613 18095 6647
rect 18429 6613 18463 6647
rect 1685 6409 1719 6443
rect 2237 6409 2271 6443
rect 11345 6409 11379 6443
rect 13277 6409 13311 6443
rect 14013 6409 14047 6443
rect 14381 6409 14415 6443
rect 14841 6409 14875 6443
rect 15209 6409 15243 6443
rect 17601 6409 17635 6443
rect 2605 6341 2639 6375
rect 5926 6341 5960 6375
rect 9996 6341 10030 6375
rect 12164 6341 12198 6375
rect 13921 6341 13955 6375
rect 17785 6341 17819 6375
rect 1777 6273 1811 6307
rect 3433 6273 3467 6307
rect 3893 6273 3927 6307
rect 4169 6273 4203 6307
rect 6193 6273 6227 6307
rect 6561 6273 6595 6307
rect 6828 6273 6862 6307
rect 8125 6273 8159 6307
rect 10241 6273 10275 6307
rect 11897 6273 11931 6307
rect 14749 6273 14783 6307
rect 15577 6273 15611 6307
rect 18245 6273 18279 6307
rect 1593 6205 1627 6239
rect 2697 6205 2731 6239
rect 2881 6205 2915 6239
rect 3525 6205 3559 6239
rect 3709 6205 3743 6239
rect 8769 6205 8803 6239
rect 10793 6205 10827 6239
rect 14105 6205 14139 6239
rect 14933 6205 14967 6239
rect 15669 6205 15703 6239
rect 15761 6205 15795 6239
rect 16681 6205 16715 6239
rect 16957 6205 16991 6239
rect 2145 6069 2179 6103
rect 3065 6069 3099 6103
rect 4813 6069 4847 6103
rect 7941 6069 7975 6103
rect 8861 6069 8895 6103
rect 13553 6069 13587 6103
rect 17969 6069 18003 6103
rect 18429 6069 18463 6103
rect 2881 5865 2915 5899
rect 5917 5865 5951 5899
rect 6193 5865 6227 5899
rect 7297 5865 7331 5899
rect 9229 5865 9263 5899
rect 10517 5865 10551 5899
rect 10885 5865 10919 5899
rect 11989 5865 12023 5899
rect 14197 5865 14231 5899
rect 15117 5865 15151 5899
rect 15485 5865 15519 5899
rect 17233 5865 17267 5899
rect 17877 5865 17911 5899
rect 2789 5797 2823 5831
rect 8309 5797 8343 5831
rect 1685 5729 1719 5763
rect 1777 5729 1811 5763
rect 3341 5729 3375 5763
rect 3525 5729 3559 5763
rect 4537 5729 4571 5763
rect 6745 5729 6779 5763
rect 9413 5729 9447 5763
rect 11345 5729 11379 5763
rect 12081 5729 12115 5763
rect 14473 5729 14507 5763
rect 15945 5729 15979 5763
rect 16037 5729 16071 5763
rect 16313 5729 16347 5763
rect 16589 5729 16623 5763
rect 17417 5729 17451 5763
rect 1869 5661 1903 5695
rect 2605 5661 2639 5695
rect 4804 5661 4838 5695
rect 6561 5661 6595 5695
rect 7573 5661 7607 5695
rect 8125 5661 8159 5695
rect 8953 5661 8987 5695
rect 9505 5661 9539 5695
rect 10241 5661 10275 5695
rect 10793 5661 10827 5695
rect 13921 5661 13955 5695
rect 14749 5661 14783 5695
rect 17601 5661 17635 5695
rect 18061 5661 18095 5695
rect 18245 5661 18279 5695
rect 3249 5593 3283 5627
rect 6653 5593 6687 5627
rect 13737 5593 13771 5627
rect 14657 5593 14691 5627
rect 15853 5593 15887 5627
rect 2237 5525 2271 5559
rect 2421 5525 2455 5559
rect 3985 5525 4019 5559
rect 7113 5525 7147 5559
rect 9689 5525 9723 5559
rect 10701 5525 10735 5559
rect 11253 5525 11287 5559
rect 15209 5525 15243 5559
rect 17785 5525 17819 5559
rect 18429 5525 18463 5559
rect 1501 5321 1535 5355
rect 1961 5321 1995 5355
rect 2421 5321 2455 5355
rect 2605 5321 2639 5355
rect 3065 5321 3099 5355
rect 3433 5321 3467 5355
rect 3893 5321 3927 5355
rect 5641 5321 5675 5355
rect 13277 5321 13311 5355
rect 13645 5321 13679 5355
rect 14013 5321 14047 5355
rect 14473 5321 14507 5355
rect 14841 5321 14875 5355
rect 15301 5321 15335 5355
rect 16497 5321 16531 5355
rect 16681 5321 16715 5355
rect 17049 5321 17083 5355
rect 3801 5253 3835 5287
rect 6929 5253 6963 5287
rect 7757 5253 7791 5287
rect 12403 5253 12437 5287
rect 13185 5253 13219 5287
rect 15761 5253 15795 5287
rect 1685 5185 1719 5219
rect 1777 5185 1811 5219
rect 2145 5185 2179 5219
rect 2973 5185 3007 5219
rect 4261 5185 4295 5219
rect 4537 5185 4571 5219
rect 5733 5185 5767 5219
rect 8217 5185 8251 5219
rect 9505 5185 9539 5219
rect 11529 5185 11563 5219
rect 12300 5185 12334 5219
rect 14105 5185 14139 5219
rect 14933 5185 14967 5219
rect 15669 5185 15703 5219
rect 16129 5185 16163 5219
rect 17601 5185 17635 5219
rect 17877 5185 17911 5219
rect 18245 5185 18279 5219
rect 3157 5117 3191 5151
rect 3985 5117 4019 5151
rect 5549 5117 5583 5151
rect 6469 5117 6503 5151
rect 7021 5117 7055 5151
rect 7113 5117 7147 5151
rect 7849 5117 7883 5151
rect 7941 5117 7975 5151
rect 11713 5117 11747 5151
rect 12173 5117 12207 5151
rect 13369 5117 13403 5151
rect 14197 5117 14231 5151
rect 15025 5117 15059 5151
rect 15853 5117 15887 5151
rect 17141 5117 17175 5151
rect 17233 5117 17267 5151
rect 2329 5049 2363 5083
rect 9045 5049 9079 5083
rect 12817 5049 12851 5083
rect 17785 5049 17819 5083
rect 18429 5049 18463 5083
rect 6101 4981 6135 5015
rect 6561 4981 6595 5015
rect 7389 4981 7423 5015
rect 8493 4981 8527 5015
rect 8677 4981 8711 5015
rect 9229 4981 9263 5015
rect 16313 4981 16347 5015
rect 18061 4981 18095 5015
rect 1501 4777 1535 4811
rect 6193 4777 6227 4811
rect 8401 4777 8435 4811
rect 10609 4777 10643 4811
rect 12817 4777 12851 4811
rect 2697 4709 2731 4743
rect 3617 4709 3651 4743
rect 14381 4709 14415 4743
rect 15669 4709 15703 4743
rect 17601 4709 17635 4743
rect 5641 4641 5675 4675
rect 6745 4641 6779 4675
rect 6929 4641 6963 4675
rect 11345 4641 11379 4675
rect 11529 4641 11563 4675
rect 12173 4641 12207 4675
rect 13461 4641 13495 4675
rect 14749 4641 14783 4675
rect 15761 4641 15795 4675
rect 15945 4641 15979 4675
rect 1685 4573 1719 4607
rect 2053 4573 2087 4607
rect 2329 4573 2363 4607
rect 2605 4573 2639 4607
rect 2881 4573 2915 4607
rect 3157 4573 3191 4607
rect 3433 4573 3467 4607
rect 4261 4573 4295 4607
rect 6653 4573 6687 4607
rect 7481 4573 7515 4607
rect 8309 4573 8343 4607
rect 10333 4573 10367 4607
rect 12357 4573 12391 4607
rect 14565 4573 14599 4607
rect 14933 4573 14967 4607
rect 15509 4573 15543 4607
rect 16589 4573 16623 4607
rect 16865 4573 16899 4607
rect 17141 4573 17175 4607
rect 17417 4573 17451 4607
rect 17693 4573 17727 4607
rect 18153 4573 18187 4607
rect 18245 4573 18279 4607
rect 3801 4505 3835 4539
rect 5825 4505 5859 4539
rect 14289 4505 14323 4539
rect 15393 4505 15427 4539
rect 1869 4437 1903 4471
rect 2145 4437 2179 4471
rect 2421 4437 2455 4471
rect 2973 4437 3007 4471
rect 3249 4437 3283 4471
rect 4077 4437 4111 4471
rect 5733 4437 5767 4471
rect 6285 4437 6319 4471
rect 8769 4437 8803 4471
rect 10793 4437 10827 4471
rect 10885 4437 10919 4471
rect 13921 4437 13955 4471
rect 16129 4437 16163 4471
rect 16405 4437 16439 4471
rect 16773 4437 16807 4471
rect 17049 4437 17083 4471
rect 17325 4437 17359 4471
rect 17877 4437 17911 4471
rect 17969 4437 18003 4471
rect 18429 4437 18463 4471
rect 6101 4233 6135 4267
rect 6469 4233 6503 4267
rect 5733 4165 5767 4199
rect 1685 4097 1719 4131
rect 2053 4097 2087 4131
rect 2329 4097 2363 4131
rect 2605 4097 2639 4131
rect 2881 4097 2915 4131
rect 3157 4097 3191 4131
rect 3341 4097 3375 4131
rect 3893 4097 3927 4131
rect 9045 4097 9079 4131
rect 9137 4097 9171 4131
rect 10333 4097 10367 4131
rect 12357 4097 12391 4131
rect 13461 4097 13495 4131
rect 14105 4097 14139 4131
rect 14448 4097 14482 4131
rect 16681 4097 16715 4131
rect 16957 4097 16991 4131
rect 17233 4097 17267 4131
rect 17601 4097 17635 4131
rect 17877 4097 17911 4131
rect 18245 4097 18279 4131
rect 5549 4029 5583 4063
rect 5641 4029 5675 4063
rect 9321 4029 9355 4063
rect 10149 4029 10183 4063
rect 10793 4029 10827 4063
rect 12541 4029 12575 4063
rect 13001 4029 13035 4063
rect 15669 4029 15703 4063
rect 16313 4029 16347 4063
rect 16497 4029 16531 4063
rect 1501 3961 1535 3995
rect 2145 3961 2179 3995
rect 3525 3961 3559 3995
rect 9781 3961 9815 3995
rect 13921 3961 13955 3995
rect 14519 3961 14553 3995
rect 16865 3961 16899 3995
rect 17785 3961 17819 3995
rect 18061 3961 18095 3995
rect 1869 3893 1903 3927
rect 2421 3893 2455 3927
rect 2697 3893 2731 3927
rect 2973 3893 3007 3927
rect 3709 3893 3743 3927
rect 8585 3893 8619 3927
rect 8861 3893 8895 3927
rect 13093 3893 13127 3927
rect 13277 3893 13311 3927
rect 13645 3893 13679 3927
rect 13829 3893 13863 3927
rect 14197 3893 14231 3927
rect 17141 3893 17175 3927
rect 17417 3893 17451 3927
rect 18429 3893 18463 3927
rect 13829 3689 13863 3723
rect 16773 3689 16807 3723
rect 3433 3621 3467 3655
rect 8309 3621 8343 3655
rect 12541 3621 12575 3655
rect 17325 3621 17359 3655
rect 3985 3553 4019 3587
rect 8493 3553 8527 3587
rect 8677 3553 8711 3587
rect 14105 3553 14139 3587
rect 15853 3553 15887 3587
rect 16221 3553 16255 3587
rect 1685 3485 1719 3519
rect 2053 3485 2087 3519
rect 2421 3485 2455 3519
rect 2513 3485 2547 3519
rect 2881 3485 2915 3519
rect 3341 3485 3375 3519
rect 3617 3485 3651 3519
rect 3801 3485 3835 3519
rect 5549 3485 5583 3519
rect 6745 3485 6779 3519
rect 6837 3485 6871 3519
rect 7640 3485 7674 3519
rect 9137 3485 9171 3519
rect 9505 3485 9539 3519
rect 9632 3485 9666 3519
rect 10057 3485 10091 3519
rect 10333 3485 10367 3519
rect 10425 3485 10459 3519
rect 10920 3485 10954 3519
rect 11345 3485 11379 3519
rect 11805 3485 11839 3519
rect 12725 3485 12759 3519
rect 12817 3485 12851 3519
rect 13128 3485 13162 3519
rect 13404 3485 13438 3519
rect 13645 3485 13679 3519
rect 16037 3485 16071 3519
rect 16957 3485 16991 3519
rect 17141 3485 17175 3519
rect 17509 3485 17543 3519
rect 17877 3485 17911 3519
rect 18245 3485 18279 3519
rect 11529 3417 11563 3451
rect 13231 3417 13265 3451
rect 14289 3417 14323 3451
rect 1501 3349 1535 3383
rect 1869 3349 1903 3383
rect 2237 3349 2271 3383
rect 2697 3349 2731 3383
rect 3065 3349 3099 3383
rect 3157 3349 3191 3383
rect 5365 3349 5399 3383
rect 6561 3349 6595 3383
rect 7021 3349 7055 3383
rect 7711 3349 7745 3383
rect 8953 3349 8987 3383
rect 9321 3349 9355 3383
rect 9735 3349 9769 3383
rect 9873 3349 9907 3383
rect 10149 3349 10183 3383
rect 10609 3349 10643 3383
rect 11023 3349 11057 3383
rect 11161 3349 11195 3383
rect 11621 3349 11655 3383
rect 12449 3349 12483 3383
rect 13001 3349 13035 3383
rect 13507 3349 13541 3383
rect 16681 3349 16715 3383
rect 17693 3349 17727 3383
rect 18061 3349 18095 3383
rect 18429 3349 18463 3383
rect 3709 3145 3743 3179
rect 4537 3145 4571 3179
rect 16405 3145 16439 3179
rect 5089 3077 5123 3111
rect 9045 3077 9079 3111
rect 10977 3077 11011 3111
rect 11529 3077 11563 3111
rect 13645 3077 13679 3111
rect 1409 3009 1443 3043
rect 2145 3009 2179 3043
rect 2513 3009 2547 3043
rect 2605 3009 2639 3043
rect 3249 3009 3283 3043
rect 3341 3009 3375 3043
rect 3893 3009 3927 3043
rect 4169 3009 4203 3043
rect 4721 3009 4755 3043
rect 4997 3009 5031 3043
rect 5549 3009 5583 3043
rect 6745 3009 6779 3043
rect 6837 3009 6871 3043
rect 7113 3009 7147 3043
rect 9229 3009 9263 3043
rect 11161 3009 11195 3043
rect 13461 3009 13495 3043
rect 15510 3009 15544 3043
rect 15761 3009 15795 3043
rect 16313 3009 16347 3043
rect 16773 3009 16807 3043
rect 17417 3009 17451 3043
rect 17509 3009 17543 3043
rect 17877 3009 17911 3043
rect 18245 3009 18279 3043
rect 1961 2941 1995 2975
rect 8217 2941 8251 2975
rect 9505 2941 9539 2975
rect 13185 2941 13219 2975
rect 13369 2941 13403 2975
rect 14657 2941 14691 2975
rect 1593 2873 1627 2907
rect 2789 2873 2823 2907
rect 5365 2873 5399 2907
rect 17233 2873 17267 2907
rect 18061 2873 18095 2907
rect 2329 2805 2363 2839
rect 3065 2805 3099 2839
rect 3525 2805 3559 2839
rect 3985 2805 4019 2839
rect 4813 2805 4847 2839
rect 6561 2805 6595 2839
rect 7021 2805 7055 2839
rect 7297 2805 7331 2839
rect 11253 2805 11287 2839
rect 15439 2805 15473 2839
rect 15945 2805 15979 2839
rect 16129 2805 16163 2839
rect 16957 2805 16991 2839
rect 17693 2805 17727 2839
rect 18429 2805 18463 2839
rect 1501 2601 1535 2635
rect 1869 2601 1903 2635
rect 5181 2601 5215 2635
rect 6193 2601 6227 2635
rect 13737 2601 13771 2635
rect 11529 2533 11563 2567
rect 17233 2533 17267 2567
rect 11805 2465 11839 2499
rect 13553 2465 13587 2499
rect 14197 2465 14231 2499
rect 14381 2465 14415 2499
rect 15301 2465 15335 2499
rect 1685 2397 1719 2431
rect 2237 2397 2271 2431
rect 2697 2397 2731 2431
rect 3157 2397 3191 2431
rect 3617 2397 3651 2431
rect 4077 2397 4111 2431
rect 4537 2397 4571 2431
rect 4997 2397 5031 2431
rect 5365 2397 5399 2431
rect 5917 2397 5951 2431
rect 6009 2397 6043 2431
rect 6377 2397 6411 2431
rect 6561 2397 6595 2431
rect 7021 2397 7055 2431
rect 7481 2397 7515 2431
rect 7941 2397 7975 2431
rect 8677 2397 8711 2431
rect 9229 2397 9263 2431
rect 9597 2397 9631 2431
rect 10057 2397 10091 2431
rect 10517 2397 10551 2431
rect 10701 2397 10735 2431
rect 11136 2397 11170 2431
rect 11713 2397 11747 2431
rect 13921 2397 13955 2431
rect 16129 2397 16163 2431
rect 16681 2397 16715 2431
rect 17049 2397 17083 2431
rect 17417 2397 17451 2431
rect 17785 2397 17819 2431
rect 18153 2397 18187 2431
rect 11989 2329 12023 2363
rect 2053 2261 2087 2295
rect 2513 2261 2547 2295
rect 2973 2261 3007 2295
rect 3433 2261 3467 2295
rect 3893 2261 3927 2295
rect 4353 2261 4387 2295
rect 4813 2261 4847 2295
rect 5457 2261 5491 2295
rect 5733 2261 5767 2295
rect 6745 2261 6779 2295
rect 7205 2261 7239 2295
rect 7665 2261 7699 2295
rect 8125 2261 8159 2295
rect 8493 2261 8527 2295
rect 9045 2261 9079 2295
rect 9413 2261 9447 2295
rect 9873 2261 9907 2295
rect 10333 2261 10367 2295
rect 10885 2261 10919 2295
rect 11207 2261 11241 2295
rect 16313 2261 16347 2295
rect 16865 2261 16899 2295
rect 17601 2261 17635 2295
rect 17969 2261 18003 2295
rect 18337 2261 18371 2295
<< metal1 >>
rect 3786 15172 3792 15224
rect 3844 15212 3850 15224
rect 4706 15212 4712 15224
rect 3844 15184 4712 15212
rect 3844 15172 3850 15184
rect 4706 15172 4712 15184
rect 4764 15172 4770 15224
rect 5902 14968 5908 15020
rect 5960 15008 5966 15020
rect 14918 15008 14924 15020
rect 5960 14980 14924 15008
rect 5960 14968 5966 14980
rect 14918 14968 14924 14980
rect 14976 14968 14982 15020
rect 2130 14900 2136 14952
rect 2188 14940 2194 14952
rect 7466 14940 7472 14952
rect 2188 14912 7472 14940
rect 2188 14900 2194 14912
rect 7466 14900 7472 14912
rect 7524 14900 7530 14952
rect 8754 14900 8760 14952
rect 8812 14940 8818 14952
rect 16390 14940 16396 14952
rect 8812 14912 16396 14940
rect 8812 14900 8818 14912
rect 16390 14900 16396 14912
rect 16448 14900 16454 14952
rect 4522 14832 4528 14884
rect 4580 14872 4586 14884
rect 4580 14844 8524 14872
rect 4580 14832 4586 14844
rect 3970 14764 3976 14816
rect 4028 14804 4034 14816
rect 7006 14804 7012 14816
rect 4028 14776 7012 14804
rect 4028 14764 4034 14776
rect 7006 14764 7012 14776
rect 7064 14764 7070 14816
rect 8496 14804 8524 14844
rect 11330 14832 11336 14884
rect 11388 14872 11394 14884
rect 18966 14872 18972 14884
rect 11388 14844 18972 14872
rect 11388 14832 11394 14844
rect 18966 14832 18972 14844
rect 19024 14832 19030 14884
rect 12434 14804 12440 14816
rect 8496 14776 12440 14804
rect 12434 14764 12440 14776
rect 12492 14764 12498 14816
rect 12618 14764 12624 14816
rect 12676 14804 12682 14816
rect 13538 14804 13544 14816
rect 12676 14776 13544 14804
rect 12676 14764 12682 14776
rect 13538 14764 13544 14776
rect 13596 14804 13602 14816
rect 18322 14804 18328 14816
rect 13596 14776 18328 14804
rect 13596 14764 13602 14776
rect 18322 14764 18328 14776
rect 18380 14764 18386 14816
rect 1104 14714 18860 14736
rect 1104 14662 3174 14714
rect 3226 14662 3238 14714
rect 3290 14662 3302 14714
rect 3354 14662 3366 14714
rect 3418 14662 3430 14714
rect 3482 14662 7622 14714
rect 7674 14662 7686 14714
rect 7738 14662 7750 14714
rect 7802 14662 7814 14714
rect 7866 14662 7878 14714
rect 7930 14662 12070 14714
rect 12122 14662 12134 14714
rect 12186 14662 12198 14714
rect 12250 14662 12262 14714
rect 12314 14662 12326 14714
rect 12378 14662 16518 14714
rect 16570 14662 16582 14714
rect 16634 14662 16646 14714
rect 16698 14662 16710 14714
rect 16762 14662 16774 14714
rect 16826 14662 18860 14714
rect 1104 14640 18860 14662
rect 3421 14603 3479 14609
rect 3421 14569 3433 14603
rect 3467 14600 3479 14603
rect 3510 14600 3516 14612
rect 3467 14572 3516 14600
rect 3467 14569 3479 14572
rect 3421 14563 3479 14569
rect 3510 14560 3516 14572
rect 3568 14560 3574 14612
rect 5534 14560 5540 14612
rect 5592 14600 5598 14612
rect 5721 14603 5779 14609
rect 5721 14600 5733 14603
rect 5592 14572 5733 14600
rect 5592 14560 5598 14572
rect 5721 14569 5733 14572
rect 5767 14569 5779 14603
rect 5721 14563 5779 14569
rect 6086 14560 6092 14612
rect 6144 14600 6150 14612
rect 6546 14600 6552 14612
rect 6144 14572 6552 14600
rect 6144 14560 6150 14572
rect 6546 14560 6552 14572
rect 6604 14600 6610 14612
rect 6641 14603 6699 14609
rect 6641 14600 6653 14603
rect 6604 14572 6653 14600
rect 6604 14560 6610 14572
rect 6641 14569 6653 14572
rect 6687 14569 6699 14603
rect 6641 14563 6699 14569
rect 6730 14560 6736 14612
rect 6788 14600 6794 14612
rect 7009 14603 7067 14609
rect 7009 14600 7021 14603
rect 6788 14572 7021 14600
rect 6788 14560 6794 14572
rect 7009 14569 7021 14572
rect 7055 14569 7067 14603
rect 7374 14600 7380 14612
rect 7335 14572 7380 14600
rect 7009 14563 7067 14569
rect 7374 14560 7380 14572
rect 7432 14560 7438 14612
rect 8662 14600 8668 14612
rect 8623 14572 8668 14600
rect 8662 14560 8668 14572
rect 8720 14560 8726 14612
rect 9306 14600 9312 14612
rect 9267 14572 9312 14600
rect 9306 14560 9312 14572
rect 9364 14560 9370 14612
rect 9950 14600 9956 14612
rect 9911 14572 9956 14600
rect 9950 14560 9956 14572
rect 10008 14560 10014 14612
rect 10594 14600 10600 14612
rect 10555 14572 10600 14600
rect 10594 14560 10600 14572
rect 10652 14560 10658 14612
rect 11238 14560 11244 14612
rect 11296 14600 11302 14612
rect 11793 14603 11851 14609
rect 11793 14600 11805 14603
rect 11296 14572 11805 14600
rect 11296 14560 11302 14572
rect 2958 14492 2964 14544
rect 3016 14532 3022 14544
rect 6822 14532 6828 14544
rect 3016 14504 6828 14532
rect 3016 14492 3022 14504
rect 3160 14473 3188 14504
rect 6822 14492 6828 14504
rect 6880 14492 6886 14544
rect 10229 14535 10287 14541
rect 10229 14501 10241 14535
rect 10275 14532 10287 14535
rect 11054 14532 11060 14544
rect 10275 14504 11060 14532
rect 10275 14501 10287 14504
rect 10229 14495 10287 14501
rect 11054 14492 11060 14504
rect 11112 14492 11118 14544
rect 3145 14467 3203 14473
rect 2746 14436 3004 14464
rect 1946 14396 1952 14408
rect 1907 14368 1952 14396
rect 1946 14356 1952 14368
rect 2004 14356 2010 14408
rect 2222 14396 2228 14408
rect 2183 14368 2228 14396
rect 2222 14356 2228 14368
rect 2280 14396 2286 14408
rect 2746 14396 2774 14436
rect 2280 14368 2774 14396
rect 2869 14399 2927 14405
rect 2280 14356 2286 14368
rect 2869 14365 2881 14399
rect 2915 14365 2927 14399
rect 2976 14396 3004 14436
rect 3145 14433 3157 14467
rect 3191 14433 3203 14467
rect 3970 14464 3976 14476
rect 3145 14427 3203 14433
rect 3436 14436 3976 14464
rect 3436 14396 3464 14436
rect 3970 14424 3976 14436
rect 4028 14424 4034 14476
rect 4154 14424 4160 14476
rect 4212 14464 4218 14476
rect 4617 14467 4675 14473
rect 4617 14464 4629 14467
rect 4212 14436 4629 14464
rect 4212 14424 4218 14436
rect 4617 14433 4629 14436
rect 4663 14464 4675 14467
rect 5997 14467 6055 14473
rect 5997 14464 6009 14467
rect 4663 14436 6009 14464
rect 4663 14433 4675 14436
rect 4617 14427 4675 14433
rect 5997 14433 6009 14436
rect 6043 14433 6055 14467
rect 5997 14427 6055 14433
rect 6178 14424 6184 14476
rect 6236 14464 6242 14476
rect 6236 14436 6684 14464
rect 6236 14424 6242 14436
rect 3602 14396 3608 14408
rect 2976 14368 3464 14396
rect 3563 14368 3608 14396
rect 2869 14359 2927 14365
rect 2884 14328 2912 14359
rect 3602 14356 3608 14368
rect 3660 14356 3666 14408
rect 4341 14399 4399 14405
rect 4341 14365 4353 14399
rect 4387 14396 4399 14399
rect 4430 14396 4436 14408
rect 4387 14368 4436 14396
rect 4387 14365 4399 14368
rect 4341 14359 4399 14365
rect 4430 14356 4436 14368
rect 4488 14356 4494 14408
rect 4706 14396 4712 14408
rect 4667 14368 4712 14396
rect 4706 14356 4712 14368
rect 4764 14356 4770 14408
rect 4982 14396 4988 14408
rect 4943 14368 4988 14396
rect 4982 14356 4988 14368
rect 5040 14356 5046 14408
rect 5902 14396 5908 14408
rect 5863 14368 5908 14396
rect 5902 14356 5908 14368
rect 5960 14356 5966 14408
rect 6546 14396 6552 14408
rect 6507 14368 6552 14396
rect 6546 14356 6552 14368
rect 6604 14356 6610 14408
rect 6656 14396 6684 14436
rect 6825 14399 6883 14405
rect 6825 14396 6837 14399
rect 6656 14368 6837 14396
rect 6825 14365 6837 14368
rect 6871 14365 6883 14399
rect 6825 14359 6883 14365
rect 7374 14356 7380 14408
rect 7432 14396 7438 14408
rect 7469 14399 7527 14405
rect 7469 14396 7481 14399
rect 7432 14368 7481 14396
rect 7432 14356 7438 14368
rect 7469 14365 7481 14368
rect 7515 14365 7527 14399
rect 7469 14359 7527 14365
rect 8662 14356 8668 14408
rect 8720 14396 8726 14408
rect 9125 14399 9183 14405
rect 9125 14396 9137 14399
rect 8720 14368 9137 14396
rect 8720 14356 8726 14368
rect 9125 14365 9137 14368
rect 9171 14365 9183 14399
rect 9125 14359 9183 14365
rect 9306 14356 9312 14408
rect 9364 14396 9370 14408
rect 9585 14399 9643 14405
rect 9585 14396 9597 14399
rect 9364 14368 9597 14396
rect 9364 14356 9370 14368
rect 9585 14365 9597 14368
rect 9631 14365 9643 14399
rect 9585 14359 9643 14365
rect 9950 14356 9956 14408
rect 10008 14396 10014 14408
rect 10045 14399 10103 14405
rect 10045 14396 10057 14399
rect 10008 14368 10057 14396
rect 10008 14356 10014 14368
rect 10045 14365 10057 14368
rect 10091 14365 10103 14399
rect 10045 14359 10103 14365
rect 10594 14356 10600 14408
rect 10652 14396 10658 14408
rect 11716 14405 11744 14572
rect 11793 14569 11805 14572
rect 11839 14569 11851 14603
rect 12526 14600 12532 14612
rect 12487 14572 12532 14600
rect 11793 14563 11851 14569
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 13170 14600 13176 14612
rect 13131 14572 13176 14600
rect 13170 14560 13176 14572
rect 13228 14560 13234 14612
rect 14277 14535 14335 14541
rect 14277 14501 14289 14535
rect 14323 14532 14335 14535
rect 15286 14532 15292 14544
rect 14323 14504 15292 14532
rect 14323 14501 14335 14504
rect 14277 14495 14335 14501
rect 15286 14492 15292 14504
rect 15344 14492 15350 14544
rect 12894 14424 12900 14476
rect 12952 14464 12958 14476
rect 14182 14464 14188 14476
rect 12952 14436 14188 14464
rect 12952 14424 12958 14436
rect 14182 14424 14188 14436
rect 14240 14424 14246 14476
rect 15105 14467 15163 14473
rect 15105 14433 15117 14467
rect 15151 14464 15163 14467
rect 16758 14464 16764 14476
rect 15151 14436 16764 14464
rect 15151 14433 15163 14436
rect 15105 14427 15163 14433
rect 16758 14424 16764 14436
rect 16816 14424 16822 14476
rect 10873 14399 10931 14405
rect 10873 14396 10885 14399
rect 10652 14368 10885 14396
rect 10652 14356 10658 14368
rect 10873 14365 10885 14368
rect 10919 14365 10931 14399
rect 10873 14359 10931 14365
rect 11701 14399 11759 14405
rect 11701 14365 11713 14399
rect 11747 14365 11759 14399
rect 11974 14396 11980 14408
rect 11935 14368 11980 14396
rect 11701 14359 11759 14365
rect 11974 14356 11980 14368
rect 12032 14396 12038 14408
rect 12253 14399 12311 14405
rect 12253 14396 12265 14399
rect 12032 14368 12265 14396
rect 12032 14356 12038 14368
rect 12253 14365 12265 14368
rect 12299 14365 12311 14399
rect 12253 14359 12311 14365
rect 12526 14356 12532 14408
rect 12584 14396 12590 14408
rect 12805 14399 12863 14405
rect 12805 14396 12817 14399
rect 12584 14368 12817 14396
rect 12584 14356 12590 14368
rect 12805 14365 12817 14368
rect 12851 14365 12863 14399
rect 12805 14359 12863 14365
rect 13170 14356 13176 14408
rect 13228 14396 13234 14408
rect 13265 14399 13323 14405
rect 13265 14396 13277 14399
rect 13228 14368 13277 14396
rect 13228 14356 13234 14368
rect 13265 14365 13277 14368
rect 13311 14365 13323 14399
rect 13265 14359 13323 14365
rect 13814 14356 13820 14408
rect 13872 14396 13878 14408
rect 14093 14399 14151 14405
rect 14093 14396 14105 14399
rect 13872 14368 14105 14396
rect 13872 14356 13878 14368
rect 14093 14365 14105 14368
rect 14139 14396 14151 14399
rect 14369 14399 14427 14405
rect 14369 14396 14381 14399
rect 14139 14368 14381 14396
rect 14139 14365 14151 14368
rect 14093 14359 14151 14365
rect 14369 14365 14381 14368
rect 14415 14365 14427 14399
rect 14369 14359 14427 14365
rect 15289 14399 15347 14405
rect 15289 14365 15301 14399
rect 15335 14396 15347 14399
rect 15470 14396 15476 14408
rect 15335 14368 15476 14396
rect 15335 14365 15347 14368
rect 15289 14359 15347 14365
rect 15470 14356 15476 14368
rect 15528 14396 15534 14408
rect 15565 14399 15623 14405
rect 15565 14396 15577 14399
rect 15528 14368 15577 14396
rect 15528 14356 15534 14368
rect 15565 14365 15577 14368
rect 15611 14365 15623 14399
rect 15565 14359 15623 14365
rect 16022 14356 16028 14408
rect 16080 14396 16086 14408
rect 16209 14399 16267 14405
rect 16209 14396 16221 14399
rect 16080 14368 16221 14396
rect 16080 14356 16086 14368
rect 16209 14365 16221 14368
rect 16255 14365 16267 14399
rect 16209 14359 16267 14365
rect 16298 14356 16304 14408
rect 16356 14396 16362 14408
rect 16485 14399 16543 14405
rect 16485 14396 16497 14399
rect 16356 14368 16497 14396
rect 16356 14356 16362 14368
rect 16485 14365 16497 14368
rect 16531 14396 16543 14399
rect 16942 14396 16948 14408
rect 16531 14368 16948 14396
rect 16531 14365 16543 14368
rect 16485 14359 16543 14365
rect 16942 14356 16948 14368
rect 17000 14356 17006 14408
rect 17037 14399 17095 14405
rect 17037 14365 17049 14399
rect 17083 14396 17095 14399
rect 17218 14396 17224 14408
rect 17083 14368 17224 14396
rect 17083 14365 17095 14368
rect 17037 14359 17095 14365
rect 17218 14356 17224 14368
rect 17276 14356 17282 14408
rect 17678 14396 17684 14408
rect 17639 14368 17684 14396
rect 17678 14356 17684 14368
rect 17736 14356 17742 14408
rect 17954 14396 17960 14408
rect 17915 14368 17960 14396
rect 17954 14356 17960 14368
rect 18012 14356 18018 14408
rect 4246 14328 4252 14340
rect 2884 14300 4252 14328
rect 4246 14288 4252 14300
rect 4304 14288 4310 14340
rect 5166 14288 5172 14340
rect 5224 14328 5230 14340
rect 13354 14328 13360 14340
rect 5224 14300 6500 14328
rect 5224 14288 5230 14300
rect 3142 14220 3148 14272
rect 3200 14260 3206 14272
rect 5810 14260 5816 14272
rect 3200 14232 5816 14260
rect 3200 14220 3206 14232
rect 5810 14220 5816 14232
rect 5868 14220 5874 14272
rect 6362 14260 6368 14272
rect 6323 14232 6368 14260
rect 6362 14220 6368 14232
rect 6420 14220 6426 14272
rect 6472 14260 6500 14300
rect 7576 14300 13360 14328
rect 7576 14260 7604 14300
rect 13354 14288 13360 14300
rect 13412 14288 13418 14340
rect 6472 14232 7604 14260
rect 7653 14263 7711 14269
rect 7653 14229 7665 14263
rect 7699 14260 7711 14263
rect 8110 14260 8116 14272
rect 7699 14232 8116 14260
rect 7699 14229 7711 14232
rect 7653 14223 7711 14229
rect 8110 14220 8116 14232
rect 8168 14220 8174 14272
rect 8662 14220 8668 14272
rect 8720 14260 8726 14272
rect 8941 14263 8999 14269
rect 8941 14260 8953 14263
rect 8720 14232 8953 14260
rect 8720 14220 8726 14232
rect 8941 14229 8953 14232
rect 8987 14229 8999 14263
rect 8941 14223 8999 14229
rect 9030 14220 9036 14272
rect 9088 14260 9094 14272
rect 9401 14263 9459 14269
rect 9401 14260 9413 14263
rect 9088 14232 9413 14260
rect 9088 14220 9094 14232
rect 9401 14229 9413 14232
rect 9447 14229 9459 14263
rect 10686 14260 10692 14272
rect 10647 14232 10692 14260
rect 9401 14223 9459 14229
rect 10686 14220 10692 14232
rect 10744 14220 10750 14272
rect 11422 14220 11428 14272
rect 11480 14260 11486 14272
rect 11517 14263 11575 14269
rect 11517 14260 11529 14263
rect 11480 14232 11529 14260
rect 11480 14220 11486 14232
rect 11517 14229 11529 14232
rect 11563 14229 11575 14263
rect 11517 14223 11575 14229
rect 11790 14220 11796 14272
rect 11848 14260 11854 14272
rect 12161 14263 12219 14269
rect 12161 14260 12173 14263
rect 11848 14232 12173 14260
rect 11848 14220 11854 14232
rect 12161 14229 12173 14232
rect 12207 14229 12219 14263
rect 12161 14223 12219 14229
rect 12621 14263 12679 14269
rect 12621 14229 12633 14263
rect 12667 14260 12679 14263
rect 12710 14260 12716 14272
rect 12667 14232 12716 14260
rect 12667 14229 12679 14232
rect 12621 14223 12679 14229
rect 12710 14220 12716 14232
rect 12768 14220 12774 14272
rect 13449 14263 13507 14269
rect 13449 14229 13461 14263
rect 13495 14260 13507 14263
rect 13722 14260 13728 14272
rect 13495 14232 13728 14260
rect 13495 14229 13507 14232
rect 13449 14223 13507 14229
rect 13722 14220 13728 14232
rect 13780 14220 13786 14272
rect 15378 14260 15384 14272
rect 15339 14232 15384 14260
rect 15378 14220 15384 14232
rect 15436 14220 15442 14272
rect 1104 14170 18860 14192
rect 1104 14118 5398 14170
rect 5450 14118 5462 14170
rect 5514 14118 5526 14170
rect 5578 14118 5590 14170
rect 5642 14118 5654 14170
rect 5706 14118 9846 14170
rect 9898 14118 9910 14170
rect 9962 14118 9974 14170
rect 10026 14118 10038 14170
rect 10090 14118 10102 14170
rect 10154 14118 14294 14170
rect 14346 14118 14358 14170
rect 14410 14118 14422 14170
rect 14474 14118 14486 14170
rect 14538 14118 14550 14170
rect 14602 14118 18860 14170
rect 1104 14096 18860 14118
rect 2774 14016 2780 14068
rect 2832 14056 2838 14068
rect 3050 14056 3056 14068
rect 2832 14028 3056 14056
rect 2832 14016 2838 14028
rect 3050 14016 3056 14028
rect 3108 14056 3114 14068
rect 3510 14056 3516 14068
rect 3108 14028 3516 14056
rect 3108 14016 3114 14028
rect 3510 14016 3516 14028
rect 3568 14016 3574 14068
rect 4338 14056 4344 14068
rect 4299 14028 4344 14056
rect 4338 14016 4344 14028
rect 4396 14016 4402 14068
rect 4706 14056 4712 14068
rect 4667 14028 4712 14056
rect 4706 14016 4712 14028
rect 4764 14016 4770 14068
rect 4798 14016 4804 14068
rect 4856 14056 4862 14068
rect 4985 14059 5043 14065
rect 4985 14056 4997 14059
rect 4856 14028 4997 14056
rect 4856 14016 4862 14028
rect 4985 14025 4997 14028
rect 5031 14025 5043 14059
rect 6270 14056 6276 14068
rect 4985 14019 5043 14025
rect 5092 14028 6276 14056
rect 2038 13948 2044 14000
rect 2096 13988 2102 14000
rect 5092 13988 5120 14028
rect 6270 14016 6276 14028
rect 6328 14016 6334 14068
rect 6454 14016 6460 14068
rect 6512 14016 6518 14068
rect 6638 14016 6644 14068
rect 6696 14056 6702 14068
rect 8113 14059 8171 14065
rect 8113 14056 8125 14059
rect 6696 14028 8125 14056
rect 6696 14016 6702 14028
rect 8113 14025 8125 14028
rect 8159 14025 8171 14059
rect 8113 14019 8171 14025
rect 8665 14059 8723 14065
rect 8665 14025 8677 14059
rect 8711 14056 8723 14059
rect 8754 14056 8760 14068
rect 8711 14028 8760 14056
rect 8711 14025 8723 14028
rect 8665 14019 8723 14025
rect 2096 13960 5120 13988
rect 2096 13948 2102 13960
rect 1949 13923 2007 13929
rect 1949 13889 1961 13923
rect 1995 13920 2007 13923
rect 2130 13920 2136 13932
rect 1995 13892 2136 13920
rect 1995 13889 2007 13892
rect 1949 13883 2007 13889
rect 2130 13880 2136 13892
rect 2188 13880 2194 13932
rect 2240 13929 2268 13960
rect 2225 13923 2283 13929
rect 2225 13889 2237 13923
rect 2271 13889 2283 13923
rect 2225 13883 2283 13889
rect 2869 13923 2927 13929
rect 2869 13889 2881 13923
rect 2915 13920 2927 13923
rect 3694 13920 3700 13932
rect 2915 13892 3700 13920
rect 2915 13889 2927 13892
rect 2869 13883 2927 13889
rect 3694 13880 3700 13892
rect 3752 13880 3758 13932
rect 4062 13920 4068 13932
rect 4023 13892 4068 13920
rect 4062 13880 4068 13892
rect 4120 13880 4126 13932
rect 4522 13920 4528 13932
rect 4483 13892 4528 13920
rect 4522 13880 4528 13892
rect 4580 13880 4586 13932
rect 5166 13920 5172 13932
rect 5127 13892 5172 13920
rect 5166 13880 5172 13892
rect 5224 13880 5230 13932
rect 5534 13920 5540 13932
rect 5495 13892 5540 13920
rect 5534 13880 5540 13892
rect 5592 13880 5598 13932
rect 5810 13920 5816 13932
rect 5771 13892 5816 13920
rect 5810 13880 5816 13892
rect 5868 13880 5874 13932
rect 5997 13923 6055 13929
rect 5997 13889 6009 13923
rect 6043 13889 6055 13923
rect 5997 13883 6055 13889
rect 6365 13923 6423 13929
rect 6365 13889 6377 13923
rect 6411 13920 6423 13923
rect 6472 13920 6500 14016
rect 6411 13892 6500 13920
rect 6411 13889 6423 13892
rect 6365 13883 6423 13889
rect 3142 13852 3148 13864
rect 3103 13824 3148 13852
rect 3142 13812 3148 13824
rect 3200 13812 3206 13864
rect 3602 13812 3608 13864
rect 3660 13852 3666 13864
rect 3789 13855 3847 13861
rect 3789 13852 3801 13855
rect 3660 13824 3801 13852
rect 3660 13812 3666 13824
rect 3789 13821 3801 13824
rect 3835 13821 3847 13855
rect 3789 13815 3847 13821
rect 4172 13824 5396 13852
rect 934 13744 940 13796
rect 992 13784 998 13796
rect 4172 13784 4200 13824
rect 5368 13793 5396 13824
rect 5442 13812 5448 13864
rect 5500 13852 5506 13864
rect 6012 13852 6040 13883
rect 6546 13880 6552 13932
rect 6604 13920 6610 13932
rect 6825 13923 6883 13929
rect 6825 13920 6837 13923
rect 6604 13892 6837 13920
rect 6604 13880 6610 13892
rect 6825 13889 6837 13892
rect 6871 13889 6883 13923
rect 7006 13920 7012 13932
rect 6967 13892 7012 13920
rect 6825 13883 6883 13889
rect 7006 13880 7012 13892
rect 7064 13880 7070 13932
rect 7469 13923 7527 13929
rect 7469 13889 7481 13923
rect 7515 13920 7527 13923
rect 8021 13923 8079 13929
rect 7515 13892 7696 13920
rect 7515 13889 7527 13892
rect 7469 13883 7527 13889
rect 5500 13824 5948 13852
rect 6012 13824 6408 13852
rect 5500 13812 5506 13824
rect 992 13756 4200 13784
rect 5353 13787 5411 13793
rect 992 13744 998 13756
rect 5353 13753 5365 13787
rect 5399 13753 5411 13787
rect 5920 13784 5948 13824
rect 6380 13796 6408 13824
rect 6472 13824 7236 13852
rect 6178 13784 6184 13796
rect 5920 13756 6040 13784
rect 6139 13756 6184 13784
rect 5353 13747 5411 13753
rect 1946 13676 1952 13728
rect 2004 13716 2010 13728
rect 3970 13716 3976 13728
rect 2004 13688 3976 13716
rect 2004 13676 2010 13688
rect 3970 13676 3976 13688
rect 4028 13676 4034 13728
rect 4062 13676 4068 13728
rect 4120 13716 4126 13728
rect 5629 13719 5687 13725
rect 5629 13716 5641 13719
rect 4120 13688 5641 13716
rect 4120 13676 4126 13688
rect 5629 13685 5641 13688
rect 5675 13685 5687 13719
rect 6012 13716 6040 13756
rect 6178 13744 6184 13756
rect 6236 13744 6242 13796
rect 6362 13744 6368 13796
rect 6420 13744 6426 13796
rect 6472 13716 6500 13824
rect 6549 13787 6607 13793
rect 6549 13753 6561 13787
rect 6595 13784 6607 13787
rect 6730 13784 6736 13796
rect 6595 13756 6736 13784
rect 6595 13753 6607 13756
rect 6549 13747 6607 13753
rect 6730 13744 6736 13756
rect 6788 13744 6794 13796
rect 7208 13784 7236 13824
rect 7208 13756 7328 13784
rect 6012 13688 6500 13716
rect 6641 13719 6699 13725
rect 5629 13679 5687 13685
rect 6641 13685 6653 13719
rect 6687 13716 6699 13719
rect 6822 13716 6828 13728
rect 6687 13688 6828 13716
rect 6687 13685 6699 13688
rect 6641 13679 6699 13685
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 7300 13725 7328 13756
rect 7668 13725 7696 13892
rect 8021 13889 8033 13923
rect 8067 13889 8079 13923
rect 8021 13883 8079 13889
rect 8297 13923 8355 13929
rect 8297 13889 8309 13923
rect 8343 13920 8355 13923
rect 8680 13920 8708 14019
rect 8754 14016 8760 14028
rect 8812 14016 8818 14068
rect 11057 14059 11115 14065
rect 11057 14025 11069 14059
rect 11103 14056 11115 14059
rect 11146 14056 11152 14068
rect 11103 14028 11152 14056
rect 11103 14025 11115 14028
rect 11057 14019 11115 14025
rect 11146 14016 11152 14028
rect 11204 14016 11210 14068
rect 11698 14056 11704 14068
rect 11348 14028 11704 14056
rect 11348 14000 11376 14028
rect 11698 14016 11704 14028
rect 11756 14016 11762 14068
rect 12434 14016 12440 14068
rect 12492 14056 12498 14068
rect 12529 14059 12587 14065
rect 12529 14056 12541 14059
rect 12492 14028 12541 14056
rect 12492 14016 12498 14028
rect 12529 14025 12541 14028
rect 12575 14025 12587 14059
rect 13262 14056 13268 14068
rect 13223 14028 13268 14056
rect 12529 14019 12587 14025
rect 13262 14016 13268 14028
rect 13320 14016 13326 14068
rect 14001 14059 14059 14065
rect 14001 14056 14013 14059
rect 13648 14028 14013 14056
rect 10229 13991 10287 13997
rect 10229 13988 10241 13991
rect 10060 13960 10241 13988
rect 10060 13929 10088 13960
rect 10229 13957 10241 13960
rect 10275 13988 10287 13991
rect 11330 13988 11336 14000
rect 10275 13960 11336 13988
rect 10275 13957 10287 13960
rect 10229 13951 10287 13957
rect 11330 13948 11336 13960
rect 11388 13948 11394 14000
rect 11609 13991 11667 13997
rect 11609 13957 11621 13991
rect 11655 13988 11667 13991
rect 12618 13988 12624 14000
rect 11655 13960 12624 13988
rect 11655 13957 11667 13960
rect 11609 13951 11667 13957
rect 8343 13892 8708 13920
rect 10045 13923 10103 13929
rect 8343 13889 8355 13892
rect 8297 13883 8355 13889
rect 10045 13889 10057 13923
rect 10091 13889 10103 13923
rect 10045 13883 10103 13889
rect 11241 13923 11299 13929
rect 11241 13889 11253 13923
rect 11287 13920 11299 13923
rect 11624 13920 11652 13951
rect 12618 13948 12624 13960
rect 12676 13948 12682 14000
rect 11287 13892 11652 13920
rect 12713 13923 12771 13929
rect 11287 13889 11299 13892
rect 11241 13883 11299 13889
rect 12713 13889 12725 13923
rect 12759 13920 12771 13923
rect 12894 13920 12900 13932
rect 12759 13892 12900 13920
rect 12759 13889 12771 13892
rect 12713 13883 12771 13889
rect 8036 13852 8064 13883
rect 12894 13880 12900 13892
rect 12952 13880 12958 13932
rect 13449 13923 13507 13929
rect 13449 13889 13461 13923
rect 13495 13920 13507 13923
rect 13648 13920 13676 14028
rect 14001 14025 14013 14028
rect 14047 14025 14059 14059
rect 14918 14056 14924 14068
rect 14879 14028 14924 14056
rect 14001 14019 14059 14025
rect 14016 13988 14044 14019
rect 14918 14016 14924 14028
rect 14976 14016 14982 14068
rect 15838 13988 15844 14000
rect 14016 13960 15844 13988
rect 15838 13948 15844 13960
rect 15896 13948 15902 14000
rect 13495 13892 13676 13920
rect 13825 13923 13883 13929
rect 13495 13889 13507 13892
rect 13449 13883 13507 13889
rect 13825 13889 13837 13923
rect 13871 13920 13883 13923
rect 15010 13920 15016 13932
rect 13871 13892 15016 13920
rect 13871 13889 13883 13892
rect 13825 13883 13883 13889
rect 15010 13880 15016 13892
rect 15068 13880 15074 13932
rect 15105 13923 15163 13929
rect 15105 13889 15117 13923
rect 15151 13920 15163 13923
rect 15746 13920 15752 13932
rect 15151 13892 15752 13920
rect 15151 13889 15163 13892
rect 15105 13883 15163 13889
rect 15746 13880 15752 13892
rect 15804 13880 15810 13932
rect 15933 13923 15991 13929
rect 15933 13889 15945 13923
rect 15979 13920 15991 13923
rect 16206 13920 16212 13932
rect 15979 13892 16212 13920
rect 15979 13889 15991 13892
rect 15933 13883 15991 13889
rect 16206 13880 16212 13892
rect 16264 13880 16270 13932
rect 16482 13920 16488 13932
rect 16443 13892 16488 13920
rect 16482 13880 16488 13892
rect 16540 13880 16546 13932
rect 17957 13923 18015 13929
rect 17957 13920 17969 13923
rect 16592 13892 17969 13920
rect 8481 13855 8539 13861
rect 8481 13852 8493 13855
rect 8036 13824 8493 13852
rect 8481 13821 8493 13824
rect 8527 13852 8539 13855
rect 9490 13852 9496 13864
rect 8527 13824 9496 13852
rect 8527 13821 8539 13824
rect 8481 13815 8539 13821
rect 9490 13812 9496 13824
rect 9548 13812 9554 13864
rect 11882 13812 11888 13864
rect 11940 13852 11946 13864
rect 16592 13852 16620 13892
rect 17957 13889 17969 13892
rect 18003 13889 18015 13923
rect 17957 13883 18015 13889
rect 16758 13852 16764 13864
rect 11940 13824 16620 13852
rect 16719 13824 16764 13852
rect 11940 13812 11946 13824
rect 16758 13812 16764 13824
rect 16816 13812 16822 13864
rect 17037 13855 17095 13861
rect 17037 13852 17049 13855
rect 16868 13824 17049 13852
rect 7834 13784 7840 13796
rect 7795 13756 7840 13784
rect 7834 13744 7840 13756
rect 7892 13744 7898 13796
rect 9674 13744 9680 13796
rect 9732 13784 9738 13796
rect 16025 13787 16083 13793
rect 16025 13784 16037 13787
rect 9732 13756 16037 13784
rect 9732 13744 9738 13756
rect 16025 13753 16037 13756
rect 16071 13753 16083 13787
rect 16025 13747 16083 13753
rect 16114 13744 16120 13796
rect 16172 13784 16178 13796
rect 16868 13784 16896 13824
rect 17037 13821 17049 13824
rect 17083 13821 17095 13855
rect 17037 13815 17095 13821
rect 17681 13855 17739 13861
rect 17681 13821 17693 13855
rect 17727 13852 17739 13855
rect 17770 13852 17776 13864
rect 17727 13824 17776 13852
rect 17727 13821 17739 13824
rect 17681 13815 17739 13821
rect 17770 13812 17776 13824
rect 17828 13812 17834 13864
rect 16172 13756 16896 13784
rect 16172 13744 16178 13756
rect 7285 13719 7343 13725
rect 7285 13685 7297 13719
rect 7331 13685 7343 13719
rect 7285 13679 7343 13685
rect 7653 13719 7711 13725
rect 7653 13685 7665 13719
rect 7699 13716 7711 13719
rect 8294 13716 8300 13728
rect 7699 13688 8300 13716
rect 7699 13685 7711 13688
rect 7653 13679 7711 13685
rect 8294 13676 8300 13688
rect 8352 13676 8358 13728
rect 9858 13716 9864 13728
rect 9819 13688 9864 13716
rect 9858 13676 9864 13688
rect 9916 13676 9922 13728
rect 13354 13676 13360 13728
rect 13412 13716 13418 13728
rect 13633 13719 13691 13725
rect 13633 13716 13645 13719
rect 13412 13688 13645 13716
rect 13412 13676 13418 13688
rect 13633 13685 13645 13688
rect 13679 13685 13691 13719
rect 16298 13716 16304 13728
rect 16259 13688 16304 13716
rect 13633 13679 13691 13685
rect 16298 13676 16304 13688
rect 16356 13676 16362 13728
rect 16758 13676 16764 13728
rect 16816 13716 16822 13728
rect 17034 13716 17040 13728
rect 16816 13688 17040 13716
rect 16816 13676 16822 13688
rect 17034 13676 17040 13688
rect 17092 13676 17098 13728
rect 1104 13626 18860 13648
rect 1104 13574 3174 13626
rect 3226 13574 3238 13626
rect 3290 13574 3302 13626
rect 3354 13574 3366 13626
rect 3418 13574 3430 13626
rect 3482 13574 7622 13626
rect 7674 13574 7686 13626
rect 7738 13574 7750 13626
rect 7802 13574 7814 13626
rect 7866 13574 7878 13626
rect 7930 13574 12070 13626
rect 12122 13574 12134 13626
rect 12186 13574 12198 13626
rect 12250 13574 12262 13626
rect 12314 13574 12326 13626
rect 12378 13574 16518 13626
rect 16570 13574 16582 13626
rect 16634 13574 16646 13626
rect 16698 13574 16710 13626
rect 16762 13574 16774 13626
rect 16826 13574 18860 13626
rect 1104 13552 18860 13574
rect 2866 13472 2872 13524
rect 2924 13512 2930 13524
rect 3329 13515 3387 13521
rect 3329 13512 3341 13515
rect 2924 13484 3341 13512
rect 2924 13472 2930 13484
rect 3329 13481 3341 13484
rect 3375 13481 3387 13515
rect 3329 13475 3387 13481
rect 3510 13472 3516 13524
rect 3568 13512 3574 13524
rect 4893 13515 4951 13521
rect 4893 13512 4905 13515
rect 3568 13484 4905 13512
rect 3568 13472 3574 13484
rect 4893 13481 4905 13484
rect 4939 13481 4951 13515
rect 7190 13512 7196 13524
rect 4893 13475 4951 13481
rect 6196 13484 7196 13512
rect 2498 13404 2504 13456
rect 2556 13444 2562 13456
rect 3881 13447 3939 13453
rect 3881 13444 3893 13447
rect 2556 13416 3893 13444
rect 2556 13404 2562 13416
rect 3881 13413 3893 13416
rect 3927 13413 3939 13447
rect 3881 13407 3939 13413
rect 4154 13404 4160 13456
rect 4212 13444 4218 13456
rect 6196 13444 6224 13484
rect 7190 13472 7196 13484
rect 7248 13512 7254 13524
rect 7248 13484 12296 13512
rect 7248 13472 7254 13484
rect 4212 13416 6224 13444
rect 4212 13404 4218 13416
rect 6270 13404 6276 13456
rect 6328 13444 6334 13456
rect 6328 13416 8524 13444
rect 6328 13404 6334 13416
rect 1946 13376 1952 13388
rect 1907 13348 1952 13376
rect 1946 13336 1952 13348
rect 2004 13336 2010 13388
rect 5442 13376 5448 13388
rect 3068 13348 4384 13376
rect 2225 13311 2283 13317
rect 2225 13277 2237 13311
rect 2271 13308 2283 13311
rect 2774 13308 2780 13320
rect 2271 13280 2780 13308
rect 2271 13277 2283 13280
rect 2225 13271 2283 13277
rect 2774 13268 2780 13280
rect 2832 13268 2838 13320
rect 2866 13268 2872 13320
rect 2924 13308 2930 13320
rect 2924 13280 2969 13308
rect 2924 13268 2930 13280
rect 290 13200 296 13252
rect 348 13240 354 13252
rect 3068 13240 3096 13348
rect 3142 13268 3148 13320
rect 3200 13308 3206 13320
rect 3510 13308 3516 13320
rect 3200 13280 3245 13308
rect 3471 13280 3516 13308
rect 3200 13268 3206 13280
rect 3510 13268 3516 13280
rect 3568 13268 3574 13320
rect 4062 13308 4068 13320
rect 4023 13280 4068 13308
rect 4062 13268 4068 13280
rect 4120 13268 4126 13320
rect 348 13212 3096 13240
rect 3252 13212 4292 13240
rect 348 13200 354 13212
rect 1578 13132 1584 13184
rect 1636 13172 1642 13184
rect 3252 13172 3280 13212
rect 1636 13144 3280 13172
rect 1636 13132 1642 13144
rect 3418 13132 3424 13184
rect 3476 13172 3482 13184
rect 4154 13172 4160 13184
rect 3476 13144 4160 13172
rect 3476 13132 3482 13144
rect 4154 13132 4160 13144
rect 4212 13132 4218 13184
rect 4264 13181 4292 13212
rect 4249 13175 4307 13181
rect 4249 13141 4261 13175
rect 4295 13141 4307 13175
rect 4356 13172 4384 13348
rect 4724 13348 5448 13376
rect 4433 13311 4491 13317
rect 4433 13277 4445 13311
rect 4479 13308 4491 13311
rect 4724 13308 4752 13348
rect 5442 13336 5448 13348
rect 5500 13336 5506 13388
rect 5718 13376 5724 13388
rect 5679 13348 5724 13376
rect 5718 13336 5724 13348
rect 5776 13336 5782 13388
rect 5994 13336 6000 13388
rect 6052 13376 6058 13388
rect 6457 13379 6515 13385
rect 6457 13376 6469 13379
rect 6052 13348 6469 13376
rect 6052 13336 6058 13348
rect 6457 13345 6469 13348
rect 6503 13345 6515 13379
rect 6457 13339 6515 13345
rect 6549 13379 6607 13385
rect 6549 13345 6561 13379
rect 6595 13376 6607 13379
rect 7469 13379 7527 13385
rect 7469 13376 7481 13379
rect 6595 13348 7481 13376
rect 6595 13345 6607 13348
rect 6549 13339 6607 13345
rect 7469 13345 7481 13348
rect 7515 13376 7527 13379
rect 7742 13376 7748 13388
rect 7515 13348 7748 13376
rect 7515 13345 7527 13348
rect 7469 13339 7527 13345
rect 7742 13336 7748 13348
rect 7800 13336 7806 13388
rect 4479 13280 4752 13308
rect 4801 13311 4859 13317
rect 4479 13277 4491 13280
rect 4433 13271 4491 13277
rect 4801 13277 4813 13311
rect 4847 13308 4859 13311
rect 6638 13308 6644 13320
rect 4847 13280 6644 13308
rect 4847 13277 4859 13280
rect 4801 13271 4859 13277
rect 6638 13268 6644 13280
rect 6696 13268 6702 13320
rect 7190 13268 7196 13320
rect 7248 13308 7254 13320
rect 7285 13311 7343 13317
rect 7285 13308 7297 13311
rect 7248 13280 7297 13308
rect 7248 13268 7254 13280
rect 7285 13277 7297 13280
rect 7331 13277 7343 13311
rect 8496 13308 8524 13416
rect 9398 13336 9404 13388
rect 9456 13376 9462 13388
rect 9769 13379 9827 13385
rect 9769 13376 9781 13379
rect 9456 13348 9781 13376
rect 9456 13336 9462 13348
rect 9769 13345 9781 13348
rect 9815 13345 9827 13379
rect 9769 13339 9827 13345
rect 11609 13379 11667 13385
rect 11609 13345 11621 13379
rect 11655 13376 11667 13379
rect 11974 13376 11980 13388
rect 11655 13348 11980 13376
rect 11655 13345 11667 13348
rect 11609 13339 11667 13345
rect 11974 13336 11980 13348
rect 12032 13336 12038 13388
rect 12161 13311 12219 13317
rect 12161 13308 12173 13311
rect 8496 13280 12173 13308
rect 7285 13271 7343 13277
rect 12161 13277 12173 13280
rect 12207 13277 12219 13311
rect 12268 13308 12296 13484
rect 12342 13472 12348 13524
rect 12400 13512 12406 13524
rect 13814 13512 13820 13524
rect 12400 13484 13820 13512
rect 12400 13472 12406 13484
rect 13814 13472 13820 13484
rect 13872 13472 13878 13524
rect 16669 13515 16727 13521
rect 16669 13481 16681 13515
rect 16715 13512 16727 13515
rect 16850 13512 16856 13524
rect 16715 13484 16856 13512
rect 16715 13481 16727 13484
rect 16669 13475 16727 13481
rect 16850 13472 16856 13484
rect 16908 13472 16914 13524
rect 16301 13447 16359 13453
rect 16301 13413 16313 13447
rect 16347 13444 16359 13447
rect 17678 13444 17684 13456
rect 16347 13416 17684 13444
rect 16347 13413 16359 13416
rect 16301 13407 16359 13413
rect 17678 13404 17684 13416
rect 17736 13404 17742 13456
rect 12434 13336 12440 13388
rect 12492 13376 12498 13388
rect 16114 13376 16120 13388
rect 12492 13348 12537 13376
rect 13648 13348 16120 13376
rect 12492 13336 12498 13348
rect 12342 13308 12348 13320
rect 12255 13280 12348 13308
rect 12161 13271 12219 13277
rect 5537 13243 5595 13249
rect 5537 13209 5549 13243
rect 5583 13240 5595 13243
rect 5583 13212 6868 13240
rect 5583 13209 5595 13212
rect 5537 13203 5595 13209
rect 4617 13175 4675 13181
rect 4617 13172 4629 13175
rect 4356 13144 4629 13172
rect 4249 13135 4307 13141
rect 4617 13141 4629 13144
rect 4663 13141 4675 13175
rect 5166 13172 5172 13184
rect 5127 13144 5172 13172
rect 4617 13135 4675 13141
rect 5166 13132 5172 13144
rect 5224 13132 5230 13184
rect 5629 13175 5687 13181
rect 5629 13141 5641 13175
rect 5675 13172 5687 13175
rect 5997 13175 6055 13181
rect 5997 13172 6009 13175
rect 5675 13144 6009 13172
rect 5675 13141 5687 13144
rect 5629 13135 5687 13141
rect 5997 13141 6009 13144
rect 6043 13141 6055 13175
rect 5997 13135 6055 13141
rect 6270 13132 6276 13184
rect 6328 13172 6334 13184
rect 6840 13181 6868 13212
rect 6914 13200 6920 13252
rect 6972 13240 6978 13252
rect 9585 13243 9643 13249
rect 6972 13212 9352 13240
rect 6972 13200 6978 13212
rect 6365 13175 6423 13181
rect 6365 13172 6377 13175
rect 6328 13144 6377 13172
rect 6328 13132 6334 13144
rect 6365 13141 6377 13144
rect 6411 13141 6423 13175
rect 6365 13135 6423 13141
rect 6825 13175 6883 13181
rect 6825 13141 6837 13175
rect 6871 13141 6883 13175
rect 7190 13172 7196 13184
rect 7151 13144 7196 13172
rect 6825 13135 6883 13141
rect 7190 13132 7196 13144
rect 7248 13132 7254 13184
rect 8386 13132 8392 13184
rect 8444 13172 8450 13184
rect 9217 13175 9275 13181
rect 9217 13172 9229 13175
rect 8444 13144 9229 13172
rect 8444 13132 8450 13144
rect 9217 13141 9229 13144
rect 9263 13141 9275 13175
rect 9324 13172 9352 13212
rect 9585 13209 9597 13243
rect 9631 13240 9643 13243
rect 10045 13243 10103 13249
rect 10045 13240 10057 13243
rect 9631 13212 10057 13240
rect 9631 13209 9643 13212
rect 9585 13203 9643 13209
rect 10045 13209 10057 13212
rect 10091 13209 10103 13243
rect 12176 13240 12204 13271
rect 12342 13268 12348 13280
rect 12400 13308 12406 13320
rect 13648 13308 13676 13348
rect 16114 13336 16120 13348
rect 16172 13336 16178 13388
rect 16853 13379 16911 13385
rect 16853 13345 16865 13379
rect 16899 13376 16911 13379
rect 16942 13376 16948 13388
rect 16899 13348 16948 13376
rect 16899 13345 16911 13348
rect 16853 13339 16911 13345
rect 16942 13336 16948 13348
rect 17000 13336 17006 13388
rect 16485 13311 16543 13317
rect 12400 13280 13676 13308
rect 13740 13280 13952 13308
rect 12400 13268 12406 13280
rect 13740 13240 13768 13280
rect 12176 13212 13768 13240
rect 13924 13240 13952 13280
rect 16485 13277 16497 13311
rect 16531 13308 16543 13311
rect 17678 13308 17684 13320
rect 16531 13280 17684 13308
rect 16531 13277 16543 13280
rect 16485 13271 16543 13277
rect 17678 13268 17684 13280
rect 17736 13268 17742 13320
rect 17957 13311 18015 13317
rect 17957 13277 17969 13311
rect 18003 13308 18015 13311
rect 18046 13308 18052 13320
rect 18003 13280 18052 13308
rect 18003 13277 18015 13280
rect 17957 13271 18015 13277
rect 18046 13268 18052 13280
rect 18104 13268 18110 13320
rect 16574 13240 16580 13252
rect 13924 13212 16580 13240
rect 10045 13203 10103 13209
rect 16574 13200 16580 13212
rect 16632 13200 16638 13252
rect 17126 13240 17132 13252
rect 17087 13212 17132 13240
rect 17126 13200 17132 13212
rect 17184 13200 17190 13252
rect 17497 13243 17555 13249
rect 17497 13209 17509 13243
rect 17543 13240 17555 13243
rect 17586 13240 17592 13252
rect 17543 13212 17592 13240
rect 17543 13209 17555 13212
rect 17497 13203 17555 13209
rect 17586 13200 17592 13212
rect 17644 13200 17650 13252
rect 9674 13172 9680 13184
rect 9324 13144 9680 13172
rect 9217 13135 9275 13141
rect 9674 13132 9680 13144
rect 9732 13132 9738 13184
rect 10965 13175 11023 13181
rect 10965 13141 10977 13175
rect 11011 13172 11023 13175
rect 11146 13172 11152 13184
rect 11011 13144 11152 13172
rect 11011 13141 11023 13144
rect 10965 13135 11023 13141
rect 11146 13132 11152 13144
rect 11204 13132 11210 13184
rect 11330 13172 11336 13184
rect 11291 13144 11336 13172
rect 11330 13132 11336 13144
rect 11388 13132 11394 13184
rect 11425 13175 11483 13181
rect 11425 13141 11437 13175
rect 11471 13172 11483 13175
rect 11793 13175 11851 13181
rect 11793 13172 11805 13175
rect 11471 13144 11805 13172
rect 11471 13141 11483 13144
rect 11425 13135 11483 13141
rect 11793 13141 11805 13144
rect 11839 13141 11851 13175
rect 11793 13135 11851 13141
rect 11882 13132 11888 13184
rect 11940 13172 11946 13184
rect 12253 13175 12311 13181
rect 12253 13172 12265 13175
rect 11940 13144 12265 13172
rect 11940 13132 11946 13144
rect 12253 13141 12265 13144
rect 12299 13141 12311 13175
rect 12618 13172 12624 13184
rect 12579 13144 12624 13172
rect 12253 13135 12311 13141
rect 12618 13132 12624 13144
rect 12676 13132 12682 13184
rect 13814 13172 13820 13184
rect 13727 13144 13820 13172
rect 13814 13132 13820 13144
rect 13872 13172 13878 13184
rect 15194 13172 15200 13184
rect 13872 13144 15200 13172
rect 13872 13132 13878 13144
rect 15194 13132 15200 13144
rect 15252 13132 15258 13184
rect 17034 13172 17040 13184
rect 16995 13144 17040 13172
rect 17034 13132 17040 13144
rect 17092 13132 17098 13184
rect 17402 13172 17408 13184
rect 17363 13144 17408 13172
rect 17402 13132 17408 13144
rect 17460 13132 17466 13184
rect 1104 13082 18860 13104
rect 1104 13030 5398 13082
rect 5450 13030 5462 13082
rect 5514 13030 5526 13082
rect 5578 13030 5590 13082
rect 5642 13030 5654 13082
rect 5706 13030 9846 13082
rect 9898 13030 9910 13082
rect 9962 13030 9974 13082
rect 10026 13030 10038 13082
rect 10090 13030 10102 13082
rect 10154 13030 14294 13082
rect 14346 13030 14358 13082
rect 14410 13030 14422 13082
rect 14474 13030 14486 13082
rect 14538 13030 14550 13082
rect 14602 13030 18860 13082
rect 1104 13008 18860 13030
rect 2866 12928 2872 12980
rect 2924 12968 2930 12980
rect 3881 12971 3939 12977
rect 2924 12940 3832 12968
rect 2924 12928 2930 12940
rect 2958 12792 2964 12844
rect 3016 12832 3022 12844
rect 3145 12835 3203 12841
rect 3145 12832 3157 12835
rect 3016 12804 3157 12832
rect 3016 12792 3022 12804
rect 3145 12801 3157 12804
rect 3191 12801 3203 12835
rect 3418 12832 3424 12844
rect 3379 12804 3424 12832
rect 3145 12795 3203 12801
rect 3418 12792 3424 12804
rect 3476 12792 3482 12844
rect 3804 12832 3832 12940
rect 3881 12937 3893 12971
rect 3927 12968 3939 12971
rect 4709 12971 4767 12977
rect 4709 12968 4721 12971
rect 3927 12940 4721 12968
rect 3927 12937 3939 12940
rect 3881 12931 3939 12937
rect 4709 12937 4721 12940
rect 4755 12968 4767 12971
rect 4982 12968 4988 12980
rect 4755 12940 4988 12968
rect 4755 12937 4767 12940
rect 4709 12931 4767 12937
rect 4982 12928 4988 12940
rect 5040 12928 5046 12980
rect 5166 12968 5172 12980
rect 5127 12940 5172 12968
rect 5166 12928 5172 12940
rect 5224 12928 5230 12980
rect 6641 12971 6699 12977
rect 5276 12940 6592 12968
rect 5276 12900 5304 12940
rect 5000 12872 5304 12900
rect 4525 12835 4583 12841
rect 3804 12804 4476 12832
rect 1949 12767 2007 12773
rect 1949 12733 1961 12767
rect 1995 12764 2007 12767
rect 2130 12764 2136 12776
rect 1995 12736 2136 12764
rect 1995 12733 2007 12736
rect 1949 12727 2007 12733
rect 2130 12724 2136 12736
rect 2188 12724 2194 12776
rect 2222 12724 2228 12776
rect 2280 12764 2286 12776
rect 2774 12764 2780 12776
rect 2280 12736 2780 12764
rect 2280 12724 2286 12736
rect 2774 12724 2780 12736
rect 2832 12724 2838 12776
rect 2869 12767 2927 12773
rect 2869 12733 2881 12767
rect 2915 12733 2927 12767
rect 2869 12727 2927 12733
rect 2884 12696 2912 12727
rect 3510 12724 3516 12776
rect 3568 12764 3574 12776
rect 3973 12767 4031 12773
rect 3973 12764 3985 12767
rect 3568 12736 3985 12764
rect 3568 12724 3574 12736
rect 3973 12733 3985 12736
rect 4019 12733 4031 12767
rect 3973 12727 4031 12733
rect 4062 12724 4068 12776
rect 4120 12764 4126 12776
rect 4448 12764 4476 12804
rect 4525 12801 4537 12835
rect 4571 12832 4583 12835
rect 5000 12832 5028 12872
rect 5350 12860 5356 12912
rect 5408 12900 5414 12912
rect 5629 12903 5687 12909
rect 5629 12900 5641 12903
rect 5408 12872 5641 12900
rect 5408 12860 5414 12872
rect 5629 12869 5641 12872
rect 5675 12869 5687 12903
rect 6564 12900 6592 12940
rect 6641 12937 6653 12971
rect 6687 12968 6699 12971
rect 7190 12968 7196 12980
rect 6687 12940 7196 12968
rect 6687 12937 6699 12940
rect 6641 12931 6699 12937
rect 7190 12928 7196 12940
rect 7248 12928 7254 12980
rect 9217 12971 9275 12977
rect 9217 12937 9229 12971
rect 9263 12968 9275 12971
rect 9585 12971 9643 12977
rect 9585 12968 9597 12971
rect 9263 12940 9597 12968
rect 9263 12937 9275 12940
rect 9217 12931 9275 12937
rect 9585 12937 9597 12940
rect 9631 12937 9643 12971
rect 9585 12931 9643 12937
rect 11330 12928 11336 12980
rect 11388 12968 11394 12980
rect 11609 12971 11667 12977
rect 11609 12968 11621 12971
rect 11388 12940 11621 12968
rect 11388 12928 11394 12940
rect 11609 12937 11621 12940
rect 11655 12937 11667 12971
rect 11609 12931 11667 12937
rect 11977 12971 12035 12977
rect 11977 12937 11989 12971
rect 12023 12968 12035 12971
rect 12618 12968 12624 12980
rect 12023 12940 12624 12968
rect 12023 12937 12035 12940
rect 11977 12931 12035 12937
rect 12618 12928 12624 12940
rect 12676 12928 12682 12980
rect 13541 12971 13599 12977
rect 13541 12937 13553 12971
rect 13587 12968 13599 12971
rect 13909 12971 13967 12977
rect 13909 12968 13921 12971
rect 13587 12940 13921 12968
rect 13587 12937 13599 12940
rect 13541 12931 13599 12937
rect 13909 12937 13921 12940
rect 13955 12937 13967 12971
rect 13909 12931 13967 12937
rect 16853 12971 16911 12977
rect 16853 12937 16865 12971
rect 16899 12968 16911 12971
rect 17770 12968 17776 12980
rect 16899 12940 17776 12968
rect 16899 12937 16911 12940
rect 16853 12931 16911 12937
rect 17770 12928 17776 12940
rect 17828 12928 17834 12980
rect 6914 12900 6920 12912
rect 6564 12872 6920 12900
rect 5629 12863 5687 12869
rect 6914 12860 6920 12872
rect 6972 12860 6978 12912
rect 7006 12860 7012 12912
rect 7064 12900 7070 12912
rect 9953 12903 10011 12909
rect 9953 12900 9965 12903
rect 7064 12872 9965 12900
rect 7064 12860 7070 12872
rect 9953 12869 9965 12872
rect 9999 12900 10011 12903
rect 10413 12903 10471 12909
rect 10413 12900 10425 12903
rect 9999 12872 10425 12900
rect 9999 12869 10011 12872
rect 9953 12863 10011 12869
rect 10413 12869 10425 12872
rect 10459 12900 10471 12903
rect 16942 12900 16948 12912
rect 10459 12872 14320 12900
rect 16903 12872 16948 12900
rect 10459 12869 10471 12872
rect 10413 12863 10471 12869
rect 6270 12832 6276 12844
rect 4571 12804 5028 12832
rect 5092 12804 6276 12832
rect 4571 12801 4583 12804
rect 4525 12795 4583 12801
rect 5092 12764 5120 12804
rect 6270 12792 6276 12804
rect 6328 12792 6334 12844
rect 9122 12832 9128 12844
rect 9083 12804 9128 12832
rect 9122 12792 9128 12804
rect 9180 12792 9186 12844
rect 10045 12835 10103 12841
rect 10045 12801 10057 12835
rect 10091 12832 10103 12835
rect 12069 12835 12127 12841
rect 10091 12804 10364 12832
rect 10091 12801 10103 12804
rect 10045 12795 10103 12801
rect 5258 12764 5264 12776
rect 4120 12736 4165 12764
rect 4448 12736 5120 12764
rect 5219 12736 5264 12764
rect 4120 12724 4126 12736
rect 5258 12724 5264 12736
rect 5316 12724 5322 12776
rect 5353 12767 5411 12773
rect 5353 12733 5365 12767
rect 5399 12733 5411 12767
rect 5353 12727 5411 12733
rect 3878 12696 3884 12708
rect 2884 12668 3884 12696
rect 3878 12656 3884 12668
rect 3936 12656 3942 12708
rect 3988 12668 4936 12696
rect 3050 12588 3056 12640
rect 3108 12628 3114 12640
rect 3237 12631 3295 12637
rect 3237 12628 3249 12631
rect 3108 12600 3249 12628
rect 3108 12588 3114 12600
rect 3237 12597 3249 12600
rect 3283 12597 3295 12631
rect 3510 12628 3516 12640
rect 3471 12600 3516 12628
rect 3237 12591 3295 12597
rect 3510 12588 3516 12600
rect 3568 12588 3574 12640
rect 3786 12588 3792 12640
rect 3844 12628 3850 12640
rect 3988 12628 4016 12668
rect 3844 12600 4016 12628
rect 3844 12588 3850 12600
rect 4154 12588 4160 12640
rect 4212 12628 4218 12640
rect 4341 12631 4399 12637
rect 4341 12628 4353 12631
rect 4212 12600 4353 12628
rect 4212 12588 4218 12600
rect 4341 12597 4353 12600
rect 4387 12597 4399 12631
rect 4341 12591 4399 12597
rect 4706 12588 4712 12640
rect 4764 12628 4770 12640
rect 4801 12631 4859 12637
rect 4801 12628 4813 12631
rect 4764 12600 4813 12628
rect 4764 12588 4770 12600
rect 4801 12597 4813 12600
rect 4847 12597 4859 12631
rect 4908 12628 4936 12668
rect 5166 12656 5172 12708
rect 5224 12696 5230 12708
rect 5368 12696 5396 12727
rect 7374 12724 7380 12776
rect 7432 12764 7438 12776
rect 7742 12764 7748 12776
rect 7432 12736 7748 12764
rect 7432 12724 7438 12736
rect 7742 12724 7748 12736
rect 7800 12764 7806 12776
rect 9309 12767 9367 12773
rect 9309 12764 9321 12767
rect 7800 12736 9321 12764
rect 7800 12724 7806 12736
rect 9309 12733 9321 12736
rect 9355 12733 9367 12767
rect 9309 12727 9367 12733
rect 5224 12668 5396 12696
rect 5224 12656 5230 12668
rect 6730 12656 6736 12708
rect 6788 12696 6794 12708
rect 6825 12699 6883 12705
rect 6825 12696 6837 12699
rect 6788 12668 6837 12696
rect 6788 12656 6794 12668
rect 6825 12665 6837 12668
rect 6871 12696 6883 12699
rect 8665 12699 8723 12705
rect 8665 12696 8677 12699
rect 6871 12668 8677 12696
rect 6871 12665 6883 12668
rect 6825 12659 6883 12665
rect 8665 12665 8677 12668
rect 8711 12696 8723 12699
rect 10060 12696 10088 12795
rect 10226 12764 10232 12776
rect 10187 12736 10232 12764
rect 10226 12724 10232 12736
rect 10284 12724 10290 12776
rect 10336 12764 10364 12804
rect 12069 12801 12081 12835
rect 12115 12832 12127 12835
rect 12342 12832 12348 12844
rect 12115 12804 12348 12832
rect 12115 12801 12127 12804
rect 12069 12795 12127 12801
rect 12342 12792 12348 12804
rect 12400 12792 12406 12844
rect 12986 12792 12992 12844
rect 13044 12832 13050 12844
rect 14292 12841 14320 12872
rect 16942 12860 16948 12872
rect 17000 12860 17006 12912
rect 17126 12860 17132 12912
rect 17184 12900 17190 12912
rect 17313 12903 17371 12909
rect 17313 12900 17325 12903
rect 17184 12872 17325 12900
rect 17184 12860 17190 12872
rect 17313 12869 17325 12872
rect 17359 12869 17371 12903
rect 17586 12900 17592 12912
rect 17547 12872 17592 12900
rect 17313 12863 17371 12869
rect 17586 12860 17592 12872
rect 17644 12860 17650 12912
rect 13449 12835 13507 12841
rect 13449 12832 13461 12835
rect 13044 12804 13461 12832
rect 13044 12792 13050 12804
rect 13449 12801 13461 12804
rect 13495 12801 13507 12835
rect 13449 12795 13507 12801
rect 14277 12835 14335 12841
rect 14277 12801 14289 12835
rect 14323 12801 14335 12835
rect 14277 12795 14335 12801
rect 14369 12835 14427 12841
rect 14369 12801 14381 12835
rect 14415 12832 14427 12835
rect 15194 12832 15200 12844
rect 14415 12804 15200 12832
rect 14415 12801 14427 12804
rect 14369 12795 14427 12801
rect 12158 12764 12164 12776
rect 10336 12736 12164 12764
rect 12158 12724 12164 12736
rect 12216 12724 12222 12776
rect 12253 12767 12311 12773
rect 12253 12733 12265 12767
rect 12299 12764 12311 12767
rect 12434 12764 12440 12776
rect 12299 12736 12440 12764
rect 12299 12733 12311 12736
rect 12253 12727 12311 12733
rect 12434 12724 12440 12736
rect 12492 12764 12498 12776
rect 13354 12764 13360 12776
rect 12492 12736 13360 12764
rect 12492 12724 12498 12736
rect 13354 12724 13360 12736
rect 13412 12764 13418 12776
rect 13633 12767 13691 12773
rect 13633 12764 13645 12767
rect 13412 12736 13645 12764
rect 13412 12724 13418 12736
rect 13633 12733 13645 12736
rect 13679 12733 13691 12767
rect 13633 12727 13691 12733
rect 8711 12668 10088 12696
rect 12713 12699 12771 12705
rect 8711 12665 8723 12668
rect 8665 12659 8723 12665
rect 12713 12665 12725 12699
rect 12759 12696 12771 12699
rect 13170 12696 13176 12708
rect 12759 12668 13176 12696
rect 12759 12665 12771 12668
rect 12713 12659 12771 12665
rect 13170 12656 13176 12668
rect 13228 12656 13234 12708
rect 5813 12631 5871 12637
rect 5813 12628 5825 12631
rect 4908 12600 5825 12628
rect 4801 12591 4859 12597
rect 5813 12597 5825 12600
rect 5859 12597 5871 12631
rect 5813 12591 5871 12597
rect 6638 12588 6644 12640
rect 6696 12628 6702 12640
rect 8757 12631 8815 12637
rect 8757 12628 8769 12631
rect 6696 12600 8769 12628
rect 6696 12588 6702 12600
rect 8757 12597 8769 12600
rect 8803 12597 8815 12631
rect 8757 12591 8815 12597
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 13081 12631 13139 12637
rect 13081 12628 13093 12631
rect 12492 12600 13093 12628
rect 12492 12588 12498 12600
rect 13081 12597 13093 12600
rect 13127 12597 13139 12631
rect 14292 12628 14320 12795
rect 15194 12792 15200 12804
rect 15252 12832 15258 12844
rect 16206 12832 16212 12844
rect 15252 12804 16212 12832
rect 15252 12792 15258 12804
rect 16206 12792 16212 12804
rect 16264 12792 16270 12844
rect 16574 12792 16580 12844
rect 16632 12832 16638 12844
rect 17494 12832 17500 12844
rect 16632 12804 17500 12832
rect 16632 12792 16638 12804
rect 17494 12792 17500 12804
rect 17552 12792 17558 12844
rect 14458 12724 14464 12776
rect 14516 12764 14522 12776
rect 17221 12767 17279 12773
rect 14516 12736 14561 12764
rect 14516 12724 14522 12736
rect 17221 12733 17233 12767
rect 17267 12764 17279 12767
rect 17681 12767 17739 12773
rect 17681 12764 17693 12767
rect 17267 12736 17693 12764
rect 17267 12733 17279 12736
rect 17221 12727 17279 12733
rect 17681 12733 17693 12736
rect 17727 12764 17739 12767
rect 17770 12764 17776 12776
rect 17727 12736 17776 12764
rect 17727 12733 17739 12736
rect 17681 12727 17739 12733
rect 17770 12724 17776 12736
rect 17828 12724 17834 12776
rect 17957 12767 18015 12773
rect 17957 12733 17969 12767
rect 18003 12764 18015 12767
rect 18230 12764 18236 12776
rect 18003 12736 18236 12764
rect 18003 12733 18015 12736
rect 17957 12727 18015 12733
rect 18230 12724 18236 12736
rect 18288 12724 18294 12776
rect 15838 12656 15844 12708
rect 15896 12696 15902 12708
rect 19610 12696 19616 12708
rect 15896 12668 19616 12696
rect 15896 12656 15902 12668
rect 19610 12656 19616 12668
rect 19668 12656 19674 12708
rect 14829 12631 14887 12637
rect 14829 12628 14841 12631
rect 14292 12600 14841 12628
rect 13081 12591 13139 12597
rect 14829 12597 14841 12600
rect 14875 12628 14887 12631
rect 16850 12628 16856 12640
rect 14875 12600 16856 12628
rect 14875 12597 14887 12600
rect 14829 12591 14887 12597
rect 16850 12588 16856 12600
rect 16908 12588 16914 12640
rect 1104 12538 18860 12560
rect 1104 12486 3174 12538
rect 3226 12486 3238 12538
rect 3290 12486 3302 12538
rect 3354 12486 3366 12538
rect 3418 12486 3430 12538
rect 3482 12486 7622 12538
rect 7674 12486 7686 12538
rect 7738 12486 7750 12538
rect 7802 12486 7814 12538
rect 7866 12486 7878 12538
rect 7930 12486 12070 12538
rect 12122 12486 12134 12538
rect 12186 12486 12198 12538
rect 12250 12486 12262 12538
rect 12314 12486 12326 12538
rect 12378 12486 16518 12538
rect 16570 12486 16582 12538
rect 16634 12486 16646 12538
rect 16698 12486 16710 12538
rect 16762 12486 16774 12538
rect 16826 12486 18860 12538
rect 1104 12464 18860 12486
rect 2958 12384 2964 12436
rect 3016 12424 3022 12436
rect 4065 12427 4123 12433
rect 4065 12424 4077 12427
rect 3016 12396 4077 12424
rect 3016 12384 3022 12396
rect 4065 12393 4077 12396
rect 4111 12393 4123 12427
rect 4065 12387 4123 12393
rect 7190 12384 7196 12436
rect 7248 12424 7254 12436
rect 7466 12424 7472 12436
rect 7248 12396 7472 12424
rect 7248 12384 7254 12396
rect 7466 12384 7472 12396
rect 7524 12384 7530 12436
rect 9122 12384 9128 12436
rect 9180 12424 9186 12436
rect 9677 12427 9735 12433
rect 9677 12424 9689 12427
rect 9180 12396 9689 12424
rect 9180 12384 9186 12396
rect 9677 12393 9689 12396
rect 9723 12393 9735 12427
rect 12802 12424 12808 12436
rect 12763 12396 12808 12424
rect 9677 12387 9735 12393
rect 12802 12384 12808 12396
rect 12860 12384 12866 12436
rect 12986 12384 12992 12436
rect 13044 12424 13050 12436
rect 14093 12427 14151 12433
rect 14093 12424 14105 12427
rect 13044 12396 14105 12424
rect 13044 12384 13050 12396
rect 14093 12393 14105 12396
rect 14139 12393 14151 12427
rect 14093 12387 14151 12393
rect 17954 12384 17960 12436
rect 18012 12424 18018 12436
rect 18138 12424 18144 12436
rect 18012 12396 18144 12424
rect 18012 12384 18018 12396
rect 18138 12384 18144 12396
rect 18196 12384 18202 12436
rect 5902 12356 5908 12368
rect 1964 12328 5908 12356
rect 1964 12297 1992 12328
rect 5902 12316 5908 12328
rect 5960 12316 5966 12368
rect 10410 12316 10416 12368
rect 10468 12356 10474 12368
rect 10873 12359 10931 12365
rect 10873 12356 10885 12359
rect 10468 12328 10885 12356
rect 10468 12316 10474 12328
rect 10873 12325 10885 12328
rect 10919 12325 10931 12359
rect 13817 12359 13875 12365
rect 13817 12356 13829 12359
rect 10873 12319 10931 12325
rect 11139 12328 13829 12356
rect 1949 12291 2007 12297
rect 1949 12257 1961 12291
rect 1995 12257 2007 12291
rect 1949 12251 2007 12257
rect 3053 12291 3111 12297
rect 3053 12257 3065 12291
rect 3099 12288 3111 12291
rect 4062 12288 4068 12300
rect 3099 12260 4068 12288
rect 3099 12257 3111 12260
rect 3053 12251 3111 12257
rect 4062 12248 4068 12260
rect 4120 12288 4126 12300
rect 4985 12291 5043 12297
rect 4985 12288 4997 12291
rect 4120 12260 4997 12288
rect 4120 12248 4126 12260
rect 4985 12257 4997 12260
rect 5031 12288 5043 12291
rect 6546 12288 6552 12300
rect 5031 12260 6552 12288
rect 5031 12257 5043 12260
rect 4985 12251 5043 12257
rect 6546 12248 6552 12260
rect 6604 12288 6610 12300
rect 6641 12291 6699 12297
rect 6641 12288 6653 12291
rect 6604 12260 6653 12288
rect 6604 12248 6610 12260
rect 6641 12257 6653 12260
rect 6687 12257 6699 12291
rect 6641 12251 6699 12257
rect 7469 12291 7527 12297
rect 7469 12257 7481 12291
rect 7515 12288 7527 12291
rect 8297 12291 8355 12297
rect 8297 12288 8309 12291
rect 7515 12260 8309 12288
rect 7515 12257 7527 12260
rect 7469 12251 7527 12257
rect 8297 12257 8309 12260
rect 8343 12257 8355 12291
rect 10226 12288 10232 12300
rect 10187 12260 10232 12288
rect 8297 12251 8355 12257
rect 2225 12223 2283 12229
rect 2225 12189 2237 12223
rect 2271 12220 2283 12223
rect 2774 12220 2780 12232
rect 2271 12192 2780 12220
rect 2271 12189 2283 12192
rect 2225 12183 2283 12189
rect 2774 12180 2780 12192
rect 2832 12220 2838 12232
rect 5261 12223 5319 12229
rect 5261 12220 5273 12223
rect 2832 12192 5273 12220
rect 2832 12180 2838 12192
rect 5261 12189 5273 12192
rect 5307 12189 5319 12223
rect 5261 12183 5319 12189
rect 7098 12180 7104 12232
rect 7156 12220 7162 12232
rect 7285 12223 7343 12229
rect 7285 12220 7297 12223
rect 7156 12192 7297 12220
rect 7156 12180 7162 12192
rect 7285 12189 7297 12192
rect 7331 12189 7343 12223
rect 7285 12183 7343 12189
rect 7374 12180 7380 12232
rect 7432 12220 7438 12232
rect 7484 12220 7512 12251
rect 10226 12248 10232 12260
rect 10284 12248 10290 12300
rect 7432 12192 7512 12220
rect 7432 12180 7438 12192
rect 2406 12152 2412 12164
rect 2367 12124 2412 12152
rect 2406 12112 2412 12124
rect 2464 12152 2470 12164
rect 2685 12155 2743 12161
rect 2685 12152 2697 12155
rect 2464 12124 2697 12152
rect 2464 12112 2470 12124
rect 2685 12121 2697 12124
rect 2731 12121 2743 12155
rect 3142 12152 3148 12164
rect 3103 12124 3148 12152
rect 2685 12115 2743 12121
rect 3142 12112 3148 12124
rect 3200 12112 3206 12164
rect 3237 12155 3295 12161
rect 3237 12121 3249 12155
rect 3283 12152 3295 12155
rect 3789 12155 3847 12161
rect 3789 12152 3801 12155
rect 3283 12124 3801 12152
rect 3283 12121 3295 12124
rect 3237 12115 3295 12121
rect 3789 12121 3801 12124
rect 3835 12121 3847 12155
rect 3789 12115 3847 12121
rect 3878 12112 3884 12164
rect 3936 12152 3942 12164
rect 4249 12155 4307 12161
rect 4249 12152 4261 12155
rect 3936 12124 4261 12152
rect 3936 12112 3942 12124
rect 4249 12121 4261 12124
rect 4295 12152 4307 12155
rect 4801 12155 4859 12161
rect 4801 12152 4813 12155
rect 4295 12124 4813 12152
rect 4295 12121 4307 12124
rect 4249 12115 4307 12121
rect 4801 12121 4813 12124
rect 4847 12152 4859 12155
rect 4982 12152 4988 12164
rect 4847 12124 4988 12152
rect 4847 12121 4859 12124
rect 4801 12115 4859 12121
rect 4982 12112 4988 12124
rect 5040 12112 5046 12164
rect 6457 12155 6515 12161
rect 6457 12121 6469 12155
rect 6503 12152 6515 12155
rect 6503 12124 7788 12152
rect 6503 12121 6515 12124
rect 6457 12115 6515 12121
rect 2498 12084 2504 12096
rect 2459 12056 2504 12084
rect 2498 12044 2504 12056
rect 2556 12044 2562 12096
rect 3326 12044 3332 12096
rect 3384 12084 3390 12096
rect 3605 12087 3663 12093
rect 3605 12084 3617 12087
rect 3384 12056 3617 12084
rect 3384 12044 3390 12056
rect 3605 12053 3617 12056
rect 3651 12053 3663 12087
rect 3605 12047 3663 12053
rect 4338 12044 4344 12096
rect 4396 12084 4402 12096
rect 4433 12087 4491 12093
rect 4433 12084 4445 12087
rect 4396 12056 4445 12084
rect 4396 12044 4402 12056
rect 4433 12053 4445 12056
rect 4479 12053 4491 12087
rect 4433 12047 4491 12053
rect 4890 12044 4896 12096
rect 4948 12084 4954 12096
rect 6086 12084 6092 12096
rect 4948 12056 4993 12084
rect 6047 12056 6092 12084
rect 4948 12044 4954 12056
rect 6086 12044 6092 12056
rect 6144 12044 6150 12096
rect 6549 12087 6607 12093
rect 6549 12053 6561 12087
rect 6595 12084 6607 12087
rect 6917 12087 6975 12093
rect 6917 12084 6929 12087
rect 6595 12056 6929 12084
rect 6595 12053 6607 12056
rect 6549 12047 6607 12053
rect 6917 12053 6929 12056
rect 6963 12053 6975 12087
rect 6917 12047 6975 12053
rect 7006 12044 7012 12096
rect 7064 12084 7070 12096
rect 7760 12093 7788 12124
rect 7926 12112 7932 12164
rect 7984 12152 7990 12164
rect 8205 12155 8263 12161
rect 8205 12152 8217 12155
rect 7984 12124 8217 12152
rect 7984 12112 7990 12124
rect 8205 12121 8217 12124
rect 8251 12152 8263 12155
rect 9493 12155 9551 12161
rect 9493 12152 9505 12155
rect 8251 12124 9505 12152
rect 8251 12121 8263 12124
rect 8205 12115 8263 12121
rect 9493 12121 9505 12124
rect 9539 12152 9551 12155
rect 10137 12155 10195 12161
rect 10137 12152 10149 12155
rect 9539 12124 10149 12152
rect 9539 12121 9551 12124
rect 9493 12115 9551 12121
rect 10137 12121 10149 12124
rect 10183 12152 10195 12155
rect 11139 12152 11167 12328
rect 13817 12325 13829 12328
rect 13863 12356 13875 12359
rect 16577 12359 16635 12365
rect 16577 12356 16589 12359
rect 13863 12328 16589 12356
rect 13863 12325 13875 12328
rect 13817 12319 13875 12325
rect 11330 12248 11336 12300
rect 11388 12288 11394 12300
rect 11425 12291 11483 12297
rect 11425 12288 11437 12291
rect 11388 12260 11437 12288
rect 11388 12248 11394 12260
rect 11425 12257 11437 12260
rect 11471 12257 11483 12291
rect 11425 12251 11483 12257
rect 12342 12248 12348 12300
rect 12400 12248 12406 12300
rect 12434 12248 12440 12300
rect 12492 12288 12498 12300
rect 12621 12291 12679 12297
rect 12492 12260 12537 12288
rect 12492 12248 12498 12260
rect 12621 12257 12633 12291
rect 12667 12257 12679 12291
rect 13354 12288 13360 12300
rect 13315 12260 13360 12288
rect 12621 12251 12679 12257
rect 11238 12220 11244 12232
rect 11199 12192 11244 12220
rect 11238 12180 11244 12192
rect 11296 12180 11302 12232
rect 12360 12220 12388 12248
rect 12636 12220 12664 12251
rect 13354 12248 13360 12260
rect 13412 12248 13418 12300
rect 14568 12297 14596 12328
rect 16577 12325 16589 12328
rect 16623 12356 16635 12359
rect 17218 12356 17224 12368
rect 16623 12328 17224 12356
rect 16623 12325 16635 12328
rect 16577 12319 16635 12325
rect 17218 12316 17224 12328
rect 17276 12316 17282 12368
rect 17589 12359 17647 12365
rect 17589 12325 17601 12359
rect 17635 12356 17647 12359
rect 18690 12356 18696 12368
rect 17635 12328 18696 12356
rect 17635 12325 17647 12328
rect 17589 12319 17647 12325
rect 18690 12316 18696 12328
rect 18748 12316 18754 12368
rect 14553 12291 14611 12297
rect 14553 12257 14565 12291
rect 14599 12257 14611 12291
rect 14553 12251 14611 12257
rect 14642 12248 14648 12300
rect 14700 12288 14706 12300
rect 16945 12291 17003 12297
rect 14700 12260 14745 12288
rect 14700 12248 14706 12260
rect 16945 12257 16957 12291
rect 16991 12288 17003 12291
rect 16991 12260 17724 12288
rect 16991 12257 17003 12260
rect 16945 12251 17003 12257
rect 12360 12192 12664 12220
rect 15194 12180 15200 12232
rect 15252 12220 15258 12232
rect 17696 12229 17724 12260
rect 17405 12223 17463 12229
rect 17405 12220 17417 12223
rect 15252 12192 17417 12220
rect 15252 12180 15258 12192
rect 17405 12189 17417 12192
rect 17451 12189 17463 12223
rect 17405 12183 17463 12189
rect 17681 12223 17739 12229
rect 17681 12189 17693 12223
rect 17727 12220 17739 12223
rect 17862 12220 17868 12232
rect 17727 12192 17868 12220
rect 17727 12189 17739 12192
rect 17681 12183 17739 12189
rect 17862 12180 17868 12192
rect 17920 12180 17926 12232
rect 17954 12180 17960 12232
rect 18012 12220 18018 12232
rect 18012 12192 18057 12220
rect 18012 12180 18018 12192
rect 12345 12155 12403 12161
rect 10183 12124 11167 12152
rect 11256 12124 12112 12152
rect 10183 12121 10195 12124
rect 10137 12115 10195 12121
rect 7377 12087 7435 12093
rect 7377 12084 7389 12087
rect 7064 12056 7389 12084
rect 7064 12044 7070 12056
rect 7377 12053 7389 12056
rect 7423 12053 7435 12087
rect 7377 12047 7435 12053
rect 7745 12087 7803 12093
rect 7745 12053 7757 12087
rect 7791 12053 7803 12087
rect 8110 12084 8116 12096
rect 8071 12056 8116 12084
rect 7745 12047 7803 12053
rect 8110 12044 8116 12056
rect 8168 12084 8174 12096
rect 8573 12087 8631 12093
rect 8573 12084 8585 12087
rect 8168 12056 8585 12084
rect 8168 12044 8174 12056
rect 8573 12053 8585 12056
rect 8619 12084 8631 12087
rect 10045 12087 10103 12093
rect 10045 12084 10057 12087
rect 8619 12056 10057 12084
rect 8619 12053 8631 12056
rect 8573 12047 8631 12053
rect 10045 12053 10057 12056
rect 10091 12084 10103 12087
rect 10505 12087 10563 12093
rect 10505 12084 10517 12087
rect 10091 12056 10517 12084
rect 10091 12053 10103 12056
rect 10045 12047 10103 12053
rect 10505 12053 10517 12056
rect 10551 12084 10563 12087
rect 11256 12084 11284 12124
rect 10551 12056 11284 12084
rect 11333 12087 11391 12093
rect 10551 12053 10563 12056
rect 10505 12047 10563 12053
rect 11333 12053 11345 12087
rect 11379 12084 11391 12087
rect 11977 12087 12035 12093
rect 11977 12084 11989 12087
rect 11379 12056 11989 12084
rect 11379 12053 11391 12056
rect 11333 12047 11391 12053
rect 11977 12053 11989 12056
rect 12023 12053 12035 12087
rect 12084 12084 12112 12124
rect 12345 12121 12357 12155
rect 12391 12152 12403 12155
rect 12802 12152 12808 12164
rect 12391 12124 12808 12152
rect 12391 12121 12403 12124
rect 12345 12115 12403 12121
rect 12802 12112 12808 12124
rect 12860 12112 12866 12164
rect 15013 12155 15071 12161
rect 15013 12152 15025 12155
rect 13004 12124 15025 12152
rect 13004 12084 13032 12124
rect 13170 12084 13176 12096
rect 12084 12056 13032 12084
rect 13131 12056 13176 12084
rect 11977 12047 12035 12053
rect 13170 12044 13176 12056
rect 13228 12044 13234 12096
rect 13262 12044 13268 12096
rect 13320 12084 13326 12096
rect 14476 12093 14504 12124
rect 15013 12121 15025 12124
rect 15059 12152 15071 12155
rect 17129 12155 17187 12161
rect 15059 12124 16528 12152
rect 15059 12121 15071 12124
rect 15013 12115 15071 12121
rect 14461 12087 14519 12093
rect 13320 12056 13365 12084
rect 13320 12044 13326 12056
rect 14461 12053 14473 12087
rect 14507 12053 14519 12087
rect 14461 12047 14519 12053
rect 15289 12087 15347 12093
rect 15289 12053 15301 12087
rect 15335 12084 15347 12087
rect 15930 12084 15936 12096
rect 15335 12056 15936 12084
rect 15335 12053 15347 12056
rect 15289 12047 15347 12053
rect 15930 12044 15936 12056
rect 15988 12044 15994 12096
rect 16022 12044 16028 12096
rect 16080 12084 16086 12096
rect 16393 12087 16451 12093
rect 16393 12084 16405 12087
rect 16080 12056 16405 12084
rect 16080 12044 16086 12056
rect 16393 12053 16405 12056
rect 16439 12053 16451 12087
rect 16500 12084 16528 12124
rect 17129 12121 17141 12155
rect 17175 12152 17187 12155
rect 17175 12124 17724 12152
rect 17175 12121 17187 12124
rect 17129 12115 17187 12121
rect 17696 12096 17724 12124
rect 17313 12087 17371 12093
rect 17313 12084 17325 12087
rect 16500 12056 17325 12084
rect 16393 12047 16451 12053
rect 17313 12053 17325 12056
rect 17359 12084 17371 12087
rect 17586 12084 17592 12096
rect 17359 12056 17592 12084
rect 17359 12053 17371 12056
rect 17313 12047 17371 12053
rect 17586 12044 17592 12056
rect 17644 12044 17650 12096
rect 17678 12044 17684 12096
rect 17736 12044 17742 12096
rect 1104 11994 18860 12016
rect 1104 11942 5398 11994
rect 5450 11942 5462 11994
rect 5514 11942 5526 11994
rect 5578 11942 5590 11994
rect 5642 11942 5654 11994
rect 5706 11942 9846 11994
rect 9898 11942 9910 11994
rect 9962 11942 9974 11994
rect 10026 11942 10038 11994
rect 10090 11942 10102 11994
rect 10154 11942 14294 11994
rect 14346 11942 14358 11994
rect 14410 11942 14422 11994
rect 14474 11942 14486 11994
rect 14538 11942 14550 11994
rect 14602 11942 18860 11994
rect 1104 11920 18860 11942
rect 2406 11840 2412 11892
rect 2464 11880 2470 11892
rect 3326 11880 3332 11892
rect 2464 11852 3188 11880
rect 3287 11852 3332 11880
rect 2464 11840 2470 11852
rect 3050 11812 3056 11824
rect 2516 11784 3056 11812
rect 2516 11753 2544 11784
rect 3050 11772 3056 11784
rect 3108 11772 3114 11824
rect 3160 11812 3188 11852
rect 3326 11840 3332 11852
rect 3384 11840 3390 11892
rect 3421 11883 3479 11889
rect 3421 11849 3433 11883
rect 3467 11880 3479 11883
rect 3510 11880 3516 11892
rect 3467 11852 3516 11880
rect 3467 11849 3479 11852
rect 3421 11843 3479 11849
rect 3510 11840 3516 11852
rect 3568 11840 3574 11892
rect 4338 11880 4344 11892
rect 4299 11852 4344 11880
rect 4338 11840 4344 11852
rect 4396 11840 4402 11892
rect 4890 11840 4896 11892
rect 4948 11880 4954 11892
rect 5445 11883 5503 11889
rect 5445 11880 5457 11883
rect 4948 11852 5457 11880
rect 4948 11840 4954 11852
rect 5445 11849 5457 11852
rect 5491 11849 5503 11883
rect 5902 11880 5908 11892
rect 5863 11852 5908 11880
rect 5445 11843 5503 11849
rect 5902 11840 5908 11852
rect 5960 11880 5966 11892
rect 8297 11883 8355 11889
rect 5960 11852 7696 11880
rect 5960 11840 5966 11852
rect 4154 11812 4160 11824
rect 3160 11784 4160 11812
rect 4154 11772 4160 11784
rect 4212 11772 4218 11824
rect 4433 11815 4491 11821
rect 4433 11781 4445 11815
rect 4479 11812 4491 11815
rect 6086 11812 6092 11824
rect 4479 11784 6092 11812
rect 4479 11781 4491 11784
rect 4433 11775 4491 11781
rect 6086 11772 6092 11784
rect 6144 11772 6150 11824
rect 6454 11812 6460 11824
rect 6415 11784 6460 11812
rect 6454 11772 6460 11784
rect 6512 11772 6518 11824
rect 6638 11772 6644 11824
rect 6696 11812 6702 11824
rect 7101 11815 7159 11821
rect 7101 11812 7113 11815
rect 6696 11784 7113 11812
rect 6696 11772 6702 11784
rect 7101 11781 7113 11784
rect 7147 11781 7159 11815
rect 7668 11812 7696 11852
rect 8297 11849 8309 11883
rect 8343 11880 8355 11883
rect 8386 11880 8392 11892
rect 8343 11852 8392 11880
rect 8343 11849 8355 11852
rect 8297 11843 8355 11849
rect 8386 11840 8392 11852
rect 8444 11840 8450 11892
rect 8478 11840 8484 11892
rect 8536 11880 8542 11892
rect 9125 11883 9183 11889
rect 9125 11880 9137 11883
rect 8536 11852 9137 11880
rect 8536 11840 8542 11852
rect 9125 11849 9137 11852
rect 9171 11849 9183 11883
rect 9125 11843 9183 11849
rect 9674 11840 9680 11892
rect 9732 11880 9738 11892
rect 9953 11883 10011 11889
rect 9953 11880 9965 11883
rect 9732 11852 9965 11880
rect 9732 11840 9738 11852
rect 9953 11849 9965 11852
rect 9999 11880 10011 11883
rect 10413 11883 10471 11889
rect 10413 11880 10425 11883
rect 9999 11852 10425 11880
rect 9999 11849 10011 11852
rect 9953 11843 10011 11849
rect 10413 11849 10425 11852
rect 10459 11880 10471 11883
rect 10962 11880 10968 11892
rect 10459 11852 10968 11880
rect 10459 11849 10471 11852
rect 10413 11843 10471 11849
rect 10962 11840 10968 11852
rect 11020 11840 11026 11892
rect 13081 11883 13139 11889
rect 13081 11849 13093 11883
rect 13127 11880 13139 11883
rect 13262 11880 13268 11892
rect 13127 11852 13268 11880
rect 13127 11849 13139 11852
rect 13081 11843 13139 11849
rect 13262 11840 13268 11852
rect 13320 11840 13326 11892
rect 13630 11840 13636 11892
rect 13688 11880 13694 11892
rect 15013 11883 15071 11889
rect 15013 11880 15025 11883
rect 13688 11852 15025 11880
rect 13688 11840 13694 11852
rect 15013 11849 15025 11852
rect 15059 11880 15071 11883
rect 16393 11883 16451 11889
rect 16393 11880 16405 11883
rect 15059 11852 16405 11880
rect 15059 11849 15071 11852
rect 15013 11843 15071 11849
rect 16393 11849 16405 11852
rect 16439 11880 16451 11883
rect 18138 11880 18144 11892
rect 16439 11852 18144 11880
rect 16439 11849 16451 11852
rect 16393 11843 16451 11849
rect 18138 11840 18144 11852
rect 18196 11840 18202 11892
rect 12621 11815 12679 11821
rect 12621 11812 12633 11815
rect 7668 11784 12633 11812
rect 7101 11775 7159 11781
rect 12621 11781 12633 11784
rect 12667 11812 12679 11815
rect 15194 11812 15200 11824
rect 12667 11784 15200 11812
rect 12667 11781 12679 11784
rect 12621 11775 12679 11781
rect 15194 11772 15200 11784
rect 15252 11772 15258 11824
rect 15930 11812 15936 11824
rect 15891 11784 15936 11812
rect 15930 11772 15936 11784
rect 15988 11772 15994 11824
rect 17218 11812 17224 11824
rect 17179 11784 17224 11812
rect 17218 11772 17224 11784
rect 17276 11772 17282 11824
rect 1949 11747 2007 11753
rect 1949 11713 1961 11747
rect 1995 11744 2007 11747
rect 2501 11747 2559 11753
rect 1995 11716 2360 11744
rect 1995 11713 2007 11716
rect 1949 11707 2007 11713
rect 2222 11676 2228 11688
rect 2183 11648 2228 11676
rect 2222 11636 2228 11648
rect 2280 11636 2286 11688
rect 2332 11676 2360 11716
rect 2501 11713 2513 11747
rect 2547 11713 2559 11747
rect 2501 11707 2559 11713
rect 2777 11747 2835 11753
rect 2777 11713 2789 11747
rect 2823 11744 2835 11747
rect 5718 11744 5724 11756
rect 2823 11716 5724 11744
rect 2823 11713 2835 11716
rect 2777 11707 2835 11713
rect 5718 11704 5724 11716
rect 5776 11704 5782 11756
rect 5813 11747 5871 11753
rect 5813 11713 5825 11747
rect 5859 11744 5871 11747
rect 6472 11744 6500 11772
rect 7006 11744 7012 11756
rect 5859 11716 6500 11744
rect 6967 11716 7012 11744
rect 5859 11713 5871 11716
rect 5813 11707 5871 11713
rect 7006 11704 7012 11716
rect 7064 11704 7070 11756
rect 7374 11744 7380 11756
rect 7116 11716 7380 11744
rect 3418 11676 3424 11688
rect 2332 11648 3424 11676
rect 3418 11636 3424 11648
rect 3476 11636 3482 11688
rect 3605 11679 3663 11685
rect 3605 11645 3617 11679
rect 3651 11676 3663 11679
rect 4522 11676 4528 11688
rect 3651 11648 4528 11676
rect 3651 11645 3663 11648
rect 3605 11639 3663 11645
rect 4522 11636 4528 11648
rect 4580 11636 4586 11688
rect 6089 11679 6147 11685
rect 6089 11645 6101 11679
rect 6135 11676 6147 11679
rect 7116 11676 7144 11716
rect 7374 11704 7380 11716
rect 7432 11704 7438 11756
rect 9217 11747 9275 11753
rect 9217 11713 9229 11747
rect 9263 11744 9275 11747
rect 9766 11744 9772 11756
rect 9263 11716 9772 11744
rect 9263 11713 9275 11716
rect 9217 11707 9275 11713
rect 9766 11704 9772 11716
rect 9824 11704 9830 11756
rect 12710 11744 12716 11756
rect 12623 11716 12716 11744
rect 12710 11704 12716 11716
rect 12768 11744 12774 11756
rect 13262 11744 13268 11756
rect 12768 11716 13268 11744
rect 12768 11704 12774 11716
rect 13262 11704 13268 11716
rect 13320 11704 13326 11756
rect 14550 11704 14556 11756
rect 14608 11744 14614 11756
rect 15105 11747 15163 11753
rect 15105 11744 15117 11747
rect 14608 11716 15117 11744
rect 14608 11704 14614 11716
rect 15105 11713 15117 11716
rect 15151 11713 15163 11747
rect 17129 11747 17187 11753
rect 15105 11707 15163 11713
rect 15212 11716 16160 11744
rect 6135 11648 7144 11676
rect 6135 11645 6147 11648
rect 6089 11639 6147 11645
rect 7190 11636 7196 11688
rect 7248 11676 7254 11688
rect 7745 11679 7803 11685
rect 7745 11676 7757 11679
rect 7248 11648 7293 11676
rect 7392 11648 7757 11676
rect 7248 11636 7254 11648
rect 2240 11608 2268 11636
rect 3789 11611 3847 11617
rect 3789 11608 3801 11611
rect 2240 11580 3801 11608
rect 3789 11577 3801 11580
rect 3835 11577 3847 11611
rect 3789 11571 3847 11577
rect 5258 11568 5264 11620
rect 5316 11608 5322 11620
rect 6641 11611 6699 11617
rect 6641 11608 6653 11611
rect 5316 11580 6653 11608
rect 5316 11568 5322 11580
rect 6641 11577 6653 11580
rect 6687 11577 6699 11611
rect 6641 11571 6699 11577
rect 7098 11568 7104 11620
rect 7156 11608 7162 11620
rect 7392 11608 7420 11648
rect 7745 11645 7757 11648
rect 7791 11645 7803 11679
rect 7745 11639 7803 11645
rect 8113 11679 8171 11685
rect 8113 11645 8125 11679
rect 8159 11645 8171 11679
rect 8113 11639 8171 11645
rect 8205 11679 8263 11685
rect 8205 11645 8217 11679
rect 8251 11676 8263 11679
rect 8251 11648 8800 11676
rect 8251 11645 8263 11648
rect 8205 11639 8263 11645
rect 7156 11580 7420 11608
rect 8128 11608 8156 11639
rect 8386 11608 8392 11620
rect 8128 11580 8392 11608
rect 7156 11568 7162 11580
rect 8386 11568 8392 11580
rect 8444 11568 8450 11620
rect 8772 11617 8800 11648
rect 9398 11636 9404 11688
rect 9456 11676 9462 11688
rect 10042 11676 10048 11688
rect 9456 11648 9549 11676
rect 10003 11648 10048 11676
rect 9456 11636 9462 11648
rect 10042 11636 10048 11648
rect 10100 11636 10106 11688
rect 10226 11676 10232 11688
rect 10187 11648 10232 11676
rect 10226 11636 10232 11648
rect 10284 11636 10290 11688
rect 12529 11679 12587 11685
rect 12529 11645 12541 11679
rect 12575 11676 12587 11679
rect 12618 11676 12624 11688
rect 12575 11648 12624 11676
rect 12575 11645 12587 11648
rect 12529 11639 12587 11645
rect 12618 11636 12624 11648
rect 12676 11676 12682 11688
rect 14642 11676 14648 11688
rect 12676 11648 14648 11676
rect 12676 11636 12682 11648
rect 14642 11636 14648 11648
rect 14700 11636 14706 11688
rect 14921 11679 14979 11685
rect 14921 11645 14933 11679
rect 14967 11645 14979 11679
rect 15212 11676 15240 11716
rect 16022 11676 16028 11688
rect 14921 11639 14979 11645
rect 15120 11648 15240 11676
rect 15983 11648 16028 11676
rect 8757 11611 8815 11617
rect 8757 11577 8769 11611
rect 8803 11577 8815 11611
rect 8757 11571 8815 11577
rect 8846 11568 8852 11620
rect 8904 11608 8910 11620
rect 9416 11608 9444 11636
rect 13078 11608 13084 11620
rect 8904 11580 9352 11608
rect 9416 11580 13084 11608
rect 8904 11568 8910 11580
rect 1854 11500 1860 11552
rect 1912 11540 1918 11552
rect 2317 11543 2375 11549
rect 2317 11540 2329 11543
rect 1912 11512 2329 11540
rect 1912 11500 1918 11512
rect 2317 11509 2329 11512
rect 2363 11509 2375 11543
rect 2590 11540 2596 11552
rect 2551 11512 2596 11540
rect 2317 11503 2375 11509
rect 2590 11500 2596 11512
rect 2648 11500 2654 11552
rect 2958 11540 2964 11552
rect 2919 11512 2964 11540
rect 2958 11500 2964 11512
rect 3016 11500 3022 11552
rect 3418 11500 3424 11552
rect 3476 11540 3482 11552
rect 3694 11540 3700 11552
rect 3476 11512 3700 11540
rect 3476 11500 3482 11512
rect 3694 11500 3700 11512
rect 3752 11500 3758 11552
rect 3970 11540 3976 11552
rect 3931 11512 3976 11540
rect 3970 11500 3976 11512
rect 4028 11500 4034 11552
rect 5442 11500 5448 11552
rect 5500 11540 5506 11552
rect 7561 11543 7619 11549
rect 7561 11540 7573 11543
rect 5500 11512 7573 11540
rect 5500 11500 5506 11512
rect 7561 11509 7573 11512
rect 7607 11540 7619 11543
rect 7926 11540 7932 11552
rect 7607 11512 7932 11540
rect 7607 11509 7619 11512
rect 7561 11503 7619 11509
rect 7926 11500 7932 11512
rect 7984 11500 7990 11552
rect 8665 11543 8723 11549
rect 8665 11509 8677 11543
rect 8711 11540 8723 11543
rect 9122 11540 9128 11552
rect 8711 11512 9128 11540
rect 8711 11509 8723 11512
rect 8665 11503 8723 11509
rect 9122 11500 9128 11512
rect 9180 11500 9186 11552
rect 9324 11540 9352 11580
rect 13078 11568 13084 11580
rect 13136 11568 13142 11620
rect 14936 11608 14964 11639
rect 15120 11608 15148 11648
rect 16022 11636 16028 11648
rect 16080 11636 16086 11688
rect 16132 11685 16160 11716
rect 17129 11713 17141 11747
rect 17175 11744 17187 11747
rect 17586 11744 17592 11756
rect 17175 11716 17592 11744
rect 17175 11713 17187 11716
rect 17129 11707 17187 11713
rect 17586 11704 17592 11716
rect 17644 11744 17650 11756
rect 18414 11744 18420 11756
rect 17644 11716 18420 11744
rect 17644 11704 17650 11716
rect 18414 11704 18420 11716
rect 18472 11704 18478 11756
rect 16117 11679 16175 11685
rect 16117 11645 16129 11679
rect 16163 11645 16175 11679
rect 16117 11639 16175 11645
rect 17310 11636 17316 11688
rect 17368 11676 17374 11688
rect 17405 11679 17463 11685
rect 17405 11676 17417 11679
rect 17368 11648 17417 11676
rect 17368 11636 17374 11648
rect 17405 11645 17417 11648
rect 17451 11645 17463 11679
rect 17678 11676 17684 11688
rect 17639 11648 17684 11676
rect 17405 11639 17463 11645
rect 17678 11636 17684 11648
rect 17736 11636 17742 11688
rect 17957 11679 18015 11685
rect 17957 11645 17969 11679
rect 18003 11676 18015 11679
rect 18874 11676 18880 11688
rect 18003 11648 18880 11676
rect 18003 11645 18015 11648
rect 17957 11639 18015 11645
rect 18874 11636 18880 11648
rect 18932 11636 18938 11688
rect 14936 11580 15148 11608
rect 15028 11552 15056 11580
rect 9585 11543 9643 11549
rect 9585 11540 9597 11543
rect 9324 11512 9597 11540
rect 9585 11509 9597 11512
rect 9631 11509 9643 11543
rect 9585 11503 9643 11509
rect 9858 11500 9864 11552
rect 9916 11540 9922 11552
rect 13170 11540 13176 11552
rect 9916 11512 13176 11540
rect 9916 11500 9922 11512
rect 13170 11500 13176 11512
rect 13228 11500 13234 11552
rect 14550 11540 14556 11552
rect 14511 11512 14556 11540
rect 14550 11500 14556 11512
rect 14608 11500 14614 11552
rect 15010 11500 15016 11552
rect 15068 11500 15074 11552
rect 15378 11500 15384 11552
rect 15436 11540 15442 11552
rect 15473 11543 15531 11549
rect 15473 11540 15485 11543
rect 15436 11512 15485 11540
rect 15436 11500 15442 11512
rect 15473 11509 15485 11512
rect 15519 11509 15531 11543
rect 15473 11503 15531 11509
rect 15562 11500 15568 11552
rect 15620 11540 15626 11552
rect 16761 11543 16819 11549
rect 15620 11512 15665 11540
rect 15620 11500 15626 11512
rect 16761 11509 16773 11543
rect 16807 11540 16819 11543
rect 16850 11540 16856 11552
rect 16807 11512 16856 11540
rect 16807 11509 16819 11512
rect 16761 11503 16819 11509
rect 16850 11500 16856 11512
rect 16908 11500 16914 11552
rect 1104 11450 18860 11472
rect 1104 11398 3174 11450
rect 3226 11398 3238 11450
rect 3290 11398 3302 11450
rect 3354 11398 3366 11450
rect 3418 11398 3430 11450
rect 3482 11398 7622 11450
rect 7674 11398 7686 11450
rect 7738 11398 7750 11450
rect 7802 11398 7814 11450
rect 7866 11398 7878 11450
rect 7930 11398 12070 11450
rect 12122 11398 12134 11450
rect 12186 11398 12198 11450
rect 12250 11398 12262 11450
rect 12314 11398 12326 11450
rect 12378 11398 16518 11450
rect 16570 11398 16582 11450
rect 16634 11398 16646 11450
rect 16698 11398 16710 11450
rect 16762 11398 16774 11450
rect 16826 11398 18860 11450
rect 1104 11376 18860 11398
rect 2866 11336 2872 11348
rect 2516 11308 2872 11336
rect 1302 11228 1308 11280
rect 1360 11268 1366 11280
rect 2317 11271 2375 11277
rect 2317 11268 2329 11271
rect 1360 11240 2329 11268
rect 1360 11228 1366 11240
rect 2317 11237 2329 11240
rect 2363 11237 2375 11271
rect 2317 11231 2375 11237
rect 1946 11200 1952 11212
rect 1907 11172 1952 11200
rect 1946 11160 1952 11172
rect 2004 11160 2010 11212
rect 2222 11132 2228 11144
rect 2183 11104 2228 11132
rect 2222 11092 2228 11104
rect 2280 11092 2286 11144
rect 2516 11141 2544 11308
rect 2866 11296 2872 11308
rect 2924 11296 2930 11348
rect 4525 11339 4583 11345
rect 4525 11336 4537 11339
rect 3252 11308 4537 11336
rect 3252 11268 3280 11308
rect 4525 11305 4537 11308
rect 4571 11336 4583 11339
rect 4798 11336 4804 11348
rect 4571 11308 4804 11336
rect 4571 11305 4583 11308
rect 4525 11299 4583 11305
rect 4798 11296 4804 11308
rect 4856 11296 4862 11348
rect 7006 11296 7012 11348
rect 7064 11336 7070 11348
rect 7745 11339 7803 11345
rect 7745 11336 7757 11339
rect 7064 11308 7757 11336
rect 7064 11296 7070 11308
rect 7745 11305 7757 11308
rect 7791 11305 7803 11339
rect 7745 11299 7803 11305
rect 8570 11296 8576 11348
rect 8628 11336 8634 11348
rect 8941 11339 8999 11345
rect 8941 11336 8953 11339
rect 8628 11308 8953 11336
rect 8628 11296 8634 11308
rect 8941 11305 8953 11308
rect 8987 11305 8999 11339
rect 14093 11339 14151 11345
rect 14093 11336 14105 11339
rect 8941 11299 8999 11305
rect 10888 11308 14105 11336
rect 2792 11240 3280 11268
rect 3329 11271 3387 11277
rect 2792 11209 2820 11240
rect 3329 11237 3341 11271
rect 3375 11268 3387 11271
rect 3602 11268 3608 11280
rect 3375 11240 3608 11268
rect 3375 11237 3387 11240
rect 3329 11231 3387 11237
rect 3602 11228 3608 11240
rect 3660 11228 3666 11280
rect 8110 11268 8116 11280
rect 7024 11240 8116 11268
rect 7024 11212 7052 11240
rect 8110 11228 8116 11240
rect 8168 11228 8174 11280
rect 8846 11268 8852 11280
rect 8220 11240 8852 11268
rect 2777 11203 2835 11209
rect 2777 11169 2789 11203
rect 2823 11169 2835 11203
rect 2777 11163 2835 11169
rect 2869 11203 2927 11209
rect 2869 11169 2881 11203
rect 2915 11200 2927 11203
rect 3970 11200 3976 11212
rect 2915 11172 3976 11200
rect 2915 11169 2927 11172
rect 2869 11163 2927 11169
rect 3970 11160 3976 11172
rect 4028 11160 4034 11212
rect 7006 11160 7012 11212
rect 7064 11160 7070 11212
rect 8220 11209 8248 11240
rect 8846 11228 8852 11240
rect 8904 11228 8910 11280
rect 9858 11268 9864 11280
rect 8956 11240 9864 11268
rect 8205 11203 8263 11209
rect 8205 11169 8217 11203
rect 8251 11169 8263 11203
rect 8205 11163 8263 11169
rect 8297 11203 8355 11209
rect 8297 11169 8309 11203
rect 8343 11169 8355 11203
rect 8297 11163 8355 11169
rect 2501 11135 2559 11141
rect 2501 11101 2513 11135
rect 2547 11101 2559 11135
rect 2958 11132 2964 11144
rect 2919 11104 2964 11132
rect 2501 11095 2559 11101
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 3142 11092 3148 11144
rect 3200 11132 3206 11144
rect 3510 11132 3516 11144
rect 3200 11104 3516 11132
rect 3200 11092 3206 11104
rect 3510 11092 3516 11104
rect 3568 11092 3574 11144
rect 3694 11092 3700 11144
rect 3752 11132 3758 11144
rect 3752 11104 4016 11132
rect 3752 11092 3758 11104
rect 2240 11064 2268 11092
rect 3988 11076 4016 11104
rect 4522 11092 4528 11144
rect 4580 11132 4586 11144
rect 5638 11135 5696 11141
rect 5638 11132 5650 11135
rect 4580 11104 5650 11132
rect 4580 11092 4586 11104
rect 5638 11101 5650 11104
rect 5684 11101 5696 11135
rect 5638 11095 5696 11101
rect 5905 11135 5963 11141
rect 5905 11101 5917 11135
rect 5951 11132 5963 11135
rect 5994 11132 6000 11144
rect 5951 11104 6000 11132
rect 5951 11101 5963 11104
rect 5905 11095 5963 11101
rect 5994 11092 6000 11104
rect 6052 11092 6058 11144
rect 7466 11092 7472 11144
rect 7524 11132 7530 11144
rect 8110 11132 8116 11144
rect 7524 11104 8116 11132
rect 7524 11092 7530 11104
rect 8110 11092 8116 11104
rect 8168 11132 8174 11144
rect 8312 11132 8340 11163
rect 8168 11104 8340 11132
rect 8168 11092 8174 11104
rect 8478 11092 8484 11144
rect 8536 11132 8542 11144
rect 8573 11135 8631 11141
rect 8573 11132 8585 11135
rect 8536 11104 8585 11132
rect 8536 11092 8542 11104
rect 8573 11101 8585 11104
rect 8619 11101 8631 11135
rect 8956 11132 8984 11240
rect 9858 11228 9864 11240
rect 9916 11228 9922 11280
rect 9214 11160 9220 11212
rect 9272 11200 9278 11212
rect 9493 11203 9551 11209
rect 9493 11200 9505 11203
rect 9272 11172 9505 11200
rect 9272 11160 9278 11172
rect 9493 11169 9505 11172
rect 9539 11169 9551 11203
rect 9766 11200 9772 11212
rect 9727 11172 9772 11200
rect 9493 11163 9551 11169
rect 9766 11160 9772 11172
rect 9824 11160 9830 11212
rect 8573 11095 8631 11101
rect 8680 11104 8984 11132
rect 3789 11067 3847 11073
rect 3789 11064 3801 11067
rect 2240 11036 3801 11064
rect 3789 11033 3801 11036
rect 3835 11033 3847 11067
rect 3789 11027 3847 11033
rect 3970 11024 3976 11076
rect 4028 11024 4034 11076
rect 7282 11024 7288 11076
rect 7340 11064 7346 11076
rect 7653 11067 7711 11073
rect 7653 11064 7665 11067
rect 7340 11036 7665 11064
rect 7340 11024 7346 11036
rect 7653 11033 7665 11036
rect 7699 11064 7711 11067
rect 8680 11064 8708 11104
rect 9122 11092 9128 11144
rect 9180 11132 9186 11144
rect 9309 11135 9367 11141
rect 9309 11132 9321 11135
rect 9180 11104 9321 11132
rect 9180 11092 9186 11104
rect 9309 11101 9321 11104
rect 9355 11101 9367 11135
rect 9309 11095 9367 11101
rect 9401 11135 9459 11141
rect 9401 11101 9413 11135
rect 9447 11132 9459 11135
rect 10888 11132 10916 11308
rect 14093 11305 14105 11308
rect 14139 11305 14151 11339
rect 14093 11299 14151 11305
rect 15470 11296 15476 11348
rect 15528 11336 15534 11348
rect 15746 11336 15752 11348
rect 15528 11308 15752 11336
rect 15528 11296 15534 11308
rect 15746 11296 15752 11308
rect 15804 11296 15810 11348
rect 16025 11339 16083 11345
rect 16025 11305 16037 11339
rect 16071 11336 16083 11339
rect 16071 11308 17724 11336
rect 16071 11305 16083 11308
rect 16025 11299 16083 11305
rect 16117 11271 16175 11277
rect 16117 11268 16129 11271
rect 14568 11240 16129 11268
rect 14568 11209 14596 11240
rect 16117 11237 16129 11240
rect 16163 11237 16175 11271
rect 16117 11231 16175 11237
rect 17034 11228 17040 11280
rect 17092 11268 17098 11280
rect 17586 11268 17592 11280
rect 17092 11240 17592 11268
rect 17092 11228 17098 11240
rect 17586 11228 17592 11240
rect 17644 11228 17650 11280
rect 14553 11203 14611 11209
rect 14553 11169 14565 11203
rect 14599 11169 14611 11203
rect 14734 11200 14740 11212
rect 14695 11172 14740 11200
rect 14553 11163 14611 11169
rect 14734 11160 14740 11172
rect 14792 11160 14798 11212
rect 15378 11200 15384 11212
rect 15339 11172 15384 11200
rect 15378 11160 15384 11172
rect 15436 11160 15442 11212
rect 15470 11160 15476 11212
rect 15528 11200 15534 11212
rect 16669 11203 16727 11209
rect 16669 11200 16681 11203
rect 15528 11172 15573 11200
rect 15672 11172 16681 11200
rect 15528 11160 15534 11172
rect 9447 11104 10916 11132
rect 9447 11101 9459 11104
rect 9401 11095 9459 11101
rect 10962 11092 10968 11144
rect 11020 11132 11026 11144
rect 11238 11132 11244 11144
rect 11020 11104 11244 11132
rect 11020 11092 11026 11104
rect 11238 11092 11244 11104
rect 11296 11092 11302 11144
rect 11514 11092 11520 11144
rect 11572 11132 11578 11144
rect 11701 11135 11759 11141
rect 11701 11132 11713 11135
rect 11572 11104 11713 11132
rect 11572 11092 11578 11104
rect 11701 11101 11713 11104
rect 11747 11101 11759 11135
rect 15194 11132 15200 11144
rect 11701 11095 11759 11101
rect 11961 11104 15200 11132
rect 7699 11036 8708 11064
rect 7699 11033 7711 11036
rect 7653 11027 7711 11033
rect 2774 10956 2780 11008
rect 2832 10996 2838 11008
rect 5442 10996 5448 11008
rect 2832 10968 5448 10996
rect 2832 10956 2838 10968
rect 5442 10956 5448 10968
rect 5500 10956 5506 11008
rect 8128 11005 8156 11036
rect 8754 11024 8760 11076
rect 8812 11064 8818 11076
rect 11961 11073 11989 11104
rect 15194 11092 15200 11104
rect 15252 11092 15258 11144
rect 15289 11135 15347 11141
rect 15289 11101 15301 11135
rect 15335 11132 15347 11135
rect 15562 11132 15568 11144
rect 15335 11104 15568 11132
rect 15335 11101 15347 11104
rect 15289 11095 15347 11101
rect 15562 11092 15568 11104
rect 15620 11092 15626 11144
rect 11946 11067 12004 11073
rect 11946 11064 11958 11067
rect 8812 11036 11958 11064
rect 8812 11024 8818 11036
rect 11946 11033 11958 11036
rect 11992 11033 12004 11067
rect 13630 11064 13636 11076
rect 11946 11027 12004 11033
rect 12406 11036 13636 11064
rect 8113 10999 8171 11005
rect 8113 10965 8125 10999
rect 8159 10965 8171 10999
rect 8113 10959 8171 10965
rect 10318 10956 10324 11008
rect 10376 10996 10382 11008
rect 12406 10996 12434 11036
rect 13630 11024 13636 11036
rect 13688 11024 13694 11076
rect 14461 11067 14519 11073
rect 14461 11033 14473 11067
rect 14507 11064 14519 11067
rect 14642 11064 14648 11076
rect 14507 11036 14648 11064
rect 14507 11033 14519 11036
rect 14461 11027 14519 11033
rect 14642 11024 14648 11036
rect 14700 11024 14706 11076
rect 15102 11064 15108 11076
rect 14752 11036 15108 11064
rect 13078 10996 13084 11008
rect 10376 10968 12434 10996
rect 12991 10968 13084 10996
rect 10376 10956 10382 10968
rect 13078 10956 13084 10968
rect 13136 10996 13142 11008
rect 14752 10996 14780 11036
rect 15102 11024 15108 11036
rect 15160 11064 15166 11076
rect 15672 11064 15700 11172
rect 16669 11169 16681 11172
rect 16715 11169 16727 11203
rect 16669 11163 16727 11169
rect 17696 11144 17724 11308
rect 16485 11135 16543 11141
rect 16485 11101 16497 11135
rect 16531 11132 16543 11135
rect 16850 11132 16856 11144
rect 16531 11104 16856 11132
rect 16531 11101 16543 11104
rect 16485 11095 16543 11101
rect 16850 11092 16856 11104
rect 16908 11092 16914 11144
rect 17037 11135 17095 11141
rect 17037 11101 17049 11135
rect 17083 11132 17095 11135
rect 17126 11132 17132 11144
rect 17083 11104 17132 11132
rect 17083 11101 17095 11104
rect 17037 11095 17095 11101
rect 17126 11092 17132 11104
rect 17184 11092 17190 11144
rect 17405 11135 17463 11141
rect 17405 11101 17417 11135
rect 17451 11132 17463 11135
rect 17494 11132 17500 11144
rect 17451 11104 17500 11132
rect 17451 11101 17463 11104
rect 17405 11095 17463 11101
rect 17494 11092 17500 11104
rect 17552 11092 17558 11144
rect 17678 11132 17684 11144
rect 17639 11104 17684 11132
rect 17678 11092 17684 11104
rect 17736 11092 17742 11144
rect 17954 11132 17960 11144
rect 17915 11104 17960 11132
rect 17954 11092 17960 11104
rect 18012 11092 18018 11144
rect 15160 11036 15700 11064
rect 15160 11024 15166 11036
rect 16390 11024 16396 11076
rect 16448 11064 16454 11076
rect 16577 11067 16635 11073
rect 16577 11064 16589 11067
rect 16448 11036 16589 11064
rect 16448 11024 16454 11036
rect 16577 11033 16589 11036
rect 16623 11033 16635 11067
rect 18598 11064 18604 11076
rect 16577 11027 16635 11033
rect 17328 11036 18604 11064
rect 14918 10996 14924 11008
rect 13136 10968 14780 10996
rect 14879 10968 14924 10996
rect 13136 10956 13142 10968
rect 14918 10956 14924 10968
rect 14976 10956 14982 11008
rect 17328 11005 17356 11036
rect 18598 11024 18604 11036
rect 18656 11024 18662 11076
rect 17313 10999 17371 11005
rect 17313 10965 17325 10999
rect 17359 10965 17371 10999
rect 17313 10959 17371 10965
rect 17589 10999 17647 11005
rect 17589 10965 17601 10999
rect 17635 10996 17647 10999
rect 18046 10996 18052 11008
rect 17635 10968 18052 10996
rect 17635 10965 17647 10968
rect 17589 10959 17647 10965
rect 18046 10956 18052 10968
rect 18104 10956 18110 11008
rect 1104 10906 18860 10928
rect 1104 10854 5398 10906
rect 5450 10854 5462 10906
rect 5514 10854 5526 10906
rect 5578 10854 5590 10906
rect 5642 10854 5654 10906
rect 5706 10854 9846 10906
rect 9898 10854 9910 10906
rect 9962 10854 9974 10906
rect 10026 10854 10038 10906
rect 10090 10854 10102 10906
rect 10154 10854 14294 10906
rect 14346 10854 14358 10906
rect 14410 10854 14422 10906
rect 14474 10854 14486 10906
rect 14538 10854 14550 10906
rect 14602 10854 18860 10906
rect 1104 10832 18860 10854
rect 1578 10752 1584 10804
rect 1636 10792 1642 10804
rect 2774 10792 2780 10804
rect 1636 10764 2780 10792
rect 1636 10752 1642 10764
rect 2774 10752 2780 10764
rect 2832 10752 2838 10804
rect 2869 10795 2927 10801
rect 2869 10761 2881 10795
rect 2915 10792 2927 10795
rect 3694 10792 3700 10804
rect 2915 10764 3700 10792
rect 2915 10761 2927 10764
rect 2869 10755 2927 10761
rect 3694 10752 3700 10764
rect 3752 10792 3758 10804
rect 4341 10795 4399 10801
rect 4341 10792 4353 10795
rect 3752 10764 4353 10792
rect 3752 10752 3758 10764
rect 4341 10761 4353 10764
rect 4387 10792 4399 10795
rect 8205 10795 8263 10801
rect 4387 10764 7972 10792
rect 4387 10761 4399 10764
rect 4341 10755 4399 10761
rect 3436 10696 3832 10724
rect 2777 10659 2835 10665
rect 2777 10625 2789 10659
rect 2823 10656 2835 10659
rect 3142 10656 3148 10668
rect 2823 10628 3148 10656
rect 2823 10625 2835 10628
rect 2777 10619 2835 10625
rect 3142 10616 3148 10628
rect 3200 10616 3206 10668
rect 1949 10591 2007 10597
rect 1949 10557 1961 10591
rect 1995 10557 2007 10591
rect 2222 10588 2228 10600
rect 2183 10560 2228 10588
rect 1949 10551 2007 10557
rect 1964 10520 1992 10551
rect 2222 10548 2228 10560
rect 2280 10548 2286 10600
rect 2961 10591 3019 10597
rect 2961 10557 2973 10591
rect 3007 10588 3019 10591
rect 3436 10588 3464 10696
rect 3510 10616 3516 10668
rect 3568 10656 3574 10668
rect 3605 10659 3663 10665
rect 3605 10656 3617 10659
rect 3568 10628 3617 10656
rect 3568 10616 3574 10628
rect 3605 10625 3617 10628
rect 3651 10625 3663 10659
rect 3605 10619 3663 10625
rect 3804 10597 3832 10696
rect 5718 10684 5724 10736
rect 5776 10724 5782 10736
rect 5914 10727 5972 10733
rect 5914 10724 5926 10727
rect 5776 10696 5926 10724
rect 5776 10684 5782 10696
rect 5914 10693 5926 10696
rect 5960 10724 5972 10727
rect 7190 10724 7196 10736
rect 5960 10696 7196 10724
rect 5960 10693 5972 10696
rect 5914 10687 5972 10693
rect 7190 10684 7196 10696
rect 7248 10684 7254 10736
rect 6086 10616 6092 10668
rect 6144 10656 6150 10668
rect 6181 10659 6239 10665
rect 6181 10656 6193 10659
rect 6144 10628 6193 10656
rect 6144 10616 6150 10628
rect 6181 10625 6193 10628
rect 6227 10656 6239 10659
rect 6825 10659 6883 10665
rect 6825 10656 6837 10659
rect 6227 10628 6837 10656
rect 6227 10625 6239 10628
rect 6181 10619 6239 10625
rect 6825 10625 6837 10628
rect 6871 10625 6883 10659
rect 7081 10659 7139 10665
rect 7081 10656 7093 10659
rect 6825 10619 6883 10625
rect 6932 10628 7093 10656
rect 3007 10560 3464 10588
rect 3697 10591 3755 10597
rect 3007 10557 3019 10560
rect 2961 10551 3019 10557
rect 3697 10557 3709 10591
rect 3743 10557 3755 10591
rect 3697 10551 3755 10557
rect 3789 10591 3847 10597
rect 3789 10557 3801 10591
rect 3835 10588 3847 10591
rect 4430 10588 4436 10600
rect 3835 10560 4436 10588
rect 3835 10557 3847 10560
rect 3789 10551 3847 10557
rect 2130 10520 2136 10532
rect 1964 10492 2136 10520
rect 2130 10480 2136 10492
rect 2188 10480 2194 10532
rect 3050 10480 3056 10532
rect 3108 10520 3114 10532
rect 3712 10520 3740 10551
rect 4430 10548 4436 10560
rect 4488 10548 4494 10600
rect 6932 10588 6960 10628
rect 7081 10625 7093 10628
rect 7127 10625 7139 10659
rect 7208 10656 7236 10684
rect 7944 10656 7972 10764
rect 8205 10761 8217 10795
rect 8251 10792 8263 10795
rect 9214 10792 9220 10804
rect 8251 10764 9220 10792
rect 8251 10761 8263 10764
rect 8205 10755 8263 10761
rect 9214 10752 9220 10764
rect 9272 10752 9278 10804
rect 11517 10795 11575 10801
rect 11517 10761 11529 10795
rect 11563 10761 11575 10795
rect 11517 10755 11575 10761
rect 8110 10684 8116 10736
rect 8168 10724 8174 10736
rect 9410 10727 9468 10733
rect 9410 10724 9422 10727
rect 8168 10696 9422 10724
rect 8168 10684 8174 10696
rect 9410 10693 9422 10696
rect 9456 10693 9468 10727
rect 10318 10724 10324 10736
rect 9410 10687 9468 10693
rect 9508 10696 10324 10724
rect 9508 10656 9536 10696
rect 10318 10684 10324 10696
rect 10376 10684 10382 10736
rect 11532 10724 11560 10755
rect 11606 10752 11612 10804
rect 11664 10792 11670 10804
rect 11974 10792 11980 10804
rect 11664 10764 11980 10792
rect 11664 10752 11670 10764
rect 11974 10752 11980 10764
rect 12032 10792 12038 10804
rect 14369 10795 14427 10801
rect 14369 10792 14381 10795
rect 12032 10764 14381 10792
rect 12032 10752 12038 10764
rect 14369 10761 14381 10764
rect 14415 10761 14427 10795
rect 14642 10792 14648 10804
rect 14603 10764 14648 10792
rect 14369 10755 14427 10761
rect 14642 10752 14648 10764
rect 14700 10752 14706 10804
rect 15105 10795 15163 10801
rect 15105 10761 15117 10795
rect 15151 10792 15163 10795
rect 16669 10795 16727 10801
rect 16669 10792 16681 10795
rect 15151 10764 16681 10792
rect 15151 10761 15163 10764
rect 15105 10755 15163 10761
rect 16669 10761 16681 10764
rect 16715 10761 16727 10795
rect 17034 10792 17040 10804
rect 16995 10764 17040 10792
rect 16669 10755 16727 10761
rect 17034 10752 17040 10764
rect 17092 10792 17098 10804
rect 17497 10795 17555 10801
rect 17497 10792 17509 10795
rect 17092 10764 17509 10792
rect 17092 10752 17098 10764
rect 17497 10761 17509 10764
rect 17543 10792 17555 10795
rect 17954 10792 17960 10804
rect 17543 10764 17960 10792
rect 17543 10761 17555 10764
rect 17497 10755 17555 10761
rect 17954 10752 17960 10764
rect 18012 10752 18018 10804
rect 13256 10727 13314 10733
rect 13256 10724 13268 10727
rect 11532 10696 13268 10724
rect 13256 10693 13268 10696
rect 13302 10724 13314 10727
rect 13354 10724 13360 10736
rect 13302 10696 13360 10724
rect 13302 10693 13314 10696
rect 13256 10687 13314 10693
rect 13354 10684 13360 10696
rect 13412 10684 13418 10736
rect 15194 10684 15200 10736
rect 15252 10684 15258 10736
rect 7208 10628 7880 10656
rect 7944 10628 9536 10656
rect 10128 10659 10186 10665
rect 7081 10619 7139 10625
rect 6840 10560 6960 10588
rect 3108 10492 3740 10520
rect 3108 10480 3114 10492
rect 2409 10455 2467 10461
rect 2409 10421 2421 10455
rect 2455 10452 2467 10455
rect 2498 10452 2504 10464
rect 2455 10424 2504 10452
rect 2455 10421 2467 10424
rect 2409 10415 2467 10421
rect 2498 10412 2504 10424
rect 2556 10412 2562 10464
rect 2682 10412 2688 10464
rect 2740 10452 2746 10464
rect 3237 10455 3295 10461
rect 3237 10452 3249 10455
rect 2740 10424 3249 10452
rect 2740 10412 2746 10424
rect 3237 10421 3249 10424
rect 3283 10421 3295 10455
rect 3712 10452 3740 10492
rect 4154 10452 4160 10464
rect 3712 10424 4160 10452
rect 3237 10415 3295 10421
rect 4154 10412 4160 10424
rect 4212 10412 4218 10464
rect 4801 10455 4859 10461
rect 4801 10421 4813 10455
rect 4847 10452 4859 10455
rect 5258 10452 5264 10464
rect 4847 10424 5264 10452
rect 4847 10421 4859 10424
rect 4801 10415 4859 10421
rect 5258 10412 5264 10424
rect 5316 10412 5322 10464
rect 6840 10452 6868 10560
rect 7852 10520 7880 10628
rect 10128 10625 10140 10659
rect 10174 10656 10186 10659
rect 11606 10656 11612 10668
rect 10174 10628 11612 10656
rect 10174 10625 10186 10628
rect 10128 10619 10186 10625
rect 11606 10616 11612 10628
rect 11664 10616 11670 10668
rect 12618 10616 12624 10668
rect 12676 10665 12682 10668
rect 12676 10656 12688 10665
rect 14458 10656 14464 10668
rect 12676 10628 12721 10656
rect 14419 10628 14464 10656
rect 12676 10619 12688 10628
rect 12676 10616 12682 10619
rect 14458 10616 14464 10628
rect 14516 10656 14522 10668
rect 15013 10659 15071 10665
rect 15013 10656 15025 10659
rect 14516 10628 15025 10656
rect 14516 10616 14522 10628
rect 15013 10625 15025 10628
rect 15059 10625 15071 10659
rect 15212 10656 15240 10684
rect 15212 10628 17264 10656
rect 15013 10619 15071 10625
rect 9674 10588 9680 10600
rect 9635 10560 9680 10588
rect 9674 10548 9680 10560
rect 9732 10588 9738 10600
rect 9861 10591 9919 10597
rect 9861 10588 9873 10591
rect 9732 10560 9873 10588
rect 9732 10548 9738 10560
rect 9861 10557 9873 10560
rect 9907 10557 9919 10591
rect 12894 10588 12900 10600
rect 12855 10560 12900 10588
rect 9861 10551 9919 10557
rect 12894 10548 12900 10560
rect 12952 10588 12958 10600
rect 12989 10591 13047 10597
rect 12989 10588 13001 10591
rect 12952 10560 13001 10588
rect 12952 10548 12958 10560
rect 12989 10557 13001 10560
rect 13035 10557 13047 10591
rect 12989 10551 13047 10557
rect 15102 10548 15108 10600
rect 15160 10588 15166 10600
rect 15197 10591 15255 10597
rect 15197 10588 15209 10591
rect 15160 10560 15209 10588
rect 15160 10548 15166 10560
rect 15197 10557 15209 10560
rect 15243 10557 15255 10591
rect 17126 10588 17132 10600
rect 15197 10551 15255 10557
rect 15856 10560 17132 10588
rect 8297 10523 8355 10529
rect 8297 10520 8309 10523
rect 7852 10492 8309 10520
rect 8297 10489 8309 10492
rect 8343 10489 8355 10523
rect 8297 10483 8355 10489
rect 10870 10480 10876 10532
rect 10928 10520 10934 10532
rect 15856 10520 15884 10560
rect 17126 10548 17132 10560
rect 17184 10548 17190 10600
rect 17236 10597 17264 10628
rect 17221 10591 17279 10597
rect 17221 10557 17233 10591
rect 17267 10588 17279 10591
rect 17310 10588 17316 10600
rect 17267 10560 17316 10588
rect 17267 10557 17279 10560
rect 17221 10551 17279 10557
rect 17310 10548 17316 10560
rect 17368 10548 17374 10600
rect 17678 10588 17684 10600
rect 17639 10560 17684 10588
rect 17678 10548 17684 10560
rect 17736 10548 17742 10600
rect 17957 10591 18015 10597
rect 17957 10557 17969 10591
rect 18003 10588 18015 10591
rect 18322 10588 18328 10600
rect 18003 10560 18328 10588
rect 18003 10557 18015 10560
rect 17957 10551 18015 10557
rect 18322 10548 18328 10560
rect 18380 10548 18386 10600
rect 10928 10492 11376 10520
rect 10928 10480 10934 10492
rect 8386 10452 8392 10464
rect 6840 10424 8392 10452
rect 8386 10412 8392 10424
rect 8444 10452 8450 10464
rect 10594 10452 10600 10464
rect 8444 10424 10600 10452
rect 8444 10412 8450 10424
rect 10594 10412 10600 10424
rect 10652 10412 10658 10464
rect 11238 10452 11244 10464
rect 11199 10424 11244 10452
rect 11238 10412 11244 10424
rect 11296 10412 11302 10464
rect 11348 10452 11376 10492
rect 14384 10492 15884 10520
rect 16485 10523 16543 10529
rect 14384 10452 14412 10492
rect 16485 10489 16497 10523
rect 16531 10520 16543 10523
rect 17696 10520 17724 10548
rect 16531 10492 17724 10520
rect 16531 10489 16543 10492
rect 16485 10483 16543 10489
rect 11348 10424 14412 10452
rect 1104 10362 18860 10384
rect 1104 10310 3174 10362
rect 3226 10310 3238 10362
rect 3290 10310 3302 10362
rect 3354 10310 3366 10362
rect 3418 10310 3430 10362
rect 3482 10310 7622 10362
rect 7674 10310 7686 10362
rect 7738 10310 7750 10362
rect 7802 10310 7814 10362
rect 7866 10310 7878 10362
rect 7930 10310 12070 10362
rect 12122 10310 12134 10362
rect 12186 10310 12198 10362
rect 12250 10310 12262 10362
rect 12314 10310 12326 10362
rect 12378 10310 16518 10362
rect 16570 10310 16582 10362
rect 16634 10310 16646 10362
rect 16698 10310 16710 10362
rect 16762 10310 16774 10362
rect 16826 10310 18860 10362
rect 1104 10288 18860 10310
rect 1578 10248 1584 10260
rect 1539 10220 1584 10248
rect 1578 10208 1584 10220
rect 1636 10208 1642 10260
rect 2222 10208 2228 10260
rect 2280 10248 2286 10260
rect 3789 10251 3847 10257
rect 3789 10248 3801 10251
rect 2280 10220 3801 10248
rect 2280 10208 2286 10220
rect 3789 10217 3801 10220
rect 3835 10217 3847 10251
rect 3789 10211 3847 10217
rect 4154 10208 4160 10260
rect 4212 10248 4218 10260
rect 4212 10220 10548 10248
rect 4212 10208 4218 10220
rect 3050 10180 3056 10192
rect 1964 10152 3056 10180
rect 1964 10056 1992 10152
rect 3050 10140 3056 10152
rect 3108 10140 3114 10192
rect 3510 10180 3516 10192
rect 3160 10152 3516 10180
rect 2498 10112 2504 10124
rect 2459 10084 2504 10112
rect 2498 10072 2504 10084
rect 2556 10072 2562 10124
rect 3160 10121 3188 10152
rect 3510 10140 3516 10152
rect 3568 10140 3574 10192
rect 6546 10180 6552 10192
rect 6507 10152 6552 10180
rect 6546 10140 6552 10152
rect 6604 10140 6610 10192
rect 8110 10140 8116 10192
rect 8168 10180 8174 10192
rect 9033 10183 9091 10189
rect 9033 10180 9045 10183
rect 8168 10152 9045 10180
rect 8168 10140 8174 10152
rect 9033 10149 9045 10152
rect 9079 10149 9091 10183
rect 9033 10143 9091 10149
rect 2593 10115 2651 10121
rect 2593 10081 2605 10115
rect 2639 10081 2651 10115
rect 2593 10075 2651 10081
rect 3145 10115 3203 10121
rect 3145 10081 3157 10115
rect 3191 10081 3203 10115
rect 3145 10075 3203 10081
rect 1486 10044 1492 10056
rect 1447 10016 1492 10044
rect 1486 10004 1492 10016
rect 1544 10004 1550 10056
rect 1946 10044 1952 10056
rect 1859 10016 1952 10044
rect 1946 10004 1952 10016
rect 2004 10004 2010 10056
rect 2608 10044 2636 10075
rect 3050 10044 3056 10056
rect 2608 10040 2728 10044
rect 2792 10040 3056 10044
rect 2608 10016 3056 10040
rect 2700 10012 2820 10016
rect 3050 10004 3056 10016
rect 3108 10004 3114 10056
rect 3234 10044 3240 10056
rect 3195 10016 3240 10044
rect 3234 10004 3240 10016
rect 3292 10044 3298 10056
rect 3513 10047 3571 10053
rect 3513 10044 3525 10047
rect 3292 10016 3525 10044
rect 3292 10004 3298 10016
rect 3513 10013 3525 10016
rect 3559 10013 3571 10047
rect 3513 10007 3571 10013
rect 4525 10047 4583 10053
rect 4525 10013 4537 10047
rect 4571 10044 4583 10047
rect 5994 10044 6000 10056
rect 4571 10016 6000 10044
rect 4571 10013 4583 10016
rect 4525 10007 4583 10013
rect 5994 10004 6000 10016
rect 6052 10004 6058 10056
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10044 7987 10047
rect 8110 10044 8116 10056
rect 7975 10016 8116 10044
rect 7975 10013 7987 10016
rect 7929 10007 7987 10013
rect 8110 10004 8116 10016
rect 8168 10044 8174 10056
rect 9674 10044 9680 10056
rect 8168 10016 9680 10044
rect 8168 10004 8174 10016
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 10146 10047 10204 10053
rect 10146 10013 10158 10047
rect 10192 10013 10204 10047
rect 10413 10047 10471 10053
rect 10413 10044 10425 10047
rect 10146 10007 10204 10013
rect 10336 10016 10425 10044
rect 1504 9976 1532 10004
rect 4798 9985 4804 9988
rect 3973 9979 4031 9985
rect 3973 9976 3985 9979
rect 1504 9948 3985 9976
rect 3973 9945 3985 9948
rect 4019 9945 4031 9979
rect 4792 9976 4804 9985
rect 4759 9948 4804 9976
rect 3973 9939 4031 9945
rect 4792 9939 4804 9948
rect 4798 9936 4804 9939
rect 4856 9936 4862 9988
rect 7190 9936 7196 9988
rect 7248 9976 7254 9988
rect 7374 9976 7380 9988
rect 7248 9948 7380 9976
rect 7248 9936 7254 9948
rect 7374 9936 7380 9948
rect 7432 9976 7438 9988
rect 7662 9979 7720 9985
rect 7662 9976 7674 9979
rect 7432 9948 7674 9976
rect 7432 9936 7438 9948
rect 7662 9945 7674 9948
rect 7708 9945 7720 9979
rect 7662 9939 7720 9945
rect 1670 9868 1676 9920
rect 1728 9908 1734 9920
rect 1765 9911 1823 9917
rect 1765 9908 1777 9911
rect 1728 9880 1777 9908
rect 1728 9868 1734 9880
rect 1765 9877 1777 9880
rect 1811 9877 1823 9911
rect 2038 9908 2044 9920
rect 1999 9880 2044 9908
rect 1765 9871 1823 9877
rect 2038 9868 2044 9880
rect 2096 9868 2102 9920
rect 2409 9911 2467 9917
rect 2409 9877 2421 9911
rect 2455 9908 2467 9911
rect 2682 9908 2688 9920
rect 2455 9880 2688 9908
rect 2455 9877 2467 9880
rect 2409 9871 2467 9877
rect 2682 9868 2688 9880
rect 2740 9868 2746 9920
rect 3421 9911 3479 9917
rect 3421 9877 3433 9911
rect 3467 9908 3479 9911
rect 3878 9908 3884 9920
rect 3467 9880 3884 9908
rect 3467 9877 3479 9880
rect 3421 9871 3479 9877
rect 3878 9868 3884 9880
rect 3936 9868 3942 9920
rect 5902 9908 5908 9920
rect 5863 9880 5908 9908
rect 5902 9868 5908 9880
rect 5960 9868 5966 9920
rect 7466 9868 7472 9920
rect 7524 9908 7530 9920
rect 8294 9908 8300 9920
rect 7524 9880 8300 9908
rect 7524 9868 7530 9880
rect 8294 9868 8300 9880
rect 8352 9868 8358 9920
rect 9692 9908 9720 10004
rect 10152 9976 10180 10007
rect 10226 9976 10232 9988
rect 10152 9948 10232 9976
rect 10226 9936 10232 9948
rect 10284 9936 10290 9988
rect 10336 9908 10364 10016
rect 10413 10013 10425 10016
rect 10459 10013 10471 10047
rect 10413 10007 10471 10013
rect 10520 9976 10548 10220
rect 10594 10208 10600 10260
rect 10652 10248 10658 10260
rect 11425 10251 11483 10257
rect 11425 10248 11437 10251
rect 10652 10220 11437 10248
rect 10652 10208 10658 10220
rect 11425 10217 11437 10220
rect 11471 10248 11483 10251
rect 14734 10248 14740 10260
rect 11471 10220 14740 10248
rect 11471 10217 11483 10220
rect 11425 10211 11483 10217
rect 14734 10208 14740 10220
rect 14792 10208 14798 10260
rect 16390 10208 16396 10260
rect 16448 10248 16454 10260
rect 16577 10251 16635 10257
rect 16577 10248 16589 10251
rect 16448 10220 16589 10248
rect 16448 10208 16454 10220
rect 16577 10217 16589 10220
rect 16623 10217 16635 10251
rect 16577 10211 16635 10217
rect 17126 10208 17132 10260
rect 17184 10208 17190 10260
rect 17218 10208 17224 10260
rect 17276 10248 17282 10260
rect 17402 10248 17408 10260
rect 17276 10220 17408 10248
rect 17276 10208 17282 10220
rect 17402 10208 17408 10220
rect 17460 10208 17466 10260
rect 18325 10251 18383 10257
rect 18325 10217 18337 10251
rect 18371 10248 18383 10251
rect 18414 10248 18420 10260
rect 18371 10220 18420 10248
rect 18371 10217 18383 10220
rect 18325 10211 18383 10217
rect 18414 10208 18420 10220
rect 18472 10208 18478 10260
rect 17144 10180 17172 10208
rect 17144 10152 17816 10180
rect 16206 10072 16212 10124
rect 16264 10112 16270 10124
rect 16393 10115 16451 10121
rect 16393 10112 16405 10115
rect 16264 10084 16405 10112
rect 16264 10072 16270 10084
rect 16393 10081 16405 10084
rect 16439 10112 16451 10115
rect 17034 10112 17040 10124
rect 16439 10084 17040 10112
rect 16439 10081 16451 10084
rect 16393 10075 16451 10081
rect 17034 10072 17040 10084
rect 17092 10072 17098 10124
rect 17221 10115 17279 10121
rect 17221 10081 17233 10115
rect 17267 10112 17279 10115
rect 17310 10112 17316 10124
rect 17267 10084 17316 10112
rect 17267 10081 17279 10084
rect 17221 10075 17279 10081
rect 17310 10072 17316 10084
rect 17368 10072 17374 10124
rect 17402 10072 17408 10124
rect 17460 10072 17466 10124
rect 17788 10112 17816 10152
rect 17788 10084 17908 10112
rect 11514 10004 11520 10056
rect 11572 10044 11578 10056
rect 11974 10044 11980 10056
rect 11572 10016 11980 10044
rect 11572 10004 11578 10016
rect 11974 10004 11980 10016
rect 12032 10044 12038 10056
rect 12805 10047 12863 10053
rect 12805 10044 12817 10047
rect 12032 10016 12817 10044
rect 12032 10004 12038 10016
rect 12805 10013 12817 10016
rect 12851 10044 12863 10047
rect 12894 10044 12900 10056
rect 12851 10016 12900 10044
rect 12851 10013 12863 10016
rect 12805 10007 12863 10013
rect 12894 10004 12900 10016
rect 12952 10004 12958 10056
rect 16942 10044 16948 10056
rect 16903 10016 16948 10044
rect 16942 10004 16948 10016
rect 17000 10004 17006 10056
rect 17420 10044 17448 10072
rect 17880 10053 17908 10084
rect 17773 10047 17831 10053
rect 17773 10044 17785 10047
rect 17420 10016 17785 10044
rect 17773 10013 17785 10016
rect 17819 10013 17831 10047
rect 17773 10007 17831 10013
rect 17865 10047 17923 10053
rect 17865 10013 17877 10047
rect 17911 10013 17923 10047
rect 17865 10007 17923 10013
rect 12560 9979 12618 9985
rect 10520 9948 12434 9976
rect 9692 9880 10364 9908
rect 12406 9908 12434 9948
rect 12560 9945 12572 9979
rect 12606 9976 12618 9979
rect 13078 9976 13084 9988
rect 12606 9948 13084 9976
rect 12606 9945 12618 9948
rect 12560 9939 12618 9945
rect 13078 9936 13084 9948
rect 13136 9936 13142 9988
rect 17126 9936 17132 9988
rect 17184 9976 17190 9988
rect 18414 9976 18420 9988
rect 17184 9948 18420 9976
rect 17184 9936 17190 9948
rect 18414 9936 18420 9948
rect 18472 9936 18478 9988
rect 16022 9908 16028 9920
rect 12406 9880 16028 9908
rect 16022 9868 16028 9880
rect 16080 9868 16086 9920
rect 17494 9868 17500 9920
rect 17552 9908 17558 9920
rect 17589 9911 17647 9917
rect 17589 9908 17601 9911
rect 17552 9880 17601 9908
rect 17552 9868 17558 9880
rect 17589 9877 17601 9880
rect 17635 9877 17647 9911
rect 17589 9871 17647 9877
rect 17954 9868 17960 9920
rect 18012 9908 18018 9920
rect 18049 9911 18107 9917
rect 18049 9908 18061 9911
rect 18012 9880 18061 9908
rect 18012 9868 18018 9880
rect 18049 9877 18061 9880
rect 18095 9877 18107 9911
rect 18049 9871 18107 9877
rect 1104 9818 18860 9840
rect 1104 9766 5398 9818
rect 5450 9766 5462 9818
rect 5514 9766 5526 9818
rect 5578 9766 5590 9818
rect 5642 9766 5654 9818
rect 5706 9766 9846 9818
rect 9898 9766 9910 9818
rect 9962 9766 9974 9818
rect 10026 9766 10038 9818
rect 10090 9766 10102 9818
rect 10154 9766 14294 9818
rect 14346 9766 14358 9818
rect 14410 9766 14422 9818
rect 14474 9766 14486 9818
rect 14538 9766 14550 9818
rect 14602 9766 18860 9818
rect 1104 9744 18860 9766
rect 1946 9664 1952 9716
rect 2004 9704 2010 9716
rect 2041 9707 2099 9713
rect 2041 9704 2053 9707
rect 2004 9676 2053 9704
rect 2004 9664 2010 9676
rect 2041 9673 2053 9676
rect 2087 9673 2099 9707
rect 3421 9707 3479 9713
rect 3421 9704 3433 9707
rect 2041 9667 2099 9673
rect 2608 9676 3433 9704
rect 2608 9636 2636 9676
rect 3421 9673 3433 9676
rect 3467 9704 3479 9707
rect 3694 9704 3700 9716
rect 3467 9676 3700 9704
rect 3467 9673 3479 9676
rect 3421 9667 3479 9673
rect 3694 9664 3700 9676
rect 3752 9664 3758 9716
rect 8496 9676 9076 9704
rect 1964 9608 2636 9636
rect 1486 9568 1492 9580
rect 1447 9540 1492 9568
rect 1486 9528 1492 9540
rect 1544 9528 1550 9580
rect 1964 9577 1992 9608
rect 2682 9596 2688 9648
rect 2740 9636 2746 9648
rect 3513 9639 3571 9645
rect 3513 9636 3525 9639
rect 2740 9608 3525 9636
rect 2740 9596 2746 9608
rect 3513 9605 3525 9608
rect 3559 9605 3571 9639
rect 3513 9599 3571 9605
rect 5568 9639 5626 9645
rect 5568 9605 5580 9639
rect 5614 9636 5626 9639
rect 6546 9636 6552 9648
rect 5614 9608 6552 9636
rect 5614 9605 5626 9608
rect 5568 9599 5626 9605
rect 6546 9596 6552 9608
rect 6604 9596 6610 9648
rect 8496 9636 8524 9676
rect 6840 9608 8524 9636
rect 1949 9571 2007 9577
rect 1949 9537 1961 9571
rect 1995 9537 2007 9571
rect 1949 9531 2007 9537
rect 2498 9528 2504 9580
rect 2556 9568 2562 9580
rect 2593 9571 2651 9577
rect 2593 9568 2605 9571
rect 2556 9540 2605 9568
rect 2556 9528 2562 9540
rect 2593 9537 2605 9540
rect 2639 9537 2651 9571
rect 6730 9568 6736 9580
rect 2593 9531 2651 9537
rect 2792 9540 6736 9568
rect 2314 9460 2320 9512
rect 2372 9500 2378 9512
rect 2685 9503 2743 9509
rect 2685 9500 2697 9503
rect 2372 9472 2697 9500
rect 2372 9460 2378 9472
rect 2685 9469 2697 9472
rect 2731 9469 2743 9503
rect 2685 9463 2743 9469
rect 1673 9435 1731 9441
rect 1673 9401 1685 9435
rect 1719 9432 1731 9435
rect 2792 9432 2820 9540
rect 6730 9528 6736 9540
rect 6788 9528 6794 9580
rect 2869 9503 2927 9509
rect 2869 9469 2881 9503
rect 2915 9469 2927 9503
rect 2869 9463 2927 9469
rect 1719 9404 2820 9432
rect 2884 9432 2912 9463
rect 2958 9460 2964 9512
rect 3016 9500 3022 9512
rect 3053 9503 3111 9509
rect 3053 9500 3065 9503
rect 3016 9472 3065 9500
rect 3016 9460 3022 9472
rect 3053 9469 3065 9472
rect 3099 9469 3111 9503
rect 3053 9463 3111 9469
rect 5813 9503 5871 9509
rect 5813 9469 5825 9503
rect 5859 9500 5871 9503
rect 5994 9500 6000 9512
rect 5859 9472 6000 9500
rect 5859 9469 5871 9472
rect 5813 9463 5871 9469
rect 5994 9460 6000 9472
rect 6052 9460 6058 9512
rect 4433 9435 4491 9441
rect 2884 9404 3004 9432
rect 1719 9401 1731 9404
rect 1673 9395 1731 9401
rect 1762 9364 1768 9376
rect 1723 9336 1768 9364
rect 1762 9324 1768 9336
rect 1820 9324 1826 9376
rect 2222 9364 2228 9376
rect 2183 9336 2228 9364
rect 2222 9324 2228 9336
rect 2280 9324 2286 9376
rect 2774 9324 2780 9376
rect 2832 9364 2838 9376
rect 2976 9364 3004 9404
rect 4433 9401 4445 9435
rect 4479 9432 4491 9435
rect 4522 9432 4528 9444
rect 4479 9404 4528 9432
rect 4479 9401 4491 9404
rect 4433 9395 4491 9401
rect 4522 9392 4528 9404
rect 4580 9392 4586 9444
rect 4614 9364 4620 9376
rect 2832 9336 4620 9364
rect 2832 9324 2838 9336
rect 4614 9324 4620 9336
rect 4672 9324 4678 9376
rect 5074 9324 5080 9376
rect 5132 9364 5138 9376
rect 6840 9364 6868 9608
rect 7282 9568 7288 9580
rect 7243 9540 7288 9568
rect 7282 9528 7288 9540
rect 7340 9568 7346 9580
rect 8018 9568 8024 9580
rect 7340 9540 8024 9568
rect 7340 9528 7346 9540
rect 8018 9528 8024 9540
rect 8076 9568 8082 9580
rect 8389 9571 8447 9577
rect 8389 9568 8401 9571
rect 8076 9540 8401 9568
rect 8076 9528 8082 9540
rect 8389 9537 8401 9540
rect 8435 9537 8447 9571
rect 8389 9531 8447 9537
rect 8478 9528 8484 9580
rect 8536 9568 8542 9580
rect 8829 9571 8887 9577
rect 8829 9568 8841 9571
rect 8536 9540 8841 9568
rect 8536 9528 8542 9540
rect 8829 9537 8841 9540
rect 8875 9537 8887 9571
rect 9048 9568 9076 9676
rect 16942 9664 16948 9716
rect 17000 9704 17006 9716
rect 17405 9707 17463 9713
rect 17405 9704 17417 9707
rect 17000 9676 17417 9704
rect 17000 9664 17006 9676
rect 17405 9673 17417 9676
rect 17451 9704 17463 9707
rect 17451 9676 18000 9704
rect 17451 9673 17463 9676
rect 17405 9667 17463 9673
rect 13020 9639 13078 9645
rect 13020 9605 13032 9639
rect 13066 9636 13078 9639
rect 15010 9636 15016 9648
rect 13066 9608 15016 9636
rect 13066 9605 13078 9608
rect 13020 9599 13078 9605
rect 15010 9596 15016 9608
rect 15068 9596 15074 9648
rect 17126 9636 17132 9648
rect 17087 9608 17132 9636
rect 17126 9596 17132 9608
rect 17184 9596 17190 9648
rect 17972 9636 18000 9676
rect 18233 9639 18291 9645
rect 18233 9636 18245 9639
rect 17420 9608 17908 9636
rect 17972 9608 18245 9636
rect 17420 9568 17448 9608
rect 17880 9577 17908 9608
rect 18233 9605 18245 9608
rect 18279 9605 18291 9639
rect 18233 9599 18291 9605
rect 9048 9540 12020 9568
rect 8829 9531 8887 9537
rect 7374 9460 7380 9512
rect 7432 9500 7438 9512
rect 7653 9503 7711 9509
rect 7653 9500 7665 9503
rect 7432 9472 7665 9500
rect 7432 9460 7438 9472
rect 7653 9469 7665 9472
rect 7699 9500 7711 9503
rect 8110 9500 8116 9512
rect 7699 9472 8116 9500
rect 7699 9469 7711 9472
rect 7653 9463 7711 9469
rect 8110 9460 8116 9472
rect 8168 9500 8174 9512
rect 8573 9503 8631 9509
rect 8573 9500 8585 9503
rect 8168 9472 8585 9500
rect 8168 9460 8174 9472
rect 8573 9469 8585 9472
rect 8619 9469 8631 9503
rect 8573 9463 8631 9469
rect 5132 9336 6868 9364
rect 5132 9324 5138 9336
rect 8938 9324 8944 9376
rect 8996 9364 9002 9376
rect 9953 9367 10011 9373
rect 9953 9364 9965 9367
rect 8996 9336 9965 9364
rect 8996 9324 9002 9336
rect 9953 9333 9965 9336
rect 9999 9333 10011 9367
rect 11882 9364 11888 9376
rect 11843 9336 11888 9364
rect 9953 9327 10011 9333
rect 11882 9324 11888 9336
rect 11940 9324 11946 9376
rect 11992 9364 12020 9540
rect 14016 9540 17448 9568
rect 17589 9571 17647 9577
rect 13262 9500 13268 9512
rect 13223 9472 13268 9500
rect 13262 9460 13268 9472
rect 13320 9460 13326 9512
rect 14016 9364 14044 9540
rect 17589 9537 17601 9571
rect 17635 9537 17647 9571
rect 17589 9531 17647 9537
rect 17865 9571 17923 9577
rect 17865 9537 17877 9571
rect 17911 9568 17923 9571
rect 18046 9568 18052 9580
rect 17911 9540 18052 9568
rect 17911 9537 17923 9540
rect 17865 9531 17923 9537
rect 16945 9503 17003 9509
rect 16945 9469 16957 9503
rect 16991 9500 17003 9503
rect 17402 9500 17408 9512
rect 16991 9472 17408 9500
rect 16991 9469 17003 9472
rect 16945 9463 17003 9469
rect 17402 9460 17408 9472
rect 17460 9460 17466 9512
rect 17604 9500 17632 9531
rect 18046 9528 18052 9540
rect 18104 9528 18110 9580
rect 18414 9568 18420 9580
rect 18375 9540 18420 9568
rect 18414 9528 18420 9540
rect 18472 9528 18478 9580
rect 17512 9472 17632 9500
rect 14090 9392 14096 9444
rect 14148 9432 14154 9444
rect 17221 9435 17279 9441
rect 17221 9432 17233 9435
rect 14148 9404 17233 9432
rect 14148 9392 14154 9404
rect 17221 9401 17233 9404
rect 17267 9432 17279 9435
rect 17512 9432 17540 9472
rect 18230 9460 18236 9512
rect 18288 9460 18294 9512
rect 18248 9432 18276 9460
rect 17267 9404 17540 9432
rect 17604 9404 18276 9432
rect 17267 9401 17279 9404
rect 17221 9395 17279 9401
rect 11992 9336 14044 9364
rect 15378 9324 15384 9376
rect 15436 9364 15442 9376
rect 17604 9364 17632 9404
rect 15436 9336 17632 9364
rect 17773 9367 17831 9373
rect 15436 9324 15442 9336
rect 17773 9333 17785 9367
rect 17819 9364 17831 9367
rect 17862 9364 17868 9376
rect 17819 9336 17868 9364
rect 17819 9333 17831 9336
rect 17773 9327 17831 9333
rect 17862 9324 17868 9336
rect 17920 9324 17926 9376
rect 18049 9367 18107 9373
rect 18049 9333 18061 9367
rect 18095 9364 18107 9367
rect 18230 9364 18236 9376
rect 18095 9336 18236 9364
rect 18095 9333 18107 9336
rect 18049 9327 18107 9333
rect 18230 9324 18236 9336
rect 18288 9324 18294 9376
rect 1104 9274 18860 9296
rect 1104 9222 3174 9274
rect 3226 9222 3238 9274
rect 3290 9222 3302 9274
rect 3354 9222 3366 9274
rect 3418 9222 3430 9274
rect 3482 9222 7622 9274
rect 7674 9222 7686 9274
rect 7738 9222 7750 9274
rect 7802 9222 7814 9274
rect 7866 9222 7878 9274
rect 7930 9222 12070 9274
rect 12122 9222 12134 9274
rect 12186 9222 12198 9274
rect 12250 9222 12262 9274
rect 12314 9222 12326 9274
rect 12378 9222 16518 9274
rect 16570 9222 16582 9274
rect 16634 9222 16646 9274
rect 16698 9222 16710 9274
rect 16762 9222 16774 9274
rect 16826 9222 18860 9274
rect 1104 9200 18860 9222
rect 2498 9160 2504 9172
rect 2459 9132 2504 9160
rect 2498 9120 2504 9132
rect 2556 9120 2562 9172
rect 3418 9160 3424 9172
rect 3331 9132 3424 9160
rect 3418 9120 3424 9132
rect 3476 9160 3482 9172
rect 6086 9160 6092 9172
rect 3476 9132 6092 9160
rect 3476 9120 3482 9132
rect 6086 9120 6092 9132
rect 6144 9120 6150 9172
rect 6825 9163 6883 9169
rect 6825 9129 6837 9163
rect 6871 9160 6883 9163
rect 7190 9160 7196 9172
rect 6871 9132 7196 9160
rect 6871 9129 6883 9132
rect 6825 9123 6883 9129
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 8754 9160 8760 9172
rect 8715 9132 8760 9160
rect 8754 9120 8760 9132
rect 8812 9120 8818 9172
rect 10137 9163 10195 9169
rect 10137 9129 10149 9163
rect 10183 9160 10195 9163
rect 10226 9160 10232 9172
rect 10183 9132 10232 9160
rect 10183 9129 10195 9132
rect 10137 9123 10195 9129
rect 10226 9120 10232 9132
rect 10284 9120 10290 9172
rect 11977 9163 12035 9169
rect 11977 9129 11989 9163
rect 12023 9160 12035 9163
rect 12618 9160 12624 9172
rect 12023 9132 12624 9160
rect 12023 9129 12035 9132
rect 11977 9123 12035 9129
rect 12618 9120 12624 9132
rect 12676 9120 12682 9172
rect 14734 9120 14740 9172
rect 14792 9160 14798 9172
rect 15289 9163 15347 9169
rect 15289 9160 15301 9163
rect 14792 9132 15301 9160
rect 14792 9120 14798 9132
rect 15289 9129 15301 9132
rect 15335 9160 15347 9163
rect 15378 9160 15384 9172
rect 15335 9132 15384 9160
rect 15335 9129 15347 9132
rect 15289 9123 15347 9129
rect 15378 9120 15384 9132
rect 15436 9120 15442 9172
rect 17310 9160 17316 9172
rect 17271 9132 17316 9160
rect 17310 9120 17316 9132
rect 17368 9120 17374 9172
rect 18325 9163 18383 9169
rect 18325 9160 18337 9163
rect 17604 9132 18337 9160
rect 17604 9092 17632 9132
rect 18325 9129 18337 9132
rect 18371 9129 18383 9163
rect 18325 9123 18383 9129
rect 16868 9064 17632 9092
rect 17681 9095 17739 9101
rect 2406 9024 2412 9036
rect 2056 8996 2412 9024
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8956 1731 8959
rect 1854 8956 1860 8968
rect 1719 8928 1860 8956
rect 1719 8925 1731 8928
rect 1673 8919 1731 8925
rect 1854 8916 1860 8928
rect 1912 8916 1918 8968
rect 2056 8965 2084 8996
rect 2406 8984 2412 8996
rect 2464 8984 2470 9036
rect 3145 9027 3203 9033
rect 3145 8993 3157 9027
rect 3191 9024 3203 9027
rect 3234 9024 3240 9036
rect 3191 8996 3240 9024
rect 3191 8993 3203 8996
rect 3145 8987 3203 8993
rect 3234 8984 3240 8996
rect 3292 8984 3298 9036
rect 14553 9027 14611 9033
rect 14553 8993 14565 9027
rect 14599 9024 14611 9027
rect 16022 9024 16028 9036
rect 14599 8996 16028 9024
rect 14599 8993 14611 8996
rect 14553 8987 14611 8993
rect 16022 8984 16028 8996
rect 16080 8984 16086 9036
rect 2041 8959 2099 8965
rect 2041 8925 2053 8959
rect 2087 8925 2099 8959
rect 2041 8919 2099 8925
rect 2133 8959 2191 8965
rect 2133 8925 2145 8959
rect 2179 8925 2191 8959
rect 2133 8919 2191 8925
rect 2869 8959 2927 8965
rect 2869 8925 2881 8959
rect 2915 8956 2927 8959
rect 2958 8956 2964 8968
rect 2915 8928 2964 8956
rect 2915 8925 2927 8928
rect 2869 8919 2927 8925
rect 1946 8848 1952 8900
rect 2004 8888 2010 8900
rect 2148 8888 2176 8919
rect 2958 8916 2964 8928
rect 3016 8916 3022 8968
rect 3050 8916 3056 8968
rect 3108 8956 3114 8968
rect 5353 8959 5411 8965
rect 5353 8956 5365 8959
rect 3108 8928 4016 8956
rect 3108 8916 3114 8928
rect 3513 8891 3571 8897
rect 3513 8888 3525 8891
rect 2004 8860 3525 8888
rect 2004 8848 2010 8860
rect 3513 8857 3525 8860
rect 3559 8857 3571 8891
rect 3513 8851 3571 8857
rect 1486 8820 1492 8832
rect 1447 8792 1492 8820
rect 1486 8780 1492 8792
rect 1544 8780 1550 8832
rect 1578 8780 1584 8832
rect 1636 8820 1642 8832
rect 1857 8823 1915 8829
rect 1857 8820 1869 8823
rect 1636 8792 1869 8820
rect 1636 8780 1642 8792
rect 1857 8789 1869 8792
rect 1903 8789 1915 8823
rect 1857 8783 1915 8789
rect 2317 8823 2375 8829
rect 2317 8789 2329 8823
rect 2363 8820 2375 8823
rect 2406 8820 2412 8832
rect 2363 8792 2412 8820
rect 2363 8789 2375 8792
rect 2317 8783 2375 8789
rect 2406 8780 2412 8792
rect 2464 8780 2470 8832
rect 2961 8823 3019 8829
rect 2961 8789 2973 8823
rect 3007 8820 3019 8823
rect 3418 8820 3424 8832
rect 3007 8792 3424 8820
rect 3007 8789 3019 8792
rect 2961 8783 3019 8789
rect 3418 8780 3424 8792
rect 3476 8780 3482 8832
rect 3988 8829 4016 8928
rect 4448 8928 5365 8956
rect 4448 8900 4476 8928
rect 5353 8925 5365 8928
rect 5399 8956 5411 8959
rect 5445 8959 5503 8965
rect 5445 8956 5457 8959
rect 5399 8928 5457 8956
rect 5399 8925 5411 8928
rect 5353 8919 5411 8925
rect 5445 8925 5457 8928
rect 5491 8956 5503 8959
rect 5994 8956 6000 8968
rect 5491 8928 6000 8956
rect 5491 8925 5503 8928
rect 5445 8919 5503 8925
rect 5994 8916 6000 8928
rect 6052 8956 6058 8968
rect 7374 8956 7380 8968
rect 6052 8928 7380 8956
rect 6052 8916 6058 8928
rect 7374 8916 7380 8928
rect 7432 8956 7438 8968
rect 7432 8928 7788 8956
rect 7432 8916 7438 8928
rect 7760 8900 7788 8928
rect 8938 8916 8944 8968
rect 8996 8956 9002 8968
rect 11250 8959 11308 8965
rect 11250 8956 11262 8959
rect 8996 8928 11262 8956
rect 8996 8916 9002 8928
rect 11250 8925 11262 8928
rect 11296 8925 11308 8959
rect 11514 8956 11520 8968
rect 11475 8928 11520 8956
rect 11250 8919 11308 8925
rect 11514 8916 11520 8928
rect 11572 8956 11578 8968
rect 11974 8956 11980 8968
rect 11572 8928 11980 8956
rect 11572 8916 11578 8928
rect 11974 8916 11980 8928
rect 12032 8916 12038 8968
rect 13262 8956 13268 8968
rect 13004 8928 13268 8956
rect 13004 8900 13032 8928
rect 13262 8916 13268 8928
rect 13320 8956 13326 8968
rect 13357 8959 13415 8965
rect 13357 8956 13369 8959
rect 13320 8928 13369 8956
rect 13320 8916 13326 8928
rect 13357 8925 13369 8928
rect 13403 8925 13415 8959
rect 13357 8919 13415 8925
rect 13906 8916 13912 8968
rect 13964 8956 13970 8968
rect 14734 8956 14740 8968
rect 13964 8928 14740 8956
rect 13964 8916 13970 8928
rect 14734 8916 14740 8928
rect 14792 8916 14798 8968
rect 15841 8959 15899 8965
rect 15841 8925 15853 8959
rect 15887 8956 15899 8959
rect 16298 8956 16304 8968
rect 15887 8928 16304 8956
rect 15887 8925 15899 8928
rect 15841 8919 15899 8925
rect 16298 8916 16304 8928
rect 16356 8956 16362 8968
rect 16868 8956 16896 9064
rect 17681 9061 17693 9095
rect 17727 9092 17739 9095
rect 18138 9092 18144 9104
rect 17727 9064 18144 9092
rect 17727 9061 17739 9064
rect 17681 9055 17739 9061
rect 18138 9052 18144 9064
rect 18196 9052 18202 9104
rect 17037 9027 17095 9033
rect 17037 8993 17049 9027
rect 17083 9024 17095 9027
rect 17083 8996 18552 9024
rect 17083 8993 17095 8996
rect 17037 8987 17095 8993
rect 18524 8968 18552 8996
rect 16356 8928 16896 8956
rect 16356 8916 16362 8928
rect 17310 8916 17316 8968
rect 17368 8956 17374 8968
rect 17497 8959 17555 8965
rect 17497 8956 17509 8959
rect 17368 8928 17509 8956
rect 17368 8916 17374 8928
rect 17497 8925 17509 8928
rect 17543 8925 17555 8959
rect 17497 8919 17555 8925
rect 17865 8959 17923 8965
rect 17865 8925 17877 8959
rect 17911 8956 17923 8959
rect 18046 8956 18052 8968
rect 17911 8928 18052 8956
rect 17911 8925 17923 8928
rect 17865 8919 17923 8925
rect 18046 8916 18052 8928
rect 18104 8916 18110 8968
rect 18233 8959 18291 8965
rect 18233 8925 18245 8959
rect 18279 8956 18291 8959
rect 18322 8956 18328 8968
rect 18279 8928 18328 8956
rect 18279 8925 18291 8928
rect 18233 8919 18291 8925
rect 4430 8848 4436 8900
rect 4488 8848 4494 8900
rect 4522 8848 4528 8900
rect 4580 8888 4586 8900
rect 5718 8897 5724 8900
rect 5086 8891 5144 8897
rect 5086 8888 5098 8891
rect 4580 8860 5098 8888
rect 4580 8848 4586 8860
rect 5086 8857 5098 8860
rect 5132 8857 5144 8891
rect 5712 8888 5724 8897
rect 5679 8860 5724 8888
rect 5086 8851 5144 8857
rect 5712 8851 5724 8860
rect 5718 8848 5724 8851
rect 5776 8848 5782 8900
rect 7190 8848 7196 8900
rect 7248 8888 7254 8900
rect 7622 8891 7680 8897
rect 7622 8888 7634 8891
rect 7248 8860 7634 8888
rect 7248 8848 7254 8860
rect 7622 8857 7634 8860
rect 7668 8857 7680 8891
rect 7622 8851 7680 8857
rect 7742 8848 7748 8900
rect 7800 8848 7806 8900
rect 12802 8888 12808 8900
rect 12406 8860 12808 8888
rect 3973 8823 4031 8829
rect 3973 8789 3985 8823
rect 4019 8820 4031 8823
rect 4062 8820 4068 8832
rect 4019 8792 4068 8820
rect 4019 8789 4031 8792
rect 3973 8783 4031 8789
rect 4062 8780 4068 8792
rect 4120 8780 4126 8832
rect 4246 8780 4252 8832
rect 4304 8820 4310 8832
rect 12406 8820 12434 8860
rect 12802 8848 12808 8860
rect 12860 8848 12866 8900
rect 12986 8848 12992 8900
rect 13044 8848 13050 8900
rect 13112 8891 13170 8897
rect 13112 8857 13124 8891
rect 13158 8888 13170 8891
rect 13446 8888 13452 8900
rect 13158 8860 13452 8888
rect 13158 8857 13170 8860
rect 13112 8851 13170 8857
rect 13446 8848 13452 8860
rect 13504 8848 13510 8900
rect 15933 8891 15991 8897
rect 15933 8857 15945 8891
rect 15979 8888 15991 8891
rect 17126 8888 17132 8900
rect 15979 8860 17132 8888
rect 15979 8857 15991 8860
rect 15933 8851 15991 8857
rect 17126 8848 17132 8860
rect 17184 8848 17190 8900
rect 17221 8891 17279 8897
rect 17221 8857 17233 8891
rect 17267 8888 17279 8891
rect 18248 8888 18276 8919
rect 18322 8916 18328 8928
rect 18380 8916 18386 8968
rect 18506 8956 18512 8968
rect 18467 8928 18512 8956
rect 18506 8916 18512 8928
rect 18564 8916 18570 8968
rect 17267 8860 18276 8888
rect 17267 8857 17279 8860
rect 17221 8851 17279 8857
rect 4304 8792 12434 8820
rect 14277 8823 14335 8829
rect 4304 8780 4310 8792
rect 14277 8789 14289 8823
rect 14323 8820 14335 8823
rect 14642 8820 14648 8832
rect 14323 8792 14648 8820
rect 14323 8789 14335 8792
rect 14277 8783 14335 8789
rect 14642 8780 14648 8792
rect 14700 8780 14706 8832
rect 15102 8820 15108 8832
rect 15063 8792 15108 8820
rect 15102 8780 15108 8792
rect 15160 8780 15166 8832
rect 15470 8820 15476 8832
rect 15431 8792 15476 8820
rect 15470 8780 15476 8792
rect 15528 8780 15534 8832
rect 16574 8780 16580 8832
rect 16632 8820 16638 8832
rect 16850 8820 16856 8832
rect 16632 8792 16856 8820
rect 16632 8780 16638 8792
rect 16850 8780 16856 8792
rect 16908 8820 16914 8832
rect 18049 8823 18107 8829
rect 18049 8820 18061 8823
rect 16908 8792 18061 8820
rect 16908 8780 16914 8792
rect 18049 8789 18061 8792
rect 18095 8789 18107 8823
rect 18049 8783 18107 8789
rect 1104 8730 18860 8752
rect 1104 8678 5398 8730
rect 5450 8678 5462 8730
rect 5514 8678 5526 8730
rect 5578 8678 5590 8730
rect 5642 8678 5654 8730
rect 5706 8678 9846 8730
rect 9898 8678 9910 8730
rect 9962 8678 9974 8730
rect 10026 8678 10038 8730
rect 10090 8678 10102 8730
rect 10154 8678 14294 8730
rect 14346 8678 14358 8730
rect 14410 8678 14422 8730
rect 14474 8678 14486 8730
rect 14538 8678 14550 8730
rect 14602 8678 18860 8730
rect 1104 8656 18860 8678
rect 2314 8616 2320 8628
rect 2275 8588 2320 8616
rect 2314 8576 2320 8588
rect 2372 8576 2378 8628
rect 8938 8616 8944 8628
rect 2424 8588 8944 8616
rect 1857 8551 1915 8557
rect 1857 8517 1869 8551
rect 1903 8548 1915 8551
rect 2222 8548 2228 8560
rect 1903 8520 2228 8548
rect 1903 8517 1915 8520
rect 1857 8511 1915 8517
rect 2222 8508 2228 8520
rect 2280 8508 2286 8560
rect 1946 8412 1952 8424
rect 1907 8384 1952 8412
rect 1946 8372 1952 8384
rect 2004 8372 2010 8424
rect 2133 8415 2191 8421
rect 2133 8381 2145 8415
rect 2179 8412 2191 8415
rect 2424 8412 2452 8588
rect 8938 8576 8944 8588
rect 8996 8576 9002 8628
rect 9214 8576 9220 8628
rect 9272 8616 9278 8628
rect 12897 8619 12955 8625
rect 9272 8588 9352 8616
rect 9272 8576 9278 8588
rect 2777 8551 2835 8557
rect 2777 8517 2789 8551
rect 2823 8548 2835 8551
rect 2958 8548 2964 8560
rect 2823 8520 2964 8548
rect 2823 8517 2835 8520
rect 2777 8511 2835 8517
rect 2958 8508 2964 8520
rect 3016 8508 3022 8560
rect 4976 8551 5034 8557
rect 4976 8517 4988 8551
rect 5022 8548 5034 8551
rect 5074 8548 5080 8560
rect 5022 8520 5080 8548
rect 5022 8517 5034 8520
rect 4976 8511 5034 8517
rect 2685 8483 2743 8489
rect 2685 8449 2697 8483
rect 2731 8449 2743 8483
rect 3510 8480 3516 8492
rect 3471 8452 3516 8480
rect 2685 8443 2743 8449
rect 2179 8384 2452 8412
rect 2179 8381 2191 8384
rect 2133 8375 2191 8381
rect 2700 8356 2728 8443
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 4991 8480 5019 8511
rect 5074 8508 5080 8520
rect 5132 8508 5138 8560
rect 5718 8508 5724 8560
rect 5776 8548 5782 8560
rect 5994 8548 6000 8560
rect 5776 8520 6000 8548
rect 5776 8508 5782 8520
rect 5994 8508 6000 8520
rect 6052 8508 6058 8560
rect 9324 8557 9352 8588
rect 12897 8585 12909 8619
rect 12943 8585 12955 8619
rect 12897 8579 12955 8585
rect 14369 8619 14427 8625
rect 14369 8585 14381 8619
rect 14415 8616 14427 8619
rect 15010 8616 15016 8628
rect 14415 8588 15016 8616
rect 14415 8585 14427 8588
rect 14369 8579 14427 8585
rect 9300 8551 9358 8557
rect 9300 8517 9312 8551
rect 9346 8517 9358 8551
rect 9300 8511 9358 8517
rect 11238 8508 11244 8560
rect 11296 8548 11302 8560
rect 11762 8551 11820 8557
rect 11762 8548 11774 8551
rect 11296 8520 11774 8548
rect 11296 8508 11302 8520
rect 11762 8517 11774 8520
rect 11808 8517 11820 8551
rect 12912 8548 12940 8579
rect 15010 8576 15016 8588
rect 15068 8576 15074 8628
rect 15749 8619 15807 8625
rect 15749 8585 15761 8619
rect 15795 8616 15807 8619
rect 16574 8616 16580 8628
rect 15795 8588 16580 8616
rect 15795 8585 15807 8588
rect 15749 8579 15807 8585
rect 16574 8576 16580 8588
rect 16632 8576 16638 8628
rect 17402 8576 17408 8628
rect 17460 8616 17466 8628
rect 17589 8619 17647 8625
rect 17589 8616 17601 8619
rect 17460 8588 17601 8616
rect 17460 8576 17466 8588
rect 17589 8585 17601 8588
rect 17635 8585 17647 8619
rect 17589 8579 17647 8585
rect 13256 8551 13314 8557
rect 13256 8548 13268 8551
rect 12912 8520 13268 8548
rect 11762 8511 11820 8517
rect 13256 8517 13268 8520
rect 13302 8548 13314 8551
rect 16022 8548 16028 8560
rect 13302 8520 16028 8548
rect 13302 8517 13314 8520
rect 13256 8511 13314 8517
rect 16022 8508 16028 8520
rect 16080 8508 16086 8560
rect 3804 8452 5019 8480
rect 2869 8415 2927 8421
rect 2869 8381 2881 8415
rect 2915 8381 2927 8415
rect 2869 8375 2927 8381
rect 1394 8304 1400 8356
rect 1452 8344 1458 8356
rect 1489 8347 1547 8353
rect 1489 8344 1501 8347
rect 1452 8316 1501 8344
rect 1452 8304 1458 8316
rect 1489 8313 1501 8316
rect 1535 8313 1547 8347
rect 1489 8307 1547 8313
rect 2682 8304 2688 8356
rect 2740 8304 2746 8356
rect 2498 8236 2504 8288
rect 2556 8276 2562 8288
rect 2884 8276 2912 8375
rect 3050 8372 3056 8424
rect 3108 8412 3114 8424
rect 3804 8421 3832 8452
rect 5258 8440 5264 8492
rect 5316 8480 5322 8492
rect 7478 8483 7536 8489
rect 7478 8480 7490 8483
rect 5316 8452 7490 8480
rect 5316 8440 5322 8452
rect 7478 8449 7490 8452
rect 7524 8449 7536 8483
rect 7742 8480 7748 8492
rect 7703 8452 7748 8480
rect 7478 8443 7536 8449
rect 7742 8440 7748 8452
rect 7800 8480 7806 8492
rect 9033 8483 9091 8489
rect 9033 8480 9045 8483
rect 7800 8452 9045 8480
rect 7800 8440 7806 8452
rect 9033 8449 9045 8452
rect 9079 8449 9091 8483
rect 12986 8480 12992 8492
rect 9033 8443 9091 8449
rect 11532 8452 12992 8480
rect 11532 8424 11560 8452
rect 12986 8440 12992 8452
rect 13044 8440 13050 8492
rect 15841 8483 15899 8489
rect 15841 8449 15853 8483
rect 15887 8480 15899 8483
rect 15930 8480 15936 8492
rect 15887 8452 15936 8480
rect 15887 8449 15899 8452
rect 15841 8443 15899 8449
rect 15930 8440 15936 8452
rect 15988 8440 15994 8492
rect 17034 8440 17040 8492
rect 17092 8480 17098 8492
rect 17405 8483 17463 8489
rect 17405 8480 17417 8483
rect 17092 8452 17417 8480
rect 17092 8440 17098 8452
rect 17405 8449 17417 8452
rect 17451 8480 17463 8483
rect 17773 8483 17831 8489
rect 17773 8480 17785 8483
rect 17451 8452 17785 8480
rect 17451 8449 17463 8452
rect 17405 8443 17463 8449
rect 17773 8449 17785 8452
rect 17819 8449 17831 8483
rect 17773 8443 17831 8449
rect 17862 8440 17868 8492
rect 17920 8480 17926 8492
rect 18230 8480 18236 8492
rect 17920 8452 17965 8480
rect 18191 8452 18236 8480
rect 17920 8440 17926 8452
rect 18230 8440 18236 8452
rect 18288 8440 18294 8492
rect 3605 8415 3663 8421
rect 3605 8412 3617 8415
rect 3108 8384 3617 8412
rect 3108 8372 3114 8384
rect 3605 8381 3617 8384
rect 3651 8381 3663 8415
rect 3605 8375 3663 8381
rect 3789 8415 3847 8421
rect 3789 8381 3801 8415
rect 3835 8381 3847 8415
rect 3789 8375 3847 8381
rect 3234 8344 3240 8356
rect 3068 8316 3240 8344
rect 3068 8276 3096 8316
rect 3234 8304 3240 8316
rect 3292 8344 3298 8356
rect 3804 8344 3832 8375
rect 4430 8372 4436 8424
rect 4488 8412 4494 8424
rect 4709 8415 4767 8421
rect 4709 8412 4721 8415
rect 4488 8384 4721 8412
rect 4488 8372 4494 8384
rect 4709 8381 4721 8384
rect 4755 8381 4767 8415
rect 4709 8375 4767 8381
rect 10318 8372 10324 8424
rect 10376 8412 10382 8424
rect 11057 8415 11115 8421
rect 11057 8412 11069 8415
rect 10376 8384 11069 8412
rect 10376 8372 10382 8384
rect 11057 8381 11069 8384
rect 11103 8381 11115 8415
rect 11514 8412 11520 8424
rect 11475 8384 11520 8412
rect 11057 8375 11115 8381
rect 11514 8372 11520 8384
rect 11572 8372 11578 8424
rect 16022 8412 16028 8424
rect 15983 8384 16028 8412
rect 16022 8372 16028 8384
rect 16080 8372 16086 8424
rect 3292 8316 3832 8344
rect 3292 8304 3298 8316
rect 5810 8304 5816 8356
rect 5868 8344 5874 8356
rect 6365 8347 6423 8353
rect 6365 8344 6377 8347
rect 5868 8316 6377 8344
rect 5868 8304 5874 8316
rect 6365 8313 6377 8316
rect 6411 8313 6423 8347
rect 6365 8307 6423 8313
rect 10413 8347 10471 8353
rect 10413 8313 10425 8347
rect 10459 8344 10471 8347
rect 10778 8344 10784 8356
rect 10459 8316 10784 8344
rect 10459 8313 10471 8316
rect 10413 8307 10471 8313
rect 10778 8304 10784 8316
rect 10836 8304 10842 8356
rect 18046 8344 18052 8356
rect 18007 8316 18052 8344
rect 18046 8304 18052 8316
rect 18104 8304 18110 8356
rect 18414 8344 18420 8356
rect 18375 8316 18420 8344
rect 18414 8304 18420 8316
rect 18472 8304 18478 8356
rect 2556 8248 3096 8276
rect 3145 8279 3203 8285
rect 2556 8236 2562 8248
rect 3145 8245 3157 8279
rect 3191 8276 3203 8279
rect 3694 8276 3700 8288
rect 3191 8248 3700 8276
rect 3191 8245 3203 8248
rect 3145 8239 3203 8245
rect 3694 8236 3700 8248
rect 3752 8236 3758 8288
rect 4065 8279 4123 8285
rect 4065 8245 4077 8279
rect 4111 8276 4123 8279
rect 4246 8276 4252 8288
rect 4111 8248 4252 8276
rect 4111 8245 4123 8248
rect 4065 8239 4123 8245
rect 4246 8236 4252 8248
rect 4304 8236 4310 8288
rect 4614 8236 4620 8288
rect 4672 8276 4678 8288
rect 6089 8279 6147 8285
rect 6089 8276 6101 8279
rect 4672 8248 6101 8276
rect 4672 8236 4678 8248
rect 6089 8245 6101 8248
rect 6135 8276 6147 8279
rect 8478 8276 8484 8288
rect 6135 8248 8484 8276
rect 6135 8245 6147 8248
rect 6089 8239 6147 8245
rect 8478 8236 8484 8248
rect 8536 8236 8542 8288
rect 10502 8276 10508 8288
rect 10463 8248 10508 8276
rect 10502 8236 10508 8248
rect 10560 8236 10566 8288
rect 15378 8276 15384 8288
rect 15339 8248 15384 8276
rect 15378 8236 15384 8248
rect 15436 8236 15442 8288
rect 1104 8186 18860 8208
rect 1104 8134 3174 8186
rect 3226 8134 3238 8186
rect 3290 8134 3302 8186
rect 3354 8134 3366 8186
rect 3418 8134 3430 8186
rect 3482 8134 7622 8186
rect 7674 8134 7686 8186
rect 7738 8134 7750 8186
rect 7802 8134 7814 8186
rect 7866 8134 7878 8186
rect 7930 8134 12070 8186
rect 12122 8134 12134 8186
rect 12186 8134 12198 8186
rect 12250 8134 12262 8186
rect 12314 8134 12326 8186
rect 12378 8134 16518 8186
rect 16570 8134 16582 8186
rect 16634 8134 16646 8186
rect 16698 8134 16710 8186
rect 16762 8134 16774 8186
rect 16826 8134 18860 8186
rect 1104 8112 18860 8134
rect 1486 8072 1492 8084
rect 1447 8044 1492 8072
rect 1486 8032 1492 8044
rect 1544 8032 1550 8084
rect 1946 8032 1952 8084
rect 2004 8072 2010 8084
rect 2133 8075 2191 8081
rect 2133 8072 2145 8075
rect 2004 8044 2145 8072
rect 2004 8032 2010 8044
rect 2133 8041 2145 8044
rect 2179 8041 2191 8075
rect 2133 8035 2191 8041
rect 2682 8032 2688 8084
rect 2740 8072 2746 8084
rect 3237 8075 3295 8081
rect 3237 8072 3249 8075
rect 2740 8044 3249 8072
rect 2740 8032 2746 8044
rect 3237 8041 3249 8044
rect 3283 8072 3295 8075
rect 4338 8072 4344 8084
rect 3283 8044 4344 8072
rect 3283 8041 3295 8044
rect 3237 8035 3295 8041
rect 4338 8032 4344 8044
rect 4396 8072 4402 8084
rect 11606 8072 11612 8084
rect 4396 8044 11612 8072
rect 4396 8032 4402 8044
rect 11606 8032 11612 8044
rect 11664 8032 11670 8084
rect 11885 8075 11943 8081
rect 11885 8041 11897 8075
rect 11931 8072 11943 8075
rect 12342 8072 12348 8084
rect 11931 8044 12348 8072
rect 11931 8041 11943 8044
rect 11885 8035 11943 8041
rect 12342 8032 12348 8044
rect 12400 8032 12406 8084
rect 16942 8072 16948 8084
rect 16903 8044 16948 8072
rect 16942 8032 16948 8044
rect 17000 8032 17006 8084
rect 17310 8032 17316 8084
rect 17368 8072 17374 8084
rect 17678 8072 17684 8084
rect 17368 8044 17684 8072
rect 17368 8032 17374 8044
rect 17678 8032 17684 8044
rect 17736 8032 17742 8084
rect 3694 8004 3700 8016
rect 2976 7976 3700 8004
rect 2774 7936 2780 7948
rect 2735 7908 2780 7936
rect 2774 7896 2780 7908
rect 2832 7896 2838 7948
rect 1670 7868 1676 7880
rect 1631 7840 1676 7868
rect 1670 7828 1676 7840
rect 1728 7828 1734 7880
rect 2041 7871 2099 7877
rect 2041 7837 2053 7871
rect 2087 7868 2099 7871
rect 2314 7868 2320 7880
rect 2087 7840 2320 7868
rect 2087 7837 2099 7840
rect 2041 7831 2099 7837
rect 2314 7828 2320 7840
rect 2372 7828 2378 7880
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7868 2651 7871
rect 2976 7868 3004 7976
rect 3694 7964 3700 7976
rect 3752 7964 3758 8016
rect 17221 8007 17279 8013
rect 17221 7973 17233 8007
rect 17267 8004 17279 8007
rect 18322 8004 18328 8016
rect 17267 7976 18328 8004
rect 17267 7973 17279 7976
rect 17221 7967 17279 7973
rect 18322 7964 18328 7976
rect 18380 7964 18386 8016
rect 3053 7939 3111 7945
rect 3053 7905 3065 7939
rect 3099 7936 3111 7939
rect 3786 7936 3792 7948
rect 3099 7908 3792 7936
rect 3099 7905 3111 7908
rect 3053 7899 3111 7905
rect 2639 7840 3004 7868
rect 2639 7837 2651 7840
rect 2593 7831 2651 7837
rect 1946 7760 1952 7812
rect 2004 7800 2010 7812
rect 3068 7800 3096 7899
rect 3786 7896 3792 7908
rect 3844 7936 3850 7948
rect 3844 7908 4660 7936
rect 3844 7896 3850 7908
rect 4430 7828 4436 7880
rect 4488 7868 4494 7880
rect 4525 7871 4583 7877
rect 4525 7868 4537 7871
rect 4488 7840 4537 7868
rect 4488 7828 4494 7840
rect 4525 7837 4537 7840
rect 4571 7837 4583 7871
rect 4632 7868 4660 7908
rect 5552 7908 7052 7936
rect 5552 7868 5580 7908
rect 4632 7840 5580 7868
rect 6181 7871 6239 7877
rect 4525 7831 4583 7837
rect 6181 7837 6193 7871
rect 6227 7837 6239 7871
rect 6181 7831 6239 7837
rect 2004 7772 3096 7800
rect 2004 7760 2010 7772
rect 3786 7760 3792 7812
rect 3844 7800 3850 7812
rect 4062 7800 4068 7812
rect 3844 7772 4068 7800
rect 3844 7760 3850 7772
rect 4062 7760 4068 7772
rect 4120 7800 4126 7812
rect 4770 7803 4828 7809
rect 4770 7800 4782 7803
rect 4120 7772 4782 7800
rect 4120 7760 4126 7772
rect 4770 7769 4782 7772
rect 4816 7769 4828 7803
rect 4770 7763 4828 7769
rect 1854 7732 1860 7744
rect 1815 7704 1860 7732
rect 1854 7692 1860 7704
rect 1912 7692 1918 7744
rect 2130 7692 2136 7744
rect 2188 7732 2194 7744
rect 2501 7735 2559 7741
rect 2501 7732 2513 7735
rect 2188 7704 2513 7732
rect 2188 7692 2194 7704
rect 2501 7701 2513 7704
rect 2547 7701 2559 7735
rect 2501 7695 2559 7701
rect 5905 7735 5963 7741
rect 5905 7701 5917 7735
rect 5951 7732 5963 7735
rect 5994 7732 6000 7744
rect 5951 7704 6000 7732
rect 5951 7701 5963 7704
rect 5905 7695 5963 7701
rect 5994 7692 6000 7704
rect 6052 7692 6058 7744
rect 6196 7732 6224 7831
rect 6270 7828 6276 7880
rect 6328 7868 6334 7880
rect 6917 7871 6975 7877
rect 6917 7868 6929 7871
rect 6328 7840 6929 7868
rect 6328 7828 6334 7840
rect 6917 7837 6929 7840
rect 6963 7837 6975 7871
rect 7024 7868 7052 7908
rect 8294 7896 8300 7948
rect 8352 7936 8358 7948
rect 8941 7939 8999 7945
rect 8941 7936 8953 7939
rect 8352 7908 8953 7936
rect 8352 7896 8358 7908
rect 8941 7905 8953 7908
rect 8987 7905 8999 7939
rect 8941 7899 8999 7905
rect 8956 7868 8984 7899
rect 11514 7896 11520 7948
rect 11572 7936 11578 7948
rect 12069 7939 12127 7945
rect 12069 7936 12081 7939
rect 11572 7908 12081 7936
rect 11572 7896 11578 7908
rect 12069 7905 12081 7908
rect 12115 7905 12127 7939
rect 15010 7936 15016 7948
rect 14971 7908 15016 7936
rect 12069 7899 12127 7905
rect 15010 7896 15016 7908
rect 15068 7896 15074 7948
rect 15105 7939 15163 7945
rect 15105 7905 15117 7939
rect 15151 7936 15163 7939
rect 15378 7936 15384 7948
rect 15151 7908 15384 7936
rect 15151 7905 15163 7908
rect 15105 7899 15163 7905
rect 15378 7896 15384 7908
rect 15436 7896 15442 7948
rect 10505 7871 10563 7877
rect 10505 7868 10517 7871
rect 7024 7840 8616 7868
rect 8956 7840 10517 7868
rect 6917 7831 6975 7837
rect 6825 7803 6883 7809
rect 6825 7769 6837 7803
rect 6871 7800 6883 7803
rect 7162 7803 7220 7809
rect 7162 7800 7174 7803
rect 6871 7772 7174 7800
rect 6871 7769 6883 7772
rect 6825 7763 6883 7769
rect 7162 7769 7174 7772
rect 7208 7769 7220 7803
rect 7162 7763 7220 7769
rect 6914 7732 6920 7744
rect 6196 7704 6920 7732
rect 6914 7692 6920 7704
rect 6972 7692 6978 7744
rect 8297 7735 8355 7741
rect 8297 7701 8309 7735
rect 8343 7732 8355 7735
rect 8478 7732 8484 7744
rect 8343 7704 8484 7732
rect 8343 7701 8355 7704
rect 8297 7695 8355 7701
rect 8478 7692 8484 7704
rect 8536 7692 8542 7744
rect 8588 7732 8616 7840
rect 10505 7837 10517 7840
rect 10551 7868 10563 7871
rect 10594 7868 10600 7880
rect 10551 7840 10600 7868
rect 10551 7837 10563 7840
rect 10505 7831 10563 7837
rect 10594 7828 10600 7840
rect 10652 7828 10658 7880
rect 10778 7877 10784 7880
rect 10772 7868 10784 7877
rect 10739 7840 10784 7868
rect 10772 7831 10784 7840
rect 10778 7828 10784 7831
rect 10836 7828 10842 7880
rect 15197 7871 15255 7877
rect 12268 7840 15148 7868
rect 9214 7809 9220 7812
rect 9208 7763 9220 7809
rect 9272 7800 9278 7812
rect 10796 7800 10824 7828
rect 12268 7800 12296 7840
rect 9272 7772 9308 7800
rect 9416 7772 10732 7800
rect 10796 7772 12296 7800
rect 12336 7803 12394 7809
rect 9214 7760 9220 7763
rect 9272 7760 9278 7772
rect 9416 7732 9444 7772
rect 10318 7732 10324 7744
rect 8588 7704 9444 7732
rect 10279 7704 10324 7732
rect 10318 7692 10324 7704
rect 10376 7692 10382 7744
rect 10704 7732 10732 7772
rect 12336 7769 12348 7803
rect 12382 7800 12394 7803
rect 13262 7800 13268 7812
rect 12382 7772 13268 7800
rect 12382 7769 12394 7772
rect 12336 7763 12394 7769
rect 13262 7760 13268 7772
rect 13320 7760 13326 7812
rect 15120 7800 15148 7840
rect 15197 7837 15209 7871
rect 15243 7868 15255 7871
rect 15470 7868 15476 7880
rect 15243 7840 15476 7868
rect 15243 7837 15255 7840
rect 15197 7831 15255 7837
rect 15470 7828 15476 7840
rect 15528 7828 15534 7880
rect 16942 7828 16948 7880
rect 17000 7868 17006 7880
rect 17037 7871 17095 7877
rect 17037 7868 17049 7871
rect 17000 7840 17049 7868
rect 17000 7828 17006 7840
rect 17037 7837 17049 7840
rect 17083 7837 17095 7871
rect 17037 7831 17095 7837
rect 17497 7871 17555 7877
rect 17497 7837 17509 7871
rect 17543 7868 17555 7871
rect 17586 7868 17592 7880
rect 17543 7840 17592 7868
rect 17543 7837 17555 7840
rect 17497 7831 17555 7837
rect 17586 7828 17592 7840
rect 17644 7828 17650 7880
rect 17770 7828 17776 7880
rect 17828 7868 17834 7880
rect 18233 7871 18291 7877
rect 18233 7868 18245 7871
rect 17828 7840 18245 7868
rect 17828 7828 17834 7840
rect 18233 7837 18245 7840
rect 18279 7837 18291 7871
rect 18233 7831 18291 7837
rect 16022 7800 16028 7812
rect 15120 7772 16028 7800
rect 16022 7760 16028 7772
rect 16080 7760 16086 7812
rect 12066 7732 12072 7744
rect 10704 7704 12072 7732
rect 12066 7692 12072 7704
rect 12124 7692 12130 7744
rect 13446 7732 13452 7744
rect 13407 7704 13452 7732
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 15378 7692 15384 7744
rect 15436 7732 15442 7744
rect 15565 7735 15623 7741
rect 15565 7732 15577 7735
rect 15436 7704 15577 7732
rect 15436 7692 15442 7704
rect 15565 7701 15577 7704
rect 15611 7701 15623 7735
rect 15565 7695 15623 7701
rect 17310 7692 17316 7744
rect 17368 7732 17374 7744
rect 17589 7735 17647 7741
rect 17589 7732 17601 7735
rect 17368 7704 17601 7732
rect 17368 7692 17374 7704
rect 17589 7701 17601 7704
rect 17635 7701 17647 7735
rect 18414 7732 18420 7744
rect 18375 7704 18420 7732
rect 17589 7695 17647 7701
rect 18414 7692 18420 7704
rect 18472 7692 18478 7744
rect 1104 7642 18860 7664
rect 1104 7590 5398 7642
rect 5450 7590 5462 7642
rect 5514 7590 5526 7642
rect 5578 7590 5590 7642
rect 5642 7590 5654 7642
rect 5706 7590 9846 7642
rect 9898 7590 9910 7642
rect 9962 7590 9974 7642
rect 10026 7590 10038 7642
rect 10090 7590 10102 7642
rect 10154 7590 14294 7642
rect 14346 7590 14358 7642
rect 14410 7590 14422 7642
rect 14474 7590 14486 7642
rect 14538 7590 14550 7642
rect 14602 7590 18860 7642
rect 1104 7568 18860 7590
rect 1765 7531 1823 7537
rect 1765 7497 1777 7531
rect 1811 7528 1823 7531
rect 1946 7528 1952 7540
rect 1811 7500 1952 7528
rect 1811 7497 1823 7500
rect 1765 7491 1823 7497
rect 1946 7488 1952 7500
rect 2004 7488 2010 7540
rect 2130 7528 2136 7540
rect 2091 7500 2136 7528
rect 2130 7488 2136 7500
rect 2188 7488 2194 7540
rect 2406 7488 2412 7540
rect 2464 7528 2470 7540
rect 2501 7531 2559 7537
rect 2501 7528 2513 7531
rect 2464 7500 2513 7528
rect 2464 7488 2470 7500
rect 2501 7497 2513 7500
rect 2547 7497 2559 7531
rect 2501 7491 2559 7497
rect 2961 7531 3019 7537
rect 2961 7497 2973 7531
rect 3007 7528 3019 7531
rect 3050 7528 3056 7540
rect 3007 7500 3056 7528
rect 3007 7497 3019 7500
rect 2961 7491 3019 7497
rect 3050 7488 3056 7500
rect 3108 7488 3114 7540
rect 4982 7488 4988 7540
rect 5040 7528 5046 7540
rect 9125 7531 9183 7537
rect 5040 7500 9076 7528
rect 5040 7488 5046 7500
rect 4430 7420 4436 7472
rect 4488 7460 4494 7472
rect 7868 7463 7926 7469
rect 4488 7432 5948 7460
rect 4488 7420 4494 7432
rect 2498 7392 2504 7404
rect 1504 7364 2504 7392
rect 1504 7333 1532 7364
rect 2498 7352 2504 7364
rect 2556 7352 2562 7404
rect 2593 7395 2651 7401
rect 2593 7361 2605 7395
rect 2639 7392 2651 7395
rect 2774 7392 2780 7404
rect 2639 7364 2780 7392
rect 2639 7361 2651 7364
rect 2593 7355 2651 7361
rect 2774 7352 2780 7364
rect 2832 7352 2838 7404
rect 4177 7395 4235 7401
rect 4177 7361 4189 7395
rect 4223 7392 4235 7395
rect 5166 7392 5172 7404
rect 4223 7364 5172 7392
rect 4223 7361 4235 7364
rect 4177 7355 4235 7361
rect 5166 7352 5172 7364
rect 5224 7352 5230 7404
rect 5649 7395 5707 7401
rect 5649 7361 5661 7395
rect 5695 7392 5707 7395
rect 5810 7392 5816 7404
rect 5695 7364 5816 7392
rect 5695 7361 5707 7364
rect 5649 7355 5707 7361
rect 5810 7352 5816 7364
rect 5868 7352 5874 7404
rect 5920 7401 5948 7432
rect 7868 7429 7880 7463
rect 7914 7460 7926 7463
rect 8018 7460 8024 7472
rect 7914 7432 8024 7460
rect 7914 7429 7926 7432
rect 7868 7423 7926 7429
rect 8018 7420 8024 7432
rect 8076 7420 8082 7472
rect 9048 7460 9076 7500
rect 9125 7497 9137 7531
rect 9171 7528 9183 7531
rect 9214 7528 9220 7540
rect 9171 7500 9220 7528
rect 9171 7497 9183 7500
rect 9125 7491 9183 7497
rect 9214 7488 9220 7500
rect 9272 7488 9278 7540
rect 14093 7531 14151 7537
rect 14093 7528 14105 7531
rect 9324 7500 14105 7528
rect 9324 7460 9352 7500
rect 14093 7497 14105 7500
rect 14139 7497 14151 7531
rect 14093 7491 14151 7497
rect 14553 7531 14611 7537
rect 14553 7497 14565 7531
rect 14599 7528 14611 7531
rect 14921 7531 14979 7537
rect 14921 7528 14933 7531
rect 14599 7500 14933 7528
rect 14599 7497 14611 7500
rect 14553 7491 14611 7497
rect 14921 7497 14933 7500
rect 14967 7497 14979 7531
rect 15378 7528 15384 7540
rect 15339 7500 15384 7528
rect 14921 7491 14979 7497
rect 15378 7488 15384 7500
rect 15436 7488 15442 7540
rect 16390 7528 16396 7540
rect 16351 7500 16396 7528
rect 16390 7488 16396 7500
rect 16448 7528 16454 7540
rect 17037 7531 17095 7537
rect 17037 7528 17049 7531
rect 16448 7500 17049 7528
rect 16448 7488 16454 7500
rect 17037 7497 17049 7500
rect 17083 7497 17095 7531
rect 17037 7491 17095 7497
rect 18049 7531 18107 7537
rect 18049 7497 18061 7531
rect 18095 7497 18107 7531
rect 18049 7491 18107 7497
rect 9048 7432 9352 7460
rect 10352 7463 10410 7469
rect 10352 7429 10364 7463
rect 10398 7460 10410 7463
rect 10502 7460 10508 7472
rect 10398 7432 10508 7460
rect 10398 7429 10410 7432
rect 10352 7423 10410 7429
rect 10502 7420 10508 7432
rect 10560 7420 10566 7472
rect 12066 7420 12072 7472
rect 12124 7460 12130 7472
rect 13078 7460 13084 7472
rect 12124 7432 13084 7460
rect 12124 7420 12130 7432
rect 13078 7420 13084 7432
rect 13136 7420 13142 7472
rect 17052 7460 17080 7491
rect 17678 7460 17684 7472
rect 17052 7432 17684 7460
rect 17678 7420 17684 7432
rect 17736 7460 17742 7472
rect 17736 7432 17908 7460
rect 17736 7420 17742 7432
rect 5905 7395 5963 7401
rect 5905 7361 5917 7395
rect 5951 7392 5963 7395
rect 6178 7392 6184 7404
rect 5951 7364 6184 7392
rect 5951 7361 5963 7364
rect 5905 7355 5963 7361
rect 6178 7352 6184 7364
rect 6236 7392 6242 7404
rect 8113 7395 8171 7401
rect 8113 7392 8125 7395
rect 6236 7364 8125 7392
rect 6236 7352 6242 7364
rect 8113 7361 8125 7364
rect 8159 7392 8171 7395
rect 8294 7392 8300 7404
rect 8159 7364 8300 7392
rect 8159 7361 8171 7364
rect 8113 7355 8171 7361
rect 8294 7352 8300 7364
rect 8352 7352 8358 7404
rect 9232 7364 10548 7392
rect 1489 7327 1547 7333
rect 1489 7293 1501 7327
rect 1535 7293 1547 7327
rect 1670 7324 1676 7336
rect 1631 7296 1676 7324
rect 1489 7287 1547 7293
rect 1670 7284 1676 7296
rect 1728 7284 1734 7336
rect 2409 7327 2467 7333
rect 2409 7293 2421 7327
rect 2455 7293 2467 7327
rect 4430 7324 4436 7336
rect 4391 7296 4436 7324
rect 2409 7287 2467 7293
rect 2424 7256 2452 7287
rect 4430 7284 4436 7296
rect 4488 7284 4494 7336
rect 8478 7324 8484 7336
rect 8439 7296 8484 7324
rect 8478 7284 8484 7296
rect 8536 7284 8542 7336
rect 9232 7268 9260 7364
rect 10520 7324 10548 7364
rect 10594 7352 10600 7404
rect 10652 7392 10658 7404
rect 10652 7364 11376 7392
rect 10652 7352 10658 7364
rect 11241 7327 11299 7333
rect 11241 7324 11253 7327
rect 10520 7296 11253 7324
rect 11241 7293 11253 7296
rect 11287 7293 11299 7327
rect 11348 7324 11376 7364
rect 11882 7352 11888 7404
rect 11940 7392 11946 7404
rect 12336 7395 12394 7401
rect 12336 7392 12348 7395
rect 11940 7364 12348 7392
rect 11940 7352 11946 7364
rect 12336 7361 12348 7364
rect 12382 7392 12394 7395
rect 13630 7392 13636 7404
rect 12382 7364 13636 7392
rect 12382 7361 12394 7364
rect 12336 7355 12394 7361
rect 13630 7352 13636 7364
rect 13688 7352 13694 7404
rect 14461 7395 14519 7401
rect 14461 7361 14473 7395
rect 14507 7392 14519 7395
rect 14918 7392 14924 7404
rect 14507 7364 14924 7392
rect 14507 7361 14519 7364
rect 14461 7355 14519 7361
rect 14918 7352 14924 7364
rect 14976 7352 14982 7404
rect 15286 7392 15292 7404
rect 15247 7364 15292 7392
rect 15286 7352 15292 7364
rect 15344 7352 15350 7404
rect 17129 7395 17187 7401
rect 17129 7392 17141 7395
rect 15488 7364 17141 7392
rect 11514 7324 11520 7336
rect 11348 7296 11520 7324
rect 11241 7287 11299 7293
rect 11514 7284 11520 7296
rect 11572 7324 11578 7336
rect 11974 7324 11980 7336
rect 11572 7296 11980 7324
rect 11572 7284 11578 7296
rect 11974 7284 11980 7296
rect 12032 7324 12038 7336
rect 12069 7327 12127 7333
rect 12069 7324 12081 7327
rect 12032 7296 12081 7324
rect 12032 7284 12038 7296
rect 12069 7293 12081 7296
rect 12115 7293 12127 7327
rect 14645 7327 14703 7333
rect 14645 7324 14657 7327
rect 12069 7287 12127 7293
rect 13464 7296 14657 7324
rect 2682 7256 2688 7268
rect 2424 7228 2688 7256
rect 2682 7216 2688 7228
rect 2740 7256 2746 7268
rect 3053 7259 3111 7265
rect 3053 7256 3065 7259
rect 2740 7228 3065 7256
rect 2740 7216 2746 7228
rect 3053 7225 3065 7228
rect 3099 7225 3111 7259
rect 9214 7256 9220 7268
rect 9127 7228 9220 7256
rect 3053 7219 3111 7225
rect 9214 7216 9220 7228
rect 9272 7216 9278 7268
rect 4522 7188 4528 7200
rect 4483 7160 4528 7188
rect 4522 7148 4528 7160
rect 4580 7148 4586 7200
rect 6733 7191 6791 7197
rect 6733 7157 6745 7191
rect 6779 7188 6791 7191
rect 6914 7188 6920 7200
rect 6779 7160 6920 7188
rect 6779 7157 6791 7160
rect 6733 7151 6791 7157
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 9582 7148 9588 7200
rect 9640 7188 9646 7200
rect 10689 7191 10747 7197
rect 10689 7188 10701 7191
rect 9640 7160 10701 7188
rect 9640 7148 9646 7160
rect 10689 7157 10701 7160
rect 10735 7157 10747 7191
rect 10689 7151 10747 7157
rect 11606 7148 11612 7200
rect 11664 7188 11670 7200
rect 13464 7197 13492 7296
rect 14645 7293 14657 7296
rect 14691 7293 14703 7327
rect 14645 7287 14703 7293
rect 15194 7284 15200 7336
rect 15252 7324 15258 7336
rect 15488 7324 15516 7364
rect 17129 7361 17141 7364
rect 17175 7392 17187 7395
rect 17310 7392 17316 7404
rect 17175 7364 17316 7392
rect 17175 7361 17187 7364
rect 17129 7355 17187 7361
rect 17310 7352 17316 7364
rect 17368 7352 17374 7404
rect 17586 7392 17592 7404
rect 17547 7364 17592 7392
rect 17586 7352 17592 7364
rect 17644 7352 17650 7404
rect 17880 7401 17908 7432
rect 17865 7395 17923 7401
rect 17865 7361 17877 7395
rect 17911 7361 17923 7395
rect 18064 7392 18092 7491
rect 18233 7395 18291 7401
rect 18233 7392 18245 7395
rect 18064 7364 18245 7392
rect 17865 7355 17923 7361
rect 18233 7361 18245 7364
rect 18279 7361 18291 7395
rect 18233 7355 18291 7361
rect 15252 7296 15516 7324
rect 15565 7327 15623 7333
rect 15252 7284 15258 7296
rect 15565 7293 15577 7327
rect 15611 7324 15623 7327
rect 15746 7324 15752 7336
rect 15611 7296 15752 7324
rect 15611 7293 15623 7296
rect 15565 7287 15623 7293
rect 13630 7216 13636 7268
rect 13688 7256 13694 7268
rect 15580 7256 15608 7287
rect 15746 7284 15752 7296
rect 15804 7284 15810 7336
rect 17218 7284 17224 7336
rect 17276 7324 17282 7336
rect 17276 7296 17321 7324
rect 17276 7284 17282 7296
rect 13688 7228 15608 7256
rect 13688 7216 13694 7228
rect 16206 7216 16212 7268
rect 16264 7256 16270 7268
rect 16669 7259 16727 7265
rect 16669 7256 16681 7259
rect 16264 7228 16681 7256
rect 16264 7216 16270 7228
rect 16669 7225 16681 7228
rect 16715 7225 16727 7259
rect 16669 7219 16727 7225
rect 13449 7191 13507 7197
rect 13449 7188 13461 7191
rect 11664 7160 13461 7188
rect 11664 7148 11670 7160
rect 13449 7157 13461 7160
rect 13495 7157 13507 7191
rect 13449 7151 13507 7157
rect 17773 7191 17831 7197
rect 17773 7157 17785 7191
rect 17819 7188 17831 7191
rect 18230 7188 18236 7200
rect 17819 7160 18236 7188
rect 17819 7157 17831 7160
rect 17773 7151 17831 7157
rect 18230 7148 18236 7160
rect 18288 7148 18294 7200
rect 18414 7188 18420 7200
rect 18375 7160 18420 7188
rect 18414 7148 18420 7160
rect 18472 7148 18478 7200
rect 1104 7098 18860 7120
rect 1104 7046 3174 7098
rect 3226 7046 3238 7098
rect 3290 7046 3302 7098
rect 3354 7046 3366 7098
rect 3418 7046 3430 7098
rect 3482 7046 7622 7098
rect 7674 7046 7686 7098
rect 7738 7046 7750 7098
rect 7802 7046 7814 7098
rect 7866 7046 7878 7098
rect 7930 7046 12070 7098
rect 12122 7046 12134 7098
rect 12186 7046 12198 7098
rect 12250 7046 12262 7098
rect 12314 7046 12326 7098
rect 12378 7046 16518 7098
rect 16570 7046 16582 7098
rect 16634 7046 16646 7098
rect 16698 7046 16710 7098
rect 16762 7046 16774 7098
rect 16826 7046 18860 7098
rect 1104 7024 18860 7046
rect 1486 6984 1492 6996
rect 1447 6956 1492 6984
rect 1486 6944 1492 6956
rect 1544 6944 1550 6996
rect 1670 6944 1676 6996
rect 1728 6984 1734 6996
rect 1949 6987 2007 6993
rect 1949 6984 1961 6987
rect 1728 6956 1961 6984
rect 1728 6944 1734 6956
rect 1949 6953 1961 6956
rect 1995 6953 2007 6987
rect 3510 6984 3516 6996
rect 1949 6947 2007 6953
rect 2332 6956 3004 6984
rect 3471 6956 3516 6984
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 2332 6780 2360 6956
rect 2406 6876 2412 6928
rect 2464 6916 2470 6928
rect 2866 6916 2872 6928
rect 2464 6888 2872 6916
rect 2464 6876 2470 6888
rect 2866 6876 2872 6888
rect 2924 6876 2930 6928
rect 2976 6916 3004 6956
rect 3510 6944 3516 6956
rect 3568 6944 3574 6996
rect 5074 6944 5080 6996
rect 5132 6984 5138 6996
rect 5813 6987 5871 6993
rect 5813 6984 5825 6987
rect 5132 6956 5825 6984
rect 5132 6944 5138 6956
rect 5813 6953 5825 6956
rect 5859 6953 5871 6987
rect 5813 6947 5871 6953
rect 11974 6944 11980 6996
rect 12032 6984 12038 6996
rect 12032 6956 12379 6984
rect 12032 6944 12038 6956
rect 4157 6919 4215 6925
rect 4157 6916 4169 6919
rect 2976 6888 4169 6916
rect 4157 6885 4169 6888
rect 4203 6885 4215 6919
rect 4157 6879 4215 6885
rect 12351 6916 12379 6956
rect 15286 6944 15292 6996
rect 15344 6984 15350 6996
rect 15381 6987 15439 6993
rect 15381 6984 15393 6987
rect 15344 6956 15393 6984
rect 15344 6944 15350 6956
rect 15381 6953 15393 6956
rect 15427 6953 15439 6987
rect 17678 6984 17684 6996
rect 17639 6956 17684 6984
rect 15381 6947 15439 6953
rect 17678 6944 17684 6956
rect 17736 6944 17742 6996
rect 17770 6944 17776 6996
rect 17828 6944 17834 6996
rect 15010 6916 15016 6928
rect 12351 6888 12480 6916
rect 2593 6851 2651 6857
rect 2593 6817 2605 6851
rect 2639 6848 2651 6851
rect 2682 6848 2688 6860
rect 2639 6820 2688 6848
rect 2639 6817 2651 6820
rect 2593 6811 2651 6817
rect 2682 6808 2688 6820
rect 2740 6848 2746 6860
rect 2961 6851 3019 6857
rect 2961 6848 2973 6851
rect 2740 6820 2973 6848
rect 2740 6808 2746 6820
rect 2961 6817 2973 6820
rect 3007 6848 3019 6851
rect 4430 6848 4436 6860
rect 3007 6820 4292 6848
rect 4391 6820 4436 6848
rect 3007 6817 3019 6820
rect 2961 6811 3019 6817
rect 1719 6752 2360 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 3694 6740 3700 6792
rect 3752 6780 3758 6792
rect 3789 6783 3847 6789
rect 3789 6780 3801 6783
rect 3752 6752 3801 6780
rect 3752 6740 3758 6752
rect 3789 6749 3801 6752
rect 3835 6749 3847 6783
rect 3789 6743 3847 6749
rect 2222 6672 2228 6724
rect 2280 6712 2286 6724
rect 2409 6715 2467 6721
rect 2409 6712 2421 6715
rect 2280 6684 2421 6712
rect 2280 6672 2286 6684
rect 2409 6681 2421 6684
rect 2455 6681 2467 6715
rect 4264 6712 4292 6820
rect 4430 6808 4436 6820
rect 4488 6808 4494 6860
rect 5997 6851 6055 6857
rect 5997 6817 6009 6851
rect 6043 6848 6055 6851
rect 6086 6848 6092 6860
rect 6043 6820 6092 6848
rect 6043 6817 6055 6820
rect 5997 6811 6055 6817
rect 4341 6783 4399 6789
rect 4341 6749 4353 6783
rect 4387 6780 4399 6783
rect 6012 6780 6040 6811
rect 6086 6808 6092 6820
rect 6144 6808 6150 6860
rect 12351 6857 12379 6888
rect 12345 6851 12403 6857
rect 12345 6817 12357 6851
rect 12391 6817 12403 6851
rect 12345 6811 12403 6817
rect 4387 6752 6040 6780
rect 4387 6749 4399 6752
rect 4341 6743 4399 6749
rect 8386 6740 8392 6792
rect 8444 6780 8450 6792
rect 8481 6783 8539 6789
rect 8481 6780 8493 6783
rect 8444 6752 8493 6780
rect 8444 6740 8450 6752
rect 8481 6749 8493 6752
rect 8527 6780 8539 6783
rect 9309 6783 9367 6789
rect 9309 6780 9321 6783
rect 8527 6752 9321 6780
rect 8527 6749 8539 6752
rect 8481 6743 8539 6749
rect 9309 6749 9321 6752
rect 9355 6780 9367 6783
rect 12452 6780 12480 6888
rect 14844 6888 15016 6916
rect 14844 6857 14872 6888
rect 15010 6876 15016 6888
rect 15068 6876 15074 6928
rect 14829 6851 14887 6857
rect 14829 6817 14841 6851
rect 14875 6817 14887 6851
rect 14829 6811 14887 6817
rect 14921 6851 14979 6857
rect 14921 6817 14933 6851
rect 14967 6848 14979 6851
rect 15102 6848 15108 6860
rect 14967 6820 15108 6848
rect 14967 6817 14979 6820
rect 14921 6811 14979 6817
rect 15102 6808 15108 6820
rect 15160 6808 15166 6860
rect 16206 6848 16212 6860
rect 16167 6820 16212 6848
rect 16206 6808 16212 6820
rect 16264 6808 16270 6860
rect 16301 6851 16359 6857
rect 16301 6817 16313 6851
rect 16347 6817 16359 6851
rect 16301 6811 16359 6817
rect 13817 6783 13875 6789
rect 13817 6780 13829 6783
rect 9355 6752 10272 6780
rect 9355 6749 9367 6752
rect 9309 6743 9367 6749
rect 10244 6724 10272 6752
rect 10336 6752 12204 6780
rect 12452 6752 13829 6780
rect 4678 6715 4736 6721
rect 4678 6712 4690 6715
rect 4264 6684 4690 6712
rect 2409 6675 2467 6681
rect 4678 6681 4690 6684
rect 4724 6681 4736 6715
rect 4678 6675 4736 6681
rect 6086 6672 6092 6724
rect 6144 6712 6150 6724
rect 9582 6721 9588 6724
rect 8225 6715 8283 6721
rect 8225 6712 8237 6715
rect 6144 6684 8237 6712
rect 6144 6672 6150 6684
rect 8225 6681 8237 6684
rect 8271 6712 8283 6715
rect 9576 6712 9588 6721
rect 8271 6684 8340 6712
rect 9543 6684 9588 6712
rect 8271 6681 8283 6684
rect 8225 6675 8283 6681
rect 1857 6647 1915 6653
rect 1857 6613 1869 6647
rect 1903 6644 1915 6647
rect 2314 6644 2320 6656
rect 1903 6616 2320 6644
rect 1903 6613 1915 6616
rect 1857 6607 1915 6613
rect 2314 6604 2320 6616
rect 2372 6604 2378 6656
rect 3050 6644 3056 6656
rect 3011 6616 3056 6644
rect 3050 6604 3056 6616
rect 3108 6604 3114 6656
rect 3142 6604 3148 6656
rect 3200 6644 3206 6656
rect 3970 6644 3976 6656
rect 3200 6616 3245 6644
rect 3931 6616 3976 6644
rect 3200 6604 3206 6616
rect 3970 6604 3976 6616
rect 4028 6604 4034 6656
rect 7101 6647 7159 6653
rect 7101 6613 7113 6647
rect 7147 6644 7159 6647
rect 7282 6644 7288 6656
rect 7147 6616 7288 6644
rect 7147 6613 7159 6616
rect 7101 6607 7159 6613
rect 7282 6604 7288 6616
rect 7340 6604 7346 6656
rect 8312 6644 8340 6684
rect 9576 6675 9588 6684
rect 9582 6672 9588 6675
rect 9640 6672 9646 6724
rect 10226 6672 10232 6724
rect 10284 6672 10290 6724
rect 10336 6644 10364 6752
rect 11330 6672 11336 6724
rect 11388 6712 11394 6724
rect 12078 6715 12136 6721
rect 12078 6712 12090 6715
rect 11388 6684 12090 6712
rect 11388 6672 11394 6684
rect 12078 6681 12090 6684
rect 12124 6681 12136 6715
rect 12176 6712 12204 6752
rect 13817 6749 13829 6752
rect 13863 6749 13875 6783
rect 13817 6743 13875 6749
rect 15378 6740 15384 6792
rect 15436 6780 15442 6792
rect 16316 6780 16344 6811
rect 16574 6808 16580 6860
rect 16632 6848 16638 6860
rect 17129 6851 17187 6857
rect 17129 6848 17141 6851
rect 16632 6820 17141 6848
rect 16632 6808 16638 6820
rect 17129 6817 17141 6820
rect 17175 6848 17187 6851
rect 17218 6848 17224 6860
rect 17175 6820 17224 6848
rect 17175 6817 17187 6820
rect 17129 6811 17187 6817
rect 17218 6808 17224 6820
rect 17276 6808 17282 6860
rect 17788 6848 17816 6944
rect 17328 6820 17816 6848
rect 17328 6792 17356 6820
rect 15436 6752 16344 6780
rect 17037 6783 17095 6789
rect 15436 6740 15442 6752
rect 17037 6749 17049 6783
rect 17083 6780 17095 6783
rect 17310 6780 17316 6792
rect 17083 6752 17316 6780
rect 17083 6749 17095 6752
rect 17037 6743 17095 6749
rect 17310 6740 17316 6752
rect 17368 6740 17374 6792
rect 17862 6780 17868 6792
rect 17823 6752 17868 6780
rect 17862 6740 17868 6752
rect 17920 6740 17926 6792
rect 18230 6780 18236 6792
rect 18191 6752 18236 6780
rect 18230 6740 18236 6752
rect 18288 6740 18294 6792
rect 12894 6712 12900 6724
rect 12176 6684 12900 6712
rect 12078 6675 12136 6681
rect 12894 6672 12900 6684
rect 12952 6672 12958 6724
rect 12986 6672 12992 6724
rect 13044 6712 13050 6724
rect 13550 6715 13608 6721
rect 13550 6712 13562 6715
rect 13044 6684 13562 6712
rect 13044 6672 13050 6684
rect 13550 6681 13562 6684
rect 13596 6681 13608 6715
rect 13550 6675 13608 6681
rect 16117 6715 16175 6721
rect 16117 6681 16129 6715
rect 16163 6712 16175 6715
rect 16945 6715 17003 6721
rect 16163 6684 16620 6712
rect 16163 6681 16175 6684
rect 16117 6675 16175 6681
rect 8312 6616 10364 6644
rect 10689 6647 10747 6653
rect 10689 6613 10701 6647
rect 10735 6644 10747 6647
rect 10870 6644 10876 6656
rect 10735 6616 10876 6644
rect 10735 6613 10747 6616
rect 10689 6607 10747 6613
rect 10870 6604 10876 6616
rect 10928 6604 10934 6656
rect 10962 6604 10968 6656
rect 11020 6644 11026 6656
rect 11020 6616 11065 6644
rect 11020 6604 11026 6616
rect 11514 6604 11520 6656
rect 11572 6644 11578 6656
rect 12437 6647 12495 6653
rect 12437 6644 12449 6647
rect 11572 6616 12449 6644
rect 11572 6604 11578 6616
rect 12437 6613 12449 6616
rect 12483 6613 12495 6647
rect 12437 6607 12495 6613
rect 14090 6604 14096 6656
rect 14148 6644 14154 6656
rect 14461 6647 14519 6653
rect 14461 6644 14473 6647
rect 14148 6616 14473 6644
rect 14148 6604 14154 6616
rect 14461 6613 14473 6616
rect 14507 6644 14519 6647
rect 15013 6647 15071 6653
rect 15013 6644 15025 6647
rect 14507 6616 15025 6644
rect 14507 6613 14519 6616
rect 14461 6607 14519 6613
rect 15013 6613 15025 6616
rect 15059 6613 15071 6647
rect 15746 6644 15752 6656
rect 15707 6616 15752 6644
rect 15013 6607 15071 6613
rect 15746 6604 15752 6616
rect 15804 6604 15810 6656
rect 16592 6653 16620 6684
rect 16945 6681 16957 6715
rect 16991 6712 17003 6715
rect 17405 6715 17463 6721
rect 17405 6712 17417 6715
rect 16991 6684 17417 6712
rect 16991 6681 17003 6684
rect 16945 6675 17003 6681
rect 17405 6681 17417 6684
rect 17451 6681 17463 6715
rect 17405 6675 17463 6681
rect 16577 6647 16635 6653
rect 16577 6613 16589 6647
rect 16623 6613 16635 6647
rect 18046 6644 18052 6656
rect 18007 6616 18052 6644
rect 16577 6607 16635 6613
rect 18046 6604 18052 6616
rect 18104 6604 18110 6656
rect 18414 6644 18420 6656
rect 18375 6616 18420 6644
rect 18414 6604 18420 6616
rect 18472 6604 18478 6656
rect 1104 6554 18860 6576
rect 1104 6502 5398 6554
rect 5450 6502 5462 6554
rect 5514 6502 5526 6554
rect 5578 6502 5590 6554
rect 5642 6502 5654 6554
rect 5706 6502 9846 6554
rect 9898 6502 9910 6554
rect 9962 6502 9974 6554
rect 10026 6502 10038 6554
rect 10090 6502 10102 6554
rect 10154 6502 14294 6554
rect 14346 6502 14358 6554
rect 14410 6502 14422 6554
rect 14474 6502 14486 6554
rect 14538 6502 14550 6554
rect 14602 6502 18860 6554
rect 1104 6480 18860 6502
rect 1673 6443 1731 6449
rect 1673 6409 1685 6443
rect 1719 6440 1731 6443
rect 2225 6443 2283 6449
rect 2225 6440 2237 6443
rect 1719 6412 2237 6440
rect 1719 6409 1731 6412
rect 1673 6403 1731 6409
rect 2225 6409 2237 6412
rect 2271 6409 2283 6443
rect 2225 6403 2283 6409
rect 3050 6400 3056 6452
rect 3108 6440 3114 6452
rect 3878 6440 3884 6452
rect 3108 6412 3884 6440
rect 3108 6400 3114 6412
rect 3878 6400 3884 6412
rect 3936 6400 3942 6452
rect 7006 6400 7012 6452
rect 7064 6440 7070 6452
rect 8110 6440 8116 6452
rect 7064 6412 8116 6440
rect 7064 6400 7070 6412
rect 8110 6400 8116 6412
rect 8168 6400 8174 6452
rect 11330 6440 11336 6452
rect 11291 6412 11336 6440
rect 11330 6400 11336 6412
rect 11388 6400 11394 6452
rect 13262 6440 13268 6452
rect 13223 6412 13268 6440
rect 13262 6400 13268 6412
rect 13320 6400 13326 6452
rect 14001 6443 14059 6449
rect 14001 6409 14013 6443
rect 14047 6440 14059 6443
rect 14369 6443 14427 6449
rect 14369 6440 14381 6443
rect 14047 6412 14381 6440
rect 14047 6409 14059 6412
rect 14001 6403 14059 6409
rect 14369 6409 14381 6412
rect 14415 6409 14427 6443
rect 14369 6403 14427 6409
rect 14829 6443 14887 6449
rect 14829 6409 14841 6443
rect 14875 6440 14887 6443
rect 15197 6443 15255 6449
rect 15197 6440 15209 6443
rect 14875 6412 15209 6440
rect 14875 6409 14887 6412
rect 14829 6403 14887 6409
rect 15197 6409 15209 6412
rect 15243 6409 15255 6443
rect 15197 6403 15255 6409
rect 16942 6400 16948 6452
rect 17000 6440 17006 6452
rect 17218 6440 17224 6452
rect 17000 6412 17224 6440
rect 17000 6400 17006 6412
rect 17218 6400 17224 6412
rect 17276 6400 17282 6452
rect 17310 6400 17316 6452
rect 17368 6440 17374 6452
rect 17589 6443 17647 6449
rect 17589 6440 17601 6443
rect 17368 6412 17601 6440
rect 17368 6400 17374 6412
rect 17589 6409 17601 6412
rect 17635 6409 17647 6443
rect 17589 6403 17647 6409
rect 2593 6375 2651 6381
rect 2593 6341 2605 6375
rect 2639 6372 2651 6375
rect 3510 6372 3516 6384
rect 2639 6344 3516 6372
rect 2639 6341 2651 6344
rect 2593 6335 2651 6341
rect 3510 6332 3516 6344
rect 3568 6332 3574 6384
rect 5810 6372 5816 6384
rect 3712 6344 5816 6372
rect 1765 6307 1823 6313
rect 1765 6273 1777 6307
rect 1811 6304 1823 6307
rect 2498 6304 2504 6316
rect 1811 6276 2504 6304
rect 1811 6273 1823 6276
rect 1765 6267 1823 6273
rect 2498 6264 2504 6276
rect 2556 6264 2562 6316
rect 3418 6304 3424 6316
rect 3379 6276 3424 6304
rect 3418 6264 3424 6276
rect 3476 6264 3482 6316
rect 3712 6248 3740 6344
rect 5810 6332 5816 6344
rect 5868 6332 5874 6384
rect 5902 6332 5908 6384
rect 5960 6381 5966 6384
rect 5960 6372 5972 6381
rect 9984 6375 10042 6381
rect 5960 6344 6005 6372
rect 5960 6335 5972 6344
rect 9984 6341 9996 6375
rect 10030 6372 10042 6375
rect 11606 6372 11612 6384
rect 10030 6344 11612 6372
rect 10030 6341 10042 6344
rect 9984 6335 10042 6341
rect 5960 6332 5966 6335
rect 11606 6332 11612 6344
rect 11664 6332 11670 6384
rect 12152 6375 12210 6381
rect 12152 6341 12164 6375
rect 12198 6372 12210 6375
rect 12342 6372 12348 6384
rect 12198 6344 12348 6372
rect 12198 6341 12210 6344
rect 12152 6335 12210 6341
rect 12342 6332 12348 6344
rect 12400 6332 12406 6384
rect 3878 6304 3884 6316
rect 3839 6276 3884 6304
rect 3878 6264 3884 6276
rect 3936 6264 3942 6316
rect 4157 6307 4215 6313
rect 4157 6273 4169 6307
rect 4203 6304 4215 6307
rect 5626 6304 5632 6316
rect 4203 6276 5632 6304
rect 4203 6273 4215 6276
rect 4157 6267 4215 6273
rect 5626 6264 5632 6276
rect 5684 6264 5690 6316
rect 6178 6304 6184 6316
rect 6139 6276 6184 6304
rect 6178 6264 6184 6276
rect 6236 6304 6242 6316
rect 6549 6307 6607 6313
rect 6549 6304 6561 6307
rect 6236 6276 6561 6304
rect 6236 6264 6242 6276
rect 6549 6273 6561 6276
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 6816 6307 6874 6313
rect 6816 6273 6828 6307
rect 6862 6304 6874 6307
rect 8113 6307 8171 6313
rect 8113 6304 8125 6307
rect 6862 6276 8125 6304
rect 6862 6273 6874 6276
rect 6816 6267 6874 6273
rect 8113 6273 8125 6276
rect 8159 6273 8171 6307
rect 10226 6304 10232 6316
rect 10139 6276 10232 6304
rect 8113 6267 8171 6273
rect 10226 6264 10232 6276
rect 10284 6304 10290 6316
rect 11885 6307 11943 6313
rect 11885 6304 11897 6307
rect 10284 6276 11897 6304
rect 10284 6264 10290 6276
rect 11885 6273 11897 6276
rect 11931 6273 11943 6307
rect 13280 6304 13308 6400
rect 13909 6375 13967 6381
rect 13909 6341 13921 6375
rect 13955 6372 13967 6375
rect 15746 6372 15752 6384
rect 13955 6344 15752 6372
rect 13955 6341 13967 6344
rect 13909 6335 13967 6341
rect 15746 6332 15752 6344
rect 15804 6332 15810 6384
rect 16206 6332 16212 6384
rect 16264 6372 16270 6384
rect 17773 6375 17831 6381
rect 17773 6372 17785 6375
rect 16264 6344 17785 6372
rect 16264 6332 16270 6344
rect 17604 6316 17632 6344
rect 17773 6341 17785 6344
rect 17819 6341 17831 6375
rect 17773 6335 17831 6341
rect 14737 6307 14795 6313
rect 13280 6276 14228 6304
rect 11885 6267 11943 6273
rect 1578 6236 1584 6248
rect 1539 6208 1584 6236
rect 1578 6196 1584 6208
rect 1636 6196 1642 6248
rect 2682 6236 2688 6248
rect 2643 6208 2688 6236
rect 2682 6196 2688 6208
rect 2740 6196 2746 6248
rect 2869 6239 2927 6245
rect 2869 6205 2881 6239
rect 2915 6236 2927 6239
rect 2958 6236 2964 6248
rect 2915 6208 2964 6236
rect 2915 6205 2927 6208
rect 2869 6199 2927 6205
rect 2958 6196 2964 6208
rect 3016 6196 3022 6248
rect 3326 6196 3332 6248
rect 3384 6236 3390 6248
rect 3513 6239 3571 6245
rect 3513 6236 3525 6239
rect 3384 6208 3525 6236
rect 3384 6196 3390 6208
rect 3513 6205 3525 6208
rect 3559 6205 3571 6239
rect 3513 6199 3571 6205
rect 3694 6196 3700 6248
rect 3752 6236 3758 6248
rect 8757 6239 8815 6245
rect 3752 6208 3845 6236
rect 3752 6196 3758 6208
rect 8757 6205 8769 6239
rect 8803 6236 8815 6239
rect 8803 6208 8892 6236
rect 8803 6205 8815 6208
rect 8757 6199 8815 6205
rect 2976 6168 3004 6196
rect 4522 6168 4528 6180
rect 2976 6140 4528 6168
rect 4522 6128 4528 6140
rect 4580 6128 4586 6180
rect 8864 6112 8892 6208
rect 10502 6196 10508 6248
rect 10560 6236 10566 6248
rect 10781 6239 10839 6245
rect 10781 6236 10793 6239
rect 10560 6208 10793 6236
rect 10560 6196 10566 6208
rect 10781 6205 10793 6208
rect 10827 6236 10839 6239
rect 11514 6236 11520 6248
rect 10827 6208 11520 6236
rect 10827 6205 10839 6208
rect 10781 6199 10839 6205
rect 11514 6196 11520 6208
rect 11572 6196 11578 6248
rect 13446 6196 13452 6248
rect 13504 6236 13510 6248
rect 14093 6239 14151 6245
rect 14093 6236 14105 6239
rect 13504 6208 14105 6236
rect 13504 6196 13510 6208
rect 14093 6205 14105 6208
rect 14139 6205 14151 6239
rect 14200 6236 14228 6276
rect 14737 6273 14749 6307
rect 14783 6304 14795 6307
rect 15102 6304 15108 6316
rect 14783 6276 15108 6304
rect 14783 6273 14795 6276
rect 14737 6267 14795 6273
rect 15102 6264 15108 6276
rect 15160 6264 15166 6316
rect 15565 6307 15623 6313
rect 15565 6273 15577 6307
rect 15611 6304 15623 6307
rect 16850 6304 16856 6316
rect 15611 6276 16856 6304
rect 15611 6273 15623 6276
rect 15565 6267 15623 6273
rect 16850 6264 16856 6276
rect 16908 6264 16914 6316
rect 17586 6264 17592 6316
rect 17644 6264 17650 6316
rect 18138 6264 18144 6316
rect 18196 6304 18202 6316
rect 18233 6307 18291 6313
rect 18233 6304 18245 6307
rect 18196 6276 18245 6304
rect 18196 6264 18202 6276
rect 18233 6273 18245 6276
rect 18279 6273 18291 6307
rect 18233 6267 18291 6273
rect 14921 6239 14979 6245
rect 14921 6236 14933 6239
rect 14200 6208 14933 6236
rect 14093 6199 14151 6205
rect 14921 6205 14933 6208
rect 14967 6236 14979 6239
rect 15378 6236 15384 6248
rect 14967 6208 15384 6236
rect 14967 6205 14979 6208
rect 14921 6199 14979 6205
rect 15378 6196 15384 6208
rect 15436 6196 15442 6248
rect 15470 6196 15476 6248
rect 15528 6236 15534 6248
rect 15657 6239 15715 6245
rect 15657 6236 15669 6239
rect 15528 6208 15669 6236
rect 15528 6196 15534 6208
rect 15657 6205 15669 6208
rect 15703 6205 15715 6239
rect 15657 6199 15715 6205
rect 15746 6196 15752 6248
rect 15804 6236 15810 6248
rect 16574 6236 16580 6248
rect 15804 6208 16580 6236
rect 15804 6196 15810 6208
rect 16574 6196 16580 6208
rect 16632 6196 16638 6248
rect 16669 6239 16727 6245
rect 16669 6205 16681 6239
rect 16715 6236 16727 6239
rect 16758 6236 16764 6248
rect 16715 6208 16764 6236
rect 16715 6205 16727 6208
rect 16669 6199 16727 6205
rect 16758 6196 16764 6208
rect 16816 6196 16822 6248
rect 16942 6236 16948 6248
rect 16903 6208 16948 6236
rect 16942 6196 16948 6208
rect 17000 6196 17006 6248
rect 10870 6128 10876 6180
rect 10928 6168 10934 6180
rect 11330 6168 11336 6180
rect 10928 6140 11336 6168
rect 10928 6128 10934 6140
rect 11330 6128 11336 6140
rect 11388 6128 11394 6180
rect 15930 6168 15936 6180
rect 12820 6140 15936 6168
rect 1762 6060 1768 6112
rect 1820 6100 1826 6112
rect 2133 6103 2191 6109
rect 2133 6100 2145 6103
rect 1820 6072 2145 6100
rect 1820 6060 1826 6072
rect 2133 6069 2145 6072
rect 2179 6069 2191 6103
rect 3050 6100 3056 6112
rect 3011 6072 3056 6100
rect 2133 6063 2191 6069
rect 3050 6060 3056 6072
rect 3108 6060 3114 6112
rect 3418 6060 3424 6112
rect 3476 6100 3482 6112
rect 3970 6100 3976 6112
rect 3476 6072 3976 6100
rect 3476 6060 3482 6072
rect 3970 6060 3976 6072
rect 4028 6060 4034 6112
rect 4798 6100 4804 6112
rect 4759 6072 4804 6100
rect 4798 6060 4804 6072
rect 4856 6060 4862 6112
rect 7929 6103 7987 6109
rect 7929 6069 7941 6103
rect 7975 6100 7987 6103
rect 8018 6100 8024 6112
rect 7975 6072 8024 6100
rect 7975 6069 7987 6072
rect 7929 6063 7987 6069
rect 8018 6060 8024 6072
rect 8076 6060 8082 6112
rect 8846 6100 8852 6112
rect 8807 6072 8852 6100
rect 8846 6060 8852 6072
rect 8904 6060 8910 6112
rect 9122 6060 9128 6112
rect 9180 6100 9186 6112
rect 12820 6100 12848 6140
rect 15930 6128 15936 6140
rect 15988 6128 15994 6180
rect 9180 6072 12848 6100
rect 9180 6060 9186 6072
rect 13078 6060 13084 6112
rect 13136 6100 13142 6112
rect 13541 6103 13599 6109
rect 13541 6100 13553 6103
rect 13136 6072 13553 6100
rect 13136 6060 13142 6072
rect 13541 6069 13553 6072
rect 13587 6069 13599 6103
rect 13541 6063 13599 6069
rect 13814 6060 13820 6112
rect 13872 6100 13878 6112
rect 16390 6100 16396 6112
rect 13872 6072 16396 6100
rect 13872 6060 13878 6072
rect 16390 6060 16396 6072
rect 16448 6060 16454 6112
rect 16776 6100 16804 6196
rect 18782 6168 18788 6180
rect 17972 6140 18788 6168
rect 17972 6112 18000 6140
rect 18782 6128 18788 6140
rect 18840 6128 18846 6180
rect 16942 6100 16948 6112
rect 16776 6072 16948 6100
rect 16942 6060 16948 6072
rect 17000 6060 17006 6112
rect 17954 6100 17960 6112
rect 17915 6072 17960 6100
rect 17954 6060 17960 6072
rect 18012 6060 18018 6112
rect 18414 6100 18420 6112
rect 18375 6072 18420 6100
rect 18414 6060 18420 6072
rect 18472 6060 18478 6112
rect 1104 6010 18860 6032
rect 1104 5958 3174 6010
rect 3226 5958 3238 6010
rect 3290 5958 3302 6010
rect 3354 5958 3366 6010
rect 3418 5958 3430 6010
rect 3482 5958 7622 6010
rect 7674 5958 7686 6010
rect 7738 5958 7750 6010
rect 7802 5958 7814 6010
rect 7866 5958 7878 6010
rect 7930 5958 12070 6010
rect 12122 5958 12134 6010
rect 12186 5958 12198 6010
rect 12250 5958 12262 6010
rect 12314 5958 12326 6010
rect 12378 5958 16518 6010
rect 16570 5958 16582 6010
rect 16634 5958 16646 6010
rect 16698 5958 16710 6010
rect 16762 5958 16774 6010
rect 16826 5958 18860 6010
rect 1104 5936 18860 5958
rect 2682 5856 2688 5908
rect 2740 5896 2746 5908
rect 2869 5899 2927 5905
rect 2869 5896 2881 5899
rect 2740 5868 2881 5896
rect 2740 5856 2746 5868
rect 2869 5865 2881 5868
rect 2915 5865 2927 5899
rect 2869 5859 2927 5865
rect 5905 5899 5963 5905
rect 5905 5865 5917 5899
rect 5951 5896 5963 5899
rect 6086 5896 6092 5908
rect 5951 5868 6092 5896
rect 5951 5865 5963 5868
rect 5905 5859 5963 5865
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 6178 5856 6184 5908
rect 6236 5896 6242 5908
rect 6236 5868 6281 5896
rect 6236 5856 6242 5868
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 7285 5899 7343 5905
rect 7285 5896 7297 5899
rect 6972 5868 7297 5896
rect 6972 5856 6978 5868
rect 7285 5865 7297 5868
rect 7331 5865 7343 5899
rect 9217 5899 9275 5905
rect 7285 5859 7343 5865
rect 7392 5868 8432 5896
rect 2777 5831 2835 5837
rect 2777 5797 2789 5831
rect 2823 5828 2835 5831
rect 4062 5828 4068 5840
rect 2823 5800 4068 5828
rect 2823 5797 2835 5800
rect 2777 5791 2835 5797
rect 4062 5788 4068 5800
rect 4120 5788 4126 5840
rect 5810 5788 5816 5840
rect 5868 5828 5874 5840
rect 7392 5828 7420 5868
rect 8294 5828 8300 5840
rect 5868 5800 7420 5828
rect 8255 5800 8300 5828
rect 5868 5788 5874 5800
rect 8294 5788 8300 5800
rect 8352 5788 8358 5840
rect 8404 5828 8432 5868
rect 9217 5865 9229 5899
rect 9263 5896 9275 5899
rect 10318 5896 10324 5908
rect 9263 5868 10324 5896
rect 9263 5865 9275 5868
rect 9217 5859 9275 5865
rect 10318 5856 10324 5868
rect 10376 5856 10382 5908
rect 10502 5896 10508 5908
rect 10463 5868 10508 5896
rect 10502 5856 10508 5868
rect 10560 5856 10566 5908
rect 10870 5896 10876 5908
rect 10831 5868 10876 5896
rect 10870 5856 10876 5868
rect 10928 5856 10934 5908
rect 11977 5899 12035 5905
rect 11977 5865 11989 5899
rect 12023 5896 12035 5899
rect 12986 5896 12992 5908
rect 12023 5868 12992 5896
rect 12023 5865 12035 5868
rect 11977 5859 12035 5865
rect 12986 5856 12992 5868
rect 13044 5856 13050 5908
rect 13170 5856 13176 5908
rect 13228 5896 13234 5908
rect 14182 5896 14188 5908
rect 13228 5868 14188 5896
rect 13228 5856 13234 5868
rect 14182 5856 14188 5868
rect 14240 5856 14246 5908
rect 15102 5896 15108 5908
rect 15063 5868 15108 5896
rect 15102 5856 15108 5868
rect 15160 5856 15166 5908
rect 15470 5896 15476 5908
rect 15431 5868 15476 5896
rect 15470 5856 15476 5868
rect 15528 5856 15534 5908
rect 16390 5856 16396 5908
rect 16448 5896 16454 5908
rect 17221 5899 17279 5905
rect 17221 5896 17233 5899
rect 16448 5868 17233 5896
rect 16448 5856 16454 5868
rect 17221 5865 17233 5868
rect 17267 5865 17279 5899
rect 17862 5896 17868 5908
rect 17823 5868 17868 5896
rect 17221 5859 17279 5865
rect 8404 5800 11054 5828
rect 1670 5760 1676 5772
rect 1631 5732 1676 5760
rect 1670 5720 1676 5732
rect 1728 5720 1734 5772
rect 1762 5720 1768 5772
rect 1820 5760 1826 5772
rect 1820 5732 1865 5760
rect 1820 5720 1826 5732
rect 2866 5720 2872 5772
rect 2924 5760 2930 5772
rect 3329 5763 3387 5769
rect 3329 5760 3341 5763
rect 2924 5732 3341 5760
rect 2924 5720 2930 5732
rect 3329 5729 3341 5732
rect 3375 5729 3387 5763
rect 3329 5723 3387 5729
rect 3513 5763 3571 5769
rect 3513 5729 3525 5763
rect 3559 5760 3571 5763
rect 3694 5760 3700 5772
rect 3559 5732 3700 5760
rect 3559 5729 3571 5732
rect 3513 5723 3571 5729
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5692 1915 5695
rect 2038 5692 2044 5704
rect 1903 5664 2044 5692
rect 1903 5661 1915 5664
rect 1857 5655 1915 5661
rect 2038 5652 2044 5664
rect 2096 5652 2102 5704
rect 2590 5692 2596 5704
rect 2551 5664 2596 5692
rect 2590 5652 2596 5664
rect 2648 5652 2654 5704
rect 3344 5692 3372 5723
rect 3694 5720 3700 5732
rect 3752 5720 3758 5772
rect 4430 5720 4436 5772
rect 4488 5760 4494 5772
rect 4525 5763 4583 5769
rect 4525 5760 4537 5763
rect 4488 5732 4537 5760
rect 4488 5720 4494 5732
rect 4525 5729 4537 5732
rect 4571 5729 4583 5763
rect 4525 5723 4583 5729
rect 5902 5720 5908 5772
rect 5960 5760 5966 5772
rect 6733 5763 6791 5769
rect 6733 5760 6745 5763
rect 5960 5732 6745 5760
rect 5960 5720 5966 5732
rect 6733 5729 6745 5732
rect 6779 5729 6791 5763
rect 6733 5723 6791 5729
rect 9401 5763 9459 5769
rect 9401 5729 9413 5763
rect 9447 5760 9459 5763
rect 9766 5760 9772 5772
rect 9447 5732 9772 5760
rect 9447 5729 9459 5732
rect 9401 5723 9459 5729
rect 9766 5720 9772 5732
rect 9824 5720 9830 5772
rect 11026 5760 11054 5800
rect 11139 5800 16620 5828
rect 11139 5760 11167 5800
rect 11330 5760 11336 5772
rect 10152 5732 10916 5760
rect 11026 5732 11167 5760
rect 11291 5732 11336 5760
rect 4246 5692 4252 5704
rect 3344 5664 4252 5692
rect 4246 5652 4252 5664
rect 4304 5652 4310 5704
rect 4798 5701 4804 5704
rect 4792 5692 4804 5701
rect 4759 5664 4804 5692
rect 4792 5655 4804 5664
rect 4798 5652 4804 5655
rect 4856 5652 4862 5704
rect 6546 5692 6552 5704
rect 4991 5664 6552 5692
rect 2240 5596 2636 5624
rect 2240 5565 2268 5596
rect 2608 5568 2636 5596
rect 2866 5584 2872 5636
rect 2924 5624 2930 5636
rect 3237 5627 3295 5633
rect 3237 5624 3249 5627
rect 2924 5596 3249 5624
rect 2924 5584 2930 5596
rect 3237 5593 3249 5596
rect 3283 5624 3295 5627
rect 4991 5624 5019 5664
rect 6546 5652 6552 5664
rect 6604 5652 6610 5704
rect 7561 5695 7619 5701
rect 7561 5661 7573 5695
rect 7607 5692 7619 5695
rect 8113 5695 8171 5701
rect 8113 5692 8125 5695
rect 7607 5664 8125 5692
rect 7607 5661 7619 5664
rect 7561 5655 7619 5661
rect 8113 5661 8125 5664
rect 8159 5692 8171 5695
rect 8202 5692 8208 5704
rect 8159 5664 8208 5692
rect 8159 5661 8171 5664
rect 8113 5655 8171 5661
rect 8202 5652 8208 5664
rect 8260 5652 8266 5704
rect 8294 5652 8300 5704
rect 8352 5692 8358 5704
rect 8941 5695 8999 5701
rect 8941 5692 8953 5695
rect 8352 5664 8953 5692
rect 8352 5652 8358 5664
rect 8941 5661 8953 5664
rect 8987 5692 8999 5695
rect 9493 5695 9551 5701
rect 9493 5692 9505 5695
rect 8987 5664 9505 5692
rect 8987 5661 8999 5664
rect 8941 5655 8999 5661
rect 9493 5661 9505 5664
rect 9539 5661 9551 5695
rect 9493 5655 9551 5661
rect 3283 5596 5019 5624
rect 3283 5593 3295 5596
rect 3237 5587 3295 5593
rect 6270 5584 6276 5636
rect 6328 5624 6334 5636
rect 6641 5627 6699 5633
rect 6641 5624 6653 5627
rect 6328 5596 6653 5624
rect 6328 5584 6334 5596
rect 6641 5593 6653 5596
rect 6687 5624 6699 5627
rect 9122 5624 9128 5636
rect 6687 5596 9128 5624
rect 6687 5593 6699 5596
rect 6641 5587 6699 5593
rect 9122 5584 9128 5596
rect 9180 5584 9186 5636
rect 10152 5624 10180 5732
rect 10229 5695 10287 5701
rect 10229 5661 10241 5695
rect 10275 5692 10287 5695
rect 10781 5695 10839 5701
rect 10781 5692 10793 5695
rect 10275 5664 10793 5692
rect 10275 5661 10287 5664
rect 10229 5655 10287 5661
rect 10781 5661 10793 5664
rect 10827 5661 10839 5695
rect 10888 5692 10916 5732
rect 11330 5720 11336 5732
rect 11388 5720 11394 5772
rect 11698 5720 11704 5772
rect 11756 5760 11762 5772
rect 12069 5763 12127 5769
rect 12069 5760 12081 5763
rect 11756 5732 12081 5760
rect 11756 5720 11762 5732
rect 12069 5729 12081 5732
rect 12115 5729 12127 5763
rect 12069 5723 12127 5729
rect 12434 5720 12440 5772
rect 12492 5760 12498 5772
rect 14461 5763 14519 5769
rect 14461 5760 14473 5763
rect 12492 5732 14473 5760
rect 12492 5720 12498 5732
rect 14461 5729 14473 5732
rect 14507 5760 14519 5763
rect 15746 5760 15752 5772
rect 14507 5732 15752 5760
rect 14507 5729 14519 5732
rect 14461 5723 14519 5729
rect 15746 5720 15752 5732
rect 15804 5720 15810 5772
rect 15930 5760 15936 5772
rect 15891 5732 15936 5760
rect 15930 5720 15936 5732
rect 15988 5720 15994 5772
rect 16022 5720 16028 5772
rect 16080 5760 16086 5772
rect 16298 5760 16304 5772
rect 16080 5732 16125 5760
rect 16259 5732 16304 5760
rect 16080 5720 16086 5732
rect 16298 5720 16304 5732
rect 16356 5720 16362 5772
rect 16592 5769 16620 5800
rect 16666 5788 16672 5840
rect 16724 5828 16730 5840
rect 17034 5828 17040 5840
rect 16724 5800 17040 5828
rect 16724 5788 16730 5800
rect 17034 5788 17040 5800
rect 17092 5788 17098 5840
rect 17236 5828 17264 5859
rect 17862 5856 17868 5868
rect 17920 5856 17926 5908
rect 17236 5800 18092 5828
rect 16577 5763 16635 5769
rect 16577 5729 16589 5763
rect 16623 5729 16635 5763
rect 16577 5723 16635 5729
rect 17310 5720 17316 5772
rect 17368 5760 17374 5772
rect 17405 5763 17463 5769
rect 17405 5760 17417 5763
rect 17368 5732 17417 5760
rect 17368 5720 17374 5732
rect 17405 5729 17417 5732
rect 17451 5729 17463 5763
rect 17405 5723 17463 5729
rect 11146 5692 11152 5704
rect 10888 5664 11152 5692
rect 10781 5655 10839 5661
rect 9508 5596 10180 5624
rect 2225 5559 2283 5565
rect 2225 5525 2237 5559
rect 2271 5525 2283 5559
rect 2406 5556 2412 5568
rect 2367 5528 2412 5556
rect 2225 5519 2283 5525
rect 2406 5516 2412 5528
rect 2464 5516 2470 5568
rect 2590 5516 2596 5568
rect 2648 5516 2654 5568
rect 3970 5556 3976 5568
rect 3931 5528 3976 5556
rect 3970 5516 3976 5528
rect 4028 5516 4034 5568
rect 7098 5556 7104 5568
rect 7059 5528 7104 5556
rect 7098 5516 7104 5528
rect 7156 5556 7162 5568
rect 9508 5556 9536 5596
rect 7156 5528 9536 5556
rect 7156 5516 7162 5528
rect 9674 5516 9680 5568
rect 9732 5556 9738 5568
rect 10244 5556 10272 5655
rect 11146 5652 11152 5664
rect 11204 5652 11210 5704
rect 13906 5652 13912 5704
rect 13964 5692 13970 5704
rect 13964 5664 14009 5692
rect 13964 5652 13970 5664
rect 14182 5652 14188 5704
rect 14240 5692 14246 5704
rect 14737 5695 14795 5701
rect 14737 5692 14749 5695
rect 14240 5664 14749 5692
rect 14240 5652 14246 5664
rect 14737 5661 14749 5664
rect 14783 5692 14795 5695
rect 16206 5692 16212 5704
rect 14783 5664 16212 5692
rect 14783 5661 14795 5664
rect 14737 5655 14795 5661
rect 16206 5652 16212 5664
rect 16264 5652 16270 5704
rect 16316 5692 16344 5720
rect 17034 5692 17040 5704
rect 16316 5664 17040 5692
rect 17034 5652 17040 5664
rect 17092 5652 17098 5704
rect 17420 5692 17448 5723
rect 18064 5701 18092 5800
rect 17589 5695 17647 5701
rect 17589 5692 17601 5695
rect 17420 5664 17601 5692
rect 17589 5661 17601 5664
rect 17635 5661 17647 5695
rect 17589 5655 17647 5661
rect 18049 5695 18107 5701
rect 18049 5661 18061 5695
rect 18095 5661 18107 5695
rect 18049 5655 18107 5661
rect 18233 5695 18291 5701
rect 18233 5661 18245 5695
rect 18279 5661 18291 5695
rect 18233 5655 18291 5661
rect 11330 5624 11336 5636
rect 10704 5596 11336 5624
rect 10704 5565 10732 5596
rect 11330 5584 11336 5596
rect 11388 5624 11394 5636
rect 11388 5596 11560 5624
rect 11388 5584 11394 5596
rect 9732 5528 10272 5556
rect 10689 5559 10747 5565
rect 9732 5516 9738 5528
rect 10689 5525 10701 5559
rect 10735 5525 10747 5559
rect 10689 5519 10747 5525
rect 11054 5516 11060 5568
rect 11112 5556 11118 5568
rect 11241 5559 11299 5565
rect 11241 5556 11253 5559
rect 11112 5528 11253 5556
rect 11112 5516 11118 5528
rect 11241 5525 11253 5528
rect 11287 5525 11299 5559
rect 11532 5556 11560 5596
rect 12158 5584 12164 5636
rect 12216 5624 12222 5636
rect 13725 5627 13783 5633
rect 13725 5624 13737 5627
rect 12216 5596 13737 5624
rect 12216 5584 12222 5596
rect 13725 5593 13737 5596
rect 13771 5593 13783 5627
rect 14550 5624 14556 5636
rect 13725 5587 13783 5593
rect 14108 5596 14556 5624
rect 14108 5556 14136 5596
rect 14550 5584 14556 5596
rect 14608 5584 14614 5636
rect 14645 5627 14703 5633
rect 14645 5593 14657 5627
rect 14691 5624 14703 5627
rect 15286 5624 15292 5636
rect 14691 5596 15292 5624
rect 14691 5593 14703 5596
rect 14645 5587 14703 5593
rect 15286 5584 15292 5596
rect 15344 5584 15350 5636
rect 15841 5627 15899 5633
rect 15841 5593 15853 5627
rect 15887 5624 15899 5627
rect 16942 5624 16948 5636
rect 15887 5596 16948 5624
rect 15887 5593 15899 5596
rect 15841 5587 15899 5593
rect 16942 5584 16948 5596
rect 17000 5584 17006 5636
rect 18248 5624 18276 5655
rect 17788 5596 18276 5624
rect 11532 5528 14136 5556
rect 11241 5519 11299 5525
rect 15194 5516 15200 5568
rect 15252 5556 15258 5568
rect 17788 5565 17816 5596
rect 17773 5559 17831 5565
rect 15252 5528 15297 5556
rect 15252 5516 15258 5528
rect 17773 5525 17785 5559
rect 17819 5525 17831 5559
rect 18414 5556 18420 5568
rect 18375 5528 18420 5556
rect 17773 5519 17831 5525
rect 18414 5516 18420 5528
rect 18472 5516 18478 5568
rect 1104 5466 18860 5488
rect 1104 5414 5398 5466
rect 5450 5414 5462 5466
rect 5514 5414 5526 5466
rect 5578 5414 5590 5466
rect 5642 5414 5654 5466
rect 5706 5414 9846 5466
rect 9898 5414 9910 5466
rect 9962 5414 9974 5466
rect 10026 5414 10038 5466
rect 10090 5414 10102 5466
rect 10154 5414 14294 5466
rect 14346 5414 14358 5466
rect 14410 5414 14422 5466
rect 14474 5414 14486 5466
rect 14538 5414 14550 5466
rect 14602 5414 18860 5466
rect 1104 5392 18860 5414
rect 1486 5352 1492 5364
rect 1447 5324 1492 5352
rect 1486 5312 1492 5324
rect 1544 5312 1550 5364
rect 1946 5352 1952 5364
rect 1907 5324 1952 5352
rect 1946 5312 1952 5324
rect 2004 5312 2010 5364
rect 2222 5312 2228 5364
rect 2280 5352 2286 5364
rect 2409 5355 2467 5361
rect 2409 5352 2421 5355
rect 2280 5324 2421 5352
rect 2280 5312 2286 5324
rect 2409 5321 2421 5324
rect 2455 5321 2467 5355
rect 2409 5315 2467 5321
rect 2498 5312 2504 5364
rect 2556 5352 2562 5364
rect 2593 5355 2651 5361
rect 2593 5352 2605 5355
rect 2556 5324 2605 5352
rect 2556 5312 2562 5324
rect 2593 5321 2605 5324
rect 2639 5321 2651 5355
rect 3050 5352 3056 5364
rect 3011 5324 3056 5352
rect 2593 5315 2651 5321
rect 3050 5312 3056 5324
rect 3108 5312 3114 5364
rect 3421 5355 3479 5361
rect 3421 5321 3433 5355
rect 3467 5352 3479 5355
rect 3510 5352 3516 5364
rect 3467 5324 3516 5352
rect 3467 5321 3479 5324
rect 3421 5315 3479 5321
rect 3510 5312 3516 5324
rect 3568 5312 3574 5364
rect 3878 5352 3884 5364
rect 3839 5324 3884 5352
rect 3878 5312 3884 5324
rect 3936 5312 3942 5364
rect 5629 5355 5687 5361
rect 5629 5321 5641 5355
rect 5675 5352 5687 5355
rect 5718 5352 5724 5364
rect 5675 5324 5724 5352
rect 5675 5321 5687 5324
rect 5629 5315 5687 5321
rect 5718 5312 5724 5324
rect 5776 5352 5782 5364
rect 13265 5355 13323 5361
rect 5776 5324 13124 5352
rect 5776 5312 5782 5324
rect 2682 5244 2688 5296
rect 2740 5284 2746 5296
rect 3789 5287 3847 5293
rect 3789 5284 3801 5287
rect 2740 5256 3801 5284
rect 2740 5244 2746 5256
rect 3789 5253 3801 5256
rect 3835 5284 3847 5287
rect 4154 5284 4160 5296
rect 3835 5256 4160 5284
rect 3835 5253 3847 5256
rect 3789 5247 3847 5253
rect 4154 5244 4160 5256
rect 4212 5284 4218 5296
rect 6917 5287 6975 5293
rect 4212 5256 5764 5284
rect 4212 5244 4218 5256
rect 1302 5176 1308 5228
rect 1360 5216 1366 5228
rect 1673 5219 1731 5225
rect 1673 5216 1685 5219
rect 1360 5188 1685 5216
rect 1360 5176 1366 5188
rect 1673 5185 1685 5188
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 1765 5219 1823 5225
rect 1765 5185 1777 5219
rect 1811 5216 1823 5219
rect 1854 5216 1860 5228
rect 1811 5188 1860 5216
rect 1811 5185 1823 5188
rect 1765 5179 1823 5185
rect 1854 5176 1860 5188
rect 1912 5176 1918 5228
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5216 2191 5219
rect 2406 5216 2412 5228
rect 2179 5188 2412 5216
rect 2179 5185 2191 5188
rect 2133 5179 2191 5185
rect 2406 5176 2412 5188
rect 2464 5176 2470 5228
rect 2961 5219 3019 5225
rect 2961 5185 2973 5219
rect 3007 5216 3019 5219
rect 3234 5216 3240 5228
rect 3007 5188 3240 5216
rect 3007 5185 3019 5188
rect 2961 5179 3019 5185
rect 3234 5176 3240 5188
rect 3292 5216 3298 5228
rect 4062 5216 4068 5228
rect 3292 5188 4068 5216
rect 3292 5176 3298 5188
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 4246 5216 4252 5228
rect 4207 5188 4252 5216
rect 4246 5176 4252 5188
rect 4304 5176 4310 5228
rect 4522 5216 4528 5228
rect 4483 5188 4528 5216
rect 4522 5176 4528 5188
rect 4580 5176 4586 5228
rect 5736 5225 5764 5256
rect 6917 5253 6929 5287
rect 6963 5284 6975 5287
rect 7466 5284 7472 5296
rect 6963 5256 7472 5284
rect 6963 5253 6975 5256
rect 6917 5247 6975 5253
rect 7466 5244 7472 5256
rect 7524 5244 7530 5296
rect 7745 5287 7803 5293
rect 7745 5253 7757 5287
rect 7791 5284 7803 5287
rect 7791 5256 10272 5284
rect 7791 5253 7803 5256
rect 7745 5247 7803 5253
rect 5721 5219 5779 5225
rect 5460 5188 5672 5216
rect 3050 5108 3056 5160
rect 3108 5148 3114 5160
rect 3145 5151 3203 5157
rect 3145 5148 3157 5151
rect 3108 5120 3157 5148
rect 3108 5108 3114 5120
rect 3145 5117 3157 5120
rect 3191 5117 3203 5151
rect 3145 5111 3203 5117
rect 3694 5108 3700 5160
rect 3752 5148 3758 5160
rect 3973 5151 4031 5157
rect 3973 5148 3985 5151
rect 3752 5120 3985 5148
rect 3752 5108 3758 5120
rect 3973 5117 3985 5120
rect 4019 5117 4031 5151
rect 3973 5111 4031 5117
rect 2317 5083 2375 5089
rect 2317 5049 2329 5083
rect 2363 5080 2375 5083
rect 3786 5080 3792 5092
rect 2363 5052 3792 5080
rect 2363 5049 2375 5052
rect 2317 5043 2375 5049
rect 3786 5040 3792 5052
rect 3844 5040 3850 5092
rect 2222 4972 2228 5024
rect 2280 5012 2286 5024
rect 5460 5012 5488 5188
rect 5537 5151 5595 5157
rect 5537 5117 5549 5151
rect 5583 5117 5595 5151
rect 5644 5148 5672 5188
rect 5721 5185 5733 5219
rect 5767 5216 5779 5219
rect 5810 5216 5816 5228
rect 5767 5188 5816 5216
rect 5767 5185 5779 5188
rect 5721 5179 5779 5185
rect 5810 5176 5816 5188
rect 5868 5176 5874 5228
rect 7282 5176 7288 5228
rect 7340 5216 7346 5228
rect 8202 5216 8208 5228
rect 7340 5188 7972 5216
rect 8163 5188 8208 5216
rect 7340 5176 7346 5188
rect 6457 5151 6515 5157
rect 6457 5148 6469 5151
rect 5644 5120 6469 5148
rect 5537 5111 5595 5117
rect 6457 5117 6469 5120
rect 6503 5148 6515 5151
rect 7006 5148 7012 5160
rect 6503 5120 7012 5148
rect 6503 5117 6515 5120
rect 6457 5111 6515 5117
rect 5552 5080 5580 5111
rect 7006 5108 7012 5120
rect 7064 5108 7070 5160
rect 7101 5151 7159 5157
rect 7101 5117 7113 5151
rect 7147 5117 7159 5151
rect 7101 5111 7159 5117
rect 5902 5080 5908 5092
rect 5552 5052 5908 5080
rect 5902 5040 5908 5052
rect 5960 5080 5966 5092
rect 7116 5080 7144 5111
rect 7190 5108 7196 5160
rect 7248 5148 7254 5160
rect 7944 5157 7972 5188
rect 8202 5176 8208 5188
rect 8260 5176 8266 5228
rect 9493 5219 9551 5225
rect 9493 5185 9505 5219
rect 9539 5216 9551 5219
rect 9674 5216 9680 5228
rect 9539 5188 9680 5216
rect 9539 5185 9551 5188
rect 9493 5179 9551 5185
rect 9674 5176 9680 5188
rect 9732 5176 9738 5228
rect 7837 5151 7895 5157
rect 7837 5148 7849 5151
rect 7248 5120 7849 5148
rect 7248 5108 7254 5120
rect 7837 5117 7849 5120
rect 7883 5117 7895 5151
rect 7837 5111 7895 5117
rect 7929 5151 7987 5157
rect 7929 5117 7941 5151
rect 7975 5117 7987 5151
rect 7929 5111 7987 5117
rect 5960 5052 7144 5080
rect 9033 5083 9091 5089
rect 5960 5040 5966 5052
rect 9033 5049 9045 5083
rect 9079 5080 9091 5083
rect 9398 5080 9404 5092
rect 9079 5052 9404 5080
rect 9079 5049 9091 5052
rect 9033 5043 9091 5049
rect 9398 5040 9404 5052
rect 9456 5040 9462 5092
rect 2280 4984 5488 5012
rect 2280 4972 2286 4984
rect 5810 4972 5816 5024
rect 5868 5012 5874 5024
rect 6089 5015 6147 5021
rect 6089 5012 6101 5015
rect 5868 4984 6101 5012
rect 5868 4972 5874 4984
rect 6089 4981 6101 4984
rect 6135 4981 6147 5015
rect 6089 4975 6147 4981
rect 6549 5015 6607 5021
rect 6549 4981 6561 5015
rect 6595 5012 6607 5015
rect 6730 5012 6736 5024
rect 6595 4984 6736 5012
rect 6595 4981 6607 4984
rect 6549 4975 6607 4981
rect 6730 4972 6736 4984
rect 6788 4972 6794 5024
rect 7374 5012 7380 5024
rect 7335 4984 7380 5012
rect 7374 4972 7380 4984
rect 7432 4972 7438 5024
rect 8478 5012 8484 5024
rect 8439 4984 8484 5012
rect 8478 4972 8484 4984
rect 8536 4972 8542 5024
rect 8665 5015 8723 5021
rect 8665 4981 8677 5015
rect 8711 5012 8723 5015
rect 8938 5012 8944 5024
rect 8711 4984 8944 5012
rect 8711 4981 8723 4984
rect 8665 4975 8723 4981
rect 8938 4972 8944 4984
rect 8996 4972 9002 5024
rect 9214 5012 9220 5024
rect 9175 4984 9220 5012
rect 9214 4972 9220 4984
rect 9272 4972 9278 5024
rect 10244 5012 10272 5256
rect 10870 5244 10876 5296
rect 10928 5284 10934 5296
rect 10928 5256 11652 5284
rect 10928 5244 10934 5256
rect 11238 5176 11244 5228
rect 11296 5216 11302 5228
rect 11517 5219 11575 5225
rect 11517 5216 11529 5219
rect 11296 5188 11529 5216
rect 11296 5176 11302 5188
rect 11517 5185 11529 5188
rect 11563 5185 11575 5219
rect 11624 5216 11652 5256
rect 12158 5244 12164 5296
rect 12216 5284 12222 5296
rect 12391 5287 12449 5293
rect 12391 5284 12403 5287
rect 12216 5256 12403 5284
rect 12216 5244 12222 5256
rect 12391 5253 12403 5256
rect 12437 5253 12449 5287
rect 12391 5247 12449 5253
rect 12288 5219 12346 5225
rect 12288 5216 12300 5219
rect 11624 5188 12300 5216
rect 11517 5179 11575 5185
rect 12288 5185 12300 5188
rect 12334 5185 12346 5219
rect 13096 5216 13124 5324
rect 13265 5321 13277 5355
rect 13311 5352 13323 5355
rect 13633 5355 13691 5361
rect 13633 5352 13645 5355
rect 13311 5324 13645 5352
rect 13311 5321 13323 5324
rect 13265 5315 13323 5321
rect 13633 5321 13645 5324
rect 13679 5321 13691 5355
rect 13633 5315 13691 5321
rect 13814 5312 13820 5364
rect 13872 5352 13878 5364
rect 14001 5355 14059 5361
rect 14001 5352 14013 5355
rect 13872 5324 14013 5352
rect 13872 5312 13878 5324
rect 14001 5321 14013 5324
rect 14047 5321 14059 5355
rect 14001 5315 14059 5321
rect 14461 5355 14519 5361
rect 14461 5321 14473 5355
rect 14507 5321 14519 5355
rect 14461 5315 14519 5321
rect 14829 5355 14887 5361
rect 14829 5321 14841 5355
rect 14875 5352 14887 5355
rect 15194 5352 15200 5364
rect 14875 5324 15200 5352
rect 14875 5321 14887 5324
rect 14829 5315 14887 5321
rect 13173 5287 13231 5293
rect 13173 5253 13185 5287
rect 13219 5284 13231 5287
rect 14476 5284 14504 5315
rect 15194 5312 15200 5324
rect 15252 5312 15258 5364
rect 15286 5312 15292 5364
rect 15344 5352 15350 5364
rect 16482 5352 16488 5364
rect 15344 5324 15389 5352
rect 15856 5324 16488 5352
rect 15344 5312 15350 5324
rect 13219 5256 14504 5284
rect 13219 5253 13231 5256
rect 13173 5247 13231 5253
rect 15010 5244 15016 5296
rect 15068 5284 15074 5296
rect 15746 5284 15752 5296
rect 15068 5256 15752 5284
rect 15068 5244 15074 5256
rect 15746 5244 15752 5256
rect 15804 5244 15810 5296
rect 13096 5188 13584 5216
rect 12288 5179 12346 5185
rect 11146 5108 11152 5160
rect 11204 5148 11210 5160
rect 11701 5151 11759 5157
rect 11701 5148 11713 5151
rect 11204 5120 11713 5148
rect 11204 5108 11210 5120
rect 11701 5117 11713 5120
rect 11747 5117 11759 5151
rect 12158 5148 12164 5160
rect 12119 5120 12164 5148
rect 11701 5111 11759 5117
rect 12158 5108 12164 5120
rect 12216 5108 12222 5160
rect 12894 5108 12900 5160
rect 12952 5148 12958 5160
rect 13357 5151 13415 5157
rect 13357 5148 13369 5151
rect 12952 5120 13369 5148
rect 12952 5108 12958 5120
rect 13357 5117 13369 5120
rect 13403 5117 13415 5151
rect 13357 5111 13415 5117
rect 12805 5083 12863 5089
rect 12805 5080 12817 5083
rect 12268 5052 12817 5080
rect 12268 5012 12296 5052
rect 12805 5049 12817 5052
rect 12851 5049 12863 5083
rect 13556 5080 13584 5188
rect 13998 5176 14004 5228
rect 14056 5216 14062 5228
rect 14093 5219 14151 5225
rect 14093 5216 14105 5219
rect 14056 5188 14105 5216
rect 14056 5176 14062 5188
rect 14093 5185 14105 5188
rect 14139 5216 14151 5219
rect 14274 5216 14280 5228
rect 14139 5188 14280 5216
rect 14139 5185 14151 5188
rect 14093 5179 14151 5185
rect 14274 5176 14280 5188
rect 14332 5176 14338 5228
rect 14918 5216 14924 5228
rect 14831 5188 14924 5216
rect 14918 5176 14924 5188
rect 14976 5216 14982 5228
rect 14976 5188 15240 5216
rect 14976 5176 14982 5188
rect 14185 5151 14243 5157
rect 14185 5117 14197 5151
rect 14231 5148 14243 5151
rect 15013 5151 15071 5157
rect 15013 5148 15025 5151
rect 14231 5120 15025 5148
rect 14231 5117 14243 5120
rect 14185 5111 14243 5117
rect 15013 5117 15025 5120
rect 15059 5117 15071 5151
rect 15212 5148 15240 5188
rect 15470 5176 15476 5228
rect 15528 5216 15534 5228
rect 15657 5219 15715 5225
rect 15657 5216 15669 5219
rect 15528 5188 15669 5216
rect 15528 5176 15534 5188
rect 15657 5185 15669 5188
rect 15703 5185 15715 5219
rect 15856 5216 15884 5324
rect 16482 5312 16488 5324
rect 16540 5312 16546 5364
rect 16669 5355 16727 5361
rect 16669 5321 16681 5355
rect 16715 5352 16727 5355
rect 16850 5352 16856 5364
rect 16715 5324 16856 5352
rect 16715 5321 16727 5324
rect 16669 5315 16727 5321
rect 16850 5312 16856 5324
rect 16908 5312 16914 5364
rect 17034 5352 17040 5364
rect 16995 5324 17040 5352
rect 17034 5312 17040 5324
rect 17092 5312 17098 5364
rect 15657 5179 15715 5185
rect 15764 5188 15884 5216
rect 15764 5148 15792 5188
rect 15930 5176 15936 5228
rect 15988 5216 15994 5228
rect 16117 5219 16175 5225
rect 16117 5216 16129 5219
rect 15988 5188 16129 5216
rect 15988 5176 15994 5188
rect 16117 5185 16129 5188
rect 16163 5185 16175 5219
rect 17586 5216 17592 5228
rect 17547 5188 17592 5216
rect 16117 5179 16175 5185
rect 17586 5176 17592 5188
rect 17644 5176 17650 5228
rect 17865 5219 17923 5225
rect 17865 5216 17877 5219
rect 17788 5188 17877 5216
rect 15212 5120 15792 5148
rect 15841 5151 15899 5157
rect 15013 5111 15071 5117
rect 15841 5117 15853 5151
rect 15887 5148 15899 5151
rect 16022 5148 16028 5160
rect 15887 5120 16028 5148
rect 15887 5117 15899 5120
rect 15841 5111 15899 5117
rect 13556 5052 13768 5080
rect 12805 5043 12863 5049
rect 10244 4984 12296 5012
rect 13740 5012 13768 5052
rect 13998 5040 14004 5092
rect 14056 5080 14062 5092
rect 14200 5080 14228 5111
rect 16022 5108 16028 5120
rect 16080 5108 16086 5160
rect 16850 5148 16856 5160
rect 16132 5120 16856 5148
rect 14056 5052 14228 5080
rect 14056 5040 14062 5052
rect 16132 5012 16160 5120
rect 16850 5108 16856 5120
rect 16908 5148 16914 5160
rect 17126 5148 17132 5160
rect 16908 5120 17132 5148
rect 16908 5108 16914 5120
rect 17126 5108 17132 5120
rect 17184 5108 17190 5160
rect 17221 5151 17279 5157
rect 17221 5117 17233 5151
rect 17267 5117 17279 5151
rect 17221 5111 17279 5117
rect 16206 5040 16212 5092
rect 16264 5080 16270 5092
rect 17236 5080 17264 5111
rect 17788 5089 17816 5188
rect 17865 5185 17877 5188
rect 17911 5185 17923 5219
rect 17865 5179 17923 5185
rect 18233 5219 18291 5225
rect 18233 5185 18245 5219
rect 18279 5216 18291 5219
rect 18598 5216 18604 5228
rect 18279 5188 18604 5216
rect 18279 5185 18291 5188
rect 18233 5179 18291 5185
rect 18598 5176 18604 5188
rect 18656 5176 18662 5228
rect 16264 5052 17264 5080
rect 17773 5083 17831 5089
rect 16264 5040 16270 5052
rect 17773 5049 17785 5083
rect 17819 5049 17831 5083
rect 18414 5080 18420 5092
rect 18375 5052 18420 5080
rect 17773 5043 17831 5049
rect 18414 5040 18420 5052
rect 18472 5040 18478 5092
rect 16298 5012 16304 5024
rect 13740 4984 16160 5012
rect 16259 4984 16304 5012
rect 16298 4972 16304 4984
rect 16356 4972 16362 5024
rect 18046 5012 18052 5024
rect 18007 4984 18052 5012
rect 18046 4972 18052 4984
rect 18104 4972 18110 5024
rect 1104 4922 18860 4944
rect 1104 4870 3174 4922
rect 3226 4870 3238 4922
rect 3290 4870 3302 4922
rect 3354 4870 3366 4922
rect 3418 4870 3430 4922
rect 3482 4870 7622 4922
rect 7674 4870 7686 4922
rect 7738 4870 7750 4922
rect 7802 4870 7814 4922
rect 7866 4870 7878 4922
rect 7930 4870 12070 4922
rect 12122 4870 12134 4922
rect 12186 4870 12198 4922
rect 12250 4870 12262 4922
rect 12314 4870 12326 4922
rect 12378 4870 16518 4922
rect 16570 4870 16582 4922
rect 16634 4870 16646 4922
rect 16698 4870 16710 4922
rect 16762 4870 16774 4922
rect 16826 4870 18860 4922
rect 1104 4848 18860 4870
rect 1486 4808 1492 4820
rect 1447 4780 1492 4808
rect 1486 4768 1492 4780
rect 1544 4768 1550 4820
rect 2314 4768 2320 4820
rect 2372 4808 2378 4820
rect 2774 4808 2780 4820
rect 2372 4780 2780 4808
rect 2372 4768 2378 4780
rect 2774 4768 2780 4780
rect 2832 4768 2838 4820
rect 6181 4811 6239 4817
rect 6181 4777 6193 4811
rect 6227 4808 6239 4811
rect 7190 4808 7196 4820
rect 6227 4780 7196 4808
rect 6227 4777 6239 4780
rect 6181 4771 6239 4777
rect 7190 4768 7196 4780
rect 7248 4768 7254 4820
rect 8018 4768 8024 4820
rect 8076 4808 8082 4820
rect 8389 4811 8447 4817
rect 8389 4808 8401 4811
rect 8076 4780 8401 4808
rect 8076 4768 8082 4780
rect 8389 4777 8401 4780
rect 8435 4777 8447 4811
rect 8389 4771 8447 4777
rect 10410 4768 10416 4820
rect 10468 4808 10474 4820
rect 10597 4811 10655 4817
rect 10597 4808 10609 4811
rect 10468 4780 10609 4808
rect 10468 4768 10474 4780
rect 10597 4777 10609 4780
rect 10643 4808 10655 4811
rect 10962 4808 10968 4820
rect 10643 4780 10968 4808
rect 10643 4777 10655 4780
rect 10597 4771 10655 4777
rect 10962 4768 10968 4780
rect 11020 4768 11026 4820
rect 12710 4808 12716 4820
rect 11808 4780 12716 4808
rect 2406 4700 2412 4752
rect 2464 4740 2470 4752
rect 2685 4743 2743 4749
rect 2685 4740 2697 4743
rect 2464 4712 2697 4740
rect 2464 4700 2470 4712
rect 2685 4709 2697 4712
rect 2731 4709 2743 4743
rect 2685 4703 2743 4709
rect 3605 4743 3663 4749
rect 3605 4709 3617 4743
rect 3651 4740 3663 4743
rect 11808 4740 11836 4780
rect 12710 4768 12716 4780
rect 12768 4768 12774 4820
rect 12805 4811 12863 4817
rect 12805 4777 12817 4811
rect 12851 4808 12863 4811
rect 12851 4780 17448 4808
rect 12851 4777 12863 4780
rect 12805 4771 12863 4777
rect 3651 4712 11836 4740
rect 3651 4709 3663 4712
rect 3605 4703 3663 4709
rect 1673 4607 1731 4613
rect 1673 4573 1685 4607
rect 1719 4573 1731 4607
rect 1673 4567 1731 4573
rect 2041 4607 2099 4613
rect 2041 4573 2053 4607
rect 2087 4604 2099 4607
rect 2087 4576 2268 4604
rect 2087 4573 2099 4576
rect 2041 4567 2099 4573
rect 1688 4536 1716 4567
rect 2240 4536 2268 4576
rect 2314 4564 2320 4616
rect 2372 4604 2378 4616
rect 2593 4607 2651 4613
rect 2372 4576 2417 4604
rect 2372 4564 2378 4576
rect 2593 4573 2605 4607
rect 2639 4604 2651 4607
rect 2682 4604 2688 4616
rect 2639 4576 2688 4604
rect 2639 4573 2651 4576
rect 2593 4567 2651 4573
rect 2682 4564 2688 4576
rect 2740 4564 2746 4616
rect 2866 4604 2872 4616
rect 2827 4576 2872 4604
rect 2866 4564 2872 4576
rect 2924 4564 2930 4616
rect 3145 4607 3203 4613
rect 3145 4573 3157 4607
rect 3191 4573 3203 4607
rect 3145 4567 3203 4573
rect 3421 4607 3479 4613
rect 3421 4573 3433 4607
rect 3467 4604 3479 4607
rect 3620 4604 3648 4703
rect 11882 4700 11888 4752
rect 11940 4740 11946 4752
rect 13998 4740 14004 4752
rect 11940 4712 14004 4740
rect 11940 4700 11946 4712
rect 13998 4700 14004 4712
rect 14056 4700 14062 4752
rect 14182 4700 14188 4752
rect 14240 4740 14246 4752
rect 14369 4743 14427 4749
rect 14369 4740 14381 4743
rect 14240 4712 14381 4740
rect 14240 4700 14246 4712
rect 14369 4709 14381 4712
rect 14415 4709 14427 4743
rect 14369 4703 14427 4709
rect 15657 4743 15715 4749
rect 15657 4709 15669 4743
rect 15703 4740 15715 4743
rect 16206 4740 16212 4752
rect 15703 4712 16212 4740
rect 15703 4709 15715 4712
rect 15657 4703 15715 4709
rect 16206 4700 16212 4712
rect 16264 4700 16270 4752
rect 16316 4712 17356 4740
rect 5629 4675 5687 4681
rect 5629 4641 5641 4675
rect 5675 4672 5687 4675
rect 6086 4672 6092 4684
rect 5675 4644 6092 4672
rect 5675 4641 5687 4644
rect 5629 4635 5687 4641
rect 6086 4632 6092 4644
rect 6144 4632 6150 4684
rect 6730 4672 6736 4684
rect 6691 4644 6736 4672
rect 6730 4632 6736 4644
rect 6788 4632 6794 4684
rect 6822 4632 6828 4684
rect 6880 4672 6886 4684
rect 6917 4675 6975 4681
rect 6917 4672 6929 4675
rect 6880 4644 6929 4672
rect 6880 4632 6886 4644
rect 6917 4641 6929 4644
rect 6963 4672 6975 4675
rect 6963 4644 9674 4672
rect 6963 4641 6975 4644
rect 6917 4635 6975 4641
rect 4246 4604 4252 4616
rect 3467 4576 3648 4604
rect 4159 4576 4252 4604
rect 3467 4573 3479 4576
rect 3421 4567 3479 4573
rect 3160 4536 3188 4567
rect 4246 4564 4252 4576
rect 4304 4604 4310 4616
rect 6638 4604 6644 4616
rect 4304 4576 6408 4604
rect 6599 4576 6644 4604
rect 4304 4564 4310 4576
rect 3786 4536 3792 4548
rect 1688 4508 2176 4536
rect 2240 4508 2774 4536
rect 3160 4508 3792 4536
rect 1854 4468 1860 4480
rect 1815 4440 1860 4468
rect 1854 4428 1860 4440
rect 1912 4428 1918 4480
rect 2148 4477 2176 4508
rect 2133 4471 2191 4477
rect 2133 4437 2145 4471
rect 2179 4437 2191 4471
rect 2133 4431 2191 4437
rect 2409 4471 2467 4477
rect 2409 4437 2421 4471
rect 2455 4468 2467 4471
rect 2498 4468 2504 4480
rect 2455 4440 2504 4468
rect 2455 4437 2467 4440
rect 2409 4431 2467 4437
rect 2498 4428 2504 4440
rect 2556 4428 2562 4480
rect 2746 4468 2774 4508
rect 3786 4496 3792 4508
rect 3844 4496 3850 4548
rect 5813 4539 5871 4545
rect 5813 4505 5825 4539
rect 5859 4536 5871 4539
rect 6380 4536 6408 4576
rect 6638 4564 6644 4576
rect 6696 4564 6702 4616
rect 7466 4604 7472 4616
rect 7427 4576 7472 4604
rect 7466 4564 7472 4576
rect 7524 4564 7530 4616
rect 8294 4604 8300 4616
rect 8255 4576 8300 4604
rect 8294 4564 8300 4576
rect 8352 4564 8358 4616
rect 9646 4604 9674 4644
rect 9766 4632 9772 4684
rect 9824 4672 9830 4684
rect 10870 4672 10876 4684
rect 9824 4644 10876 4672
rect 9824 4632 9830 4644
rect 10870 4632 10876 4644
rect 10928 4672 10934 4684
rect 11333 4675 11391 4681
rect 11333 4672 11345 4675
rect 10928 4644 11345 4672
rect 10928 4632 10934 4644
rect 11333 4641 11345 4644
rect 11379 4641 11391 4675
rect 11333 4635 11391 4641
rect 11422 4632 11428 4684
rect 11480 4672 11486 4684
rect 11517 4675 11575 4681
rect 11517 4672 11529 4675
rect 11480 4644 11529 4672
rect 11480 4632 11486 4644
rect 11517 4641 11529 4644
rect 11563 4641 11575 4675
rect 11517 4635 11575 4641
rect 12161 4675 12219 4681
rect 12161 4641 12173 4675
rect 12207 4672 12219 4675
rect 12526 4672 12532 4684
rect 12207 4644 12532 4672
rect 12207 4641 12219 4644
rect 12161 4635 12219 4641
rect 12526 4632 12532 4644
rect 12584 4632 12590 4684
rect 12802 4632 12808 4684
rect 12860 4672 12866 4684
rect 13449 4675 13507 4681
rect 13449 4672 13461 4675
rect 12860 4644 13461 4672
rect 12860 4632 12866 4644
rect 13449 4641 13461 4644
rect 13495 4641 13507 4675
rect 13449 4635 13507 4641
rect 10042 4604 10048 4616
rect 9646 4576 10048 4604
rect 10042 4564 10048 4576
rect 10100 4564 10106 4616
rect 10321 4607 10379 4613
rect 10321 4604 10333 4607
rect 10244 4576 10333 4604
rect 10134 4536 10140 4548
rect 5859 4508 6316 4536
rect 6380 4508 10140 4536
rect 5859 4505 5871 4508
rect 5813 4499 5871 4505
rect 2961 4471 3019 4477
rect 2961 4468 2973 4471
rect 2746 4440 2973 4468
rect 2961 4437 2973 4440
rect 3007 4437 3019 4471
rect 3234 4468 3240 4480
rect 3195 4440 3240 4468
rect 2961 4431 3019 4437
rect 3234 4428 3240 4440
rect 3292 4428 3298 4480
rect 4062 4468 4068 4480
rect 4023 4440 4068 4468
rect 4062 4428 4068 4440
rect 4120 4428 4126 4480
rect 5721 4471 5779 4477
rect 5721 4437 5733 4471
rect 5767 4468 5779 4471
rect 6086 4468 6092 4480
rect 5767 4440 6092 4468
rect 5767 4437 5779 4440
rect 5721 4431 5779 4437
rect 6086 4428 6092 4440
rect 6144 4428 6150 4480
rect 6288 4477 6316 4508
rect 10134 4496 10140 4508
rect 10192 4496 10198 4548
rect 6273 4471 6331 4477
rect 6273 4437 6285 4471
rect 6319 4437 6331 4471
rect 6273 4431 6331 4437
rect 8757 4471 8815 4477
rect 8757 4437 8769 4471
rect 8803 4468 8815 4471
rect 9582 4468 9588 4480
rect 8803 4440 9588 4468
rect 8803 4437 8815 4440
rect 8757 4431 8815 4437
rect 9582 4428 9588 4440
rect 9640 4428 9646 4480
rect 9674 4428 9680 4480
rect 9732 4468 9738 4480
rect 10244 4468 10272 4576
rect 10321 4573 10333 4576
rect 10367 4573 10379 4607
rect 10321 4567 10379 4573
rect 12345 4607 12403 4613
rect 12345 4573 12357 4607
rect 12391 4604 12403 4607
rect 13354 4604 13360 4616
rect 12391 4576 13360 4604
rect 12391 4573 12403 4576
rect 12345 4567 12403 4573
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 13464 4604 13492 4635
rect 13722 4632 13728 4684
rect 13780 4672 13786 4684
rect 14737 4675 14795 4681
rect 14737 4672 14749 4675
rect 13780 4644 14749 4672
rect 13780 4632 13786 4644
rect 14737 4641 14749 4644
rect 14783 4641 14795 4675
rect 14737 4635 14795 4641
rect 15010 4632 15016 4684
rect 15068 4672 15074 4684
rect 15746 4672 15752 4684
rect 15068 4644 15541 4672
rect 15707 4644 15752 4672
rect 15068 4632 15074 4644
rect 13814 4604 13820 4616
rect 13464 4576 13820 4604
rect 13814 4564 13820 4576
rect 13872 4564 13878 4616
rect 14553 4607 14611 4613
rect 14553 4604 14565 4607
rect 14108 4576 14565 4604
rect 14108 4480 14136 4576
rect 14553 4573 14565 4576
rect 14599 4573 14611 4607
rect 14553 4567 14611 4573
rect 14642 4564 14648 4616
rect 14700 4604 14706 4616
rect 14918 4604 14924 4616
rect 14700 4576 14924 4604
rect 14700 4564 14706 4576
rect 14918 4564 14924 4576
rect 14976 4564 14982 4616
rect 15513 4613 15541 4644
rect 15746 4632 15752 4644
rect 15804 4672 15810 4684
rect 15933 4675 15991 4681
rect 15933 4672 15945 4675
rect 15804 4644 15945 4672
rect 15804 4632 15810 4644
rect 15933 4641 15945 4644
rect 15979 4672 15991 4675
rect 16316 4672 16344 4712
rect 15979 4644 16344 4672
rect 15979 4641 15991 4644
rect 15933 4635 15991 4641
rect 16390 4632 16396 4684
rect 16448 4672 16454 4684
rect 16448 4644 16896 4672
rect 16448 4632 16454 4644
rect 15497 4607 15555 4613
rect 15497 4573 15509 4607
rect 15543 4573 15555 4607
rect 15497 4567 15555 4573
rect 16577 4607 16635 4613
rect 16577 4573 16589 4607
rect 16623 4604 16635 4607
rect 16758 4604 16764 4616
rect 16623 4576 16764 4604
rect 16623 4573 16635 4576
rect 16577 4567 16635 4573
rect 16758 4564 16764 4576
rect 16816 4564 16822 4616
rect 16868 4613 16896 4644
rect 16853 4607 16911 4613
rect 16853 4573 16865 4607
rect 16899 4573 16911 4607
rect 16853 4567 16911 4573
rect 17129 4607 17187 4613
rect 17129 4573 17141 4607
rect 17175 4573 17187 4607
rect 17129 4567 17187 4573
rect 14274 4536 14280 4548
rect 14235 4508 14280 4536
rect 14274 4496 14280 4508
rect 14332 4496 14338 4548
rect 15381 4539 15439 4545
rect 15381 4505 15393 4539
rect 15427 4505 15439 4539
rect 17144 4536 17172 4567
rect 15381 4499 15439 4505
rect 15948 4508 17172 4536
rect 17328 4536 17356 4712
rect 17420 4613 17448 4780
rect 17589 4743 17647 4749
rect 17589 4709 17601 4743
rect 17635 4740 17647 4743
rect 18138 4740 18144 4752
rect 17635 4712 18144 4740
rect 17635 4709 17647 4712
rect 17589 4703 17647 4709
rect 18138 4700 18144 4712
rect 18196 4700 18202 4752
rect 17405 4607 17463 4613
rect 17405 4573 17417 4607
rect 17451 4573 17463 4607
rect 17405 4567 17463 4573
rect 17681 4607 17739 4613
rect 17681 4573 17693 4607
rect 17727 4573 17739 4607
rect 17681 4567 17739 4573
rect 17696 4536 17724 4567
rect 18046 4564 18052 4616
rect 18104 4604 18110 4616
rect 18141 4607 18199 4613
rect 18141 4604 18153 4607
rect 18104 4576 18153 4604
rect 18104 4564 18110 4576
rect 18141 4573 18153 4576
rect 18187 4573 18199 4607
rect 18141 4567 18199 4573
rect 18233 4607 18291 4613
rect 18233 4573 18245 4607
rect 18279 4604 18291 4607
rect 18322 4604 18328 4616
rect 18279 4576 18328 4604
rect 18279 4573 18291 4576
rect 18233 4567 18291 4573
rect 18322 4564 18328 4576
rect 18380 4564 18386 4616
rect 17328 4508 17724 4536
rect 10778 4468 10784 4480
rect 9732 4440 10272 4468
rect 10739 4440 10784 4468
rect 9732 4428 9738 4440
rect 10778 4428 10784 4440
rect 10836 4428 10842 4480
rect 10870 4428 10876 4480
rect 10928 4468 10934 4480
rect 13909 4471 13967 4477
rect 10928 4440 10973 4468
rect 10928 4428 10934 4440
rect 13909 4437 13921 4471
rect 13955 4468 13967 4471
rect 14090 4468 14096 4480
rect 13955 4440 14096 4468
rect 13955 4437 13967 4440
rect 13909 4431 13967 4437
rect 14090 4428 14096 4440
rect 14148 4428 14154 4480
rect 15396 4468 15424 4499
rect 15948 4468 15976 4508
rect 16114 4468 16120 4480
rect 15396 4440 15976 4468
rect 16075 4440 16120 4468
rect 16114 4428 16120 4440
rect 16172 4428 16178 4480
rect 16390 4468 16396 4480
rect 16351 4440 16396 4468
rect 16390 4428 16396 4440
rect 16448 4428 16454 4480
rect 16761 4471 16819 4477
rect 16761 4437 16773 4471
rect 16807 4468 16819 4471
rect 16850 4468 16856 4480
rect 16807 4440 16856 4468
rect 16807 4437 16819 4440
rect 16761 4431 16819 4437
rect 16850 4428 16856 4440
rect 16908 4428 16914 4480
rect 17037 4471 17095 4477
rect 17037 4437 17049 4471
rect 17083 4468 17095 4471
rect 17218 4468 17224 4480
rect 17083 4440 17224 4468
rect 17083 4437 17095 4440
rect 17037 4431 17095 4437
rect 17218 4428 17224 4440
rect 17276 4428 17282 4480
rect 17310 4428 17316 4480
rect 17368 4468 17374 4480
rect 17862 4468 17868 4480
rect 17368 4440 17413 4468
rect 17823 4440 17868 4468
rect 17368 4428 17374 4440
rect 17862 4428 17868 4440
rect 17920 4428 17926 4480
rect 17954 4428 17960 4480
rect 18012 4468 18018 4480
rect 18414 4468 18420 4480
rect 18012 4440 18057 4468
rect 18375 4440 18420 4468
rect 18012 4428 18018 4440
rect 18414 4428 18420 4440
rect 18472 4428 18478 4480
rect 1104 4378 18860 4400
rect 1104 4326 5398 4378
rect 5450 4326 5462 4378
rect 5514 4326 5526 4378
rect 5578 4326 5590 4378
rect 5642 4326 5654 4378
rect 5706 4326 9846 4378
rect 9898 4326 9910 4378
rect 9962 4326 9974 4378
rect 10026 4326 10038 4378
rect 10090 4326 10102 4378
rect 10154 4326 14294 4378
rect 14346 4326 14358 4378
rect 14410 4326 14422 4378
rect 14474 4326 14486 4378
rect 14538 4326 14550 4378
rect 14602 4326 18860 4378
rect 1104 4304 18860 4326
rect 4798 4224 4804 4276
rect 4856 4264 4862 4276
rect 5534 4264 5540 4276
rect 4856 4236 5540 4264
rect 4856 4224 4862 4236
rect 5534 4224 5540 4236
rect 5592 4264 5598 4276
rect 6086 4264 6092 4276
rect 5592 4236 5948 4264
rect 6047 4236 6092 4264
rect 5592 4224 5598 4236
rect 3234 4196 3240 4208
rect 1964 4168 3240 4196
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4128 1731 4131
rect 1964 4128 1992 4168
rect 3234 4156 3240 4168
rect 3292 4156 3298 4208
rect 5721 4199 5779 4205
rect 5721 4165 5733 4199
rect 5767 4196 5779 4199
rect 5810 4196 5816 4208
rect 5767 4168 5816 4196
rect 5767 4165 5779 4168
rect 5721 4159 5779 4165
rect 5810 4156 5816 4168
rect 5868 4156 5874 4208
rect 5920 4196 5948 4236
rect 6086 4224 6092 4236
rect 6144 4224 6150 4276
rect 6457 4267 6515 4273
rect 6457 4233 6469 4267
rect 6503 4264 6515 4267
rect 6638 4264 6644 4276
rect 6503 4236 6644 4264
rect 6503 4233 6515 4236
rect 6457 4227 6515 4233
rect 6638 4224 6644 4236
rect 6696 4224 6702 4276
rect 7006 4224 7012 4276
rect 7064 4264 7070 4276
rect 16390 4264 16396 4276
rect 7064 4236 16396 4264
rect 7064 4224 7070 4236
rect 16390 4224 16396 4236
rect 16448 4224 16454 4276
rect 6822 4196 6828 4208
rect 5920 4168 6828 4196
rect 6822 4156 6828 4168
rect 6880 4156 6886 4208
rect 8938 4156 8944 4208
rect 8996 4196 9002 4208
rect 8996 4168 9628 4196
rect 8996 4156 9002 4168
rect 1719 4100 1992 4128
rect 2041 4131 2099 4137
rect 1719 4097 1731 4100
rect 1673 4091 1731 4097
rect 2041 4097 2053 4131
rect 2087 4128 2099 4131
rect 2317 4131 2375 4137
rect 2087 4100 2176 4128
rect 2087 4097 2099 4100
rect 2041 4091 2099 4097
rect 1486 3992 1492 4004
rect 1447 3964 1492 3992
rect 1486 3952 1492 3964
rect 1544 3952 1550 4004
rect 2148 4001 2176 4100
rect 2317 4097 2329 4131
rect 2363 4097 2375 4131
rect 2590 4128 2596 4140
rect 2551 4100 2596 4128
rect 2317 4091 2375 4097
rect 2133 3995 2191 4001
rect 2133 3961 2145 3995
rect 2179 3961 2191 3995
rect 2332 3992 2360 4091
rect 2590 4088 2596 4100
rect 2648 4088 2654 4140
rect 2866 4128 2872 4140
rect 2827 4100 2872 4128
rect 2866 4088 2872 4100
rect 2924 4088 2930 4140
rect 3145 4131 3203 4137
rect 3145 4097 3157 4131
rect 3191 4097 3203 4131
rect 3145 4091 3203 4097
rect 3329 4131 3387 4137
rect 3329 4097 3341 4131
rect 3375 4128 3387 4131
rect 3510 4128 3516 4140
rect 3375 4100 3516 4128
rect 3375 4097 3387 4100
rect 3329 4091 3387 4097
rect 2682 4020 2688 4072
rect 2740 4060 2746 4072
rect 3160 4060 3188 4091
rect 3510 4088 3516 4100
rect 3568 4088 3574 4140
rect 3878 4128 3884 4140
rect 3791 4100 3884 4128
rect 3878 4088 3884 4100
rect 3936 4128 3942 4140
rect 6454 4128 6460 4140
rect 3936 4100 6460 4128
rect 3936 4088 3942 4100
rect 6454 4088 6460 4100
rect 6512 4088 6518 4140
rect 8294 4088 8300 4140
rect 8352 4128 8358 4140
rect 9033 4131 9091 4137
rect 9033 4128 9045 4131
rect 8352 4100 9045 4128
rect 8352 4088 8358 4100
rect 9033 4097 9045 4100
rect 9079 4097 9091 4131
rect 9033 4091 9091 4097
rect 9122 4088 9128 4140
rect 9180 4128 9186 4140
rect 9600 4128 9628 4168
rect 10778 4156 10784 4208
rect 10836 4196 10842 4208
rect 10836 4168 14479 4196
rect 10836 4156 10842 4168
rect 14451 4140 14479 4168
rect 15120 4168 16528 4196
rect 10321 4131 10379 4137
rect 10321 4128 10333 4131
rect 9180 4100 9225 4128
rect 9600 4100 10333 4128
rect 9180 4088 9186 4100
rect 10321 4097 10333 4100
rect 10367 4097 10379 4131
rect 10321 4091 10379 4097
rect 11790 4088 11796 4140
rect 11848 4128 11854 4140
rect 12345 4131 12403 4137
rect 12345 4128 12357 4131
rect 11848 4100 12357 4128
rect 11848 4088 11854 4100
rect 12345 4097 12357 4100
rect 12391 4097 12403 4131
rect 12345 4091 12403 4097
rect 13262 4088 13268 4140
rect 13320 4128 13326 4140
rect 13449 4131 13507 4137
rect 13449 4128 13461 4131
rect 13320 4100 13461 4128
rect 13320 4088 13326 4100
rect 13449 4097 13461 4100
rect 13495 4097 13507 4131
rect 13449 4091 13507 4097
rect 13814 4088 13820 4140
rect 13872 4128 13878 4140
rect 14451 4137 14464 4140
rect 14093 4131 14151 4137
rect 14093 4128 14105 4131
rect 13872 4100 14105 4128
rect 13872 4088 13878 4100
rect 14093 4097 14105 4100
rect 14139 4097 14151 4131
rect 14093 4091 14151 4097
rect 14436 4131 14464 4137
rect 14436 4097 14448 4131
rect 14436 4091 14464 4097
rect 14458 4088 14464 4091
rect 14516 4088 14522 4140
rect 15120 4128 15148 4168
rect 14568 4100 15148 4128
rect 16500 4128 16528 4168
rect 16669 4131 16727 4137
rect 16669 4128 16681 4131
rect 16500 4100 16681 4128
rect 2740 4032 3188 4060
rect 2740 4020 2746 4032
rect 4154 4020 4160 4072
rect 4212 4060 4218 4072
rect 4706 4060 4712 4072
rect 4212 4032 4712 4060
rect 4212 4020 4218 4032
rect 4706 4020 4712 4032
rect 4764 4020 4770 4072
rect 5534 4060 5540 4072
rect 5495 4032 5540 4060
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 5629 4063 5687 4069
rect 5629 4029 5641 4063
rect 5675 4060 5687 4063
rect 6178 4060 6184 4072
rect 5675 4032 6184 4060
rect 5675 4029 5687 4032
rect 5629 4023 5687 4029
rect 6178 4020 6184 4032
rect 6236 4020 6242 4072
rect 7466 4060 7472 4072
rect 6288 4032 7472 4060
rect 2774 3992 2780 4004
rect 2332 3964 2780 3992
rect 2133 3955 2191 3961
rect 2774 3952 2780 3964
rect 2832 3952 2838 4004
rect 2866 3952 2872 4004
rect 2924 3992 2930 4004
rect 3513 3995 3571 4001
rect 3513 3992 3525 3995
rect 2924 3964 3525 3992
rect 2924 3952 2930 3964
rect 3513 3961 3525 3964
rect 3559 3992 3571 3995
rect 6288 3992 6316 4032
rect 7466 4020 7472 4032
rect 7524 4020 7530 4072
rect 9309 4063 9367 4069
rect 9309 4029 9321 4063
rect 9355 4060 9367 4063
rect 9582 4060 9588 4072
rect 9355 4032 9588 4060
rect 9355 4029 9367 4032
rect 9309 4023 9367 4029
rect 9582 4020 9588 4032
rect 9640 4020 9646 4072
rect 10137 4063 10195 4069
rect 10137 4029 10149 4063
rect 10183 4060 10195 4063
rect 10686 4060 10692 4072
rect 10183 4032 10692 4060
rect 10183 4029 10195 4032
rect 10137 4023 10195 4029
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 10781 4063 10839 4069
rect 10781 4029 10793 4063
rect 10827 4060 10839 4063
rect 12529 4063 12587 4069
rect 10827 4032 11652 4060
rect 10827 4029 10839 4032
rect 10781 4023 10839 4029
rect 9769 3995 9827 4001
rect 3559 3964 6316 3992
rect 6932 3964 8984 3992
rect 3559 3961 3571 3964
rect 3513 3955 3571 3961
rect 1854 3924 1860 3936
rect 1815 3896 1860 3924
rect 1854 3884 1860 3896
rect 1912 3884 1918 3936
rect 1946 3884 1952 3936
rect 2004 3924 2010 3936
rect 2409 3927 2467 3933
rect 2409 3924 2421 3927
rect 2004 3896 2421 3924
rect 2004 3884 2010 3896
rect 2409 3893 2421 3896
rect 2455 3893 2467 3927
rect 2682 3924 2688 3936
rect 2643 3896 2688 3924
rect 2409 3887 2467 3893
rect 2682 3884 2688 3896
rect 2740 3884 2746 3936
rect 2958 3924 2964 3936
rect 2919 3896 2964 3924
rect 2958 3884 2964 3896
rect 3016 3884 3022 3936
rect 3694 3924 3700 3936
rect 3655 3896 3700 3924
rect 3694 3884 3700 3896
rect 3752 3884 3758 3936
rect 6730 3884 6736 3936
rect 6788 3924 6794 3936
rect 6932 3924 6960 3964
rect 6788 3896 6960 3924
rect 6788 3884 6794 3896
rect 8478 3884 8484 3936
rect 8536 3924 8542 3936
rect 8573 3927 8631 3933
rect 8573 3924 8585 3927
rect 8536 3896 8585 3924
rect 8536 3884 8542 3896
rect 8573 3893 8585 3896
rect 8619 3893 8631 3927
rect 8846 3924 8852 3936
rect 8807 3896 8852 3924
rect 8573 3887 8631 3893
rect 8846 3884 8852 3896
rect 8904 3884 8910 3936
rect 8956 3924 8984 3964
rect 9769 3961 9781 3995
rect 9815 3992 9827 3995
rect 11624 3992 11652 4032
rect 12529 4029 12541 4063
rect 12575 4060 12587 4063
rect 12618 4060 12624 4072
rect 12575 4032 12624 4060
rect 12575 4029 12587 4032
rect 12529 4023 12587 4029
rect 12618 4020 12624 4032
rect 12676 4020 12682 4072
rect 12989 4063 13047 4069
rect 12989 4029 13001 4063
rect 13035 4060 13047 4063
rect 13170 4060 13176 4072
rect 13035 4032 13176 4060
rect 13035 4029 13047 4032
rect 12989 4023 13047 4029
rect 13170 4020 13176 4032
rect 13228 4020 13234 4072
rect 14568 4060 14596 4100
rect 16669 4097 16681 4100
rect 16715 4097 16727 4131
rect 16669 4091 16727 4097
rect 16945 4131 17003 4137
rect 16945 4097 16957 4131
rect 16991 4097 17003 4131
rect 16945 4091 17003 4097
rect 15654 4060 15660 4072
rect 13372 4032 14596 4060
rect 15615 4032 15660 4060
rect 13372 3992 13400 4032
rect 15654 4020 15660 4032
rect 15712 4020 15718 4072
rect 16301 4063 16359 4069
rect 16301 4029 16313 4063
rect 16347 4029 16359 4063
rect 16301 4023 16359 4029
rect 16485 4063 16543 4069
rect 16485 4029 16497 4063
rect 16531 4029 16543 4063
rect 16960 4060 16988 4091
rect 17034 4088 17040 4140
rect 17092 4128 17098 4140
rect 17221 4131 17279 4137
rect 17221 4128 17233 4131
rect 17092 4100 17233 4128
rect 17092 4088 17098 4100
rect 17221 4097 17233 4100
rect 17267 4097 17279 4131
rect 17586 4128 17592 4140
rect 17547 4100 17592 4128
rect 17221 4091 17279 4097
rect 17586 4088 17592 4100
rect 17644 4128 17650 4140
rect 17770 4128 17776 4140
rect 17644 4100 17776 4128
rect 17644 4088 17650 4100
rect 17770 4088 17776 4100
rect 17828 4088 17834 4140
rect 17865 4131 17923 4137
rect 17865 4097 17877 4131
rect 17911 4128 17923 4131
rect 17954 4128 17960 4140
rect 17911 4100 17960 4128
rect 17911 4097 17923 4100
rect 17865 4091 17923 4097
rect 17954 4088 17960 4100
rect 18012 4088 18018 4140
rect 18233 4131 18291 4137
rect 18233 4097 18245 4131
rect 18279 4097 18291 4131
rect 18233 4091 18291 4097
rect 18248 4060 18276 4091
rect 16485 4023 16543 4029
rect 16592 4032 16988 4060
rect 17788 4032 18276 4060
rect 9815 3964 11100 3992
rect 11624 3964 13400 3992
rect 9815 3961 9827 3964
rect 9769 3955 9827 3961
rect 10318 3924 10324 3936
rect 8956 3896 10324 3924
rect 10318 3884 10324 3896
rect 10376 3884 10382 3936
rect 11072 3924 11100 3964
rect 13446 3952 13452 4004
rect 13504 3992 13510 4004
rect 13909 3995 13967 4001
rect 13909 3992 13921 3995
rect 13504 3964 13921 3992
rect 13504 3952 13510 3964
rect 13909 3961 13921 3964
rect 13955 3961 13967 3995
rect 13909 3955 13967 3961
rect 14507 3995 14565 4001
rect 14507 3961 14519 3995
rect 14553 3992 14565 3995
rect 16316 3992 16344 4023
rect 14553 3964 16344 3992
rect 14553 3961 14565 3964
rect 14507 3955 14565 3961
rect 16390 3952 16396 4004
rect 16448 3992 16454 4004
rect 16500 3992 16528 4023
rect 16448 3964 16528 3992
rect 16448 3952 16454 3964
rect 12802 3924 12808 3936
rect 11072 3896 12808 3924
rect 12802 3884 12808 3896
rect 12860 3884 12866 3936
rect 13078 3884 13084 3936
rect 13136 3924 13142 3936
rect 13136 3896 13181 3924
rect 13136 3884 13142 3896
rect 13262 3884 13268 3936
rect 13320 3924 13326 3936
rect 13630 3924 13636 3936
rect 13320 3896 13365 3924
rect 13591 3896 13636 3924
rect 13320 3884 13326 3896
rect 13630 3884 13636 3896
rect 13688 3884 13694 3936
rect 13814 3924 13820 3936
rect 13775 3896 13820 3924
rect 13814 3884 13820 3896
rect 13872 3884 13878 3936
rect 13998 3884 14004 3936
rect 14056 3924 14062 3936
rect 14185 3927 14243 3933
rect 14185 3924 14197 3927
rect 14056 3896 14197 3924
rect 14056 3884 14062 3896
rect 14185 3893 14197 3896
rect 14231 3893 14243 3927
rect 14185 3887 14243 3893
rect 14642 3884 14648 3936
rect 14700 3924 14706 3936
rect 16592 3924 16620 4032
rect 16853 3995 16911 4001
rect 16853 3961 16865 3995
rect 16899 3992 16911 3995
rect 17034 3992 17040 4004
rect 16899 3964 17040 3992
rect 16899 3961 16911 3964
rect 16853 3955 16911 3961
rect 17034 3952 17040 3964
rect 17092 3952 17098 4004
rect 17788 4001 17816 4032
rect 17773 3995 17831 4001
rect 17773 3961 17785 3995
rect 17819 3961 17831 3995
rect 17773 3955 17831 3961
rect 18049 3995 18107 4001
rect 18049 3961 18061 3995
rect 18095 3992 18107 3995
rect 18874 3992 18880 4004
rect 18095 3964 18880 3992
rect 18095 3961 18107 3964
rect 18049 3955 18107 3961
rect 18874 3952 18880 3964
rect 18932 3952 18938 4004
rect 17126 3924 17132 3936
rect 14700 3896 16620 3924
rect 17087 3896 17132 3924
rect 14700 3884 14706 3896
rect 17126 3884 17132 3896
rect 17184 3884 17190 3936
rect 17405 3927 17463 3933
rect 17405 3893 17417 3927
rect 17451 3924 17463 3927
rect 17678 3924 17684 3936
rect 17451 3896 17684 3924
rect 17451 3893 17463 3896
rect 17405 3887 17463 3893
rect 17678 3884 17684 3896
rect 17736 3884 17742 3936
rect 18414 3924 18420 3936
rect 18375 3896 18420 3924
rect 18414 3884 18420 3896
rect 18472 3884 18478 3936
rect 1104 3834 18860 3856
rect 1104 3782 3174 3834
rect 3226 3782 3238 3834
rect 3290 3782 3302 3834
rect 3354 3782 3366 3834
rect 3418 3782 3430 3834
rect 3482 3782 7622 3834
rect 7674 3782 7686 3834
rect 7738 3782 7750 3834
rect 7802 3782 7814 3834
rect 7866 3782 7878 3834
rect 7930 3782 12070 3834
rect 12122 3782 12134 3834
rect 12186 3782 12198 3834
rect 12250 3782 12262 3834
rect 12314 3782 12326 3834
rect 12378 3782 16518 3834
rect 16570 3782 16582 3834
rect 16634 3782 16646 3834
rect 16698 3782 16710 3834
rect 16762 3782 16774 3834
rect 16826 3782 18860 3834
rect 1104 3760 18860 3782
rect 2590 3680 2596 3732
rect 2648 3720 2654 3732
rect 3694 3720 3700 3732
rect 2648 3692 3700 3720
rect 2648 3680 2654 3692
rect 3694 3680 3700 3692
rect 3752 3680 3758 3732
rect 9398 3680 9404 3732
rect 9456 3720 9462 3732
rect 10042 3720 10048 3732
rect 9456 3692 10048 3720
rect 9456 3680 9462 3692
rect 10042 3680 10048 3692
rect 10100 3720 10106 3732
rect 12618 3720 12624 3732
rect 10100 3692 12624 3720
rect 10100 3680 10106 3692
rect 12618 3680 12624 3692
rect 12676 3680 12682 3732
rect 13170 3680 13176 3732
rect 13228 3720 13234 3732
rect 13817 3723 13875 3729
rect 13228 3692 13768 3720
rect 13228 3680 13234 3692
rect 2774 3612 2780 3664
rect 2832 3652 2838 3664
rect 3421 3655 3479 3661
rect 3421 3652 3433 3655
rect 2832 3624 3433 3652
rect 2832 3612 2838 3624
rect 3421 3621 3433 3624
rect 3467 3621 3479 3655
rect 8110 3652 8116 3664
rect 3421 3615 3479 3621
rect 3988 3624 8116 3652
rect 2682 3584 2688 3596
rect 2056 3556 2688 3584
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3516 1731 3519
rect 1946 3516 1952 3528
rect 1719 3488 1952 3516
rect 1719 3485 1731 3488
rect 1673 3479 1731 3485
rect 1946 3476 1952 3488
rect 2004 3476 2010 3528
rect 2056 3525 2084 3556
rect 2682 3544 2688 3556
rect 2740 3544 2746 3596
rect 3988 3593 4016 3624
rect 8110 3612 8116 3624
rect 8168 3612 8174 3664
rect 8297 3655 8355 3661
rect 8297 3621 8309 3655
rect 8343 3652 8355 3655
rect 10318 3652 10324 3664
rect 8343 3624 10324 3652
rect 8343 3621 8355 3624
rect 8297 3615 8355 3621
rect 10318 3612 10324 3624
rect 10376 3612 10382 3664
rect 12526 3652 12532 3664
rect 12487 3624 12532 3652
rect 12526 3612 12532 3624
rect 12584 3612 12590 3664
rect 13630 3612 13636 3664
rect 13688 3612 13694 3664
rect 13740 3652 13768 3692
rect 13817 3689 13829 3723
rect 13863 3720 13875 3723
rect 13906 3720 13912 3732
rect 13863 3692 13912 3720
rect 13863 3689 13875 3692
rect 13817 3683 13875 3689
rect 13906 3680 13912 3692
rect 13964 3680 13970 3732
rect 16390 3680 16396 3732
rect 16448 3720 16454 3732
rect 16761 3723 16819 3729
rect 16761 3720 16773 3723
rect 16448 3692 16773 3720
rect 16448 3680 16454 3692
rect 16761 3689 16773 3692
rect 16807 3689 16819 3723
rect 16761 3683 16819 3689
rect 16942 3652 16948 3664
rect 13740 3624 16948 3652
rect 16942 3612 16948 3624
rect 17000 3612 17006 3664
rect 17313 3655 17371 3661
rect 17313 3621 17325 3655
rect 17359 3652 17371 3655
rect 18506 3652 18512 3664
rect 17359 3624 18512 3652
rect 17359 3621 17371 3624
rect 17313 3615 17371 3621
rect 18506 3612 18512 3624
rect 18564 3612 18570 3664
rect 3973 3587 4031 3593
rect 3973 3584 3985 3587
rect 2884 3556 3985 3584
rect 2041 3519 2099 3525
rect 2041 3485 2053 3519
rect 2087 3485 2099 3519
rect 2406 3516 2412 3528
rect 2367 3488 2412 3516
rect 2041 3479 2099 3485
rect 2406 3476 2412 3488
rect 2464 3476 2470 3528
rect 2498 3476 2504 3528
rect 2556 3516 2562 3528
rect 2884 3525 2912 3556
rect 3973 3553 3985 3556
rect 4019 3553 4031 3587
rect 7374 3584 7380 3596
rect 3973 3547 4031 3553
rect 5552 3556 7380 3584
rect 2869 3519 2927 3525
rect 2556 3488 2601 3516
rect 2556 3476 2562 3488
rect 2869 3485 2881 3519
rect 2915 3485 2927 3519
rect 2869 3479 2927 3485
rect 3329 3519 3387 3525
rect 3329 3485 3341 3519
rect 3375 3516 3387 3519
rect 3510 3516 3516 3528
rect 3375 3488 3516 3516
rect 3375 3485 3387 3488
rect 3329 3479 3387 3485
rect 3510 3476 3516 3488
rect 3568 3476 3574 3528
rect 3605 3519 3663 3525
rect 3605 3485 3617 3519
rect 3651 3516 3663 3519
rect 3786 3516 3792 3528
rect 3651 3488 3792 3516
rect 3651 3485 3663 3488
rect 3605 3479 3663 3485
rect 3786 3476 3792 3488
rect 3844 3476 3850 3528
rect 5552 3525 5580 3556
rect 7374 3544 7380 3556
rect 7432 3544 7438 3596
rect 8478 3584 8484 3596
rect 8439 3556 8484 3584
rect 8478 3544 8484 3556
rect 8536 3544 8542 3596
rect 8662 3584 8668 3596
rect 8623 3556 8668 3584
rect 8662 3544 8668 3556
rect 8720 3544 8726 3596
rect 11054 3584 11060 3596
rect 9140 3556 10916 3584
rect 5537 3519 5595 3525
rect 5537 3485 5549 3519
rect 5583 3485 5595 3519
rect 6730 3516 6736 3528
rect 6691 3488 6736 3516
rect 5537 3479 5595 3485
rect 6730 3476 6736 3488
rect 6788 3476 6794 3528
rect 6825 3519 6883 3525
rect 6825 3485 6837 3519
rect 6871 3516 6883 3519
rect 7628 3519 7686 3525
rect 7628 3516 7640 3519
rect 6871 3488 7640 3516
rect 6871 3485 6883 3488
rect 6825 3479 6883 3485
rect 7628 3485 7640 3488
rect 7674 3516 7686 3519
rect 8496 3516 8524 3544
rect 7674 3488 8524 3516
rect 7674 3485 7686 3488
rect 7628 3479 7686 3485
rect 8938 3476 8944 3528
rect 8996 3516 9002 3528
rect 9140 3525 9168 3556
rect 9125 3519 9183 3525
rect 9125 3516 9137 3519
rect 8996 3488 9137 3516
rect 8996 3476 9002 3488
rect 9125 3485 9137 3488
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 9493 3519 9551 3525
rect 9493 3485 9505 3519
rect 9539 3485 9551 3519
rect 9493 3479 9551 3485
rect 8570 3448 8576 3460
rect 3068 3420 3372 3448
rect 1486 3380 1492 3392
rect 1447 3352 1492 3380
rect 1486 3340 1492 3352
rect 1544 3340 1550 3392
rect 1854 3380 1860 3392
rect 1815 3352 1860 3380
rect 1854 3340 1860 3352
rect 1912 3340 1918 3392
rect 2222 3380 2228 3392
rect 2183 3352 2228 3380
rect 2222 3340 2228 3352
rect 2280 3340 2286 3392
rect 2682 3380 2688 3392
rect 2643 3352 2688 3380
rect 2682 3340 2688 3352
rect 2740 3340 2746 3392
rect 3068 3389 3096 3420
rect 3344 3392 3372 3420
rect 6840 3420 8576 3448
rect 3053 3383 3111 3389
rect 3053 3349 3065 3383
rect 3099 3349 3111 3383
rect 3053 3343 3111 3349
rect 3142 3340 3148 3392
rect 3200 3380 3206 3392
rect 3200 3352 3245 3380
rect 3200 3340 3206 3352
rect 3326 3340 3332 3392
rect 3384 3340 3390 3392
rect 4246 3340 4252 3392
rect 4304 3380 4310 3392
rect 5353 3383 5411 3389
rect 5353 3380 5365 3383
rect 4304 3352 5365 3380
rect 4304 3340 4310 3352
rect 5353 3349 5365 3352
rect 5399 3349 5411 3383
rect 5353 3343 5411 3349
rect 5810 3340 5816 3392
rect 5868 3380 5874 3392
rect 6549 3383 6607 3389
rect 6549 3380 6561 3383
rect 5868 3352 6561 3380
rect 5868 3340 5874 3352
rect 6549 3349 6561 3352
rect 6595 3349 6607 3383
rect 6549 3343 6607 3349
rect 6730 3340 6736 3392
rect 6788 3380 6794 3392
rect 6840 3380 6868 3420
rect 8570 3408 8576 3420
rect 8628 3408 8634 3460
rect 9508 3448 9536 3479
rect 9582 3476 9588 3528
rect 9640 3525 9646 3528
rect 9640 3519 9678 3525
rect 9666 3485 9678 3519
rect 9640 3479 9678 3485
rect 9640 3476 9646 3479
rect 9766 3476 9772 3528
rect 9824 3476 9830 3528
rect 10042 3516 10048 3528
rect 10003 3488 10048 3516
rect 10042 3476 10048 3488
rect 10100 3476 10106 3528
rect 10321 3519 10379 3525
rect 10321 3485 10333 3519
rect 10367 3485 10379 3519
rect 10321 3479 10379 3485
rect 10413 3519 10471 3525
rect 10413 3485 10425 3519
rect 10459 3516 10471 3519
rect 10778 3516 10784 3528
rect 10459 3488 10784 3516
rect 10459 3485 10471 3488
rect 10413 3479 10471 3485
rect 9784 3448 9812 3476
rect 9508 3420 9812 3448
rect 10336 3448 10364 3479
rect 10778 3476 10784 3488
rect 10836 3476 10842 3528
rect 10888 3525 10916 3556
rect 11026 3544 11060 3584
rect 11112 3584 11118 3596
rect 13648 3584 13676 3612
rect 14093 3587 14151 3593
rect 14093 3584 14105 3587
rect 11112 3556 13400 3584
rect 13648 3556 14105 3584
rect 11112 3544 11118 3556
rect 10888 3519 10966 3525
rect 10888 3488 10920 3519
rect 10908 3485 10920 3488
rect 10954 3485 10966 3519
rect 10908 3479 10966 3485
rect 11026 3448 11054 3544
rect 13372 3528 13400 3556
rect 14093 3553 14105 3556
rect 14139 3553 14151 3587
rect 14093 3547 14151 3553
rect 14458 3544 14464 3596
rect 14516 3584 14522 3596
rect 15838 3584 15844 3596
rect 14516 3556 15516 3584
rect 15799 3556 15844 3584
rect 14516 3544 14522 3556
rect 11330 3516 11336 3528
rect 11291 3488 11336 3516
rect 11330 3476 11336 3488
rect 11388 3476 11394 3528
rect 11793 3519 11851 3525
rect 11793 3516 11805 3519
rect 11532 3488 11805 3516
rect 11532 3460 11560 3488
rect 11793 3485 11805 3488
rect 11839 3485 11851 3519
rect 12713 3519 12771 3525
rect 12713 3516 12725 3519
rect 11793 3479 11851 3485
rect 12452 3488 12725 3516
rect 11514 3448 11520 3460
rect 10336 3420 11054 3448
rect 11475 3420 11520 3448
rect 11514 3408 11520 3420
rect 11572 3408 11578 3460
rect 12452 3392 12480 3488
rect 12713 3485 12725 3488
rect 12759 3485 12771 3519
rect 12713 3479 12771 3485
rect 12802 3476 12808 3528
rect 12860 3516 12866 3528
rect 13116 3519 13174 3525
rect 13116 3516 13128 3519
rect 12860 3488 12905 3516
rect 13004 3488 13128 3516
rect 12860 3476 12866 3488
rect 12618 3408 12624 3460
rect 12676 3448 12682 3460
rect 13004 3448 13032 3488
rect 13116 3485 13128 3488
rect 13162 3485 13174 3519
rect 13116 3479 13174 3485
rect 13354 3476 13360 3528
rect 13412 3525 13418 3528
rect 13412 3519 13450 3525
rect 13438 3485 13450 3519
rect 13412 3479 13450 3485
rect 13633 3519 13691 3525
rect 13633 3485 13645 3519
rect 13679 3516 13691 3519
rect 13722 3516 13728 3528
rect 13679 3488 13728 3516
rect 13679 3485 13691 3488
rect 13633 3479 13691 3485
rect 13412 3476 13418 3479
rect 13722 3476 13728 3488
rect 13780 3516 13786 3528
rect 13998 3516 14004 3528
rect 13780 3488 14004 3516
rect 13780 3476 13786 3488
rect 13998 3476 14004 3488
rect 14056 3476 14062 3528
rect 15488 3516 15516 3556
rect 15838 3544 15844 3556
rect 15896 3544 15902 3596
rect 16209 3587 16267 3593
rect 16209 3584 16221 3587
rect 15948 3556 16221 3584
rect 15948 3516 15976 3556
rect 16209 3553 16221 3556
rect 16255 3553 16267 3587
rect 16209 3547 16267 3553
rect 15488 3488 15976 3516
rect 16025 3519 16083 3525
rect 16025 3485 16037 3519
rect 16071 3485 16083 3519
rect 16942 3516 16948 3528
rect 16903 3488 16948 3516
rect 16025 3479 16083 3485
rect 12676 3420 13032 3448
rect 13219 3451 13277 3457
rect 12676 3408 12682 3420
rect 13219 3417 13231 3451
rect 13265 3448 13277 3451
rect 14277 3451 14335 3457
rect 14277 3448 14289 3451
rect 13265 3420 14289 3448
rect 13265 3417 13277 3420
rect 13219 3411 13277 3417
rect 14277 3417 14289 3420
rect 14323 3417 14335 3451
rect 14277 3411 14335 3417
rect 15562 3408 15568 3460
rect 15620 3448 15626 3460
rect 16040 3448 16068 3479
rect 16942 3476 16948 3488
rect 17000 3476 17006 3528
rect 17129 3519 17187 3525
rect 17129 3485 17141 3519
rect 17175 3485 17187 3519
rect 17494 3516 17500 3528
rect 17455 3488 17500 3516
rect 17129 3479 17187 3485
rect 15620 3420 16068 3448
rect 15620 3408 15626 3420
rect 16298 3408 16304 3460
rect 16356 3448 16362 3460
rect 17144 3448 17172 3479
rect 17494 3476 17500 3488
rect 17552 3476 17558 3528
rect 17862 3516 17868 3528
rect 17823 3488 17868 3516
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 18046 3476 18052 3528
rect 18104 3476 18110 3528
rect 18233 3519 18291 3525
rect 18233 3485 18245 3519
rect 18279 3516 18291 3519
rect 18690 3516 18696 3528
rect 18279 3488 18696 3516
rect 18279 3485 18291 3488
rect 18233 3479 18291 3485
rect 18690 3476 18696 3488
rect 18748 3476 18754 3528
rect 18064 3448 18092 3476
rect 16356 3420 17172 3448
rect 17328 3420 18092 3448
rect 16356 3408 16362 3420
rect 7006 3380 7012 3392
rect 6788 3352 6868 3380
rect 6967 3352 7012 3380
rect 6788 3340 6794 3352
rect 7006 3340 7012 3352
rect 7064 3340 7070 3392
rect 7699 3383 7757 3389
rect 7699 3349 7711 3383
rect 7745 3380 7757 3383
rect 7834 3380 7840 3392
rect 7745 3352 7840 3380
rect 7745 3349 7757 3352
rect 7699 3343 7757 3349
rect 7834 3340 7840 3352
rect 7892 3340 7898 3392
rect 8662 3340 8668 3392
rect 8720 3380 8726 3392
rect 8941 3383 8999 3389
rect 8941 3380 8953 3383
rect 8720 3352 8953 3380
rect 8720 3340 8726 3352
rect 8941 3349 8953 3352
rect 8987 3349 8999 3383
rect 8941 3343 8999 3349
rect 9214 3340 9220 3392
rect 9272 3380 9278 3392
rect 9309 3383 9367 3389
rect 9309 3380 9321 3383
rect 9272 3352 9321 3380
rect 9272 3340 9278 3352
rect 9309 3349 9321 3352
rect 9355 3349 9367 3383
rect 9309 3343 9367 3349
rect 9674 3340 9680 3392
rect 9732 3389 9738 3392
rect 9732 3383 9781 3389
rect 9732 3349 9735 3383
rect 9769 3349 9781 3383
rect 9732 3343 9781 3349
rect 9732 3340 9738 3343
rect 9858 3340 9864 3392
rect 9916 3380 9922 3392
rect 10137 3383 10195 3389
rect 9916 3352 9961 3380
rect 9916 3340 9922 3352
rect 10137 3349 10149 3383
rect 10183 3380 10195 3383
rect 10226 3380 10232 3392
rect 10183 3352 10232 3380
rect 10183 3349 10195 3352
rect 10137 3343 10195 3349
rect 10226 3340 10232 3352
rect 10284 3340 10290 3392
rect 10597 3383 10655 3389
rect 10597 3349 10609 3383
rect 10643 3380 10655 3383
rect 10686 3380 10692 3392
rect 10643 3352 10692 3380
rect 10643 3349 10655 3352
rect 10597 3343 10655 3349
rect 10686 3340 10692 3352
rect 10744 3340 10750 3392
rect 10962 3340 10968 3392
rect 11020 3389 11026 3392
rect 11020 3383 11069 3389
rect 11020 3349 11023 3383
rect 11057 3349 11069 3383
rect 11020 3343 11069 3349
rect 11020 3340 11026 3343
rect 11146 3340 11152 3392
rect 11204 3380 11210 3392
rect 11606 3380 11612 3392
rect 11204 3352 11249 3380
rect 11567 3352 11612 3380
rect 11204 3340 11210 3352
rect 11606 3340 11612 3352
rect 11664 3340 11670 3392
rect 12434 3340 12440 3392
rect 12492 3380 12498 3392
rect 12986 3380 12992 3392
rect 12492 3352 12537 3380
rect 12947 3352 12992 3380
rect 12492 3340 12498 3352
rect 12986 3340 12992 3352
rect 13044 3340 13050 3392
rect 13495 3383 13553 3389
rect 13495 3349 13507 3383
rect 13541 3380 13553 3383
rect 13630 3380 13636 3392
rect 13541 3352 13636 3380
rect 13541 3349 13553 3352
rect 13495 3343 13553 3349
rect 13630 3340 13636 3352
rect 13688 3340 13694 3392
rect 16669 3383 16727 3389
rect 16669 3349 16681 3383
rect 16715 3380 16727 3383
rect 17328 3380 17356 3420
rect 16715 3352 17356 3380
rect 16715 3349 16727 3352
rect 16669 3343 16727 3349
rect 17586 3340 17592 3392
rect 17644 3380 17650 3392
rect 17681 3383 17739 3389
rect 17681 3380 17693 3383
rect 17644 3352 17693 3380
rect 17644 3340 17650 3352
rect 17681 3349 17693 3352
rect 17727 3349 17739 3383
rect 18046 3380 18052 3392
rect 18007 3352 18052 3380
rect 17681 3343 17739 3349
rect 18046 3340 18052 3352
rect 18104 3340 18110 3392
rect 18414 3380 18420 3392
rect 18375 3352 18420 3380
rect 18414 3340 18420 3352
rect 18472 3340 18478 3392
rect 1104 3290 18860 3312
rect 1104 3238 5398 3290
rect 5450 3238 5462 3290
rect 5514 3238 5526 3290
rect 5578 3238 5590 3290
rect 5642 3238 5654 3290
rect 5706 3238 9846 3290
rect 9898 3238 9910 3290
rect 9962 3238 9974 3290
rect 10026 3238 10038 3290
rect 10090 3238 10102 3290
rect 10154 3238 14294 3290
rect 14346 3238 14358 3290
rect 14410 3238 14422 3290
rect 14474 3238 14486 3290
rect 14538 3238 14550 3290
rect 14602 3238 18860 3290
rect 1104 3216 18860 3238
rect 3697 3179 3755 3185
rect 3697 3176 3709 3179
rect 2516 3148 3709 3176
rect 934 3068 940 3120
rect 992 3108 998 3120
rect 2406 3108 2412 3120
rect 992 3080 2412 3108
rect 992 3068 998 3080
rect 2406 3068 2412 3080
rect 2464 3068 2470 3120
rect 1394 3040 1400 3052
rect 1355 3012 1400 3040
rect 1394 3000 1400 3012
rect 1452 3000 1458 3052
rect 2130 3040 2136 3052
rect 2091 3012 2136 3040
rect 2130 3000 2136 3012
rect 2188 3000 2194 3052
rect 2516 3049 2544 3148
rect 3697 3145 3709 3148
rect 3743 3145 3755 3179
rect 3697 3139 3755 3145
rect 4525 3179 4583 3185
rect 4525 3145 4537 3179
rect 4571 3145 4583 3179
rect 9582 3176 9588 3188
rect 4525 3139 4583 3145
rect 6840 3148 9588 3176
rect 4540 3108 4568 3139
rect 5077 3111 5135 3117
rect 5077 3108 5089 3111
rect 3252 3080 4568 3108
rect 4724 3080 5089 3108
rect 2501 3043 2559 3049
rect 2501 3009 2513 3043
rect 2547 3009 2559 3043
rect 2501 3003 2559 3009
rect 2590 3000 2596 3052
rect 2648 3040 2654 3052
rect 3252 3049 3280 3080
rect 3237 3043 3295 3049
rect 2648 3012 2693 3040
rect 2648 3000 2654 3012
rect 3237 3009 3249 3043
rect 3283 3009 3295 3043
rect 3237 3003 3295 3009
rect 3326 3000 3332 3052
rect 3384 3040 3390 3052
rect 3881 3043 3939 3049
rect 3384 3012 3429 3040
rect 3384 3000 3390 3012
rect 3881 3009 3893 3043
rect 3927 3040 3939 3043
rect 4062 3040 4068 3052
rect 3927 3012 4068 3040
rect 3927 3009 3939 3012
rect 3881 3003 3939 3009
rect 4062 3000 4068 3012
rect 4120 3000 4126 3052
rect 4724 3049 4752 3080
rect 5077 3077 5089 3080
rect 5123 3108 5135 3111
rect 5123 3080 6592 3108
rect 5123 3077 5135 3080
rect 5077 3071 5135 3077
rect 4157 3043 4215 3049
rect 4157 3009 4169 3043
rect 4203 3009 4215 3043
rect 4157 3003 4215 3009
rect 4709 3043 4767 3049
rect 4709 3009 4721 3043
rect 4755 3009 4767 3043
rect 4982 3040 4988 3052
rect 4943 3012 4988 3040
rect 4709 3003 4767 3009
rect 1949 2975 2007 2981
rect 1949 2941 1961 2975
rect 1995 2972 2007 2975
rect 4172 2972 4200 3003
rect 4982 3000 4988 3012
rect 5040 3000 5046 3052
rect 5537 3043 5595 3049
rect 5537 3009 5549 3043
rect 5583 3009 5595 3043
rect 5537 3003 5595 3009
rect 1995 2944 4200 2972
rect 1995 2941 2007 2944
rect 1949 2935 2007 2941
rect 1581 2907 1639 2913
rect 1581 2873 1593 2907
rect 1627 2904 1639 2907
rect 2590 2904 2596 2916
rect 1627 2876 2596 2904
rect 1627 2873 1639 2876
rect 1581 2867 1639 2873
rect 2590 2864 2596 2876
rect 2648 2864 2654 2916
rect 2777 2907 2835 2913
rect 2777 2904 2789 2907
rect 2700 2876 2789 2904
rect 1394 2796 1400 2848
rect 1452 2836 1458 2848
rect 2317 2839 2375 2845
rect 2317 2836 2329 2839
rect 1452 2808 2329 2836
rect 1452 2796 1458 2808
rect 2317 2805 2329 2808
rect 2363 2805 2375 2839
rect 2317 2799 2375 2805
rect 2406 2796 2412 2848
rect 2464 2836 2470 2848
rect 2700 2836 2728 2876
rect 2777 2873 2789 2876
rect 2823 2873 2835 2907
rect 2777 2867 2835 2873
rect 4154 2864 4160 2916
rect 4212 2904 4218 2916
rect 5353 2907 5411 2913
rect 5353 2904 5365 2907
rect 4212 2876 5365 2904
rect 4212 2864 4218 2876
rect 5353 2873 5365 2876
rect 5399 2873 5411 2907
rect 5552 2904 5580 3003
rect 6564 2972 6592 3080
rect 6730 3040 6736 3052
rect 6691 3012 6736 3040
rect 6730 3000 6736 3012
rect 6788 3000 6794 3052
rect 6840 3049 6868 3148
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 10870 3136 10876 3188
rect 10928 3176 10934 3188
rect 11698 3176 11704 3188
rect 10928 3148 11704 3176
rect 10928 3136 10934 3148
rect 7834 3068 7840 3120
rect 7892 3108 7898 3120
rect 9033 3111 9091 3117
rect 9033 3108 9045 3111
rect 7892 3080 9045 3108
rect 7892 3068 7898 3080
rect 9033 3077 9045 3080
rect 9079 3077 9091 3111
rect 9033 3071 9091 3077
rect 9674 3068 9680 3120
rect 9732 3108 9738 3120
rect 11532 3117 11560 3148
rect 11698 3136 11704 3148
rect 11756 3136 11762 3188
rect 12894 3136 12900 3188
rect 12952 3176 12958 3188
rect 13722 3176 13728 3188
rect 12952 3148 13728 3176
rect 12952 3136 12958 3148
rect 13722 3136 13728 3148
rect 13780 3136 13786 3188
rect 14734 3136 14740 3188
rect 14792 3176 14798 3188
rect 16393 3179 16451 3185
rect 16393 3176 16405 3179
rect 14792 3148 16405 3176
rect 14792 3136 14798 3148
rect 16393 3145 16405 3148
rect 16439 3176 16451 3179
rect 16942 3176 16948 3188
rect 16439 3148 16948 3176
rect 16439 3145 16451 3148
rect 16393 3139 16451 3145
rect 16942 3136 16948 3148
rect 17000 3136 17006 3188
rect 10965 3111 11023 3117
rect 10965 3108 10977 3111
rect 9732 3080 10977 3108
rect 9732 3068 9738 3080
rect 10965 3077 10977 3080
rect 11011 3077 11023 3111
rect 10965 3071 11023 3077
rect 11517 3111 11575 3117
rect 11517 3077 11529 3111
rect 11563 3077 11575 3111
rect 13630 3108 13636 3120
rect 13591 3080 13636 3108
rect 11517 3071 11575 3077
rect 13630 3068 13636 3080
rect 13688 3068 13694 3120
rect 14366 3068 14372 3120
rect 14424 3108 14430 3120
rect 14424 3080 16344 3108
rect 14424 3068 14430 3080
rect 6825 3043 6883 3049
rect 6825 3009 6837 3043
rect 6871 3009 6883 3043
rect 7098 3040 7104 3052
rect 7059 3012 7104 3040
rect 6825 3003 6883 3009
rect 7098 3000 7104 3012
rect 7156 3000 7162 3052
rect 9217 3043 9275 3049
rect 9217 3009 9229 3043
rect 9263 3040 9275 3043
rect 11149 3043 11207 3049
rect 9263 3012 9812 3040
rect 9263 3009 9275 3012
rect 9217 3003 9275 3009
rect 6914 2972 6920 2984
rect 6564 2944 6920 2972
rect 6914 2932 6920 2944
rect 6972 2932 6978 2984
rect 8202 2972 8208 2984
rect 8163 2944 8208 2972
rect 8202 2932 8208 2944
rect 8260 2932 8266 2984
rect 9490 2972 9496 2984
rect 9451 2944 9496 2972
rect 9490 2932 9496 2944
rect 9548 2932 9554 2984
rect 9784 2972 9812 3012
rect 11149 3009 11161 3043
rect 11195 3040 11207 3043
rect 11606 3040 11612 3052
rect 11195 3012 11612 3040
rect 11195 3009 11207 3012
rect 11149 3003 11207 3009
rect 11606 3000 11612 3012
rect 11664 3000 11670 3052
rect 13446 3040 13452 3052
rect 13407 3012 13452 3040
rect 13446 3000 13452 3012
rect 13504 3000 13510 3052
rect 14918 3000 14924 3052
rect 14976 3040 14982 3052
rect 16316 3049 16344 3080
rect 17218 3068 17224 3120
rect 17276 3108 17282 3120
rect 17276 3080 17540 3108
rect 17276 3068 17282 3080
rect 15498 3043 15556 3049
rect 15498 3040 15510 3043
rect 14976 3012 15510 3040
rect 14976 3000 14982 3012
rect 15498 3009 15510 3012
rect 15544 3009 15556 3043
rect 15498 3003 15556 3009
rect 15749 3043 15807 3049
rect 15749 3009 15761 3043
rect 15795 3009 15807 3043
rect 15749 3003 15807 3009
rect 16301 3043 16359 3049
rect 16301 3009 16313 3043
rect 16347 3009 16359 3043
rect 16301 3003 16359 3009
rect 16761 3043 16819 3049
rect 16761 3009 16773 3043
rect 16807 3040 16819 3043
rect 16850 3040 16856 3052
rect 16807 3012 16856 3040
rect 16807 3009 16819 3012
rect 16761 3003 16819 3009
rect 11422 2972 11428 2984
rect 9784 2944 11428 2972
rect 11422 2932 11428 2944
rect 11480 2932 11486 2984
rect 13170 2972 13176 2984
rect 13131 2944 13176 2972
rect 13170 2932 13176 2944
rect 13228 2932 13234 2984
rect 13354 2972 13360 2984
rect 13315 2944 13360 2972
rect 13354 2932 13360 2944
rect 13412 2932 13418 2984
rect 14642 2972 14648 2984
rect 14603 2944 14648 2972
rect 14642 2932 14648 2944
rect 14700 2932 14706 2984
rect 12802 2904 12808 2916
rect 5552 2876 12808 2904
rect 5353 2867 5411 2873
rect 12802 2864 12808 2876
rect 12860 2864 12866 2916
rect 12986 2864 12992 2916
rect 13044 2904 13050 2916
rect 15764 2904 15792 3003
rect 16850 3000 16856 3012
rect 16908 3000 16914 3052
rect 17402 3040 17408 3052
rect 17363 3012 17408 3040
rect 17402 3000 17408 3012
rect 17460 3000 17466 3052
rect 17512 3049 17540 3080
rect 17497 3043 17555 3049
rect 17497 3009 17509 3043
rect 17543 3009 17555 3043
rect 17497 3003 17555 3009
rect 17865 3043 17923 3049
rect 17865 3009 17877 3043
rect 17911 3009 17923 3043
rect 18230 3040 18236 3052
rect 18191 3012 18236 3040
rect 17865 3003 17923 3009
rect 17310 2932 17316 2984
rect 17368 2972 17374 2984
rect 17880 2972 17908 3003
rect 18230 3000 18236 3012
rect 18288 3000 18294 3052
rect 17368 2944 17908 2972
rect 17368 2932 17374 2944
rect 13044 2876 15792 2904
rect 13044 2864 13050 2876
rect 16298 2864 16304 2916
rect 16356 2904 16362 2916
rect 17221 2907 17279 2913
rect 17221 2904 17233 2907
rect 16356 2876 17233 2904
rect 16356 2864 16362 2876
rect 17221 2873 17233 2876
rect 17267 2873 17279 2907
rect 17221 2867 17279 2873
rect 18049 2907 18107 2913
rect 18049 2873 18061 2907
rect 18095 2904 18107 2907
rect 18322 2904 18328 2916
rect 18095 2876 18328 2904
rect 18095 2873 18107 2876
rect 18049 2867 18107 2873
rect 18322 2864 18328 2876
rect 18380 2864 18386 2916
rect 2464 2808 2728 2836
rect 2464 2796 2470 2808
rect 2866 2796 2872 2848
rect 2924 2836 2930 2848
rect 3053 2839 3111 2845
rect 3053 2836 3065 2839
rect 2924 2808 3065 2836
rect 2924 2796 2930 2808
rect 3053 2805 3065 2808
rect 3099 2805 3111 2839
rect 3510 2836 3516 2848
rect 3471 2808 3516 2836
rect 3053 2799 3111 2805
rect 3510 2796 3516 2808
rect 3568 2796 3574 2848
rect 3970 2836 3976 2848
rect 3931 2808 3976 2836
rect 3970 2796 3976 2808
rect 4028 2796 4034 2848
rect 4801 2839 4859 2845
rect 4801 2805 4813 2839
rect 4847 2836 4859 2839
rect 4982 2836 4988 2848
rect 4847 2808 4988 2836
rect 4847 2805 4859 2808
rect 4801 2799 4859 2805
rect 4982 2796 4988 2808
rect 5040 2796 5046 2848
rect 5534 2796 5540 2848
rect 5592 2836 5598 2848
rect 6549 2839 6607 2845
rect 6549 2836 6561 2839
rect 5592 2808 6561 2836
rect 5592 2796 5598 2808
rect 6549 2805 6561 2808
rect 6595 2805 6607 2839
rect 6549 2799 6607 2805
rect 7009 2839 7067 2845
rect 7009 2805 7021 2839
rect 7055 2836 7067 2839
rect 7098 2836 7104 2848
rect 7055 2808 7104 2836
rect 7055 2805 7067 2808
rect 7009 2799 7067 2805
rect 7098 2796 7104 2808
rect 7156 2796 7162 2848
rect 7282 2836 7288 2848
rect 7243 2808 7288 2836
rect 7282 2796 7288 2808
rect 7340 2796 7346 2848
rect 7374 2796 7380 2848
rect 7432 2836 7438 2848
rect 10870 2836 10876 2848
rect 7432 2808 10876 2836
rect 7432 2796 7438 2808
rect 10870 2796 10876 2808
rect 10928 2796 10934 2848
rect 11054 2796 11060 2848
rect 11112 2836 11118 2848
rect 11241 2839 11299 2845
rect 11241 2836 11253 2839
rect 11112 2808 11253 2836
rect 11112 2796 11118 2808
rect 11241 2805 11253 2808
rect 11287 2805 11299 2839
rect 11241 2799 11299 2805
rect 15194 2796 15200 2848
rect 15252 2836 15258 2848
rect 15427 2839 15485 2845
rect 15427 2836 15439 2839
rect 15252 2808 15439 2836
rect 15252 2796 15258 2808
rect 15427 2805 15439 2808
rect 15473 2805 15485 2839
rect 15427 2799 15485 2805
rect 15654 2796 15660 2848
rect 15712 2836 15718 2848
rect 15933 2839 15991 2845
rect 15933 2836 15945 2839
rect 15712 2808 15945 2836
rect 15712 2796 15718 2808
rect 15933 2805 15945 2808
rect 15979 2805 15991 2839
rect 16114 2836 16120 2848
rect 16075 2808 16120 2836
rect 15933 2799 15991 2805
rect 16114 2796 16120 2808
rect 16172 2796 16178 2848
rect 16942 2836 16948 2848
rect 16903 2808 16948 2836
rect 16942 2796 16948 2808
rect 17000 2796 17006 2848
rect 17681 2839 17739 2845
rect 17681 2805 17693 2839
rect 17727 2836 17739 2839
rect 17862 2836 17868 2848
rect 17727 2808 17868 2836
rect 17727 2805 17739 2808
rect 17681 2799 17739 2805
rect 17862 2796 17868 2808
rect 17920 2796 17926 2848
rect 18414 2836 18420 2848
rect 18375 2808 18420 2836
rect 18414 2796 18420 2808
rect 18472 2796 18478 2848
rect 1104 2746 18860 2768
rect 1104 2694 3174 2746
rect 3226 2694 3238 2746
rect 3290 2694 3302 2746
rect 3354 2694 3366 2746
rect 3418 2694 3430 2746
rect 3482 2694 7622 2746
rect 7674 2694 7686 2746
rect 7738 2694 7750 2746
rect 7802 2694 7814 2746
rect 7866 2694 7878 2746
rect 7930 2694 12070 2746
rect 12122 2694 12134 2746
rect 12186 2694 12198 2746
rect 12250 2694 12262 2746
rect 12314 2694 12326 2746
rect 12378 2694 16518 2746
rect 16570 2694 16582 2746
rect 16634 2694 16646 2746
rect 16698 2694 16710 2746
rect 16762 2694 16774 2746
rect 16826 2694 18860 2746
rect 1104 2672 18860 2694
rect 1486 2632 1492 2644
rect 1447 2604 1492 2632
rect 1486 2592 1492 2604
rect 1544 2592 1550 2644
rect 1857 2635 1915 2641
rect 1857 2601 1869 2635
rect 1903 2632 1915 2635
rect 2130 2632 2136 2644
rect 1903 2604 2136 2632
rect 1903 2601 1915 2604
rect 1857 2595 1915 2601
rect 2130 2592 2136 2604
rect 2188 2592 2194 2644
rect 5166 2632 5172 2644
rect 5127 2604 5172 2632
rect 5166 2592 5172 2604
rect 5224 2592 5230 2644
rect 6181 2635 6239 2641
rect 6181 2601 6193 2635
rect 6227 2632 6239 2635
rect 6362 2632 6368 2644
rect 6227 2604 6368 2632
rect 6227 2601 6239 2604
rect 6181 2595 6239 2601
rect 6362 2592 6368 2604
rect 6420 2592 6426 2644
rect 10962 2592 10968 2644
rect 11020 2632 11026 2644
rect 11974 2632 11980 2644
rect 11020 2604 11980 2632
rect 11020 2592 11026 2604
rect 11974 2592 11980 2604
rect 12032 2592 12038 2644
rect 13354 2592 13360 2644
rect 13412 2632 13418 2644
rect 13725 2635 13783 2641
rect 13725 2632 13737 2635
rect 13412 2604 13737 2632
rect 13412 2592 13418 2604
rect 13725 2601 13737 2604
rect 13771 2601 13783 2635
rect 13725 2595 13783 2601
rect 2774 2564 2780 2576
rect 1688 2536 2780 2564
rect 1688 2437 1716 2536
rect 2774 2524 2780 2536
rect 2832 2524 2838 2576
rect 10318 2564 10324 2576
rect 5920 2536 10324 2564
rect 2958 2496 2964 2508
rect 2240 2468 2964 2496
rect 2240 2437 2268 2468
rect 2958 2456 2964 2468
rect 3016 2456 3022 2508
rect 5534 2496 5540 2508
rect 3620 2468 5540 2496
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2397 1731 2431
rect 1673 2391 1731 2397
rect 2225 2431 2283 2437
rect 2225 2397 2237 2431
rect 2271 2397 2283 2431
rect 2225 2391 2283 2397
rect 2685 2431 2743 2437
rect 2685 2397 2697 2431
rect 2731 2428 2743 2431
rect 3050 2428 3056 2440
rect 2731 2400 3056 2428
rect 2731 2397 2743 2400
rect 2685 2391 2743 2397
rect 3050 2388 3056 2400
rect 3108 2388 3114 2440
rect 3620 2437 3648 2468
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 3145 2431 3203 2437
rect 3145 2397 3157 2431
rect 3191 2397 3203 2431
rect 3145 2391 3203 2397
rect 3605 2431 3663 2437
rect 3605 2397 3617 2431
rect 3651 2397 3663 2431
rect 3605 2391 3663 2397
rect 4065 2431 4123 2437
rect 4065 2397 4077 2431
rect 4111 2428 4123 2431
rect 4154 2428 4160 2440
rect 4111 2400 4160 2428
rect 4111 2397 4123 2400
rect 4065 2391 4123 2397
rect 3160 2360 3188 2391
rect 4154 2388 4160 2400
rect 4212 2388 4218 2440
rect 4525 2431 4583 2437
rect 4525 2397 4537 2431
rect 4571 2397 4583 2431
rect 4982 2428 4988 2440
rect 4943 2400 4988 2428
rect 4525 2391 4583 2397
rect 4246 2360 4252 2372
rect 3160 2332 4252 2360
rect 4246 2320 4252 2332
rect 4304 2320 4310 2372
rect 4540 2360 4568 2391
rect 4982 2388 4988 2400
rect 5040 2388 5046 2440
rect 5074 2388 5080 2440
rect 5132 2428 5138 2440
rect 5920 2437 5948 2536
rect 10318 2524 10324 2536
rect 10376 2524 10382 2576
rect 11146 2524 11152 2576
rect 11204 2524 11210 2576
rect 11422 2524 11428 2576
rect 11480 2564 11486 2576
rect 11517 2567 11575 2573
rect 11517 2564 11529 2567
rect 11480 2536 11529 2564
rect 11480 2524 11486 2536
rect 11517 2533 11529 2536
rect 11563 2533 11575 2567
rect 11517 2527 11575 2533
rect 14826 2524 14832 2576
rect 14884 2564 14890 2576
rect 14884 2536 15332 2564
rect 14884 2524 14890 2536
rect 7282 2456 7288 2508
rect 7340 2496 7346 2508
rect 11164 2496 11192 2524
rect 7340 2468 7972 2496
rect 7340 2456 7346 2468
rect 5353 2431 5411 2437
rect 5353 2428 5365 2431
rect 5132 2400 5365 2428
rect 5132 2388 5138 2400
rect 5353 2397 5365 2400
rect 5399 2397 5411 2431
rect 5353 2391 5411 2397
rect 5905 2431 5963 2437
rect 5905 2397 5917 2431
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 5994 2388 6000 2440
rect 6052 2428 6058 2440
rect 6365 2431 6423 2437
rect 6365 2428 6377 2431
rect 6052 2400 6377 2428
rect 6052 2388 6058 2400
rect 6365 2397 6377 2400
rect 6411 2397 6423 2431
rect 6546 2428 6552 2440
rect 6507 2400 6552 2428
rect 6365 2391 6423 2397
rect 6546 2388 6552 2400
rect 6604 2388 6610 2440
rect 7006 2428 7012 2440
rect 6967 2400 7012 2428
rect 7006 2388 7012 2400
rect 7064 2388 7070 2440
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 7944 2437 7972 2468
rect 10520 2468 11192 2496
rect 11793 2499 11851 2505
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 7156 2400 7481 2428
rect 7156 2388 7162 2400
rect 7469 2397 7481 2400
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 7929 2431 7987 2437
rect 7929 2397 7941 2431
rect 7975 2397 7987 2431
rect 8662 2428 8668 2440
rect 8623 2400 8668 2428
rect 7929 2391 7987 2397
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 9214 2428 9220 2440
rect 9175 2400 9220 2428
rect 9214 2388 9220 2400
rect 9272 2388 9278 2440
rect 9585 2431 9643 2437
rect 9585 2397 9597 2431
rect 9631 2428 9643 2431
rect 9766 2428 9772 2440
rect 9631 2400 9772 2428
rect 9631 2397 9643 2400
rect 9585 2391 9643 2397
rect 9766 2388 9772 2400
rect 9824 2388 9830 2440
rect 10045 2431 10103 2437
rect 10045 2397 10057 2431
rect 10091 2428 10103 2431
rect 10226 2428 10232 2440
rect 10091 2400 10232 2428
rect 10091 2397 10103 2400
rect 10045 2391 10103 2397
rect 10226 2388 10232 2400
rect 10284 2388 10290 2440
rect 10520 2437 10548 2468
rect 11793 2465 11805 2499
rect 11839 2496 11851 2499
rect 12526 2496 12532 2508
rect 11839 2468 12532 2496
rect 11839 2465 11851 2468
rect 11793 2459 11851 2465
rect 12526 2456 12532 2468
rect 12584 2456 12590 2508
rect 13538 2496 13544 2508
rect 13499 2468 13544 2496
rect 13538 2456 13544 2468
rect 13596 2456 13602 2508
rect 14182 2496 14188 2508
rect 14143 2468 14188 2496
rect 14182 2456 14188 2468
rect 14240 2456 14246 2508
rect 14369 2499 14427 2505
rect 14369 2465 14381 2499
rect 14415 2496 14427 2499
rect 15194 2496 15200 2508
rect 14415 2468 15200 2496
rect 14415 2465 14427 2468
rect 14369 2459 14427 2465
rect 15194 2456 15200 2468
rect 15252 2456 15258 2508
rect 15304 2505 15332 2536
rect 16574 2524 16580 2576
rect 16632 2564 16638 2576
rect 17221 2567 17279 2573
rect 17221 2564 17233 2567
rect 16632 2536 17233 2564
rect 16632 2524 16638 2536
rect 17221 2533 17233 2536
rect 17267 2533 17279 2567
rect 17221 2527 17279 2533
rect 15289 2499 15347 2505
rect 15289 2465 15301 2499
rect 15335 2465 15347 2499
rect 15289 2459 15347 2465
rect 10505 2431 10563 2437
rect 10505 2397 10517 2431
rect 10551 2397 10563 2431
rect 10686 2428 10692 2440
rect 10647 2400 10692 2428
rect 10505 2391 10563 2397
rect 10686 2388 10692 2400
rect 10744 2388 10750 2440
rect 11124 2431 11182 2437
rect 11124 2397 11136 2431
rect 11170 2428 11182 2431
rect 11170 2397 11192 2428
rect 11124 2391 11192 2397
rect 5810 2360 5816 2372
rect 4540 2332 5816 2360
rect 5810 2320 5816 2332
rect 5868 2320 5874 2372
rect 11164 2360 11192 2391
rect 11238 2388 11244 2440
rect 11296 2428 11302 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11296 2400 11713 2428
rect 11296 2388 11302 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 13909 2431 13967 2437
rect 13909 2397 13921 2431
rect 13955 2397 13967 2431
rect 16114 2428 16120 2440
rect 16075 2400 16120 2428
rect 13909 2391 13967 2397
rect 11330 2360 11336 2372
rect 11164 2332 11336 2360
rect 11330 2320 11336 2332
rect 11388 2320 11394 2372
rect 11440 2332 11928 2360
rect 1854 2252 1860 2304
rect 1912 2292 1918 2304
rect 2041 2295 2099 2301
rect 2041 2292 2053 2295
rect 1912 2264 2053 2292
rect 1912 2252 1918 2264
rect 2041 2261 2053 2264
rect 2087 2261 2099 2295
rect 2041 2255 2099 2261
rect 2314 2252 2320 2304
rect 2372 2292 2378 2304
rect 2501 2295 2559 2301
rect 2501 2292 2513 2295
rect 2372 2264 2513 2292
rect 2372 2252 2378 2264
rect 2501 2261 2513 2264
rect 2547 2261 2559 2295
rect 2501 2255 2559 2261
rect 2774 2252 2780 2304
rect 2832 2292 2838 2304
rect 2961 2295 3019 2301
rect 2961 2292 2973 2295
rect 2832 2264 2973 2292
rect 2832 2252 2838 2264
rect 2961 2261 2973 2264
rect 3007 2261 3019 2295
rect 2961 2255 3019 2261
rect 3234 2252 3240 2304
rect 3292 2292 3298 2304
rect 3421 2295 3479 2301
rect 3421 2292 3433 2295
rect 3292 2264 3433 2292
rect 3292 2252 3298 2264
rect 3421 2261 3433 2264
rect 3467 2261 3479 2295
rect 3421 2255 3479 2261
rect 3694 2252 3700 2304
rect 3752 2292 3758 2304
rect 3881 2295 3939 2301
rect 3881 2292 3893 2295
rect 3752 2264 3893 2292
rect 3752 2252 3758 2264
rect 3881 2261 3893 2264
rect 3927 2261 3939 2295
rect 3881 2255 3939 2261
rect 4154 2252 4160 2304
rect 4212 2292 4218 2304
rect 4341 2295 4399 2301
rect 4341 2292 4353 2295
rect 4212 2264 4353 2292
rect 4212 2252 4218 2264
rect 4341 2261 4353 2264
rect 4387 2261 4399 2295
rect 4341 2255 4399 2261
rect 4614 2252 4620 2304
rect 4672 2292 4678 2304
rect 4801 2295 4859 2301
rect 4801 2292 4813 2295
rect 4672 2264 4813 2292
rect 4672 2252 4678 2264
rect 4801 2261 4813 2264
rect 4847 2261 4859 2295
rect 4801 2255 4859 2261
rect 5074 2252 5080 2304
rect 5132 2292 5138 2304
rect 5445 2295 5503 2301
rect 5445 2292 5457 2295
rect 5132 2264 5457 2292
rect 5132 2252 5138 2264
rect 5445 2261 5457 2264
rect 5491 2261 5503 2295
rect 5718 2292 5724 2304
rect 5679 2264 5724 2292
rect 5445 2255 5503 2261
rect 5718 2252 5724 2264
rect 5776 2252 5782 2304
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6733 2295 6791 2301
rect 6733 2292 6745 2295
rect 6512 2264 6745 2292
rect 6512 2252 6518 2264
rect 6733 2261 6745 2264
rect 6779 2261 6791 2295
rect 6733 2255 6791 2261
rect 6914 2252 6920 2304
rect 6972 2292 6978 2304
rect 7193 2295 7251 2301
rect 7193 2292 7205 2295
rect 6972 2264 7205 2292
rect 6972 2252 6978 2264
rect 7193 2261 7205 2264
rect 7239 2261 7251 2295
rect 7193 2255 7251 2261
rect 7374 2252 7380 2304
rect 7432 2292 7438 2304
rect 7653 2295 7711 2301
rect 7653 2292 7665 2295
rect 7432 2264 7665 2292
rect 7432 2252 7438 2264
rect 7653 2261 7665 2264
rect 7699 2261 7711 2295
rect 7653 2255 7711 2261
rect 7834 2252 7840 2304
rect 7892 2292 7898 2304
rect 8113 2295 8171 2301
rect 8113 2292 8125 2295
rect 7892 2264 8125 2292
rect 7892 2252 7898 2264
rect 8113 2261 8125 2264
rect 8159 2261 8171 2295
rect 8113 2255 8171 2261
rect 8294 2252 8300 2304
rect 8352 2292 8358 2304
rect 8481 2295 8539 2301
rect 8481 2292 8493 2295
rect 8352 2264 8493 2292
rect 8352 2252 8358 2264
rect 8481 2261 8493 2264
rect 8527 2261 8539 2295
rect 8481 2255 8539 2261
rect 8754 2252 8760 2304
rect 8812 2292 8818 2304
rect 9033 2295 9091 2301
rect 9033 2292 9045 2295
rect 8812 2264 9045 2292
rect 8812 2252 8818 2264
rect 9033 2261 9045 2264
rect 9079 2261 9091 2295
rect 9033 2255 9091 2261
rect 9214 2252 9220 2304
rect 9272 2292 9278 2304
rect 9401 2295 9459 2301
rect 9401 2292 9413 2295
rect 9272 2264 9413 2292
rect 9272 2252 9278 2264
rect 9401 2261 9413 2264
rect 9447 2261 9459 2295
rect 9401 2255 9459 2261
rect 9674 2252 9680 2304
rect 9732 2292 9738 2304
rect 9861 2295 9919 2301
rect 9861 2292 9873 2295
rect 9732 2264 9873 2292
rect 9732 2252 9738 2264
rect 9861 2261 9873 2264
rect 9907 2261 9919 2295
rect 9861 2255 9919 2261
rect 10226 2252 10232 2304
rect 10284 2292 10290 2304
rect 10321 2295 10379 2301
rect 10321 2292 10333 2295
rect 10284 2264 10333 2292
rect 10284 2252 10290 2264
rect 10321 2261 10333 2264
rect 10367 2261 10379 2295
rect 10321 2255 10379 2261
rect 10594 2252 10600 2304
rect 10652 2292 10658 2304
rect 10873 2295 10931 2301
rect 10873 2292 10885 2295
rect 10652 2264 10885 2292
rect 10652 2252 10658 2264
rect 10873 2261 10885 2264
rect 10919 2261 10931 2295
rect 10873 2255 10931 2261
rect 11195 2295 11253 2301
rect 11195 2261 11207 2295
rect 11241 2292 11253 2295
rect 11440 2292 11468 2332
rect 11241 2264 11468 2292
rect 11900 2292 11928 2332
rect 11974 2320 11980 2372
rect 12032 2360 12038 2372
rect 12032 2332 12077 2360
rect 12032 2320 12038 2332
rect 12250 2320 12256 2372
rect 12308 2360 12314 2372
rect 12986 2360 12992 2372
rect 12308 2332 12992 2360
rect 12308 2320 12314 2332
rect 12986 2320 12992 2332
rect 13044 2360 13050 2372
rect 13924 2360 13952 2391
rect 16114 2388 16120 2400
rect 16172 2388 16178 2440
rect 16206 2388 16212 2440
rect 16264 2428 16270 2440
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 16264 2400 16681 2428
rect 16264 2388 16270 2400
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 17034 2428 17040 2440
rect 16995 2400 17040 2428
rect 16669 2391 16727 2397
rect 17034 2388 17040 2400
rect 17092 2388 17098 2440
rect 17126 2388 17132 2440
rect 17184 2428 17190 2440
rect 17405 2431 17463 2437
rect 17405 2428 17417 2431
rect 17184 2400 17417 2428
rect 17184 2388 17190 2400
rect 17405 2397 17417 2400
rect 17451 2397 17463 2431
rect 17405 2391 17463 2397
rect 17678 2388 17684 2440
rect 17736 2428 17742 2440
rect 17773 2431 17831 2437
rect 17773 2428 17785 2431
rect 17736 2400 17785 2428
rect 17736 2388 17742 2400
rect 17773 2397 17785 2400
rect 17819 2397 17831 2431
rect 18138 2428 18144 2440
rect 18099 2400 18144 2428
rect 17773 2391 17831 2397
rect 18138 2388 18144 2400
rect 18196 2388 18202 2440
rect 13044 2332 13952 2360
rect 17052 2332 17632 2360
rect 13044 2320 13050 2332
rect 17052 2304 17080 2332
rect 13170 2292 13176 2304
rect 11900 2264 13176 2292
rect 11241 2261 11253 2264
rect 11195 2255 11253 2261
rect 13170 2252 13176 2264
rect 13228 2252 13234 2304
rect 15194 2252 15200 2304
rect 15252 2292 15258 2304
rect 16301 2295 16359 2301
rect 16301 2292 16313 2295
rect 15252 2264 16313 2292
rect 15252 2252 15258 2264
rect 16301 2261 16313 2264
rect 16347 2261 16359 2295
rect 16301 2255 16359 2261
rect 16390 2252 16396 2304
rect 16448 2292 16454 2304
rect 16853 2295 16911 2301
rect 16853 2292 16865 2295
rect 16448 2264 16865 2292
rect 16448 2252 16454 2264
rect 16853 2261 16865 2264
rect 16899 2261 16911 2295
rect 16853 2255 16911 2261
rect 17034 2252 17040 2304
rect 17092 2252 17098 2304
rect 17604 2301 17632 2332
rect 17589 2295 17647 2301
rect 17589 2261 17601 2295
rect 17635 2261 17647 2295
rect 17589 2255 17647 2261
rect 17770 2252 17776 2304
rect 17828 2292 17834 2304
rect 17957 2295 18015 2301
rect 17957 2292 17969 2295
rect 17828 2264 17969 2292
rect 17828 2252 17834 2264
rect 17957 2261 17969 2264
rect 18003 2261 18015 2295
rect 17957 2255 18015 2261
rect 18046 2252 18052 2304
rect 18104 2292 18110 2304
rect 18325 2295 18383 2301
rect 18325 2292 18337 2295
rect 18104 2264 18337 2292
rect 18104 2252 18110 2264
rect 18325 2261 18337 2264
rect 18371 2261 18383 2295
rect 18325 2255 18383 2261
rect 1104 2202 18860 2224
rect 1104 2150 5398 2202
rect 5450 2150 5462 2202
rect 5514 2150 5526 2202
rect 5578 2150 5590 2202
rect 5642 2150 5654 2202
rect 5706 2150 9846 2202
rect 9898 2150 9910 2202
rect 9962 2150 9974 2202
rect 10026 2150 10038 2202
rect 10090 2150 10102 2202
rect 10154 2150 14294 2202
rect 14346 2150 14358 2202
rect 14410 2150 14422 2202
rect 14474 2150 14486 2202
rect 14538 2150 14550 2202
rect 14602 2150 18860 2202
rect 1104 2128 18860 2150
<< via1 >>
rect 3792 15172 3844 15224
rect 4712 15172 4764 15224
rect 5908 14968 5960 15020
rect 14924 14968 14976 15020
rect 2136 14900 2188 14952
rect 7472 14900 7524 14952
rect 8760 14900 8812 14952
rect 16396 14900 16448 14952
rect 4528 14832 4580 14884
rect 3976 14764 4028 14816
rect 7012 14764 7064 14816
rect 11336 14832 11388 14884
rect 18972 14832 19024 14884
rect 12440 14764 12492 14816
rect 12624 14764 12676 14816
rect 13544 14764 13596 14816
rect 18328 14764 18380 14816
rect 3174 14662 3226 14714
rect 3238 14662 3290 14714
rect 3302 14662 3354 14714
rect 3366 14662 3418 14714
rect 3430 14662 3482 14714
rect 7622 14662 7674 14714
rect 7686 14662 7738 14714
rect 7750 14662 7802 14714
rect 7814 14662 7866 14714
rect 7878 14662 7930 14714
rect 12070 14662 12122 14714
rect 12134 14662 12186 14714
rect 12198 14662 12250 14714
rect 12262 14662 12314 14714
rect 12326 14662 12378 14714
rect 16518 14662 16570 14714
rect 16582 14662 16634 14714
rect 16646 14662 16698 14714
rect 16710 14662 16762 14714
rect 16774 14662 16826 14714
rect 3516 14560 3568 14612
rect 5540 14560 5592 14612
rect 6092 14560 6144 14612
rect 6552 14560 6604 14612
rect 6736 14560 6788 14612
rect 7380 14603 7432 14612
rect 7380 14569 7389 14603
rect 7389 14569 7423 14603
rect 7423 14569 7432 14603
rect 7380 14560 7432 14569
rect 8668 14603 8720 14612
rect 8668 14569 8677 14603
rect 8677 14569 8711 14603
rect 8711 14569 8720 14603
rect 8668 14560 8720 14569
rect 9312 14603 9364 14612
rect 9312 14569 9321 14603
rect 9321 14569 9355 14603
rect 9355 14569 9364 14603
rect 9312 14560 9364 14569
rect 9956 14603 10008 14612
rect 9956 14569 9965 14603
rect 9965 14569 9999 14603
rect 9999 14569 10008 14603
rect 9956 14560 10008 14569
rect 10600 14603 10652 14612
rect 10600 14569 10609 14603
rect 10609 14569 10643 14603
rect 10643 14569 10652 14603
rect 10600 14560 10652 14569
rect 11244 14560 11296 14612
rect 2964 14492 3016 14544
rect 6828 14492 6880 14544
rect 11060 14492 11112 14544
rect 1952 14399 2004 14408
rect 1952 14365 1961 14399
rect 1961 14365 1995 14399
rect 1995 14365 2004 14399
rect 1952 14356 2004 14365
rect 2228 14399 2280 14408
rect 2228 14365 2237 14399
rect 2237 14365 2271 14399
rect 2271 14365 2280 14399
rect 2228 14356 2280 14365
rect 3976 14424 4028 14476
rect 4160 14424 4212 14476
rect 6184 14424 6236 14476
rect 3608 14399 3660 14408
rect 3608 14365 3617 14399
rect 3617 14365 3651 14399
rect 3651 14365 3660 14399
rect 3608 14356 3660 14365
rect 4436 14356 4488 14408
rect 4712 14399 4764 14408
rect 4712 14365 4721 14399
rect 4721 14365 4755 14399
rect 4755 14365 4764 14399
rect 4712 14356 4764 14365
rect 4988 14399 5040 14408
rect 4988 14365 4997 14399
rect 4997 14365 5031 14399
rect 5031 14365 5040 14399
rect 4988 14356 5040 14365
rect 5908 14399 5960 14408
rect 5908 14365 5917 14399
rect 5917 14365 5951 14399
rect 5951 14365 5960 14399
rect 5908 14356 5960 14365
rect 6552 14399 6604 14408
rect 6552 14365 6561 14399
rect 6561 14365 6595 14399
rect 6595 14365 6604 14399
rect 6552 14356 6604 14365
rect 7380 14356 7432 14408
rect 8668 14356 8720 14408
rect 9312 14356 9364 14408
rect 9956 14356 10008 14408
rect 10600 14356 10652 14408
rect 12532 14603 12584 14612
rect 12532 14569 12541 14603
rect 12541 14569 12575 14603
rect 12575 14569 12584 14603
rect 12532 14560 12584 14569
rect 13176 14603 13228 14612
rect 13176 14569 13185 14603
rect 13185 14569 13219 14603
rect 13219 14569 13228 14603
rect 13176 14560 13228 14569
rect 15292 14492 15344 14544
rect 12900 14424 12952 14476
rect 14188 14424 14240 14476
rect 16764 14467 16816 14476
rect 16764 14433 16773 14467
rect 16773 14433 16807 14467
rect 16807 14433 16816 14467
rect 16764 14424 16816 14433
rect 11980 14399 12032 14408
rect 11980 14365 11989 14399
rect 11989 14365 12023 14399
rect 12023 14365 12032 14399
rect 11980 14356 12032 14365
rect 12532 14356 12584 14408
rect 13176 14356 13228 14408
rect 13820 14356 13872 14408
rect 15476 14356 15528 14408
rect 16028 14356 16080 14408
rect 16304 14356 16356 14408
rect 16948 14356 17000 14408
rect 17224 14356 17276 14408
rect 17684 14399 17736 14408
rect 17684 14365 17693 14399
rect 17693 14365 17727 14399
rect 17727 14365 17736 14399
rect 17684 14356 17736 14365
rect 17960 14399 18012 14408
rect 17960 14365 17969 14399
rect 17969 14365 18003 14399
rect 18003 14365 18012 14399
rect 17960 14356 18012 14365
rect 4252 14288 4304 14340
rect 5172 14288 5224 14340
rect 3148 14220 3200 14272
rect 5816 14220 5868 14272
rect 6368 14263 6420 14272
rect 6368 14229 6377 14263
rect 6377 14229 6411 14263
rect 6411 14229 6420 14263
rect 6368 14220 6420 14229
rect 13360 14288 13412 14340
rect 8116 14220 8168 14272
rect 8668 14220 8720 14272
rect 9036 14220 9088 14272
rect 10692 14263 10744 14272
rect 10692 14229 10701 14263
rect 10701 14229 10735 14263
rect 10735 14229 10744 14263
rect 10692 14220 10744 14229
rect 11428 14220 11480 14272
rect 11796 14220 11848 14272
rect 12716 14220 12768 14272
rect 13728 14220 13780 14272
rect 15384 14263 15436 14272
rect 15384 14229 15393 14263
rect 15393 14229 15427 14263
rect 15427 14229 15436 14263
rect 15384 14220 15436 14229
rect 5398 14118 5450 14170
rect 5462 14118 5514 14170
rect 5526 14118 5578 14170
rect 5590 14118 5642 14170
rect 5654 14118 5706 14170
rect 9846 14118 9898 14170
rect 9910 14118 9962 14170
rect 9974 14118 10026 14170
rect 10038 14118 10090 14170
rect 10102 14118 10154 14170
rect 14294 14118 14346 14170
rect 14358 14118 14410 14170
rect 14422 14118 14474 14170
rect 14486 14118 14538 14170
rect 14550 14118 14602 14170
rect 2780 14016 2832 14068
rect 3056 14016 3108 14068
rect 3516 14016 3568 14068
rect 4344 14059 4396 14068
rect 4344 14025 4353 14059
rect 4353 14025 4387 14059
rect 4387 14025 4396 14059
rect 4344 14016 4396 14025
rect 4712 14059 4764 14068
rect 4712 14025 4721 14059
rect 4721 14025 4755 14059
rect 4755 14025 4764 14059
rect 4712 14016 4764 14025
rect 4804 14016 4856 14068
rect 2044 13948 2096 14000
rect 6276 14016 6328 14068
rect 6460 14016 6512 14068
rect 6644 14016 6696 14068
rect 2136 13880 2188 13932
rect 3700 13880 3752 13932
rect 4068 13923 4120 13932
rect 4068 13889 4077 13923
rect 4077 13889 4111 13923
rect 4111 13889 4120 13923
rect 4068 13880 4120 13889
rect 4528 13923 4580 13932
rect 4528 13889 4537 13923
rect 4537 13889 4571 13923
rect 4571 13889 4580 13923
rect 4528 13880 4580 13889
rect 5172 13923 5224 13932
rect 5172 13889 5181 13923
rect 5181 13889 5215 13923
rect 5215 13889 5224 13923
rect 5172 13880 5224 13889
rect 5540 13923 5592 13932
rect 5540 13889 5549 13923
rect 5549 13889 5583 13923
rect 5583 13889 5592 13923
rect 5540 13880 5592 13889
rect 5816 13923 5868 13932
rect 5816 13889 5825 13923
rect 5825 13889 5859 13923
rect 5859 13889 5868 13923
rect 5816 13880 5868 13889
rect 3148 13855 3200 13864
rect 3148 13821 3157 13855
rect 3157 13821 3191 13855
rect 3191 13821 3200 13855
rect 3148 13812 3200 13821
rect 3608 13812 3660 13864
rect 940 13744 992 13796
rect 5448 13812 5500 13864
rect 6552 13880 6604 13932
rect 7012 13923 7064 13932
rect 7012 13889 7021 13923
rect 7021 13889 7055 13923
rect 7055 13889 7064 13923
rect 7012 13880 7064 13889
rect 6184 13787 6236 13796
rect 1952 13676 2004 13728
rect 3976 13676 4028 13728
rect 4068 13676 4120 13728
rect 6184 13753 6193 13787
rect 6193 13753 6227 13787
rect 6227 13753 6236 13787
rect 6184 13744 6236 13753
rect 6368 13744 6420 13796
rect 6736 13744 6788 13796
rect 6828 13676 6880 13728
rect 8760 14016 8812 14068
rect 11152 14016 11204 14068
rect 11704 14016 11756 14068
rect 12440 14016 12492 14068
rect 13268 14059 13320 14068
rect 13268 14025 13277 14059
rect 13277 14025 13311 14059
rect 13311 14025 13320 14059
rect 13268 14016 13320 14025
rect 11336 13948 11388 14000
rect 12624 13948 12676 14000
rect 12900 13880 12952 13932
rect 14924 14059 14976 14068
rect 14924 14025 14933 14059
rect 14933 14025 14967 14059
rect 14967 14025 14976 14059
rect 14924 14016 14976 14025
rect 15844 13948 15896 14000
rect 15016 13880 15068 13932
rect 15752 13880 15804 13932
rect 16212 13923 16264 13932
rect 16212 13889 16221 13923
rect 16221 13889 16255 13923
rect 16255 13889 16264 13923
rect 16212 13880 16264 13889
rect 16488 13923 16540 13932
rect 16488 13889 16497 13923
rect 16497 13889 16531 13923
rect 16531 13889 16540 13923
rect 16488 13880 16540 13889
rect 9496 13812 9548 13864
rect 11888 13812 11940 13864
rect 16764 13855 16816 13864
rect 16764 13821 16773 13855
rect 16773 13821 16807 13855
rect 16807 13821 16816 13855
rect 16764 13812 16816 13821
rect 7840 13787 7892 13796
rect 7840 13753 7849 13787
rect 7849 13753 7883 13787
rect 7883 13753 7892 13787
rect 7840 13744 7892 13753
rect 9680 13744 9732 13796
rect 16120 13744 16172 13796
rect 17776 13812 17828 13864
rect 8300 13676 8352 13728
rect 9864 13719 9916 13728
rect 9864 13685 9873 13719
rect 9873 13685 9907 13719
rect 9907 13685 9916 13719
rect 9864 13676 9916 13685
rect 13360 13676 13412 13728
rect 16304 13719 16356 13728
rect 16304 13685 16313 13719
rect 16313 13685 16347 13719
rect 16347 13685 16356 13719
rect 16304 13676 16356 13685
rect 16764 13676 16816 13728
rect 17040 13676 17092 13728
rect 3174 13574 3226 13626
rect 3238 13574 3290 13626
rect 3302 13574 3354 13626
rect 3366 13574 3418 13626
rect 3430 13574 3482 13626
rect 7622 13574 7674 13626
rect 7686 13574 7738 13626
rect 7750 13574 7802 13626
rect 7814 13574 7866 13626
rect 7878 13574 7930 13626
rect 12070 13574 12122 13626
rect 12134 13574 12186 13626
rect 12198 13574 12250 13626
rect 12262 13574 12314 13626
rect 12326 13574 12378 13626
rect 16518 13574 16570 13626
rect 16582 13574 16634 13626
rect 16646 13574 16698 13626
rect 16710 13574 16762 13626
rect 16774 13574 16826 13626
rect 2872 13472 2924 13524
rect 3516 13472 3568 13524
rect 2504 13404 2556 13456
rect 4160 13404 4212 13456
rect 7196 13472 7248 13524
rect 6276 13404 6328 13456
rect 1952 13379 2004 13388
rect 1952 13345 1961 13379
rect 1961 13345 1995 13379
rect 1995 13345 2004 13379
rect 1952 13336 2004 13345
rect 2780 13268 2832 13320
rect 2872 13311 2924 13320
rect 2872 13277 2881 13311
rect 2881 13277 2915 13311
rect 2915 13277 2924 13311
rect 2872 13268 2924 13277
rect 296 13200 348 13252
rect 3148 13311 3200 13320
rect 3148 13277 3157 13311
rect 3157 13277 3191 13311
rect 3191 13277 3200 13311
rect 3516 13311 3568 13320
rect 3148 13268 3200 13277
rect 3516 13277 3525 13311
rect 3525 13277 3559 13311
rect 3559 13277 3568 13311
rect 3516 13268 3568 13277
rect 4068 13311 4120 13320
rect 4068 13277 4077 13311
rect 4077 13277 4111 13311
rect 4111 13277 4120 13311
rect 4068 13268 4120 13277
rect 1584 13132 1636 13184
rect 3424 13132 3476 13184
rect 4160 13132 4212 13184
rect 5448 13336 5500 13388
rect 5724 13379 5776 13388
rect 5724 13345 5733 13379
rect 5733 13345 5767 13379
rect 5767 13345 5776 13379
rect 5724 13336 5776 13345
rect 6000 13336 6052 13388
rect 7748 13336 7800 13388
rect 6644 13268 6696 13320
rect 7196 13268 7248 13320
rect 9404 13336 9456 13388
rect 11980 13336 12032 13388
rect 12348 13472 12400 13524
rect 13820 13472 13872 13524
rect 16856 13472 16908 13524
rect 17684 13404 17736 13456
rect 12440 13379 12492 13388
rect 12440 13345 12449 13379
rect 12449 13345 12483 13379
rect 12483 13345 12492 13379
rect 12440 13336 12492 13345
rect 5172 13175 5224 13184
rect 5172 13141 5181 13175
rect 5181 13141 5215 13175
rect 5215 13141 5224 13175
rect 5172 13132 5224 13141
rect 6276 13132 6328 13184
rect 6920 13200 6972 13252
rect 7196 13175 7248 13184
rect 7196 13141 7205 13175
rect 7205 13141 7239 13175
rect 7239 13141 7248 13175
rect 7196 13132 7248 13141
rect 8392 13132 8444 13184
rect 12348 13268 12400 13320
rect 16120 13336 16172 13388
rect 16948 13336 17000 13388
rect 17684 13311 17736 13320
rect 17684 13277 17693 13311
rect 17693 13277 17727 13311
rect 17727 13277 17736 13311
rect 17684 13268 17736 13277
rect 18052 13268 18104 13320
rect 16580 13200 16632 13252
rect 17132 13243 17184 13252
rect 17132 13209 17141 13243
rect 17141 13209 17175 13243
rect 17175 13209 17184 13243
rect 17132 13200 17184 13209
rect 17592 13200 17644 13252
rect 9680 13175 9732 13184
rect 9680 13141 9689 13175
rect 9689 13141 9723 13175
rect 9723 13141 9732 13175
rect 9680 13132 9732 13141
rect 11152 13132 11204 13184
rect 11336 13175 11388 13184
rect 11336 13141 11345 13175
rect 11345 13141 11379 13175
rect 11379 13141 11388 13175
rect 11336 13132 11388 13141
rect 11888 13132 11940 13184
rect 12624 13175 12676 13184
rect 12624 13141 12633 13175
rect 12633 13141 12667 13175
rect 12667 13141 12676 13175
rect 12624 13132 12676 13141
rect 13820 13175 13872 13184
rect 13820 13141 13829 13175
rect 13829 13141 13863 13175
rect 13863 13141 13872 13175
rect 13820 13132 13872 13141
rect 15200 13132 15252 13184
rect 17040 13175 17092 13184
rect 17040 13141 17049 13175
rect 17049 13141 17083 13175
rect 17083 13141 17092 13175
rect 17040 13132 17092 13141
rect 17408 13175 17460 13184
rect 17408 13141 17417 13175
rect 17417 13141 17451 13175
rect 17451 13141 17460 13175
rect 17408 13132 17460 13141
rect 5398 13030 5450 13082
rect 5462 13030 5514 13082
rect 5526 13030 5578 13082
rect 5590 13030 5642 13082
rect 5654 13030 5706 13082
rect 9846 13030 9898 13082
rect 9910 13030 9962 13082
rect 9974 13030 10026 13082
rect 10038 13030 10090 13082
rect 10102 13030 10154 13082
rect 14294 13030 14346 13082
rect 14358 13030 14410 13082
rect 14422 13030 14474 13082
rect 14486 13030 14538 13082
rect 14550 13030 14602 13082
rect 2872 12928 2924 12980
rect 2964 12792 3016 12844
rect 3424 12835 3476 12844
rect 3424 12801 3433 12835
rect 3433 12801 3467 12835
rect 3467 12801 3476 12835
rect 3424 12792 3476 12801
rect 4988 12928 5040 12980
rect 5172 12971 5224 12980
rect 5172 12937 5181 12971
rect 5181 12937 5215 12971
rect 5215 12937 5224 12971
rect 5172 12928 5224 12937
rect 2136 12724 2188 12776
rect 2228 12767 2280 12776
rect 2228 12733 2237 12767
rect 2237 12733 2271 12767
rect 2271 12733 2280 12767
rect 2228 12724 2280 12733
rect 2780 12724 2832 12776
rect 3516 12724 3568 12776
rect 4068 12767 4120 12776
rect 4068 12733 4077 12767
rect 4077 12733 4111 12767
rect 4111 12733 4120 12767
rect 5356 12860 5408 12912
rect 7196 12928 7248 12980
rect 11336 12928 11388 12980
rect 12624 12928 12676 12980
rect 17776 12928 17828 12980
rect 6920 12860 6972 12912
rect 7012 12860 7064 12912
rect 16948 12903 17000 12912
rect 6276 12792 6328 12844
rect 9128 12835 9180 12844
rect 9128 12801 9137 12835
rect 9137 12801 9171 12835
rect 9171 12801 9180 12835
rect 9128 12792 9180 12801
rect 5264 12767 5316 12776
rect 4068 12724 4120 12733
rect 5264 12733 5273 12767
rect 5273 12733 5307 12767
rect 5307 12733 5316 12767
rect 5264 12724 5316 12733
rect 3884 12656 3936 12708
rect 3056 12588 3108 12640
rect 3516 12631 3568 12640
rect 3516 12597 3525 12631
rect 3525 12597 3559 12631
rect 3559 12597 3568 12631
rect 3516 12588 3568 12597
rect 3792 12588 3844 12640
rect 4160 12588 4212 12640
rect 4712 12588 4764 12640
rect 5172 12656 5224 12708
rect 7380 12724 7432 12776
rect 7748 12724 7800 12776
rect 6736 12656 6788 12708
rect 10232 12767 10284 12776
rect 10232 12733 10241 12767
rect 10241 12733 10275 12767
rect 10275 12733 10284 12767
rect 10232 12724 10284 12733
rect 12348 12792 12400 12844
rect 12992 12792 13044 12844
rect 16948 12869 16957 12903
rect 16957 12869 16991 12903
rect 16991 12869 17000 12903
rect 16948 12860 17000 12869
rect 17132 12860 17184 12912
rect 17592 12903 17644 12912
rect 17592 12869 17601 12903
rect 17601 12869 17635 12903
rect 17635 12869 17644 12903
rect 17592 12860 17644 12869
rect 12164 12724 12216 12776
rect 12440 12724 12492 12776
rect 13360 12724 13412 12776
rect 13176 12656 13228 12708
rect 6644 12588 6696 12640
rect 12440 12588 12492 12640
rect 15200 12792 15252 12844
rect 16212 12792 16264 12844
rect 16580 12792 16632 12844
rect 17500 12792 17552 12844
rect 14464 12767 14516 12776
rect 14464 12733 14473 12767
rect 14473 12733 14507 12767
rect 14507 12733 14516 12767
rect 14464 12724 14516 12733
rect 17776 12724 17828 12776
rect 18236 12724 18288 12776
rect 15844 12656 15896 12708
rect 19616 12656 19668 12708
rect 16856 12588 16908 12640
rect 3174 12486 3226 12538
rect 3238 12486 3290 12538
rect 3302 12486 3354 12538
rect 3366 12486 3418 12538
rect 3430 12486 3482 12538
rect 7622 12486 7674 12538
rect 7686 12486 7738 12538
rect 7750 12486 7802 12538
rect 7814 12486 7866 12538
rect 7878 12486 7930 12538
rect 12070 12486 12122 12538
rect 12134 12486 12186 12538
rect 12198 12486 12250 12538
rect 12262 12486 12314 12538
rect 12326 12486 12378 12538
rect 16518 12486 16570 12538
rect 16582 12486 16634 12538
rect 16646 12486 16698 12538
rect 16710 12486 16762 12538
rect 16774 12486 16826 12538
rect 2964 12384 3016 12436
rect 7196 12384 7248 12436
rect 7472 12384 7524 12436
rect 9128 12384 9180 12436
rect 12808 12427 12860 12436
rect 12808 12393 12817 12427
rect 12817 12393 12851 12427
rect 12851 12393 12860 12427
rect 12808 12384 12860 12393
rect 12992 12384 13044 12436
rect 17960 12384 18012 12436
rect 18144 12384 18196 12436
rect 5908 12316 5960 12368
rect 10416 12316 10468 12368
rect 4068 12248 4120 12300
rect 6552 12248 6604 12300
rect 10232 12291 10284 12300
rect 2780 12180 2832 12232
rect 7104 12180 7156 12232
rect 7380 12180 7432 12232
rect 10232 12257 10241 12291
rect 10241 12257 10275 12291
rect 10275 12257 10284 12291
rect 10232 12248 10284 12257
rect 2412 12155 2464 12164
rect 2412 12121 2421 12155
rect 2421 12121 2455 12155
rect 2455 12121 2464 12155
rect 2412 12112 2464 12121
rect 3148 12155 3200 12164
rect 3148 12121 3157 12155
rect 3157 12121 3191 12155
rect 3191 12121 3200 12155
rect 3148 12112 3200 12121
rect 3884 12112 3936 12164
rect 4988 12112 5040 12164
rect 2504 12087 2556 12096
rect 2504 12053 2513 12087
rect 2513 12053 2547 12087
rect 2547 12053 2556 12087
rect 2504 12044 2556 12053
rect 3332 12044 3384 12096
rect 4344 12044 4396 12096
rect 4896 12087 4948 12096
rect 4896 12053 4905 12087
rect 4905 12053 4939 12087
rect 4939 12053 4948 12087
rect 6092 12087 6144 12096
rect 4896 12044 4948 12053
rect 6092 12053 6101 12087
rect 6101 12053 6135 12087
rect 6135 12053 6144 12087
rect 6092 12044 6144 12053
rect 7012 12044 7064 12096
rect 7932 12112 7984 12164
rect 11336 12248 11388 12300
rect 12348 12248 12400 12300
rect 12440 12291 12492 12300
rect 12440 12257 12449 12291
rect 12449 12257 12483 12291
rect 12483 12257 12492 12291
rect 12440 12248 12492 12257
rect 13360 12291 13412 12300
rect 11244 12223 11296 12232
rect 11244 12189 11253 12223
rect 11253 12189 11287 12223
rect 11287 12189 11296 12223
rect 11244 12180 11296 12189
rect 13360 12257 13369 12291
rect 13369 12257 13403 12291
rect 13403 12257 13412 12291
rect 13360 12248 13412 12257
rect 17224 12316 17276 12368
rect 18696 12316 18748 12368
rect 14648 12291 14700 12300
rect 14648 12257 14657 12291
rect 14657 12257 14691 12291
rect 14691 12257 14700 12291
rect 14648 12248 14700 12257
rect 15200 12180 15252 12232
rect 17868 12180 17920 12232
rect 17960 12223 18012 12232
rect 17960 12189 17969 12223
rect 17969 12189 18003 12223
rect 18003 12189 18012 12223
rect 17960 12180 18012 12189
rect 8116 12087 8168 12096
rect 8116 12053 8125 12087
rect 8125 12053 8159 12087
rect 8159 12053 8168 12087
rect 8116 12044 8168 12053
rect 12808 12112 12860 12164
rect 13176 12087 13228 12096
rect 13176 12053 13185 12087
rect 13185 12053 13219 12087
rect 13219 12053 13228 12087
rect 13176 12044 13228 12053
rect 13268 12087 13320 12096
rect 13268 12053 13277 12087
rect 13277 12053 13311 12087
rect 13311 12053 13320 12087
rect 13268 12044 13320 12053
rect 15936 12044 15988 12096
rect 16028 12044 16080 12096
rect 17592 12044 17644 12096
rect 17684 12044 17736 12096
rect 5398 11942 5450 11994
rect 5462 11942 5514 11994
rect 5526 11942 5578 11994
rect 5590 11942 5642 11994
rect 5654 11942 5706 11994
rect 9846 11942 9898 11994
rect 9910 11942 9962 11994
rect 9974 11942 10026 11994
rect 10038 11942 10090 11994
rect 10102 11942 10154 11994
rect 14294 11942 14346 11994
rect 14358 11942 14410 11994
rect 14422 11942 14474 11994
rect 14486 11942 14538 11994
rect 14550 11942 14602 11994
rect 2412 11840 2464 11892
rect 3332 11883 3384 11892
rect 3056 11772 3108 11824
rect 3332 11849 3341 11883
rect 3341 11849 3375 11883
rect 3375 11849 3384 11883
rect 3332 11840 3384 11849
rect 3516 11840 3568 11892
rect 4344 11883 4396 11892
rect 4344 11849 4353 11883
rect 4353 11849 4387 11883
rect 4387 11849 4396 11883
rect 4344 11840 4396 11849
rect 4896 11840 4948 11892
rect 5908 11883 5960 11892
rect 5908 11849 5917 11883
rect 5917 11849 5951 11883
rect 5951 11849 5960 11883
rect 5908 11840 5960 11849
rect 4160 11772 4212 11824
rect 6092 11772 6144 11824
rect 6460 11815 6512 11824
rect 6460 11781 6469 11815
rect 6469 11781 6503 11815
rect 6503 11781 6512 11815
rect 6460 11772 6512 11781
rect 6644 11772 6696 11824
rect 8392 11840 8444 11892
rect 8484 11840 8536 11892
rect 9680 11840 9732 11892
rect 10968 11840 11020 11892
rect 13268 11840 13320 11892
rect 13636 11840 13688 11892
rect 18144 11840 18196 11892
rect 15200 11772 15252 11824
rect 15936 11815 15988 11824
rect 15936 11781 15945 11815
rect 15945 11781 15979 11815
rect 15979 11781 15988 11815
rect 15936 11772 15988 11781
rect 17224 11815 17276 11824
rect 17224 11781 17233 11815
rect 17233 11781 17267 11815
rect 17267 11781 17276 11815
rect 17224 11772 17276 11781
rect 2228 11679 2280 11688
rect 2228 11645 2237 11679
rect 2237 11645 2271 11679
rect 2271 11645 2280 11679
rect 2228 11636 2280 11645
rect 5724 11704 5776 11756
rect 7012 11747 7064 11756
rect 7012 11713 7021 11747
rect 7021 11713 7055 11747
rect 7055 11713 7064 11747
rect 7012 11704 7064 11713
rect 3424 11636 3476 11688
rect 4528 11679 4580 11688
rect 4528 11645 4537 11679
rect 4537 11645 4571 11679
rect 4571 11645 4580 11679
rect 4528 11636 4580 11645
rect 7380 11704 7432 11756
rect 9772 11704 9824 11756
rect 12716 11747 12768 11756
rect 12716 11713 12725 11747
rect 12725 11713 12759 11747
rect 12759 11713 12768 11747
rect 13268 11747 13320 11756
rect 12716 11704 12768 11713
rect 13268 11713 13277 11747
rect 13277 11713 13311 11747
rect 13311 11713 13320 11747
rect 13268 11704 13320 11713
rect 14556 11704 14608 11756
rect 7196 11679 7248 11688
rect 7196 11645 7205 11679
rect 7205 11645 7239 11679
rect 7239 11645 7248 11679
rect 7196 11636 7248 11645
rect 5264 11568 5316 11620
rect 7104 11568 7156 11620
rect 8392 11568 8444 11620
rect 9404 11679 9456 11688
rect 9404 11645 9413 11679
rect 9413 11645 9447 11679
rect 9447 11645 9456 11679
rect 10048 11679 10100 11688
rect 9404 11636 9456 11645
rect 10048 11645 10057 11679
rect 10057 11645 10091 11679
rect 10091 11645 10100 11679
rect 10048 11636 10100 11645
rect 10232 11679 10284 11688
rect 10232 11645 10241 11679
rect 10241 11645 10275 11679
rect 10275 11645 10284 11679
rect 10232 11636 10284 11645
rect 12624 11636 12676 11688
rect 14648 11636 14700 11688
rect 16028 11679 16080 11688
rect 8852 11568 8904 11620
rect 1860 11500 1912 11552
rect 2596 11543 2648 11552
rect 2596 11509 2605 11543
rect 2605 11509 2639 11543
rect 2639 11509 2648 11543
rect 2596 11500 2648 11509
rect 2964 11543 3016 11552
rect 2964 11509 2973 11543
rect 2973 11509 3007 11543
rect 3007 11509 3016 11543
rect 2964 11500 3016 11509
rect 3424 11500 3476 11552
rect 3700 11500 3752 11552
rect 3976 11543 4028 11552
rect 3976 11509 3985 11543
rect 3985 11509 4019 11543
rect 4019 11509 4028 11543
rect 3976 11500 4028 11509
rect 5448 11500 5500 11552
rect 7932 11500 7984 11552
rect 9128 11500 9180 11552
rect 13084 11568 13136 11620
rect 16028 11645 16037 11679
rect 16037 11645 16071 11679
rect 16071 11645 16080 11679
rect 16028 11636 16080 11645
rect 17592 11704 17644 11756
rect 18420 11704 18472 11756
rect 17316 11636 17368 11688
rect 17684 11679 17736 11688
rect 17684 11645 17693 11679
rect 17693 11645 17727 11679
rect 17727 11645 17736 11679
rect 17684 11636 17736 11645
rect 18880 11636 18932 11688
rect 9864 11500 9916 11552
rect 13176 11500 13228 11552
rect 14556 11543 14608 11552
rect 14556 11509 14565 11543
rect 14565 11509 14599 11543
rect 14599 11509 14608 11543
rect 14556 11500 14608 11509
rect 15016 11500 15068 11552
rect 15384 11500 15436 11552
rect 15568 11543 15620 11552
rect 15568 11509 15577 11543
rect 15577 11509 15611 11543
rect 15611 11509 15620 11543
rect 15568 11500 15620 11509
rect 16856 11500 16908 11552
rect 3174 11398 3226 11450
rect 3238 11398 3290 11450
rect 3302 11398 3354 11450
rect 3366 11398 3418 11450
rect 3430 11398 3482 11450
rect 7622 11398 7674 11450
rect 7686 11398 7738 11450
rect 7750 11398 7802 11450
rect 7814 11398 7866 11450
rect 7878 11398 7930 11450
rect 12070 11398 12122 11450
rect 12134 11398 12186 11450
rect 12198 11398 12250 11450
rect 12262 11398 12314 11450
rect 12326 11398 12378 11450
rect 16518 11398 16570 11450
rect 16582 11398 16634 11450
rect 16646 11398 16698 11450
rect 16710 11398 16762 11450
rect 16774 11398 16826 11450
rect 1308 11228 1360 11280
rect 1952 11203 2004 11212
rect 1952 11169 1961 11203
rect 1961 11169 1995 11203
rect 1995 11169 2004 11203
rect 1952 11160 2004 11169
rect 2228 11135 2280 11144
rect 2228 11101 2237 11135
rect 2237 11101 2271 11135
rect 2271 11101 2280 11135
rect 2228 11092 2280 11101
rect 2872 11296 2924 11348
rect 4804 11296 4856 11348
rect 7012 11296 7064 11348
rect 8576 11296 8628 11348
rect 3608 11228 3660 11280
rect 8116 11228 8168 11280
rect 3976 11160 4028 11212
rect 7012 11160 7064 11212
rect 8852 11228 8904 11280
rect 2964 11135 3016 11144
rect 2964 11101 2973 11135
rect 2973 11101 3007 11135
rect 3007 11101 3016 11135
rect 2964 11092 3016 11101
rect 3148 11092 3200 11144
rect 3516 11135 3568 11144
rect 3516 11101 3525 11135
rect 3525 11101 3559 11135
rect 3559 11101 3568 11135
rect 3516 11092 3568 11101
rect 3700 11092 3752 11144
rect 4528 11092 4580 11144
rect 6000 11092 6052 11144
rect 7472 11092 7524 11144
rect 8116 11092 8168 11144
rect 8484 11092 8536 11144
rect 9864 11228 9916 11280
rect 9220 11160 9272 11212
rect 9772 11203 9824 11212
rect 9772 11169 9781 11203
rect 9781 11169 9815 11203
rect 9815 11169 9824 11203
rect 9772 11160 9824 11169
rect 3976 11024 4028 11076
rect 7288 11024 7340 11076
rect 9128 11092 9180 11144
rect 15476 11296 15528 11348
rect 15752 11296 15804 11348
rect 17040 11228 17092 11280
rect 17592 11228 17644 11280
rect 14740 11203 14792 11212
rect 14740 11169 14749 11203
rect 14749 11169 14783 11203
rect 14783 11169 14792 11203
rect 14740 11160 14792 11169
rect 15384 11203 15436 11212
rect 15384 11169 15393 11203
rect 15393 11169 15427 11203
rect 15427 11169 15436 11203
rect 15384 11160 15436 11169
rect 15476 11203 15528 11212
rect 15476 11169 15485 11203
rect 15485 11169 15519 11203
rect 15519 11169 15528 11203
rect 15476 11160 15528 11169
rect 10968 11092 11020 11144
rect 11244 11092 11296 11144
rect 11520 11092 11572 11144
rect 2780 10956 2832 11008
rect 5448 10956 5500 11008
rect 8760 11024 8812 11076
rect 15200 11092 15252 11144
rect 15568 11092 15620 11144
rect 10324 10956 10376 11008
rect 13636 11024 13688 11076
rect 14648 11024 14700 11076
rect 13084 10999 13136 11008
rect 13084 10965 13093 10999
rect 13093 10965 13127 10999
rect 13127 10965 13136 10999
rect 15108 11024 15160 11076
rect 16856 11092 16908 11144
rect 17132 11135 17184 11144
rect 17132 11101 17141 11135
rect 17141 11101 17175 11135
rect 17175 11101 17184 11135
rect 17132 11092 17184 11101
rect 17500 11092 17552 11144
rect 17684 11135 17736 11144
rect 17684 11101 17693 11135
rect 17693 11101 17727 11135
rect 17727 11101 17736 11135
rect 17684 11092 17736 11101
rect 17960 11135 18012 11144
rect 17960 11101 17969 11135
rect 17969 11101 18003 11135
rect 18003 11101 18012 11135
rect 17960 11092 18012 11101
rect 16396 11024 16448 11076
rect 14924 10999 14976 11008
rect 13084 10956 13136 10965
rect 14924 10965 14933 10999
rect 14933 10965 14967 10999
rect 14967 10965 14976 10999
rect 14924 10956 14976 10965
rect 18604 11024 18656 11076
rect 18052 10956 18104 11008
rect 5398 10854 5450 10906
rect 5462 10854 5514 10906
rect 5526 10854 5578 10906
rect 5590 10854 5642 10906
rect 5654 10854 5706 10906
rect 9846 10854 9898 10906
rect 9910 10854 9962 10906
rect 9974 10854 10026 10906
rect 10038 10854 10090 10906
rect 10102 10854 10154 10906
rect 14294 10854 14346 10906
rect 14358 10854 14410 10906
rect 14422 10854 14474 10906
rect 14486 10854 14538 10906
rect 14550 10854 14602 10906
rect 1584 10752 1636 10804
rect 2780 10752 2832 10804
rect 3700 10752 3752 10804
rect 3148 10616 3200 10668
rect 2228 10591 2280 10600
rect 2228 10557 2237 10591
rect 2237 10557 2271 10591
rect 2271 10557 2280 10591
rect 2228 10548 2280 10557
rect 3516 10616 3568 10668
rect 5724 10684 5776 10736
rect 7196 10684 7248 10736
rect 6092 10616 6144 10668
rect 2136 10480 2188 10532
rect 3056 10480 3108 10532
rect 4436 10548 4488 10600
rect 9220 10752 9272 10804
rect 8116 10684 8168 10736
rect 10324 10684 10376 10736
rect 11612 10752 11664 10804
rect 11980 10752 12032 10804
rect 14648 10795 14700 10804
rect 14648 10761 14657 10795
rect 14657 10761 14691 10795
rect 14691 10761 14700 10795
rect 14648 10752 14700 10761
rect 17040 10795 17092 10804
rect 17040 10761 17049 10795
rect 17049 10761 17083 10795
rect 17083 10761 17092 10795
rect 17040 10752 17092 10761
rect 17960 10752 18012 10804
rect 13360 10684 13412 10736
rect 15200 10684 15252 10736
rect 2504 10412 2556 10464
rect 2688 10412 2740 10464
rect 4160 10455 4212 10464
rect 4160 10421 4169 10455
rect 4169 10421 4203 10455
rect 4203 10421 4212 10455
rect 4160 10412 4212 10421
rect 5264 10412 5316 10464
rect 11612 10616 11664 10668
rect 12624 10659 12676 10668
rect 12624 10625 12642 10659
rect 12642 10625 12676 10659
rect 14464 10659 14516 10668
rect 12624 10616 12676 10625
rect 14464 10625 14473 10659
rect 14473 10625 14507 10659
rect 14507 10625 14516 10659
rect 14464 10616 14516 10625
rect 9680 10591 9732 10600
rect 9680 10557 9689 10591
rect 9689 10557 9723 10591
rect 9723 10557 9732 10591
rect 9680 10548 9732 10557
rect 12900 10591 12952 10600
rect 12900 10557 12909 10591
rect 12909 10557 12943 10591
rect 12943 10557 12952 10591
rect 12900 10548 12952 10557
rect 15108 10548 15160 10600
rect 17132 10591 17184 10600
rect 10876 10480 10928 10532
rect 17132 10557 17141 10591
rect 17141 10557 17175 10591
rect 17175 10557 17184 10591
rect 17132 10548 17184 10557
rect 17316 10548 17368 10600
rect 17684 10591 17736 10600
rect 17684 10557 17693 10591
rect 17693 10557 17727 10591
rect 17727 10557 17736 10591
rect 17684 10548 17736 10557
rect 18328 10548 18380 10600
rect 8392 10412 8444 10464
rect 10600 10412 10652 10464
rect 11244 10455 11296 10464
rect 11244 10421 11253 10455
rect 11253 10421 11287 10455
rect 11287 10421 11296 10455
rect 11244 10412 11296 10421
rect 3174 10310 3226 10362
rect 3238 10310 3290 10362
rect 3302 10310 3354 10362
rect 3366 10310 3418 10362
rect 3430 10310 3482 10362
rect 7622 10310 7674 10362
rect 7686 10310 7738 10362
rect 7750 10310 7802 10362
rect 7814 10310 7866 10362
rect 7878 10310 7930 10362
rect 12070 10310 12122 10362
rect 12134 10310 12186 10362
rect 12198 10310 12250 10362
rect 12262 10310 12314 10362
rect 12326 10310 12378 10362
rect 16518 10310 16570 10362
rect 16582 10310 16634 10362
rect 16646 10310 16698 10362
rect 16710 10310 16762 10362
rect 16774 10310 16826 10362
rect 1584 10251 1636 10260
rect 1584 10217 1593 10251
rect 1593 10217 1627 10251
rect 1627 10217 1636 10251
rect 1584 10208 1636 10217
rect 2228 10208 2280 10260
rect 4160 10208 4212 10260
rect 3056 10140 3108 10192
rect 2504 10115 2556 10124
rect 2504 10081 2513 10115
rect 2513 10081 2547 10115
rect 2547 10081 2556 10115
rect 2504 10072 2556 10081
rect 3516 10140 3568 10192
rect 6552 10183 6604 10192
rect 6552 10149 6561 10183
rect 6561 10149 6595 10183
rect 6595 10149 6604 10183
rect 6552 10140 6604 10149
rect 8116 10140 8168 10192
rect 1492 10047 1544 10056
rect 1492 10013 1501 10047
rect 1501 10013 1535 10047
rect 1535 10013 1544 10047
rect 1492 10004 1544 10013
rect 1952 10047 2004 10056
rect 1952 10013 1961 10047
rect 1961 10013 1995 10047
rect 1995 10013 2004 10047
rect 1952 10004 2004 10013
rect 3056 10004 3108 10056
rect 3240 10047 3292 10056
rect 3240 10013 3249 10047
rect 3249 10013 3283 10047
rect 3283 10013 3292 10047
rect 3240 10004 3292 10013
rect 6000 10004 6052 10056
rect 8116 10004 8168 10056
rect 9680 10004 9732 10056
rect 4804 9979 4856 9988
rect 4804 9945 4838 9979
rect 4838 9945 4856 9979
rect 4804 9936 4856 9945
rect 7196 9936 7248 9988
rect 7380 9936 7432 9988
rect 1676 9868 1728 9920
rect 2044 9911 2096 9920
rect 2044 9877 2053 9911
rect 2053 9877 2087 9911
rect 2087 9877 2096 9911
rect 2044 9868 2096 9877
rect 2688 9868 2740 9920
rect 3884 9868 3936 9920
rect 5908 9911 5960 9920
rect 5908 9877 5917 9911
rect 5917 9877 5951 9911
rect 5951 9877 5960 9911
rect 5908 9868 5960 9877
rect 7472 9868 7524 9920
rect 8300 9868 8352 9920
rect 10232 9936 10284 9988
rect 10600 10208 10652 10260
rect 14740 10208 14792 10260
rect 16396 10208 16448 10260
rect 17132 10208 17184 10260
rect 17224 10208 17276 10260
rect 17408 10251 17460 10260
rect 17408 10217 17417 10251
rect 17417 10217 17451 10251
rect 17451 10217 17460 10251
rect 17408 10208 17460 10217
rect 18420 10208 18472 10260
rect 16212 10072 16264 10124
rect 17040 10115 17092 10124
rect 17040 10081 17049 10115
rect 17049 10081 17083 10115
rect 17083 10081 17092 10115
rect 17040 10072 17092 10081
rect 17316 10072 17368 10124
rect 17408 10072 17460 10124
rect 11520 10004 11572 10056
rect 11980 10004 12032 10056
rect 12900 10004 12952 10056
rect 16948 10047 17000 10056
rect 16948 10013 16957 10047
rect 16957 10013 16991 10047
rect 16991 10013 17000 10047
rect 16948 10004 17000 10013
rect 13084 9936 13136 9988
rect 17132 9936 17184 9988
rect 18420 9979 18472 9988
rect 18420 9945 18429 9979
rect 18429 9945 18463 9979
rect 18463 9945 18472 9979
rect 18420 9936 18472 9945
rect 16028 9868 16080 9920
rect 17500 9868 17552 9920
rect 17960 9868 18012 9920
rect 5398 9766 5450 9818
rect 5462 9766 5514 9818
rect 5526 9766 5578 9818
rect 5590 9766 5642 9818
rect 5654 9766 5706 9818
rect 9846 9766 9898 9818
rect 9910 9766 9962 9818
rect 9974 9766 10026 9818
rect 10038 9766 10090 9818
rect 10102 9766 10154 9818
rect 14294 9766 14346 9818
rect 14358 9766 14410 9818
rect 14422 9766 14474 9818
rect 14486 9766 14538 9818
rect 14550 9766 14602 9818
rect 1952 9664 2004 9716
rect 3700 9664 3752 9716
rect 1492 9571 1544 9580
rect 1492 9537 1501 9571
rect 1501 9537 1535 9571
rect 1535 9537 1544 9571
rect 1492 9528 1544 9537
rect 2688 9596 2740 9648
rect 6552 9596 6604 9648
rect 2504 9528 2556 9580
rect 2320 9460 2372 9512
rect 6736 9528 6788 9580
rect 2964 9460 3016 9512
rect 6000 9460 6052 9512
rect 1768 9367 1820 9376
rect 1768 9333 1777 9367
rect 1777 9333 1811 9367
rect 1811 9333 1820 9367
rect 1768 9324 1820 9333
rect 2228 9367 2280 9376
rect 2228 9333 2237 9367
rect 2237 9333 2271 9367
rect 2271 9333 2280 9367
rect 2228 9324 2280 9333
rect 2780 9324 2832 9376
rect 4528 9392 4580 9444
rect 4620 9324 4672 9376
rect 5080 9324 5132 9376
rect 7288 9571 7340 9580
rect 7288 9537 7297 9571
rect 7297 9537 7331 9571
rect 7331 9537 7340 9571
rect 7288 9528 7340 9537
rect 8024 9528 8076 9580
rect 8484 9528 8536 9580
rect 16948 9664 17000 9716
rect 15016 9596 15068 9648
rect 17132 9639 17184 9648
rect 17132 9605 17141 9639
rect 17141 9605 17175 9639
rect 17175 9605 17184 9639
rect 17132 9596 17184 9605
rect 7380 9460 7432 9512
rect 8116 9460 8168 9512
rect 8944 9324 8996 9376
rect 11888 9367 11940 9376
rect 11888 9333 11897 9367
rect 11897 9333 11931 9367
rect 11931 9333 11940 9367
rect 11888 9324 11940 9333
rect 13268 9503 13320 9512
rect 13268 9469 13277 9503
rect 13277 9469 13311 9503
rect 13311 9469 13320 9503
rect 13268 9460 13320 9469
rect 17408 9460 17460 9512
rect 18052 9528 18104 9580
rect 18420 9571 18472 9580
rect 18420 9537 18429 9571
rect 18429 9537 18463 9571
rect 18463 9537 18472 9571
rect 18420 9528 18472 9537
rect 14096 9392 14148 9444
rect 18236 9460 18288 9512
rect 15384 9324 15436 9376
rect 17868 9324 17920 9376
rect 18236 9324 18288 9376
rect 3174 9222 3226 9274
rect 3238 9222 3290 9274
rect 3302 9222 3354 9274
rect 3366 9222 3418 9274
rect 3430 9222 3482 9274
rect 7622 9222 7674 9274
rect 7686 9222 7738 9274
rect 7750 9222 7802 9274
rect 7814 9222 7866 9274
rect 7878 9222 7930 9274
rect 12070 9222 12122 9274
rect 12134 9222 12186 9274
rect 12198 9222 12250 9274
rect 12262 9222 12314 9274
rect 12326 9222 12378 9274
rect 16518 9222 16570 9274
rect 16582 9222 16634 9274
rect 16646 9222 16698 9274
rect 16710 9222 16762 9274
rect 16774 9222 16826 9274
rect 2504 9163 2556 9172
rect 2504 9129 2513 9163
rect 2513 9129 2547 9163
rect 2547 9129 2556 9163
rect 2504 9120 2556 9129
rect 3424 9163 3476 9172
rect 3424 9129 3433 9163
rect 3433 9129 3467 9163
rect 3467 9129 3476 9163
rect 3424 9120 3476 9129
rect 6092 9120 6144 9172
rect 7196 9120 7248 9172
rect 8760 9163 8812 9172
rect 8760 9129 8769 9163
rect 8769 9129 8803 9163
rect 8803 9129 8812 9163
rect 8760 9120 8812 9129
rect 10232 9120 10284 9172
rect 12624 9120 12676 9172
rect 14740 9120 14792 9172
rect 15384 9120 15436 9172
rect 17316 9163 17368 9172
rect 17316 9129 17325 9163
rect 17325 9129 17359 9163
rect 17359 9129 17368 9163
rect 17316 9120 17368 9129
rect 1860 8916 1912 8968
rect 2412 8984 2464 9036
rect 3240 8984 3292 9036
rect 16028 9027 16080 9036
rect 16028 8993 16037 9027
rect 16037 8993 16071 9027
rect 16071 8993 16080 9027
rect 16028 8984 16080 8993
rect 1952 8848 2004 8900
rect 2964 8916 3016 8968
rect 3056 8916 3108 8968
rect 1492 8823 1544 8832
rect 1492 8789 1501 8823
rect 1501 8789 1535 8823
rect 1535 8789 1544 8823
rect 1492 8780 1544 8789
rect 1584 8780 1636 8832
rect 2412 8780 2464 8832
rect 3424 8780 3476 8832
rect 6000 8916 6052 8968
rect 7380 8959 7432 8968
rect 7380 8925 7389 8959
rect 7389 8925 7423 8959
rect 7423 8925 7432 8959
rect 7380 8916 7432 8925
rect 8944 8916 8996 8968
rect 11520 8959 11572 8968
rect 11520 8925 11529 8959
rect 11529 8925 11563 8959
rect 11563 8925 11572 8959
rect 11520 8916 11572 8925
rect 11980 8916 12032 8968
rect 13268 8916 13320 8968
rect 13912 8916 13964 8968
rect 14740 8959 14792 8968
rect 14740 8925 14749 8959
rect 14749 8925 14783 8959
rect 14783 8925 14792 8959
rect 14740 8916 14792 8925
rect 16304 8916 16356 8968
rect 18144 9052 18196 9104
rect 17316 8916 17368 8968
rect 18052 8916 18104 8968
rect 4436 8848 4488 8900
rect 4528 8848 4580 8900
rect 5724 8891 5776 8900
rect 5724 8857 5758 8891
rect 5758 8857 5776 8891
rect 5724 8848 5776 8857
rect 7196 8848 7248 8900
rect 7748 8848 7800 8900
rect 4068 8780 4120 8832
rect 4252 8780 4304 8832
rect 12808 8848 12860 8900
rect 12992 8848 13044 8900
rect 13452 8848 13504 8900
rect 17132 8848 17184 8900
rect 18328 8916 18380 8968
rect 18512 8959 18564 8968
rect 18512 8925 18521 8959
rect 18521 8925 18555 8959
rect 18555 8925 18564 8959
rect 18512 8916 18564 8925
rect 14648 8823 14700 8832
rect 14648 8789 14657 8823
rect 14657 8789 14691 8823
rect 14691 8789 14700 8823
rect 14648 8780 14700 8789
rect 15108 8823 15160 8832
rect 15108 8789 15117 8823
rect 15117 8789 15151 8823
rect 15151 8789 15160 8823
rect 15108 8780 15160 8789
rect 15476 8823 15528 8832
rect 15476 8789 15485 8823
rect 15485 8789 15519 8823
rect 15519 8789 15528 8823
rect 15476 8780 15528 8789
rect 16580 8780 16632 8832
rect 16856 8780 16908 8832
rect 5398 8678 5450 8730
rect 5462 8678 5514 8730
rect 5526 8678 5578 8730
rect 5590 8678 5642 8730
rect 5654 8678 5706 8730
rect 9846 8678 9898 8730
rect 9910 8678 9962 8730
rect 9974 8678 10026 8730
rect 10038 8678 10090 8730
rect 10102 8678 10154 8730
rect 14294 8678 14346 8730
rect 14358 8678 14410 8730
rect 14422 8678 14474 8730
rect 14486 8678 14538 8730
rect 14550 8678 14602 8730
rect 2320 8619 2372 8628
rect 2320 8585 2329 8619
rect 2329 8585 2363 8619
rect 2363 8585 2372 8619
rect 2320 8576 2372 8585
rect 2228 8508 2280 8560
rect 1952 8415 2004 8424
rect 1952 8381 1961 8415
rect 1961 8381 1995 8415
rect 1995 8381 2004 8415
rect 1952 8372 2004 8381
rect 8944 8576 8996 8628
rect 9220 8576 9272 8628
rect 2964 8508 3016 8560
rect 3516 8483 3568 8492
rect 3516 8449 3525 8483
rect 3525 8449 3559 8483
rect 3559 8449 3568 8483
rect 3516 8440 3568 8449
rect 5080 8508 5132 8560
rect 5724 8508 5776 8560
rect 6000 8508 6052 8560
rect 11244 8508 11296 8560
rect 15016 8576 15068 8628
rect 16580 8576 16632 8628
rect 17408 8576 17460 8628
rect 16028 8508 16080 8560
rect 1400 8304 1452 8356
rect 2688 8304 2740 8356
rect 2504 8236 2556 8288
rect 3056 8372 3108 8424
rect 5264 8440 5316 8492
rect 7748 8483 7800 8492
rect 7748 8449 7757 8483
rect 7757 8449 7791 8483
rect 7791 8449 7800 8483
rect 7748 8440 7800 8449
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 15936 8440 15988 8492
rect 17040 8440 17092 8492
rect 17868 8483 17920 8492
rect 17868 8449 17877 8483
rect 17877 8449 17911 8483
rect 17911 8449 17920 8483
rect 18236 8483 18288 8492
rect 17868 8440 17920 8449
rect 18236 8449 18245 8483
rect 18245 8449 18279 8483
rect 18279 8449 18288 8483
rect 18236 8440 18288 8449
rect 3240 8304 3292 8356
rect 4436 8372 4488 8424
rect 10324 8372 10376 8424
rect 11520 8415 11572 8424
rect 11520 8381 11529 8415
rect 11529 8381 11563 8415
rect 11563 8381 11572 8415
rect 11520 8372 11572 8381
rect 16028 8415 16080 8424
rect 16028 8381 16037 8415
rect 16037 8381 16071 8415
rect 16071 8381 16080 8415
rect 16028 8372 16080 8381
rect 5816 8304 5868 8356
rect 10784 8304 10836 8356
rect 18052 8347 18104 8356
rect 18052 8313 18061 8347
rect 18061 8313 18095 8347
rect 18095 8313 18104 8347
rect 18052 8304 18104 8313
rect 18420 8347 18472 8356
rect 18420 8313 18429 8347
rect 18429 8313 18463 8347
rect 18463 8313 18472 8347
rect 18420 8304 18472 8313
rect 3700 8236 3752 8288
rect 4252 8236 4304 8288
rect 4620 8236 4672 8288
rect 8484 8236 8536 8288
rect 10508 8279 10560 8288
rect 10508 8245 10517 8279
rect 10517 8245 10551 8279
rect 10551 8245 10560 8279
rect 10508 8236 10560 8245
rect 15384 8279 15436 8288
rect 15384 8245 15393 8279
rect 15393 8245 15427 8279
rect 15427 8245 15436 8279
rect 15384 8236 15436 8245
rect 3174 8134 3226 8186
rect 3238 8134 3290 8186
rect 3302 8134 3354 8186
rect 3366 8134 3418 8186
rect 3430 8134 3482 8186
rect 7622 8134 7674 8186
rect 7686 8134 7738 8186
rect 7750 8134 7802 8186
rect 7814 8134 7866 8186
rect 7878 8134 7930 8186
rect 12070 8134 12122 8186
rect 12134 8134 12186 8186
rect 12198 8134 12250 8186
rect 12262 8134 12314 8186
rect 12326 8134 12378 8186
rect 16518 8134 16570 8186
rect 16582 8134 16634 8186
rect 16646 8134 16698 8186
rect 16710 8134 16762 8186
rect 16774 8134 16826 8186
rect 1492 8075 1544 8084
rect 1492 8041 1501 8075
rect 1501 8041 1535 8075
rect 1535 8041 1544 8075
rect 1492 8032 1544 8041
rect 1952 8032 2004 8084
rect 2688 8032 2740 8084
rect 4344 8032 4396 8084
rect 11612 8032 11664 8084
rect 12348 8032 12400 8084
rect 16948 8075 17000 8084
rect 16948 8041 16957 8075
rect 16957 8041 16991 8075
rect 16991 8041 17000 8075
rect 16948 8032 17000 8041
rect 17316 8032 17368 8084
rect 17684 8032 17736 8084
rect 2780 7939 2832 7948
rect 2780 7905 2789 7939
rect 2789 7905 2823 7939
rect 2823 7905 2832 7939
rect 2780 7896 2832 7905
rect 1676 7871 1728 7880
rect 1676 7837 1685 7871
rect 1685 7837 1719 7871
rect 1719 7837 1728 7871
rect 1676 7828 1728 7837
rect 2320 7828 2372 7880
rect 3700 7964 3752 8016
rect 18328 7964 18380 8016
rect 1952 7760 2004 7812
rect 3792 7896 3844 7948
rect 4436 7828 4488 7880
rect 3792 7760 3844 7812
rect 4068 7760 4120 7812
rect 1860 7735 1912 7744
rect 1860 7701 1869 7735
rect 1869 7701 1903 7735
rect 1903 7701 1912 7735
rect 1860 7692 1912 7701
rect 2136 7692 2188 7744
rect 6000 7692 6052 7744
rect 6276 7828 6328 7880
rect 8300 7896 8352 7948
rect 11520 7896 11572 7948
rect 15016 7939 15068 7948
rect 15016 7905 15025 7939
rect 15025 7905 15059 7939
rect 15059 7905 15068 7939
rect 15016 7896 15068 7905
rect 15384 7896 15436 7948
rect 6920 7692 6972 7744
rect 8484 7692 8536 7744
rect 10600 7828 10652 7880
rect 10784 7871 10836 7880
rect 10784 7837 10818 7871
rect 10818 7837 10836 7871
rect 10784 7828 10836 7837
rect 9220 7803 9272 7812
rect 9220 7769 9254 7803
rect 9254 7769 9272 7803
rect 9220 7760 9272 7769
rect 10324 7735 10376 7744
rect 10324 7701 10333 7735
rect 10333 7701 10367 7735
rect 10367 7701 10376 7735
rect 10324 7692 10376 7701
rect 13268 7760 13320 7812
rect 15476 7828 15528 7880
rect 16948 7828 17000 7880
rect 17592 7828 17644 7880
rect 17776 7828 17828 7880
rect 16028 7760 16080 7812
rect 12072 7692 12124 7744
rect 13452 7735 13504 7744
rect 13452 7701 13461 7735
rect 13461 7701 13495 7735
rect 13495 7701 13504 7735
rect 13452 7692 13504 7701
rect 15384 7692 15436 7744
rect 17316 7692 17368 7744
rect 18420 7735 18472 7744
rect 18420 7701 18429 7735
rect 18429 7701 18463 7735
rect 18463 7701 18472 7735
rect 18420 7692 18472 7701
rect 5398 7590 5450 7642
rect 5462 7590 5514 7642
rect 5526 7590 5578 7642
rect 5590 7590 5642 7642
rect 5654 7590 5706 7642
rect 9846 7590 9898 7642
rect 9910 7590 9962 7642
rect 9974 7590 10026 7642
rect 10038 7590 10090 7642
rect 10102 7590 10154 7642
rect 14294 7590 14346 7642
rect 14358 7590 14410 7642
rect 14422 7590 14474 7642
rect 14486 7590 14538 7642
rect 14550 7590 14602 7642
rect 1952 7488 2004 7540
rect 2136 7531 2188 7540
rect 2136 7497 2145 7531
rect 2145 7497 2179 7531
rect 2179 7497 2188 7531
rect 2136 7488 2188 7497
rect 2412 7488 2464 7540
rect 3056 7488 3108 7540
rect 4988 7488 5040 7540
rect 4436 7420 4488 7472
rect 2504 7352 2556 7404
rect 2780 7352 2832 7404
rect 5172 7352 5224 7404
rect 5816 7352 5868 7404
rect 8024 7420 8076 7472
rect 9220 7488 9272 7540
rect 15384 7531 15436 7540
rect 15384 7497 15393 7531
rect 15393 7497 15427 7531
rect 15427 7497 15436 7531
rect 15384 7488 15436 7497
rect 16396 7531 16448 7540
rect 16396 7497 16405 7531
rect 16405 7497 16439 7531
rect 16439 7497 16448 7531
rect 16396 7488 16448 7497
rect 10508 7420 10560 7472
rect 12072 7420 12124 7472
rect 13084 7420 13136 7472
rect 17684 7420 17736 7472
rect 6184 7352 6236 7404
rect 8300 7352 8352 7404
rect 1676 7327 1728 7336
rect 1676 7293 1685 7327
rect 1685 7293 1719 7327
rect 1719 7293 1728 7327
rect 1676 7284 1728 7293
rect 4436 7327 4488 7336
rect 4436 7293 4445 7327
rect 4445 7293 4479 7327
rect 4479 7293 4488 7327
rect 4436 7284 4488 7293
rect 8484 7327 8536 7336
rect 8484 7293 8493 7327
rect 8493 7293 8527 7327
rect 8527 7293 8536 7327
rect 8484 7284 8536 7293
rect 10600 7395 10652 7404
rect 10600 7361 10609 7395
rect 10609 7361 10643 7395
rect 10643 7361 10652 7395
rect 10600 7352 10652 7361
rect 11888 7352 11940 7404
rect 13636 7352 13688 7404
rect 14924 7352 14976 7404
rect 15292 7395 15344 7404
rect 15292 7361 15301 7395
rect 15301 7361 15335 7395
rect 15335 7361 15344 7395
rect 15292 7352 15344 7361
rect 11520 7284 11572 7336
rect 11980 7284 12032 7336
rect 2688 7216 2740 7268
rect 9220 7259 9272 7268
rect 9220 7225 9229 7259
rect 9229 7225 9263 7259
rect 9263 7225 9272 7259
rect 9220 7216 9272 7225
rect 4528 7191 4580 7200
rect 4528 7157 4537 7191
rect 4537 7157 4571 7191
rect 4571 7157 4580 7191
rect 4528 7148 4580 7157
rect 6920 7148 6972 7200
rect 9588 7148 9640 7200
rect 11612 7148 11664 7200
rect 15200 7284 15252 7336
rect 17316 7352 17368 7404
rect 17592 7395 17644 7404
rect 17592 7361 17601 7395
rect 17601 7361 17635 7395
rect 17635 7361 17644 7395
rect 17592 7352 17644 7361
rect 13636 7216 13688 7268
rect 15752 7284 15804 7336
rect 17224 7327 17276 7336
rect 17224 7293 17233 7327
rect 17233 7293 17267 7327
rect 17267 7293 17276 7327
rect 17224 7284 17276 7293
rect 16212 7216 16264 7268
rect 18236 7148 18288 7200
rect 18420 7191 18472 7200
rect 18420 7157 18429 7191
rect 18429 7157 18463 7191
rect 18463 7157 18472 7191
rect 18420 7148 18472 7157
rect 3174 7046 3226 7098
rect 3238 7046 3290 7098
rect 3302 7046 3354 7098
rect 3366 7046 3418 7098
rect 3430 7046 3482 7098
rect 7622 7046 7674 7098
rect 7686 7046 7738 7098
rect 7750 7046 7802 7098
rect 7814 7046 7866 7098
rect 7878 7046 7930 7098
rect 12070 7046 12122 7098
rect 12134 7046 12186 7098
rect 12198 7046 12250 7098
rect 12262 7046 12314 7098
rect 12326 7046 12378 7098
rect 16518 7046 16570 7098
rect 16582 7046 16634 7098
rect 16646 7046 16698 7098
rect 16710 7046 16762 7098
rect 16774 7046 16826 7098
rect 1492 6987 1544 6996
rect 1492 6953 1501 6987
rect 1501 6953 1535 6987
rect 1535 6953 1544 6987
rect 1492 6944 1544 6953
rect 1676 6944 1728 6996
rect 3516 6987 3568 6996
rect 2412 6876 2464 6928
rect 2872 6876 2924 6928
rect 3516 6953 3525 6987
rect 3525 6953 3559 6987
rect 3559 6953 3568 6987
rect 3516 6944 3568 6953
rect 5080 6944 5132 6996
rect 11980 6944 12032 6996
rect 15292 6944 15344 6996
rect 17684 6987 17736 6996
rect 17684 6953 17693 6987
rect 17693 6953 17727 6987
rect 17727 6953 17736 6987
rect 17684 6944 17736 6953
rect 17776 6944 17828 6996
rect 2688 6808 2740 6860
rect 4436 6851 4488 6860
rect 3700 6740 3752 6792
rect 2228 6672 2280 6724
rect 4436 6817 4445 6851
rect 4445 6817 4479 6851
rect 4479 6817 4488 6851
rect 4436 6808 4488 6817
rect 6092 6808 6144 6860
rect 8392 6740 8444 6792
rect 15016 6876 15068 6928
rect 15108 6808 15160 6860
rect 16212 6851 16264 6860
rect 16212 6817 16221 6851
rect 16221 6817 16255 6851
rect 16255 6817 16264 6851
rect 16212 6808 16264 6817
rect 6092 6672 6144 6724
rect 9588 6715 9640 6724
rect 2320 6647 2372 6656
rect 2320 6613 2329 6647
rect 2329 6613 2363 6647
rect 2363 6613 2372 6647
rect 2320 6604 2372 6613
rect 3056 6647 3108 6656
rect 3056 6613 3065 6647
rect 3065 6613 3099 6647
rect 3099 6613 3108 6647
rect 3056 6604 3108 6613
rect 3148 6647 3200 6656
rect 3148 6613 3157 6647
rect 3157 6613 3191 6647
rect 3191 6613 3200 6647
rect 3976 6647 4028 6656
rect 3148 6604 3200 6613
rect 3976 6613 3985 6647
rect 3985 6613 4019 6647
rect 4019 6613 4028 6647
rect 3976 6604 4028 6613
rect 7288 6604 7340 6656
rect 9588 6681 9622 6715
rect 9622 6681 9640 6715
rect 9588 6672 9640 6681
rect 10232 6672 10284 6724
rect 11336 6672 11388 6724
rect 15384 6740 15436 6792
rect 16580 6808 16632 6860
rect 17224 6808 17276 6860
rect 17316 6740 17368 6792
rect 17868 6783 17920 6792
rect 17868 6749 17877 6783
rect 17877 6749 17911 6783
rect 17911 6749 17920 6783
rect 17868 6740 17920 6749
rect 18236 6783 18288 6792
rect 18236 6749 18245 6783
rect 18245 6749 18279 6783
rect 18279 6749 18288 6783
rect 18236 6740 18288 6749
rect 12900 6672 12952 6724
rect 12992 6672 13044 6724
rect 10876 6604 10928 6656
rect 10968 6647 11020 6656
rect 10968 6613 10977 6647
rect 10977 6613 11011 6647
rect 11011 6613 11020 6647
rect 10968 6604 11020 6613
rect 11520 6604 11572 6656
rect 14096 6604 14148 6656
rect 15752 6647 15804 6656
rect 15752 6613 15761 6647
rect 15761 6613 15795 6647
rect 15795 6613 15804 6647
rect 15752 6604 15804 6613
rect 18052 6647 18104 6656
rect 18052 6613 18061 6647
rect 18061 6613 18095 6647
rect 18095 6613 18104 6647
rect 18052 6604 18104 6613
rect 18420 6647 18472 6656
rect 18420 6613 18429 6647
rect 18429 6613 18463 6647
rect 18463 6613 18472 6647
rect 18420 6604 18472 6613
rect 5398 6502 5450 6554
rect 5462 6502 5514 6554
rect 5526 6502 5578 6554
rect 5590 6502 5642 6554
rect 5654 6502 5706 6554
rect 9846 6502 9898 6554
rect 9910 6502 9962 6554
rect 9974 6502 10026 6554
rect 10038 6502 10090 6554
rect 10102 6502 10154 6554
rect 14294 6502 14346 6554
rect 14358 6502 14410 6554
rect 14422 6502 14474 6554
rect 14486 6502 14538 6554
rect 14550 6502 14602 6554
rect 3056 6400 3108 6452
rect 3884 6400 3936 6452
rect 7012 6400 7064 6452
rect 8116 6400 8168 6452
rect 11336 6443 11388 6452
rect 11336 6409 11345 6443
rect 11345 6409 11379 6443
rect 11379 6409 11388 6443
rect 11336 6400 11388 6409
rect 13268 6443 13320 6452
rect 13268 6409 13277 6443
rect 13277 6409 13311 6443
rect 13311 6409 13320 6443
rect 13268 6400 13320 6409
rect 16948 6400 17000 6452
rect 17224 6400 17276 6452
rect 17316 6400 17368 6452
rect 3516 6332 3568 6384
rect 2504 6264 2556 6316
rect 3424 6307 3476 6316
rect 3424 6273 3433 6307
rect 3433 6273 3467 6307
rect 3467 6273 3476 6307
rect 3424 6264 3476 6273
rect 5816 6332 5868 6384
rect 5908 6375 5960 6384
rect 5908 6341 5926 6375
rect 5926 6341 5960 6375
rect 5908 6332 5960 6341
rect 11612 6332 11664 6384
rect 12348 6332 12400 6384
rect 3884 6307 3936 6316
rect 3884 6273 3893 6307
rect 3893 6273 3927 6307
rect 3927 6273 3936 6307
rect 3884 6264 3936 6273
rect 5632 6264 5684 6316
rect 6184 6307 6236 6316
rect 6184 6273 6193 6307
rect 6193 6273 6227 6307
rect 6227 6273 6236 6307
rect 6184 6264 6236 6273
rect 10232 6307 10284 6316
rect 10232 6273 10241 6307
rect 10241 6273 10275 6307
rect 10275 6273 10284 6307
rect 10232 6264 10284 6273
rect 15752 6332 15804 6384
rect 16212 6332 16264 6384
rect 1584 6239 1636 6248
rect 1584 6205 1593 6239
rect 1593 6205 1627 6239
rect 1627 6205 1636 6239
rect 1584 6196 1636 6205
rect 2688 6239 2740 6248
rect 2688 6205 2697 6239
rect 2697 6205 2731 6239
rect 2731 6205 2740 6239
rect 2688 6196 2740 6205
rect 2964 6196 3016 6248
rect 3332 6196 3384 6248
rect 3700 6239 3752 6248
rect 3700 6205 3709 6239
rect 3709 6205 3743 6239
rect 3743 6205 3752 6239
rect 3700 6196 3752 6205
rect 4528 6128 4580 6180
rect 10508 6196 10560 6248
rect 11520 6196 11572 6248
rect 13452 6196 13504 6248
rect 15108 6264 15160 6316
rect 16856 6264 16908 6316
rect 17592 6264 17644 6316
rect 18144 6264 18196 6316
rect 15384 6196 15436 6248
rect 15476 6196 15528 6248
rect 15752 6239 15804 6248
rect 15752 6205 15761 6239
rect 15761 6205 15795 6239
rect 15795 6205 15804 6239
rect 15752 6196 15804 6205
rect 16580 6196 16632 6248
rect 16764 6196 16816 6248
rect 16948 6239 17000 6248
rect 16948 6205 16957 6239
rect 16957 6205 16991 6239
rect 16991 6205 17000 6239
rect 16948 6196 17000 6205
rect 10876 6128 10928 6180
rect 11336 6128 11388 6180
rect 1768 6060 1820 6112
rect 3056 6103 3108 6112
rect 3056 6069 3065 6103
rect 3065 6069 3099 6103
rect 3099 6069 3108 6103
rect 3056 6060 3108 6069
rect 3424 6060 3476 6112
rect 3976 6060 4028 6112
rect 4804 6103 4856 6112
rect 4804 6069 4813 6103
rect 4813 6069 4847 6103
rect 4847 6069 4856 6103
rect 4804 6060 4856 6069
rect 8024 6060 8076 6112
rect 8852 6103 8904 6112
rect 8852 6069 8861 6103
rect 8861 6069 8895 6103
rect 8895 6069 8904 6103
rect 8852 6060 8904 6069
rect 9128 6060 9180 6112
rect 15936 6128 15988 6180
rect 13084 6060 13136 6112
rect 13820 6060 13872 6112
rect 16396 6060 16448 6112
rect 18788 6128 18840 6180
rect 16948 6060 17000 6112
rect 17960 6103 18012 6112
rect 17960 6069 17969 6103
rect 17969 6069 18003 6103
rect 18003 6069 18012 6103
rect 17960 6060 18012 6069
rect 18420 6103 18472 6112
rect 18420 6069 18429 6103
rect 18429 6069 18463 6103
rect 18463 6069 18472 6103
rect 18420 6060 18472 6069
rect 3174 5958 3226 6010
rect 3238 5958 3290 6010
rect 3302 5958 3354 6010
rect 3366 5958 3418 6010
rect 3430 5958 3482 6010
rect 7622 5958 7674 6010
rect 7686 5958 7738 6010
rect 7750 5958 7802 6010
rect 7814 5958 7866 6010
rect 7878 5958 7930 6010
rect 12070 5958 12122 6010
rect 12134 5958 12186 6010
rect 12198 5958 12250 6010
rect 12262 5958 12314 6010
rect 12326 5958 12378 6010
rect 16518 5958 16570 6010
rect 16582 5958 16634 6010
rect 16646 5958 16698 6010
rect 16710 5958 16762 6010
rect 16774 5958 16826 6010
rect 2688 5856 2740 5908
rect 6092 5856 6144 5908
rect 6184 5899 6236 5908
rect 6184 5865 6193 5899
rect 6193 5865 6227 5899
rect 6227 5865 6236 5899
rect 6184 5856 6236 5865
rect 6920 5856 6972 5908
rect 4068 5788 4120 5840
rect 5816 5788 5868 5840
rect 8300 5831 8352 5840
rect 8300 5797 8309 5831
rect 8309 5797 8343 5831
rect 8343 5797 8352 5831
rect 8300 5788 8352 5797
rect 10324 5856 10376 5908
rect 10508 5899 10560 5908
rect 10508 5865 10517 5899
rect 10517 5865 10551 5899
rect 10551 5865 10560 5899
rect 10508 5856 10560 5865
rect 10876 5899 10928 5908
rect 10876 5865 10885 5899
rect 10885 5865 10919 5899
rect 10919 5865 10928 5899
rect 10876 5856 10928 5865
rect 12992 5856 13044 5908
rect 13176 5856 13228 5908
rect 14188 5899 14240 5908
rect 14188 5865 14197 5899
rect 14197 5865 14231 5899
rect 14231 5865 14240 5899
rect 14188 5856 14240 5865
rect 15108 5899 15160 5908
rect 15108 5865 15117 5899
rect 15117 5865 15151 5899
rect 15151 5865 15160 5899
rect 15108 5856 15160 5865
rect 15476 5899 15528 5908
rect 15476 5865 15485 5899
rect 15485 5865 15519 5899
rect 15519 5865 15528 5899
rect 15476 5856 15528 5865
rect 16396 5856 16448 5908
rect 17868 5899 17920 5908
rect 1676 5763 1728 5772
rect 1676 5729 1685 5763
rect 1685 5729 1719 5763
rect 1719 5729 1728 5763
rect 1676 5720 1728 5729
rect 1768 5763 1820 5772
rect 1768 5729 1777 5763
rect 1777 5729 1811 5763
rect 1811 5729 1820 5763
rect 1768 5720 1820 5729
rect 2872 5720 2924 5772
rect 2044 5652 2096 5704
rect 2596 5695 2648 5704
rect 2596 5661 2605 5695
rect 2605 5661 2639 5695
rect 2639 5661 2648 5695
rect 2596 5652 2648 5661
rect 3700 5720 3752 5772
rect 4436 5720 4488 5772
rect 5908 5720 5960 5772
rect 9772 5720 9824 5772
rect 11336 5763 11388 5772
rect 4252 5652 4304 5704
rect 4804 5695 4856 5704
rect 4804 5661 4838 5695
rect 4838 5661 4856 5695
rect 4804 5652 4856 5661
rect 6552 5695 6604 5704
rect 2872 5584 2924 5636
rect 6552 5661 6561 5695
rect 6561 5661 6595 5695
rect 6595 5661 6604 5695
rect 6552 5652 6604 5661
rect 8208 5652 8260 5704
rect 8300 5652 8352 5704
rect 6276 5584 6328 5636
rect 9128 5584 9180 5636
rect 11336 5729 11345 5763
rect 11345 5729 11379 5763
rect 11379 5729 11388 5763
rect 11336 5720 11388 5729
rect 11704 5720 11756 5772
rect 12440 5720 12492 5772
rect 15752 5720 15804 5772
rect 15936 5763 15988 5772
rect 15936 5729 15945 5763
rect 15945 5729 15979 5763
rect 15979 5729 15988 5763
rect 15936 5720 15988 5729
rect 16028 5763 16080 5772
rect 16028 5729 16037 5763
rect 16037 5729 16071 5763
rect 16071 5729 16080 5763
rect 16304 5763 16356 5772
rect 16028 5720 16080 5729
rect 16304 5729 16313 5763
rect 16313 5729 16347 5763
rect 16347 5729 16356 5763
rect 16304 5720 16356 5729
rect 16672 5788 16724 5840
rect 17040 5788 17092 5840
rect 17868 5865 17877 5899
rect 17877 5865 17911 5899
rect 17911 5865 17920 5899
rect 17868 5856 17920 5865
rect 17316 5720 17368 5772
rect 2412 5559 2464 5568
rect 2412 5525 2421 5559
rect 2421 5525 2455 5559
rect 2455 5525 2464 5559
rect 2412 5516 2464 5525
rect 2596 5516 2648 5568
rect 3976 5559 4028 5568
rect 3976 5525 3985 5559
rect 3985 5525 4019 5559
rect 4019 5525 4028 5559
rect 3976 5516 4028 5525
rect 7104 5559 7156 5568
rect 7104 5525 7113 5559
rect 7113 5525 7147 5559
rect 7147 5525 7156 5559
rect 7104 5516 7156 5525
rect 9680 5559 9732 5568
rect 9680 5525 9689 5559
rect 9689 5525 9723 5559
rect 9723 5525 9732 5559
rect 11152 5652 11204 5704
rect 13912 5695 13964 5704
rect 13912 5661 13921 5695
rect 13921 5661 13955 5695
rect 13955 5661 13964 5695
rect 13912 5652 13964 5661
rect 14188 5652 14240 5704
rect 16212 5652 16264 5704
rect 17040 5652 17092 5704
rect 11336 5584 11388 5636
rect 9680 5516 9732 5525
rect 11060 5516 11112 5568
rect 12164 5584 12216 5636
rect 14556 5584 14608 5636
rect 15292 5584 15344 5636
rect 16948 5584 17000 5636
rect 15200 5559 15252 5568
rect 15200 5525 15209 5559
rect 15209 5525 15243 5559
rect 15243 5525 15252 5559
rect 15200 5516 15252 5525
rect 18420 5559 18472 5568
rect 18420 5525 18429 5559
rect 18429 5525 18463 5559
rect 18463 5525 18472 5559
rect 18420 5516 18472 5525
rect 5398 5414 5450 5466
rect 5462 5414 5514 5466
rect 5526 5414 5578 5466
rect 5590 5414 5642 5466
rect 5654 5414 5706 5466
rect 9846 5414 9898 5466
rect 9910 5414 9962 5466
rect 9974 5414 10026 5466
rect 10038 5414 10090 5466
rect 10102 5414 10154 5466
rect 14294 5414 14346 5466
rect 14358 5414 14410 5466
rect 14422 5414 14474 5466
rect 14486 5414 14538 5466
rect 14550 5414 14602 5466
rect 1492 5355 1544 5364
rect 1492 5321 1501 5355
rect 1501 5321 1535 5355
rect 1535 5321 1544 5355
rect 1492 5312 1544 5321
rect 1952 5355 2004 5364
rect 1952 5321 1961 5355
rect 1961 5321 1995 5355
rect 1995 5321 2004 5355
rect 1952 5312 2004 5321
rect 2228 5312 2280 5364
rect 2504 5312 2556 5364
rect 3056 5355 3108 5364
rect 3056 5321 3065 5355
rect 3065 5321 3099 5355
rect 3099 5321 3108 5355
rect 3056 5312 3108 5321
rect 3516 5312 3568 5364
rect 3884 5355 3936 5364
rect 3884 5321 3893 5355
rect 3893 5321 3927 5355
rect 3927 5321 3936 5355
rect 3884 5312 3936 5321
rect 5724 5312 5776 5364
rect 2688 5244 2740 5296
rect 4160 5244 4212 5296
rect 1308 5176 1360 5228
rect 1860 5176 1912 5228
rect 2412 5176 2464 5228
rect 3240 5176 3292 5228
rect 4068 5176 4120 5228
rect 4252 5219 4304 5228
rect 4252 5185 4261 5219
rect 4261 5185 4295 5219
rect 4295 5185 4304 5219
rect 4252 5176 4304 5185
rect 4528 5219 4580 5228
rect 4528 5185 4537 5219
rect 4537 5185 4571 5219
rect 4571 5185 4580 5219
rect 4528 5176 4580 5185
rect 7472 5244 7524 5296
rect 3056 5108 3108 5160
rect 3700 5108 3752 5160
rect 3792 5040 3844 5092
rect 2228 4972 2280 5024
rect 5816 5176 5868 5228
rect 7288 5176 7340 5228
rect 8208 5219 8260 5228
rect 7012 5151 7064 5160
rect 7012 5117 7021 5151
rect 7021 5117 7055 5151
rect 7055 5117 7064 5151
rect 7012 5108 7064 5117
rect 5908 5040 5960 5092
rect 7196 5108 7248 5160
rect 8208 5185 8217 5219
rect 8217 5185 8251 5219
rect 8251 5185 8260 5219
rect 8208 5176 8260 5185
rect 9680 5176 9732 5228
rect 9404 5040 9456 5092
rect 5816 4972 5868 5024
rect 6736 4972 6788 5024
rect 7380 5015 7432 5024
rect 7380 4981 7389 5015
rect 7389 4981 7423 5015
rect 7423 4981 7432 5015
rect 7380 4972 7432 4981
rect 8484 5015 8536 5024
rect 8484 4981 8493 5015
rect 8493 4981 8527 5015
rect 8527 4981 8536 5015
rect 8484 4972 8536 4981
rect 8944 4972 8996 5024
rect 9220 5015 9272 5024
rect 9220 4981 9229 5015
rect 9229 4981 9263 5015
rect 9263 4981 9272 5015
rect 9220 4972 9272 4981
rect 10876 5244 10928 5296
rect 11244 5176 11296 5228
rect 12164 5244 12216 5296
rect 13820 5312 13872 5364
rect 15200 5312 15252 5364
rect 15292 5355 15344 5364
rect 15292 5321 15301 5355
rect 15301 5321 15335 5355
rect 15335 5321 15344 5355
rect 16488 5355 16540 5364
rect 15292 5312 15344 5321
rect 15016 5244 15068 5296
rect 15752 5287 15804 5296
rect 15752 5253 15761 5287
rect 15761 5253 15795 5287
rect 15795 5253 15804 5287
rect 15752 5244 15804 5253
rect 11152 5108 11204 5160
rect 12164 5151 12216 5160
rect 12164 5117 12173 5151
rect 12173 5117 12207 5151
rect 12207 5117 12216 5151
rect 12164 5108 12216 5117
rect 12900 5108 12952 5160
rect 14004 5176 14056 5228
rect 14280 5176 14332 5228
rect 14924 5219 14976 5228
rect 14924 5185 14933 5219
rect 14933 5185 14967 5219
rect 14967 5185 14976 5219
rect 14924 5176 14976 5185
rect 15476 5176 15528 5228
rect 16488 5321 16497 5355
rect 16497 5321 16531 5355
rect 16531 5321 16540 5355
rect 16488 5312 16540 5321
rect 16856 5312 16908 5364
rect 17040 5355 17092 5364
rect 17040 5321 17049 5355
rect 17049 5321 17083 5355
rect 17083 5321 17092 5355
rect 17040 5312 17092 5321
rect 15936 5176 15988 5228
rect 17592 5219 17644 5228
rect 17592 5185 17601 5219
rect 17601 5185 17635 5219
rect 17635 5185 17644 5219
rect 17592 5176 17644 5185
rect 14004 5040 14056 5092
rect 16028 5108 16080 5160
rect 16856 5108 16908 5160
rect 17132 5151 17184 5160
rect 17132 5117 17141 5151
rect 17141 5117 17175 5151
rect 17175 5117 17184 5151
rect 17132 5108 17184 5117
rect 16212 5040 16264 5092
rect 18604 5176 18656 5228
rect 18420 5083 18472 5092
rect 18420 5049 18429 5083
rect 18429 5049 18463 5083
rect 18463 5049 18472 5083
rect 18420 5040 18472 5049
rect 16304 5015 16356 5024
rect 16304 4981 16313 5015
rect 16313 4981 16347 5015
rect 16347 4981 16356 5015
rect 16304 4972 16356 4981
rect 18052 5015 18104 5024
rect 18052 4981 18061 5015
rect 18061 4981 18095 5015
rect 18095 4981 18104 5015
rect 18052 4972 18104 4981
rect 3174 4870 3226 4922
rect 3238 4870 3290 4922
rect 3302 4870 3354 4922
rect 3366 4870 3418 4922
rect 3430 4870 3482 4922
rect 7622 4870 7674 4922
rect 7686 4870 7738 4922
rect 7750 4870 7802 4922
rect 7814 4870 7866 4922
rect 7878 4870 7930 4922
rect 12070 4870 12122 4922
rect 12134 4870 12186 4922
rect 12198 4870 12250 4922
rect 12262 4870 12314 4922
rect 12326 4870 12378 4922
rect 16518 4870 16570 4922
rect 16582 4870 16634 4922
rect 16646 4870 16698 4922
rect 16710 4870 16762 4922
rect 16774 4870 16826 4922
rect 1492 4811 1544 4820
rect 1492 4777 1501 4811
rect 1501 4777 1535 4811
rect 1535 4777 1544 4811
rect 1492 4768 1544 4777
rect 2320 4768 2372 4820
rect 2780 4768 2832 4820
rect 7196 4768 7248 4820
rect 8024 4768 8076 4820
rect 10416 4768 10468 4820
rect 10968 4768 11020 4820
rect 2412 4700 2464 4752
rect 12716 4768 12768 4820
rect 2320 4607 2372 4616
rect 2320 4573 2329 4607
rect 2329 4573 2363 4607
rect 2363 4573 2372 4607
rect 2320 4564 2372 4573
rect 2688 4564 2740 4616
rect 2872 4607 2924 4616
rect 2872 4573 2881 4607
rect 2881 4573 2915 4607
rect 2915 4573 2924 4607
rect 2872 4564 2924 4573
rect 11888 4700 11940 4752
rect 14004 4700 14056 4752
rect 14188 4700 14240 4752
rect 16212 4700 16264 4752
rect 6092 4632 6144 4684
rect 6736 4675 6788 4684
rect 6736 4641 6745 4675
rect 6745 4641 6779 4675
rect 6779 4641 6788 4675
rect 6736 4632 6788 4641
rect 6828 4632 6880 4684
rect 4252 4607 4304 4616
rect 4252 4573 4261 4607
rect 4261 4573 4295 4607
rect 4295 4573 4304 4607
rect 6644 4607 6696 4616
rect 4252 4564 4304 4573
rect 3792 4539 3844 4548
rect 1860 4471 1912 4480
rect 1860 4437 1869 4471
rect 1869 4437 1903 4471
rect 1903 4437 1912 4471
rect 1860 4428 1912 4437
rect 2504 4428 2556 4480
rect 3792 4505 3801 4539
rect 3801 4505 3835 4539
rect 3835 4505 3844 4539
rect 3792 4496 3844 4505
rect 6644 4573 6653 4607
rect 6653 4573 6687 4607
rect 6687 4573 6696 4607
rect 6644 4564 6696 4573
rect 7472 4607 7524 4616
rect 7472 4573 7481 4607
rect 7481 4573 7515 4607
rect 7515 4573 7524 4607
rect 7472 4564 7524 4573
rect 8300 4607 8352 4616
rect 8300 4573 8309 4607
rect 8309 4573 8343 4607
rect 8343 4573 8352 4607
rect 8300 4564 8352 4573
rect 9772 4632 9824 4684
rect 10876 4632 10928 4684
rect 11428 4632 11480 4684
rect 12532 4632 12584 4684
rect 12808 4632 12860 4684
rect 10048 4564 10100 4616
rect 3240 4471 3292 4480
rect 3240 4437 3249 4471
rect 3249 4437 3283 4471
rect 3283 4437 3292 4471
rect 3240 4428 3292 4437
rect 4068 4471 4120 4480
rect 4068 4437 4077 4471
rect 4077 4437 4111 4471
rect 4111 4437 4120 4471
rect 4068 4428 4120 4437
rect 6092 4428 6144 4480
rect 10140 4496 10192 4548
rect 9588 4428 9640 4480
rect 9680 4428 9732 4480
rect 13360 4564 13412 4616
rect 13728 4632 13780 4684
rect 15016 4632 15068 4684
rect 15752 4675 15804 4684
rect 13820 4564 13872 4616
rect 14648 4564 14700 4616
rect 14924 4607 14976 4616
rect 14924 4573 14933 4607
rect 14933 4573 14967 4607
rect 14967 4573 14976 4607
rect 14924 4564 14976 4573
rect 15752 4641 15761 4675
rect 15761 4641 15795 4675
rect 15795 4641 15804 4675
rect 15752 4632 15804 4641
rect 16396 4632 16448 4684
rect 16764 4564 16816 4616
rect 14280 4539 14332 4548
rect 14280 4505 14289 4539
rect 14289 4505 14323 4539
rect 14323 4505 14332 4539
rect 14280 4496 14332 4505
rect 18144 4700 18196 4752
rect 18052 4564 18104 4616
rect 18328 4564 18380 4616
rect 10784 4471 10836 4480
rect 10784 4437 10793 4471
rect 10793 4437 10827 4471
rect 10827 4437 10836 4471
rect 10784 4428 10836 4437
rect 10876 4471 10928 4480
rect 10876 4437 10885 4471
rect 10885 4437 10919 4471
rect 10919 4437 10928 4471
rect 10876 4428 10928 4437
rect 14096 4428 14148 4480
rect 16120 4471 16172 4480
rect 16120 4437 16129 4471
rect 16129 4437 16163 4471
rect 16163 4437 16172 4471
rect 16120 4428 16172 4437
rect 16396 4471 16448 4480
rect 16396 4437 16405 4471
rect 16405 4437 16439 4471
rect 16439 4437 16448 4471
rect 16396 4428 16448 4437
rect 16856 4428 16908 4480
rect 17224 4428 17276 4480
rect 17316 4471 17368 4480
rect 17316 4437 17325 4471
rect 17325 4437 17359 4471
rect 17359 4437 17368 4471
rect 17868 4471 17920 4480
rect 17316 4428 17368 4437
rect 17868 4437 17877 4471
rect 17877 4437 17911 4471
rect 17911 4437 17920 4471
rect 17868 4428 17920 4437
rect 17960 4471 18012 4480
rect 17960 4437 17969 4471
rect 17969 4437 18003 4471
rect 18003 4437 18012 4471
rect 18420 4471 18472 4480
rect 17960 4428 18012 4437
rect 18420 4437 18429 4471
rect 18429 4437 18463 4471
rect 18463 4437 18472 4471
rect 18420 4428 18472 4437
rect 5398 4326 5450 4378
rect 5462 4326 5514 4378
rect 5526 4326 5578 4378
rect 5590 4326 5642 4378
rect 5654 4326 5706 4378
rect 9846 4326 9898 4378
rect 9910 4326 9962 4378
rect 9974 4326 10026 4378
rect 10038 4326 10090 4378
rect 10102 4326 10154 4378
rect 14294 4326 14346 4378
rect 14358 4326 14410 4378
rect 14422 4326 14474 4378
rect 14486 4326 14538 4378
rect 14550 4326 14602 4378
rect 4804 4224 4856 4276
rect 5540 4224 5592 4276
rect 6092 4267 6144 4276
rect 3240 4156 3292 4208
rect 5816 4156 5868 4208
rect 6092 4233 6101 4267
rect 6101 4233 6135 4267
rect 6135 4233 6144 4267
rect 6092 4224 6144 4233
rect 6644 4224 6696 4276
rect 7012 4224 7064 4276
rect 16396 4224 16448 4276
rect 6828 4156 6880 4208
rect 8944 4156 8996 4208
rect 1492 3995 1544 4004
rect 1492 3961 1501 3995
rect 1501 3961 1535 3995
rect 1535 3961 1544 3995
rect 1492 3952 1544 3961
rect 2596 4131 2648 4140
rect 2596 4097 2605 4131
rect 2605 4097 2639 4131
rect 2639 4097 2648 4131
rect 2596 4088 2648 4097
rect 2872 4131 2924 4140
rect 2872 4097 2881 4131
rect 2881 4097 2915 4131
rect 2915 4097 2924 4131
rect 2872 4088 2924 4097
rect 2688 4020 2740 4072
rect 3516 4088 3568 4140
rect 3884 4131 3936 4140
rect 3884 4097 3893 4131
rect 3893 4097 3927 4131
rect 3927 4097 3936 4131
rect 3884 4088 3936 4097
rect 6460 4088 6512 4140
rect 8300 4088 8352 4140
rect 9128 4131 9180 4140
rect 9128 4097 9137 4131
rect 9137 4097 9171 4131
rect 9171 4097 9180 4131
rect 10784 4156 10836 4208
rect 9128 4088 9180 4097
rect 11796 4088 11848 4140
rect 13268 4088 13320 4140
rect 13820 4088 13872 4140
rect 14464 4131 14516 4140
rect 14464 4097 14482 4131
rect 14482 4097 14516 4131
rect 14464 4088 14516 4097
rect 4160 4020 4212 4072
rect 4712 4020 4764 4072
rect 5540 4063 5592 4072
rect 5540 4029 5549 4063
rect 5549 4029 5583 4063
rect 5583 4029 5592 4063
rect 5540 4020 5592 4029
rect 6184 4020 6236 4072
rect 2780 3952 2832 4004
rect 2872 3952 2924 4004
rect 7472 4020 7524 4072
rect 9588 4020 9640 4072
rect 10692 4020 10744 4072
rect 1860 3927 1912 3936
rect 1860 3893 1869 3927
rect 1869 3893 1903 3927
rect 1903 3893 1912 3927
rect 1860 3884 1912 3893
rect 1952 3884 2004 3936
rect 2688 3927 2740 3936
rect 2688 3893 2697 3927
rect 2697 3893 2731 3927
rect 2731 3893 2740 3927
rect 2688 3884 2740 3893
rect 2964 3927 3016 3936
rect 2964 3893 2973 3927
rect 2973 3893 3007 3927
rect 3007 3893 3016 3927
rect 2964 3884 3016 3893
rect 3700 3927 3752 3936
rect 3700 3893 3709 3927
rect 3709 3893 3743 3927
rect 3743 3893 3752 3927
rect 3700 3884 3752 3893
rect 6736 3884 6788 3936
rect 8484 3884 8536 3936
rect 8852 3927 8904 3936
rect 8852 3893 8861 3927
rect 8861 3893 8895 3927
rect 8895 3893 8904 3927
rect 8852 3884 8904 3893
rect 12624 4020 12676 4072
rect 13176 4020 13228 4072
rect 15660 4063 15712 4072
rect 15660 4029 15669 4063
rect 15669 4029 15703 4063
rect 15703 4029 15712 4063
rect 15660 4020 15712 4029
rect 17040 4088 17092 4140
rect 17592 4131 17644 4140
rect 17592 4097 17601 4131
rect 17601 4097 17635 4131
rect 17635 4097 17644 4131
rect 17592 4088 17644 4097
rect 17776 4088 17828 4140
rect 17960 4088 18012 4140
rect 10324 3884 10376 3936
rect 13452 3952 13504 4004
rect 16396 3952 16448 4004
rect 12808 3884 12860 3936
rect 13084 3927 13136 3936
rect 13084 3893 13093 3927
rect 13093 3893 13127 3927
rect 13127 3893 13136 3927
rect 13084 3884 13136 3893
rect 13268 3927 13320 3936
rect 13268 3893 13277 3927
rect 13277 3893 13311 3927
rect 13311 3893 13320 3927
rect 13636 3927 13688 3936
rect 13268 3884 13320 3893
rect 13636 3893 13645 3927
rect 13645 3893 13679 3927
rect 13679 3893 13688 3927
rect 13636 3884 13688 3893
rect 13820 3927 13872 3936
rect 13820 3893 13829 3927
rect 13829 3893 13863 3927
rect 13863 3893 13872 3927
rect 13820 3884 13872 3893
rect 14004 3884 14056 3936
rect 14648 3884 14700 3936
rect 17040 3952 17092 4004
rect 18880 3952 18932 4004
rect 17132 3927 17184 3936
rect 17132 3893 17141 3927
rect 17141 3893 17175 3927
rect 17175 3893 17184 3927
rect 17132 3884 17184 3893
rect 17684 3884 17736 3936
rect 18420 3927 18472 3936
rect 18420 3893 18429 3927
rect 18429 3893 18463 3927
rect 18463 3893 18472 3927
rect 18420 3884 18472 3893
rect 3174 3782 3226 3834
rect 3238 3782 3290 3834
rect 3302 3782 3354 3834
rect 3366 3782 3418 3834
rect 3430 3782 3482 3834
rect 7622 3782 7674 3834
rect 7686 3782 7738 3834
rect 7750 3782 7802 3834
rect 7814 3782 7866 3834
rect 7878 3782 7930 3834
rect 12070 3782 12122 3834
rect 12134 3782 12186 3834
rect 12198 3782 12250 3834
rect 12262 3782 12314 3834
rect 12326 3782 12378 3834
rect 16518 3782 16570 3834
rect 16582 3782 16634 3834
rect 16646 3782 16698 3834
rect 16710 3782 16762 3834
rect 16774 3782 16826 3834
rect 2596 3680 2648 3732
rect 3700 3680 3752 3732
rect 9404 3680 9456 3732
rect 10048 3680 10100 3732
rect 12624 3680 12676 3732
rect 13176 3680 13228 3732
rect 2780 3612 2832 3664
rect 1952 3476 2004 3528
rect 2688 3544 2740 3596
rect 8116 3612 8168 3664
rect 10324 3612 10376 3664
rect 12532 3655 12584 3664
rect 12532 3621 12541 3655
rect 12541 3621 12575 3655
rect 12575 3621 12584 3655
rect 12532 3612 12584 3621
rect 13636 3612 13688 3664
rect 13912 3680 13964 3732
rect 16396 3680 16448 3732
rect 16948 3612 17000 3664
rect 18512 3612 18564 3664
rect 2412 3519 2464 3528
rect 2412 3485 2421 3519
rect 2421 3485 2455 3519
rect 2455 3485 2464 3519
rect 2412 3476 2464 3485
rect 2504 3519 2556 3528
rect 2504 3485 2513 3519
rect 2513 3485 2547 3519
rect 2547 3485 2556 3519
rect 2504 3476 2556 3485
rect 3516 3476 3568 3528
rect 3792 3519 3844 3528
rect 3792 3485 3801 3519
rect 3801 3485 3835 3519
rect 3835 3485 3844 3519
rect 3792 3476 3844 3485
rect 7380 3544 7432 3596
rect 8484 3587 8536 3596
rect 8484 3553 8493 3587
rect 8493 3553 8527 3587
rect 8527 3553 8536 3587
rect 8484 3544 8536 3553
rect 8668 3587 8720 3596
rect 8668 3553 8677 3587
rect 8677 3553 8711 3587
rect 8711 3553 8720 3587
rect 8668 3544 8720 3553
rect 6736 3519 6788 3528
rect 6736 3485 6745 3519
rect 6745 3485 6779 3519
rect 6779 3485 6788 3519
rect 6736 3476 6788 3485
rect 8944 3476 8996 3528
rect 1492 3383 1544 3392
rect 1492 3349 1501 3383
rect 1501 3349 1535 3383
rect 1535 3349 1544 3383
rect 1492 3340 1544 3349
rect 1860 3383 1912 3392
rect 1860 3349 1869 3383
rect 1869 3349 1903 3383
rect 1903 3349 1912 3383
rect 1860 3340 1912 3349
rect 2228 3383 2280 3392
rect 2228 3349 2237 3383
rect 2237 3349 2271 3383
rect 2271 3349 2280 3383
rect 2228 3340 2280 3349
rect 2688 3383 2740 3392
rect 2688 3349 2697 3383
rect 2697 3349 2731 3383
rect 2731 3349 2740 3383
rect 2688 3340 2740 3349
rect 3148 3383 3200 3392
rect 3148 3349 3157 3383
rect 3157 3349 3191 3383
rect 3191 3349 3200 3383
rect 3148 3340 3200 3349
rect 3332 3340 3384 3392
rect 4252 3340 4304 3392
rect 5816 3340 5868 3392
rect 6736 3340 6788 3392
rect 8576 3408 8628 3460
rect 9588 3519 9640 3528
rect 9588 3485 9632 3519
rect 9632 3485 9640 3519
rect 9588 3476 9640 3485
rect 9772 3476 9824 3528
rect 10048 3519 10100 3528
rect 10048 3485 10057 3519
rect 10057 3485 10091 3519
rect 10091 3485 10100 3519
rect 10048 3476 10100 3485
rect 10784 3476 10836 3528
rect 11060 3544 11112 3596
rect 14464 3544 14516 3596
rect 15844 3587 15896 3596
rect 11336 3519 11388 3528
rect 11336 3485 11345 3519
rect 11345 3485 11379 3519
rect 11379 3485 11388 3519
rect 11336 3476 11388 3485
rect 11520 3451 11572 3460
rect 11520 3417 11529 3451
rect 11529 3417 11563 3451
rect 11563 3417 11572 3451
rect 11520 3408 11572 3417
rect 12808 3519 12860 3528
rect 12808 3485 12817 3519
rect 12817 3485 12851 3519
rect 12851 3485 12860 3519
rect 12808 3476 12860 3485
rect 12624 3408 12676 3460
rect 13360 3519 13412 3528
rect 13360 3485 13404 3519
rect 13404 3485 13412 3519
rect 13360 3476 13412 3485
rect 13728 3476 13780 3528
rect 14004 3476 14056 3528
rect 15844 3553 15853 3587
rect 15853 3553 15887 3587
rect 15887 3553 15896 3587
rect 15844 3544 15896 3553
rect 16948 3519 17000 3528
rect 15568 3408 15620 3460
rect 16948 3485 16957 3519
rect 16957 3485 16991 3519
rect 16991 3485 17000 3519
rect 16948 3476 17000 3485
rect 17500 3519 17552 3528
rect 16304 3408 16356 3460
rect 17500 3485 17509 3519
rect 17509 3485 17543 3519
rect 17543 3485 17552 3519
rect 17500 3476 17552 3485
rect 17868 3519 17920 3528
rect 17868 3485 17877 3519
rect 17877 3485 17911 3519
rect 17911 3485 17920 3519
rect 17868 3476 17920 3485
rect 18052 3476 18104 3528
rect 18696 3476 18748 3528
rect 7012 3383 7064 3392
rect 7012 3349 7021 3383
rect 7021 3349 7055 3383
rect 7055 3349 7064 3383
rect 7012 3340 7064 3349
rect 7840 3340 7892 3392
rect 8668 3340 8720 3392
rect 9220 3340 9272 3392
rect 9680 3340 9732 3392
rect 9864 3383 9916 3392
rect 9864 3349 9873 3383
rect 9873 3349 9907 3383
rect 9907 3349 9916 3383
rect 9864 3340 9916 3349
rect 10232 3340 10284 3392
rect 10692 3340 10744 3392
rect 10968 3340 11020 3392
rect 11152 3383 11204 3392
rect 11152 3349 11161 3383
rect 11161 3349 11195 3383
rect 11195 3349 11204 3383
rect 11612 3383 11664 3392
rect 11152 3340 11204 3349
rect 11612 3349 11621 3383
rect 11621 3349 11655 3383
rect 11655 3349 11664 3383
rect 11612 3340 11664 3349
rect 12440 3383 12492 3392
rect 12440 3349 12449 3383
rect 12449 3349 12483 3383
rect 12483 3349 12492 3383
rect 12992 3383 13044 3392
rect 12440 3340 12492 3349
rect 12992 3349 13001 3383
rect 13001 3349 13035 3383
rect 13035 3349 13044 3383
rect 12992 3340 13044 3349
rect 13636 3340 13688 3392
rect 17592 3340 17644 3392
rect 18052 3383 18104 3392
rect 18052 3349 18061 3383
rect 18061 3349 18095 3383
rect 18095 3349 18104 3383
rect 18052 3340 18104 3349
rect 18420 3383 18472 3392
rect 18420 3349 18429 3383
rect 18429 3349 18463 3383
rect 18463 3349 18472 3383
rect 18420 3340 18472 3349
rect 5398 3238 5450 3290
rect 5462 3238 5514 3290
rect 5526 3238 5578 3290
rect 5590 3238 5642 3290
rect 5654 3238 5706 3290
rect 9846 3238 9898 3290
rect 9910 3238 9962 3290
rect 9974 3238 10026 3290
rect 10038 3238 10090 3290
rect 10102 3238 10154 3290
rect 14294 3238 14346 3290
rect 14358 3238 14410 3290
rect 14422 3238 14474 3290
rect 14486 3238 14538 3290
rect 14550 3238 14602 3290
rect 940 3068 992 3120
rect 2412 3068 2464 3120
rect 1400 3043 1452 3052
rect 1400 3009 1409 3043
rect 1409 3009 1443 3043
rect 1443 3009 1452 3043
rect 1400 3000 1452 3009
rect 2136 3043 2188 3052
rect 2136 3009 2145 3043
rect 2145 3009 2179 3043
rect 2179 3009 2188 3043
rect 2136 3000 2188 3009
rect 2596 3043 2648 3052
rect 2596 3009 2605 3043
rect 2605 3009 2639 3043
rect 2639 3009 2648 3043
rect 2596 3000 2648 3009
rect 3332 3043 3384 3052
rect 3332 3009 3341 3043
rect 3341 3009 3375 3043
rect 3375 3009 3384 3043
rect 3332 3000 3384 3009
rect 4068 3000 4120 3052
rect 4988 3043 5040 3052
rect 4988 3009 4997 3043
rect 4997 3009 5031 3043
rect 5031 3009 5040 3043
rect 4988 3000 5040 3009
rect 2596 2864 2648 2916
rect 1400 2796 1452 2848
rect 2412 2796 2464 2848
rect 4160 2864 4212 2916
rect 6736 3043 6788 3052
rect 6736 3009 6745 3043
rect 6745 3009 6779 3043
rect 6779 3009 6788 3043
rect 6736 3000 6788 3009
rect 9588 3136 9640 3188
rect 10876 3136 10928 3188
rect 7840 3068 7892 3120
rect 9680 3068 9732 3120
rect 11704 3136 11756 3188
rect 12900 3136 12952 3188
rect 13728 3136 13780 3188
rect 14740 3136 14792 3188
rect 16948 3136 17000 3188
rect 13636 3111 13688 3120
rect 13636 3077 13645 3111
rect 13645 3077 13679 3111
rect 13679 3077 13688 3111
rect 13636 3068 13688 3077
rect 14372 3068 14424 3120
rect 7104 3043 7156 3052
rect 7104 3009 7113 3043
rect 7113 3009 7147 3043
rect 7147 3009 7156 3043
rect 7104 3000 7156 3009
rect 6920 2932 6972 2984
rect 8208 2975 8260 2984
rect 8208 2941 8217 2975
rect 8217 2941 8251 2975
rect 8251 2941 8260 2975
rect 8208 2932 8260 2941
rect 9496 2975 9548 2984
rect 9496 2941 9505 2975
rect 9505 2941 9539 2975
rect 9539 2941 9548 2975
rect 9496 2932 9548 2941
rect 11612 3000 11664 3052
rect 13452 3043 13504 3052
rect 13452 3009 13461 3043
rect 13461 3009 13495 3043
rect 13495 3009 13504 3043
rect 13452 3000 13504 3009
rect 14924 3000 14976 3052
rect 17224 3068 17276 3120
rect 11428 2932 11480 2984
rect 13176 2975 13228 2984
rect 13176 2941 13185 2975
rect 13185 2941 13219 2975
rect 13219 2941 13228 2975
rect 13176 2932 13228 2941
rect 13360 2975 13412 2984
rect 13360 2941 13369 2975
rect 13369 2941 13403 2975
rect 13403 2941 13412 2975
rect 13360 2932 13412 2941
rect 14648 2975 14700 2984
rect 14648 2941 14657 2975
rect 14657 2941 14691 2975
rect 14691 2941 14700 2975
rect 14648 2932 14700 2941
rect 12808 2864 12860 2916
rect 12992 2864 13044 2916
rect 16856 3000 16908 3052
rect 17408 3043 17460 3052
rect 17408 3009 17417 3043
rect 17417 3009 17451 3043
rect 17451 3009 17460 3043
rect 17408 3000 17460 3009
rect 18236 3043 18288 3052
rect 17316 2932 17368 2984
rect 18236 3009 18245 3043
rect 18245 3009 18279 3043
rect 18279 3009 18288 3043
rect 18236 3000 18288 3009
rect 16304 2864 16356 2916
rect 18328 2864 18380 2916
rect 2872 2796 2924 2848
rect 3516 2839 3568 2848
rect 3516 2805 3525 2839
rect 3525 2805 3559 2839
rect 3559 2805 3568 2839
rect 3516 2796 3568 2805
rect 3976 2839 4028 2848
rect 3976 2805 3985 2839
rect 3985 2805 4019 2839
rect 4019 2805 4028 2839
rect 3976 2796 4028 2805
rect 4988 2796 5040 2848
rect 5540 2796 5592 2848
rect 7104 2796 7156 2848
rect 7288 2839 7340 2848
rect 7288 2805 7297 2839
rect 7297 2805 7331 2839
rect 7331 2805 7340 2839
rect 7288 2796 7340 2805
rect 7380 2796 7432 2848
rect 10876 2796 10928 2848
rect 11060 2796 11112 2848
rect 15200 2796 15252 2848
rect 15660 2796 15712 2848
rect 16120 2839 16172 2848
rect 16120 2805 16129 2839
rect 16129 2805 16163 2839
rect 16163 2805 16172 2839
rect 16120 2796 16172 2805
rect 16948 2839 17000 2848
rect 16948 2805 16957 2839
rect 16957 2805 16991 2839
rect 16991 2805 17000 2839
rect 16948 2796 17000 2805
rect 17868 2796 17920 2848
rect 18420 2839 18472 2848
rect 18420 2805 18429 2839
rect 18429 2805 18463 2839
rect 18463 2805 18472 2839
rect 18420 2796 18472 2805
rect 3174 2694 3226 2746
rect 3238 2694 3290 2746
rect 3302 2694 3354 2746
rect 3366 2694 3418 2746
rect 3430 2694 3482 2746
rect 7622 2694 7674 2746
rect 7686 2694 7738 2746
rect 7750 2694 7802 2746
rect 7814 2694 7866 2746
rect 7878 2694 7930 2746
rect 12070 2694 12122 2746
rect 12134 2694 12186 2746
rect 12198 2694 12250 2746
rect 12262 2694 12314 2746
rect 12326 2694 12378 2746
rect 16518 2694 16570 2746
rect 16582 2694 16634 2746
rect 16646 2694 16698 2746
rect 16710 2694 16762 2746
rect 16774 2694 16826 2746
rect 1492 2635 1544 2644
rect 1492 2601 1501 2635
rect 1501 2601 1535 2635
rect 1535 2601 1544 2635
rect 1492 2592 1544 2601
rect 2136 2592 2188 2644
rect 5172 2635 5224 2644
rect 5172 2601 5181 2635
rect 5181 2601 5215 2635
rect 5215 2601 5224 2635
rect 5172 2592 5224 2601
rect 6368 2592 6420 2644
rect 10968 2592 11020 2644
rect 11980 2592 12032 2644
rect 13360 2592 13412 2644
rect 2780 2524 2832 2576
rect 2964 2456 3016 2508
rect 3056 2388 3108 2440
rect 5540 2456 5592 2508
rect 4160 2388 4212 2440
rect 4988 2431 5040 2440
rect 4252 2320 4304 2372
rect 4988 2397 4997 2431
rect 4997 2397 5031 2431
rect 5031 2397 5040 2431
rect 4988 2388 5040 2397
rect 5080 2388 5132 2440
rect 10324 2524 10376 2576
rect 11152 2524 11204 2576
rect 11428 2524 11480 2576
rect 14832 2524 14884 2576
rect 7288 2456 7340 2508
rect 6000 2431 6052 2440
rect 6000 2397 6009 2431
rect 6009 2397 6043 2431
rect 6043 2397 6052 2431
rect 6000 2388 6052 2397
rect 6552 2431 6604 2440
rect 6552 2397 6561 2431
rect 6561 2397 6595 2431
rect 6595 2397 6604 2431
rect 6552 2388 6604 2397
rect 7012 2431 7064 2440
rect 7012 2397 7021 2431
rect 7021 2397 7055 2431
rect 7055 2397 7064 2431
rect 7012 2388 7064 2397
rect 7104 2388 7156 2440
rect 8668 2431 8720 2440
rect 8668 2397 8677 2431
rect 8677 2397 8711 2431
rect 8711 2397 8720 2431
rect 8668 2388 8720 2397
rect 9220 2431 9272 2440
rect 9220 2397 9229 2431
rect 9229 2397 9263 2431
rect 9263 2397 9272 2431
rect 9220 2388 9272 2397
rect 9772 2388 9824 2440
rect 10232 2388 10284 2440
rect 12532 2456 12584 2508
rect 13544 2499 13596 2508
rect 13544 2465 13553 2499
rect 13553 2465 13587 2499
rect 13587 2465 13596 2499
rect 13544 2456 13596 2465
rect 14188 2499 14240 2508
rect 14188 2465 14197 2499
rect 14197 2465 14231 2499
rect 14231 2465 14240 2499
rect 14188 2456 14240 2465
rect 15200 2456 15252 2508
rect 16580 2524 16632 2576
rect 10692 2431 10744 2440
rect 10692 2397 10701 2431
rect 10701 2397 10735 2431
rect 10735 2397 10744 2431
rect 10692 2388 10744 2397
rect 5816 2320 5868 2372
rect 11244 2388 11296 2440
rect 16120 2431 16172 2440
rect 11336 2320 11388 2372
rect 1860 2252 1912 2304
rect 2320 2252 2372 2304
rect 2780 2252 2832 2304
rect 3240 2252 3292 2304
rect 3700 2252 3752 2304
rect 4160 2252 4212 2304
rect 4620 2252 4672 2304
rect 5080 2252 5132 2304
rect 5724 2295 5776 2304
rect 5724 2261 5733 2295
rect 5733 2261 5767 2295
rect 5767 2261 5776 2295
rect 5724 2252 5776 2261
rect 6460 2252 6512 2304
rect 6920 2252 6972 2304
rect 7380 2252 7432 2304
rect 7840 2252 7892 2304
rect 8300 2252 8352 2304
rect 8760 2252 8812 2304
rect 9220 2252 9272 2304
rect 9680 2252 9732 2304
rect 10232 2252 10284 2304
rect 10600 2252 10652 2304
rect 11980 2363 12032 2372
rect 11980 2329 11989 2363
rect 11989 2329 12023 2363
rect 12023 2329 12032 2363
rect 11980 2320 12032 2329
rect 12256 2320 12308 2372
rect 12992 2320 13044 2372
rect 16120 2397 16129 2431
rect 16129 2397 16163 2431
rect 16163 2397 16172 2431
rect 16120 2388 16172 2397
rect 16212 2388 16264 2440
rect 17040 2431 17092 2440
rect 17040 2397 17049 2431
rect 17049 2397 17083 2431
rect 17083 2397 17092 2431
rect 17040 2388 17092 2397
rect 17132 2388 17184 2440
rect 17684 2388 17736 2440
rect 18144 2431 18196 2440
rect 18144 2397 18153 2431
rect 18153 2397 18187 2431
rect 18187 2397 18196 2431
rect 18144 2388 18196 2397
rect 13176 2252 13228 2304
rect 15200 2252 15252 2304
rect 16396 2252 16448 2304
rect 17040 2252 17092 2304
rect 17776 2252 17828 2304
rect 18052 2252 18104 2304
rect 5398 2150 5450 2202
rect 5462 2150 5514 2202
rect 5526 2150 5578 2202
rect 5590 2150 5642 2202
rect 5654 2150 5706 2202
rect 9846 2150 9898 2202
rect 9910 2150 9962 2202
rect 9974 2150 10026 2202
rect 10038 2150 10090 2202
rect 10102 2150 10154 2202
rect 14294 2150 14346 2202
rect 14358 2150 14410 2202
rect 14422 2150 14474 2202
rect 14486 2150 14538 2202
rect 14550 2150 14602 2202
<< metal2 >>
rect 294 16400 350 17200
rect 938 16400 994 17200
rect 1582 16400 1638 17200
rect 2226 16538 2282 17200
rect 2226 16510 2544 16538
rect 2226 16400 2282 16510
rect 308 13258 336 16400
rect 952 13802 980 16400
rect 940 13796 992 13802
rect 940 13738 992 13744
rect 296 13252 348 13258
rect 296 13194 348 13200
rect 1596 13190 1624 16400
rect 2136 14952 2188 14958
rect 2136 14894 2188 14900
rect 1952 14408 2004 14414
rect 1950 14376 1952 14385
rect 2004 14376 2006 14385
rect 1950 14311 2006 14320
rect 2044 14000 2096 14006
rect 2044 13942 2096 13948
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1964 13394 1992 13670
rect 2056 13433 2084 13942
rect 2148 13938 2176 14894
rect 2228 14408 2280 14414
rect 2228 14350 2280 14356
rect 2136 13932 2188 13938
rect 2136 13874 2188 13880
rect 2240 13841 2268 14350
rect 2226 13832 2282 13841
rect 2226 13767 2282 13776
rect 2516 13462 2544 16510
rect 2870 16400 2926 17200
rect 3514 16400 3570 17200
rect 3790 16688 3846 16697
rect 3790 16623 3846 16632
rect 2778 15872 2834 15881
rect 2778 15807 2834 15816
rect 2792 14074 2820 15807
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 2884 13530 2912 16400
rect 3054 15056 3110 15065
rect 3054 14991 3110 15000
rect 2962 14648 3018 14657
rect 2962 14583 3018 14592
rect 2976 14550 3004 14583
rect 2964 14544 3016 14550
rect 2964 14486 3016 14492
rect 3068 14260 3096 14991
rect 3174 14716 3482 14725
rect 3174 14714 3180 14716
rect 3236 14714 3260 14716
rect 3316 14714 3340 14716
rect 3396 14714 3420 14716
rect 3476 14714 3482 14716
rect 3236 14662 3238 14714
rect 3418 14662 3420 14714
rect 3174 14660 3180 14662
rect 3236 14660 3260 14662
rect 3316 14660 3340 14662
rect 3396 14660 3420 14662
rect 3476 14660 3482 14662
rect 3174 14651 3482 14660
rect 3528 14618 3556 16400
rect 3804 15230 3832 16623
rect 4158 16538 4214 17200
rect 4158 16510 4384 16538
rect 4158 16400 4214 16510
rect 4066 16280 4122 16289
rect 4066 16215 4122 16224
rect 3792 15224 3844 15230
rect 3792 15166 3844 15172
rect 3976 14816 4028 14822
rect 3976 14758 4028 14764
rect 3516 14612 3568 14618
rect 3516 14554 3568 14560
rect 3606 14512 3662 14521
rect 3988 14482 4016 14758
rect 3606 14447 3662 14456
rect 3976 14476 4028 14482
rect 3620 14414 3648 14447
rect 3976 14418 4028 14424
rect 3608 14408 3660 14414
rect 3608 14350 3660 14356
rect 3148 14272 3200 14278
rect 2962 14240 3018 14249
rect 3068 14232 3148 14260
rect 3148 14214 3200 14220
rect 2962 14175 3018 14184
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2504 13456 2556 13462
rect 2042 13424 2098 13433
rect 1952 13388 2004 13394
rect 2504 13398 2556 13404
rect 2042 13359 2098 13368
rect 1952 13330 2004 13336
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 2872 13320 2924 13326
rect 2872 13262 2924 13268
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 2792 13025 2820 13262
rect 2778 13016 2834 13025
rect 2884 12986 2912 13262
rect 2778 12951 2834 12960
rect 2872 12980 2924 12986
rect 2872 12922 2924 12928
rect 2778 12880 2834 12889
rect 2976 12850 3004 14175
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 3068 13444 3096 14010
rect 3160 13870 3188 14214
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 3148 13864 3200 13870
rect 3148 13806 3200 13812
rect 3174 13628 3482 13637
rect 3174 13626 3180 13628
rect 3236 13626 3260 13628
rect 3316 13626 3340 13628
rect 3396 13626 3420 13628
rect 3476 13626 3482 13628
rect 3236 13574 3238 13626
rect 3418 13574 3420 13626
rect 3174 13572 3180 13574
rect 3236 13572 3260 13574
rect 3316 13572 3340 13574
rect 3396 13572 3420 13574
rect 3476 13572 3482 13574
rect 3174 13563 3482 13572
rect 3528 13530 3556 14010
rect 4080 13938 4108 16215
rect 4158 15464 4214 15473
rect 4158 15399 4214 15408
rect 4172 14482 4200 15399
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 4252 14340 4304 14346
rect 4252 14282 4304 14288
rect 3700 13932 3752 13938
rect 3700 13874 3752 13880
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 3608 13864 3660 13870
rect 3608 13806 3660 13812
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3068 13416 3188 13444
rect 3160 13326 3188 13416
rect 3514 13424 3570 13433
rect 3514 13359 3570 13368
rect 3528 13326 3556 13359
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 3436 12850 3464 13126
rect 2778 12815 2834 12824
rect 2964 12844 3016 12850
rect 2792 12782 2820 12815
rect 2964 12786 3016 12792
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 2136 12776 2188 12782
rect 2136 12718 2188 12724
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 2870 12744 2926 12753
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1308 11280 1360 11286
rect 1308 11222 1360 11228
rect 1320 5234 1348 11222
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1596 10266 1624 10746
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 1490 10160 1546 10169
rect 1490 10095 1546 10104
rect 1504 10062 1532 10095
rect 1492 10056 1544 10062
rect 1492 9998 1544 10004
rect 1676 9920 1728 9926
rect 1676 9862 1728 9868
rect 1490 9616 1546 9625
rect 1490 9551 1492 9560
rect 1544 9551 1546 9560
rect 1492 9522 1544 9528
rect 1504 9353 1532 9522
rect 1490 9344 1546 9353
rect 1490 9279 1546 9288
rect 1492 8832 1544 8838
rect 1492 8774 1544 8780
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 1504 8537 1532 8774
rect 1490 8528 1546 8537
rect 1490 8463 1546 8472
rect 1400 8356 1452 8362
rect 1400 8298 1452 8304
rect 1308 5228 1360 5234
rect 1308 5170 1360 5176
rect 940 3120 992 3126
rect 940 3062 992 3068
rect 952 800 980 3062
rect 1412 3058 1440 8298
rect 1490 8120 1546 8129
rect 1490 8055 1492 8064
rect 1544 8055 1546 8064
rect 1492 8026 1544 8032
rect 1490 7304 1546 7313
rect 1490 7239 1546 7248
rect 1504 7002 1532 7239
rect 1492 6996 1544 7002
rect 1492 6938 1544 6944
rect 1596 6905 1624 8774
rect 1688 7886 1716 9862
rect 1768 9376 1820 9382
rect 1768 9318 1820 9324
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 1676 7336 1728 7342
rect 1676 7278 1728 7284
rect 1688 7002 1716 7278
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 1582 6760 1638 6769
rect 1582 6695 1638 6704
rect 1596 6254 1624 6695
rect 1584 6248 1636 6254
rect 1584 6190 1636 6196
rect 1780 6202 1808 9318
rect 1872 8974 1900 11494
rect 1950 11248 2006 11257
rect 1950 11183 1952 11192
rect 2004 11183 2006 11192
rect 1952 11154 2004 11160
rect 2148 10713 2176 12718
rect 2240 12617 2268 12718
rect 2870 12679 2926 12688
rect 2226 12608 2282 12617
rect 2226 12543 2282 12552
rect 2780 12232 2832 12238
rect 2410 12200 2466 12209
rect 2780 12174 2832 12180
rect 2410 12135 2412 12144
rect 2464 12135 2466 12144
rect 2412 12106 2464 12112
rect 2504 12096 2556 12102
rect 2504 12038 2556 12044
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2228 11688 2280 11694
rect 2228 11630 2280 11636
rect 2240 11393 2268 11630
rect 2226 11384 2282 11393
rect 2226 11319 2282 11328
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2240 10985 2268 11086
rect 2226 10976 2282 10985
rect 2226 10911 2282 10920
rect 2134 10704 2190 10713
rect 2134 10639 2190 10648
rect 2228 10600 2280 10606
rect 2226 10568 2228 10577
rect 2280 10568 2282 10577
rect 2136 10532 2188 10538
rect 2226 10503 2282 10512
rect 2136 10474 2188 10480
rect 1952 10056 2004 10062
rect 1952 9998 2004 10004
rect 1964 9722 1992 9998
rect 2044 9920 2096 9926
rect 2044 9862 2096 9868
rect 1952 9716 2004 9722
rect 1952 9658 2004 9664
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 1950 8936 2006 8945
rect 1950 8871 1952 8880
rect 2004 8871 2006 8880
rect 1952 8842 2004 8848
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 1964 8090 1992 8366
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 1952 7812 2004 7818
rect 1952 7754 2004 7760
rect 1860 7744 1912 7750
rect 1858 7712 1860 7721
rect 1912 7712 1914 7721
rect 1858 7647 1914 7656
rect 1964 7546 1992 7754
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 1780 6174 1900 6202
rect 1768 6112 1820 6118
rect 1490 6080 1546 6089
rect 1768 6054 1820 6060
rect 1490 6015 1546 6024
rect 1504 5370 1532 6015
rect 1674 5808 1730 5817
rect 1780 5778 1808 6054
rect 1674 5743 1676 5752
rect 1728 5743 1730 5752
rect 1768 5772 1820 5778
rect 1676 5714 1728 5720
rect 1768 5714 1820 5720
rect 1492 5364 1544 5370
rect 1492 5306 1544 5312
rect 1872 5234 1900 6174
rect 2056 5710 2084 9862
rect 2148 7834 2176 10474
rect 2240 10266 2268 10503
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2240 8566 2268 9318
rect 2332 8634 2360 9454
rect 2424 9042 2452 11834
rect 2516 11665 2544 12038
rect 2792 11801 2820 12174
rect 2778 11792 2834 11801
rect 2778 11727 2834 11736
rect 2502 11656 2558 11665
rect 2502 11591 2558 11600
rect 2596 11552 2648 11558
rect 2596 11494 2648 11500
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2516 10130 2544 10406
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 2516 9178 2544 9522
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2412 9036 2464 9042
rect 2412 8978 2464 8984
rect 2412 8832 2464 8838
rect 2412 8774 2464 8780
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2228 8560 2280 8566
rect 2228 8502 2280 8508
rect 2318 8528 2374 8537
rect 2318 8463 2374 8472
rect 2332 7886 2360 8463
rect 2320 7880 2372 7886
rect 2148 7806 2268 7834
rect 2320 7822 2372 7828
rect 2136 7744 2188 7750
rect 2136 7686 2188 7692
rect 2148 7546 2176 7686
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 2134 6896 2190 6905
rect 2134 6831 2190 6840
rect 2044 5704 2096 5710
rect 1950 5672 2006 5681
rect 2044 5646 2096 5652
rect 1950 5607 2006 5616
rect 1964 5370 1992 5607
rect 1952 5364 2004 5370
rect 1952 5306 2004 5312
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 1490 4856 1546 4865
rect 1490 4791 1492 4800
rect 1544 4791 1546 4800
rect 1492 4762 1544 4768
rect 1860 4480 1912 4486
rect 1858 4448 1860 4457
rect 1912 4448 1914 4457
rect 1858 4383 1914 4392
rect 1490 4040 1546 4049
rect 1490 3975 1492 3984
rect 1544 3975 1546 3984
rect 1492 3946 1544 3952
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 1872 3641 1900 3878
rect 1858 3632 1914 3641
rect 1858 3567 1914 3576
rect 1964 3534 1992 3878
rect 1952 3528 2004 3534
rect 1952 3470 2004 3476
rect 1492 3392 1544 3398
rect 1492 3334 1544 3340
rect 1860 3392 1912 3398
rect 1860 3334 1912 3340
rect 1504 3233 1532 3334
rect 1490 3224 1546 3233
rect 1490 3159 1546 3168
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1400 2848 1452 2854
rect 1400 2790 1452 2796
rect 1490 2816 1546 2825
rect 1412 800 1440 2790
rect 1490 2751 1546 2760
rect 1504 2650 1532 2751
rect 1492 2644 1544 2650
rect 1492 2586 1544 2592
rect 1872 2417 1900 3334
rect 2148 3058 2176 6831
rect 2240 6730 2268 7806
rect 2424 7546 2452 8774
rect 2504 8288 2556 8294
rect 2504 8230 2556 8236
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2424 6934 2452 7482
rect 2516 7410 2544 8230
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2412 6928 2464 6934
rect 2412 6870 2464 6876
rect 2228 6724 2280 6730
rect 2228 6666 2280 6672
rect 2240 5370 2268 6666
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 2228 5364 2280 5370
rect 2228 5306 2280 5312
rect 2240 5030 2268 5306
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 2332 4826 2360 6598
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2424 5409 2452 5510
rect 2410 5400 2466 5409
rect 2516 5370 2544 6258
rect 2608 5710 2636 11494
rect 2884 11354 2912 12679
rect 2976 12442 3004 12786
rect 3516 12776 3568 12782
rect 3514 12744 3516 12753
rect 3568 12744 3570 12753
rect 3514 12679 3570 12688
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 2964 12436 3016 12442
rect 2964 12378 3016 12384
rect 3068 12288 3096 12582
rect 3174 12540 3482 12549
rect 3174 12538 3180 12540
rect 3236 12538 3260 12540
rect 3316 12538 3340 12540
rect 3396 12538 3420 12540
rect 3476 12538 3482 12540
rect 3236 12486 3238 12538
rect 3418 12486 3420 12538
rect 3174 12484 3180 12486
rect 3236 12484 3260 12486
rect 3316 12484 3340 12486
rect 3396 12484 3420 12486
rect 3476 12484 3482 12486
rect 3174 12475 3482 12484
rect 2976 12260 3096 12288
rect 2976 11642 3004 12260
rect 3146 12200 3202 12209
rect 3068 12144 3146 12152
rect 3068 12124 3148 12144
rect 3068 11830 3096 12124
rect 3200 12135 3202 12144
rect 3148 12106 3200 12112
rect 3332 12096 3384 12102
rect 3332 12038 3384 12044
rect 3344 11898 3372 12038
rect 3528 11898 3556 12582
rect 3332 11892 3384 11898
rect 3332 11834 3384 11840
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3056 11824 3108 11830
rect 3056 11766 3108 11772
rect 3424 11688 3476 11694
rect 2976 11614 3096 11642
rect 3620 11665 3648 13806
rect 3712 12345 3740 13874
rect 4080 13734 4108 13874
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 3790 13016 3846 13025
rect 3790 12951 3846 12960
rect 3804 12646 3832 12951
rect 3884 12708 3936 12714
rect 3884 12650 3936 12656
rect 3792 12640 3844 12646
rect 3792 12582 3844 12588
rect 3698 12336 3754 12345
rect 3698 12271 3754 12280
rect 3896 12170 3924 12650
rect 3884 12164 3936 12170
rect 3884 12106 3936 12112
rect 3606 11656 3662 11665
rect 3424 11630 3476 11636
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 2976 11150 3004 11494
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2780 11008 2832 11014
rect 2780 10950 2832 10956
rect 2792 10810 2820 10950
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 3068 10656 3096 11614
rect 3436 11558 3464 11630
rect 3528 11614 3606 11642
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3174 11452 3482 11461
rect 3174 11450 3180 11452
rect 3236 11450 3260 11452
rect 3316 11450 3340 11452
rect 3396 11450 3420 11452
rect 3476 11450 3482 11452
rect 3236 11398 3238 11450
rect 3418 11398 3420 11450
rect 3174 11396 3180 11398
rect 3236 11396 3260 11398
rect 3316 11396 3340 11398
rect 3396 11396 3420 11398
rect 3476 11396 3482 11398
rect 3174 11387 3482 11396
rect 3528 11150 3556 11614
rect 3988 11642 4016 13670
rect 4160 13456 4212 13462
rect 4160 13398 4212 13404
rect 4068 13320 4120 13326
rect 4066 13288 4068 13297
rect 4120 13288 4122 13297
rect 4066 13223 4122 13232
rect 4172 13190 4200 13398
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 4068 12776 4120 12782
rect 4068 12718 4120 12724
rect 4080 12306 4108 12718
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 4172 11830 4200 12582
rect 4160 11824 4212 11830
rect 4160 11766 4212 11772
rect 3606 11591 3662 11600
rect 3804 11614 4016 11642
rect 3700 11552 3752 11558
rect 3700 11494 3752 11500
rect 3608 11280 3660 11286
rect 3608 11222 3660 11228
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 3516 11144 3568 11150
rect 3516 11086 3568 11092
rect 3160 10674 3188 11086
rect 2884 10628 3096 10656
rect 3148 10668 3200 10674
rect 2688 10464 2740 10470
rect 2688 10406 2740 10412
rect 2700 9926 2728 10406
rect 2688 9920 2740 9926
rect 2688 9862 2740 9868
rect 2688 9648 2740 9654
rect 2686 9616 2688 9625
rect 2740 9616 2742 9625
rect 2686 9551 2742 9560
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2700 8090 2728 8298
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2792 7954 2820 9318
rect 2884 8673 2912 10628
rect 3148 10610 3200 10616
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3056 10532 3108 10538
rect 3056 10474 3108 10480
rect 3068 10198 3096 10474
rect 3174 10364 3482 10373
rect 3174 10362 3180 10364
rect 3236 10362 3260 10364
rect 3316 10362 3340 10364
rect 3396 10362 3420 10364
rect 3476 10362 3482 10364
rect 3236 10310 3238 10362
rect 3418 10310 3420 10362
rect 3174 10308 3180 10310
rect 3236 10308 3260 10310
rect 3316 10308 3340 10310
rect 3396 10308 3420 10310
rect 3476 10308 3482 10310
rect 3174 10299 3482 10308
rect 3528 10198 3556 10610
rect 3056 10192 3108 10198
rect 3056 10134 3108 10140
rect 3516 10192 3568 10198
rect 3516 10134 3568 10140
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 2976 8974 3004 9454
rect 3068 8974 3096 9998
rect 3252 9761 3280 9998
rect 3238 9752 3294 9761
rect 3238 9687 3294 9696
rect 3174 9276 3482 9285
rect 3174 9274 3180 9276
rect 3236 9274 3260 9276
rect 3316 9274 3340 9276
rect 3396 9274 3420 9276
rect 3476 9274 3482 9276
rect 3236 9222 3238 9274
rect 3418 9222 3420 9274
rect 3174 9220 3180 9222
rect 3236 9220 3260 9222
rect 3316 9220 3340 9222
rect 3396 9220 3420 9222
rect 3476 9220 3482 9222
rect 3174 9211 3482 9220
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3240 9036 3292 9042
rect 3240 8978 3292 8984
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 2870 8664 2926 8673
rect 2870 8599 2926 8608
rect 2964 8560 3016 8566
rect 2964 8502 3016 8508
rect 2976 8401 3004 8502
rect 3056 8424 3108 8430
rect 2962 8392 3018 8401
rect 3056 8366 3108 8372
rect 2962 8327 3018 8336
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 3068 7546 3096 8366
rect 3252 8362 3280 8978
rect 3436 8838 3464 9114
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3240 8356 3292 8362
rect 3240 8298 3292 8304
rect 3174 8188 3482 8197
rect 3174 8186 3180 8188
rect 3236 8186 3260 8188
rect 3316 8186 3340 8188
rect 3396 8186 3420 8188
rect 3476 8186 3482 8188
rect 3236 8134 3238 8186
rect 3418 8134 3420 8186
rect 3174 8132 3180 8134
rect 3236 8132 3260 8134
rect 3316 8132 3340 8134
rect 3396 8132 3420 8134
rect 3476 8132 3482 8134
rect 3174 8123 3482 8132
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2688 7268 2740 7274
rect 2688 7210 2740 7216
rect 2700 6866 2728 7210
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 2688 6248 2740 6254
rect 2688 6190 2740 6196
rect 2700 5914 2728 6190
rect 2688 5908 2740 5914
rect 2688 5850 2740 5856
rect 2596 5704 2648 5710
rect 2596 5646 2648 5652
rect 2792 5624 2820 7346
rect 3174 7100 3482 7109
rect 3174 7098 3180 7100
rect 3236 7098 3260 7100
rect 3316 7098 3340 7100
rect 3396 7098 3420 7100
rect 3476 7098 3482 7100
rect 3236 7046 3238 7098
rect 3418 7046 3420 7098
rect 3174 7044 3180 7046
rect 3236 7044 3260 7046
rect 3316 7044 3340 7046
rect 3396 7044 3420 7046
rect 3476 7044 3482 7046
rect 3174 7035 3482 7044
rect 3528 7002 3556 8434
rect 3516 6996 3568 7002
rect 3516 6938 3568 6944
rect 2872 6928 2924 6934
rect 2872 6870 2924 6876
rect 2884 5778 2912 6870
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3330 6624 3386 6633
rect 3068 6458 3096 6598
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 3160 6361 3188 6598
rect 3330 6559 3386 6568
rect 3146 6352 3202 6361
rect 3146 6287 3202 6296
rect 3344 6254 3372 6559
rect 3516 6384 3568 6390
rect 3516 6326 3568 6332
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 2964 6248 3016 6254
rect 2964 6190 3016 6196
rect 3332 6248 3384 6254
rect 3332 6190 3384 6196
rect 2872 5772 2924 5778
rect 2872 5714 2924 5720
rect 2872 5636 2924 5642
rect 2792 5596 2872 5624
rect 2872 5578 2924 5584
rect 2596 5568 2648 5574
rect 2596 5510 2648 5516
rect 2410 5335 2466 5344
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 2410 5264 2466 5273
rect 2410 5199 2412 5208
rect 2464 5199 2466 5208
rect 2412 5170 2464 5176
rect 2320 4820 2372 4826
rect 2320 4762 2372 4768
rect 2412 4752 2464 4758
rect 2412 4694 2464 4700
rect 2320 4616 2372 4622
rect 2318 4584 2320 4593
rect 2372 4584 2374 4593
rect 2318 4519 2374 4528
rect 2424 3534 2452 4694
rect 2504 4480 2556 4486
rect 2504 4422 2556 4428
rect 2516 3534 2544 4422
rect 2608 4298 2636 5510
rect 2688 5296 2740 5302
rect 2688 5238 2740 5244
rect 2700 4622 2728 5238
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2688 4616 2740 4622
rect 2688 4558 2740 4564
rect 2608 4270 2728 4298
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 2608 3738 2636 4082
rect 2700 4078 2728 4270
rect 2792 4128 2820 4762
rect 2884 4622 2912 5578
rect 2976 5250 3004 6190
rect 3436 6118 3464 6258
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3068 5370 3096 6054
rect 3174 6012 3482 6021
rect 3174 6010 3180 6012
rect 3236 6010 3260 6012
rect 3316 6010 3340 6012
rect 3396 6010 3420 6012
rect 3476 6010 3482 6012
rect 3236 5958 3238 6010
rect 3418 5958 3420 6010
rect 3174 5956 3180 5958
rect 3236 5956 3260 5958
rect 3316 5956 3340 5958
rect 3396 5956 3420 5958
rect 3476 5956 3482 5958
rect 3174 5947 3482 5956
rect 3238 5536 3294 5545
rect 3238 5471 3294 5480
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 2976 5222 3096 5250
rect 3252 5234 3280 5471
rect 3528 5370 3556 6326
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 3514 5264 3570 5273
rect 3068 5166 3096 5222
rect 3240 5228 3292 5234
rect 3514 5199 3570 5208
rect 3240 5170 3292 5176
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 3174 4924 3482 4933
rect 3174 4922 3180 4924
rect 3236 4922 3260 4924
rect 3316 4922 3340 4924
rect 3396 4922 3420 4924
rect 3476 4922 3482 4924
rect 3236 4870 3238 4922
rect 3418 4870 3420 4922
rect 3174 4868 3180 4870
rect 3236 4868 3260 4870
rect 3316 4868 3340 4870
rect 3396 4868 3420 4870
rect 3476 4868 3482 4870
rect 3174 4859 3482 4868
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3252 4214 3280 4422
rect 3240 4208 3292 4214
rect 3240 4150 3292 4156
rect 3528 4146 3556 5199
rect 2872 4140 2924 4146
rect 2792 4100 2872 4128
rect 2872 4082 2924 4088
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 2778 4040 2834 4049
rect 2884 4010 2912 4082
rect 2778 3975 2780 3984
rect 2832 3975 2834 3984
rect 2872 4004 2924 4010
rect 2780 3946 2832 3952
rect 2872 3946 2924 3952
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 2596 3732 2648 3738
rect 2596 3674 2648 3680
rect 2700 3602 2728 3878
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 2688 3596 2740 3602
rect 2688 3538 2740 3544
rect 2412 3528 2464 3534
rect 2412 3470 2464 3476
rect 2504 3528 2556 3534
rect 2504 3470 2556 3476
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 2688 3392 2740 3398
rect 2688 3334 2740 3340
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 2148 2650 2176 2994
rect 2136 2644 2188 2650
rect 2136 2586 2188 2592
rect 1858 2408 1914 2417
rect 1858 2343 1914 2352
rect 1860 2304 1912 2310
rect 1860 2246 1912 2252
rect 1872 800 1900 2246
rect 2240 921 2268 3334
rect 2412 3120 2464 3126
rect 2412 3062 2464 3068
rect 2424 2854 2452 3062
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 2608 2922 2636 2994
rect 2596 2916 2648 2922
rect 2596 2858 2648 2864
rect 2412 2848 2464 2854
rect 2412 2790 2464 2796
rect 2320 2304 2372 2310
rect 2320 2246 2372 2252
rect 2226 912 2282 921
rect 2226 847 2282 856
rect 2332 800 2360 2246
rect 2700 1601 2728 3334
rect 2792 2582 2820 3606
rect 2872 2848 2924 2854
rect 2872 2790 2924 2796
rect 2780 2576 2832 2582
rect 2780 2518 2832 2524
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 2686 1592 2742 1601
rect 2686 1527 2742 1536
rect 2792 800 2820 2246
rect 2884 1193 2912 2790
rect 2976 2514 3004 3878
rect 3174 3836 3482 3845
rect 3174 3834 3180 3836
rect 3236 3834 3260 3836
rect 3316 3834 3340 3836
rect 3396 3834 3420 3836
rect 3476 3834 3482 3836
rect 3236 3782 3238 3834
rect 3418 3782 3420 3834
rect 3174 3780 3180 3782
rect 3236 3780 3260 3782
rect 3316 3780 3340 3782
rect 3396 3780 3420 3782
rect 3476 3780 3482 3782
rect 3174 3771 3482 3780
rect 3516 3528 3568 3534
rect 3620 3516 3648 11222
rect 3712 11150 3740 11494
rect 3700 11144 3752 11150
rect 3700 11086 3752 11092
rect 3700 10804 3752 10810
rect 3700 10746 3752 10752
rect 3712 9722 3740 10746
rect 3700 9716 3752 9722
rect 3700 9658 3752 9664
rect 3700 8288 3752 8294
rect 3700 8230 3752 8236
rect 3712 8022 3740 8230
rect 3700 8016 3752 8022
rect 3700 7958 3752 7964
rect 3804 7954 3832 11614
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3988 11218 4016 11494
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 3976 11076 4028 11082
rect 3976 11018 4028 11024
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3792 7948 3844 7954
rect 3792 7890 3844 7896
rect 3792 7812 3844 7818
rect 3792 7754 3844 7760
rect 3700 6792 3752 6798
rect 3804 6769 3832 7754
rect 3700 6734 3752 6740
rect 3790 6760 3846 6769
rect 3712 6338 3740 6734
rect 3790 6695 3846 6704
rect 3896 6458 3924 9862
rect 3988 6746 4016 11018
rect 4160 10464 4212 10470
rect 4160 10406 4212 10412
rect 4172 10266 4200 10406
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 4264 8838 4292 14282
rect 4356 14074 4384 16510
rect 4802 16400 4858 17200
rect 5446 16400 5502 17200
rect 6090 16400 6146 17200
rect 6734 16400 6790 17200
rect 7378 16400 7434 17200
rect 8022 16400 8078 17200
rect 8666 16400 8722 17200
rect 9310 16400 9366 17200
rect 9954 16400 10010 17200
rect 10598 16400 10654 17200
rect 11242 16400 11298 17200
rect 11886 16538 11942 17200
rect 11886 16510 12020 16538
rect 11886 16400 11942 16510
rect 4712 15224 4764 15230
rect 4712 15166 4764 15172
rect 4528 14884 4580 14890
rect 4528 14826 4580 14832
rect 4436 14408 4488 14414
rect 4436 14350 4488 14356
rect 4344 14068 4396 14074
rect 4344 14010 4396 14016
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4356 11898 4384 12038
rect 4344 11892 4396 11898
rect 4344 11834 4396 11840
rect 4448 10690 4476 14350
rect 4540 13938 4568 14826
rect 4724 14414 4752 15166
rect 4712 14408 4764 14414
rect 4712 14350 4764 14356
rect 4724 14074 4752 14350
rect 4816 14074 4844 16400
rect 5460 14600 5488 16400
rect 5908 15020 5960 15026
rect 5908 14962 5960 14968
rect 5540 14612 5592 14618
rect 5460 14572 5540 14600
rect 5540 14554 5592 14560
rect 5920 14414 5948 14962
rect 6104 14618 6132 16400
rect 6748 14618 6776 16400
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 6092 14612 6144 14618
rect 6092 14554 6144 14560
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 6736 14612 6788 14618
rect 6736 14554 6788 14560
rect 6184 14476 6236 14482
rect 6184 14418 6236 14424
rect 4988 14408 5040 14414
rect 4988 14350 5040 14356
rect 5908 14408 5960 14414
rect 5908 14350 5960 14356
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 5000 12986 5028 14350
rect 5172 14340 5224 14346
rect 5172 14282 5224 14288
rect 5184 13938 5212 14282
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5398 14172 5706 14181
rect 5398 14170 5404 14172
rect 5460 14170 5484 14172
rect 5540 14170 5564 14172
rect 5620 14170 5644 14172
rect 5700 14170 5706 14172
rect 5460 14118 5462 14170
rect 5642 14118 5644 14170
rect 5398 14116 5404 14118
rect 5460 14116 5484 14118
rect 5540 14116 5564 14118
rect 5620 14116 5644 14118
rect 5700 14116 5706 14118
rect 5398 14107 5706 14116
rect 5538 13968 5594 13977
rect 5172 13932 5224 13938
rect 5828 13938 5856 14214
rect 5538 13903 5540 13912
rect 5172 13874 5224 13880
rect 5592 13903 5594 13912
rect 5816 13932 5868 13938
rect 5540 13874 5592 13880
rect 5816 13874 5868 13880
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 5460 13394 5488 13806
rect 6196 13802 6224 14418
rect 6564 14414 6592 14554
rect 6828 14544 6880 14550
rect 6828 14486 6880 14492
rect 6552 14408 6604 14414
rect 6552 14350 6604 14356
rect 6368 14272 6420 14278
rect 6420 14232 6500 14260
rect 6368 14214 6420 14220
rect 6472 14074 6500 14232
rect 6276 14068 6328 14074
rect 6276 14010 6328 14016
rect 6460 14068 6512 14074
rect 6460 14010 6512 14016
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6288 13920 6316 14010
rect 6552 13932 6604 13938
rect 6288 13892 6552 13920
rect 6552 13874 6604 13880
rect 6184 13796 6236 13802
rect 6184 13738 6236 13744
rect 6368 13796 6420 13802
rect 6368 13738 6420 13744
rect 5998 13696 6054 13705
rect 5998 13631 6054 13640
rect 6012 13394 6040 13631
rect 6276 13456 6328 13462
rect 6276 13398 6328 13404
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5724 13388 5776 13394
rect 5724 13330 5776 13336
rect 6000 13388 6052 13394
rect 6000 13330 6052 13336
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 5184 12986 5212 13126
rect 5398 13084 5706 13093
rect 5398 13082 5404 13084
rect 5460 13082 5484 13084
rect 5540 13082 5564 13084
rect 5620 13082 5644 13084
rect 5700 13082 5706 13084
rect 5460 13030 5462 13082
rect 5642 13030 5644 13082
rect 5398 13028 5404 13030
rect 5460 13028 5484 13030
rect 5540 13028 5564 13030
rect 5620 13028 5644 13030
rect 5700 13028 5706 13030
rect 5398 13019 5706 13028
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4528 11688 4580 11694
rect 4528 11630 4580 11636
rect 4540 11150 4568 11630
rect 4528 11144 4580 11150
rect 4528 11086 4580 11092
rect 4356 10662 4476 10690
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4080 7818 4108 8774
rect 4250 8392 4306 8401
rect 4250 8327 4306 8336
rect 4264 8294 4292 8327
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 4264 7970 4292 8230
rect 4356 8090 4384 10662
rect 4436 10600 4488 10606
rect 4436 10542 4488 10548
rect 4448 9330 4476 10542
rect 4540 9450 4568 11086
rect 4528 9444 4580 9450
rect 4528 9386 4580 9392
rect 4620 9376 4672 9382
rect 4448 9302 4568 9330
rect 4620 9318 4672 9324
rect 4540 8906 4568 9302
rect 4436 8900 4488 8906
rect 4436 8842 4488 8848
rect 4528 8900 4580 8906
rect 4528 8842 4580 8848
rect 4448 8430 4476 8842
rect 4436 8424 4488 8430
rect 4436 8366 4488 8372
rect 4344 8084 4396 8090
rect 4344 8026 4396 8032
rect 4264 7942 4384 7970
rect 4068 7812 4120 7818
rect 4068 7754 4120 7760
rect 3988 6718 4108 6746
rect 3976 6656 4028 6662
rect 4080 6633 4108 6718
rect 3976 6598 4028 6604
rect 4066 6624 4122 6633
rect 3988 6497 4016 6598
rect 4066 6559 4122 6568
rect 3974 6488 4030 6497
rect 3884 6452 3936 6458
rect 3974 6423 4030 6432
rect 3884 6394 3936 6400
rect 3712 6310 3832 6338
rect 3896 6322 3924 6394
rect 3700 6248 3752 6254
rect 3700 6190 3752 6196
rect 3712 5778 3740 6190
rect 3700 5772 3752 5778
rect 3700 5714 3752 5720
rect 3712 5166 3740 5714
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 3804 5098 3832 6310
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 3896 5370 3924 6258
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3988 5574 4016 6054
rect 4080 5846 4108 6559
rect 4158 6352 4214 6361
rect 4158 6287 4214 6296
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 3792 5092 3844 5098
rect 3792 5034 3844 5040
rect 3790 4720 3846 4729
rect 3790 4655 3846 4664
rect 3804 4554 3832 4655
rect 3792 4548 3844 4554
rect 3792 4490 3844 4496
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3896 4049 3924 4082
rect 3882 4040 3938 4049
rect 3882 3975 3938 3984
rect 3700 3936 3752 3942
rect 3988 3924 4016 5510
rect 4172 5302 4200 6287
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 4160 5296 4212 5302
rect 4160 5238 4212 5244
rect 4264 5234 4292 5646
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 4252 5228 4304 5234
rect 4252 5170 4304 5176
rect 4080 4486 4108 5170
rect 4252 4616 4304 4622
rect 4250 4584 4252 4593
rect 4356 4604 4384 7942
rect 4448 7886 4476 8366
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4448 7478 4476 7822
rect 4436 7472 4488 7478
rect 4436 7414 4488 7420
rect 4448 7342 4476 7414
rect 4436 7336 4488 7342
rect 4436 7278 4488 7284
rect 4448 6866 4476 7278
rect 4540 7206 4568 8842
rect 4632 8294 4660 9318
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 4436 6860 4488 6866
rect 4436 6802 4488 6808
rect 4448 5778 4476 6802
rect 4540 6186 4568 7142
rect 4528 6180 4580 6186
rect 4528 6122 4580 6128
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 4526 5672 4582 5681
rect 4526 5607 4582 5616
rect 4540 5234 4568 5607
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 4304 4584 4384 4604
rect 4306 4576 4384 4584
rect 4250 4519 4306 4528
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 4080 4185 4108 4422
rect 4066 4176 4122 4185
rect 4066 4111 4122 4120
rect 4724 4078 4752 12582
rect 5000 12434 5028 12922
rect 5356 12912 5408 12918
rect 5354 12880 5356 12889
rect 5408 12880 5410 12889
rect 5354 12815 5410 12824
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 5172 12708 5224 12714
rect 5172 12650 5224 12656
rect 5000 12406 5120 12434
rect 4988 12164 5040 12170
rect 4988 12106 5040 12112
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4908 11898 4936 12038
rect 4896 11892 4948 11898
rect 4896 11834 4948 11840
rect 4804 11348 4856 11354
rect 4804 11290 4856 11296
rect 4816 9994 4844 11290
rect 4804 9988 4856 9994
rect 4804 9930 4856 9936
rect 5000 9489 5028 12106
rect 4986 9480 5042 9489
rect 4986 9415 5042 9424
rect 5092 9382 5120 12406
rect 5184 10452 5212 12650
rect 5276 11626 5304 12718
rect 5398 11996 5706 12005
rect 5398 11994 5404 11996
rect 5460 11994 5484 11996
rect 5540 11994 5564 11996
rect 5620 11994 5644 11996
rect 5700 11994 5706 11996
rect 5460 11942 5462 11994
rect 5642 11942 5644 11994
rect 5398 11940 5404 11942
rect 5460 11940 5484 11942
rect 5540 11940 5564 11942
rect 5620 11940 5644 11942
rect 5700 11940 5706 11942
rect 5398 11931 5706 11940
rect 5736 11880 5764 13330
rect 5908 12368 5960 12374
rect 5908 12310 5960 12316
rect 5920 11898 5948 12310
rect 5644 11852 5764 11880
rect 5908 11892 5960 11898
rect 5264 11620 5316 11626
rect 5264 11562 5316 11568
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5460 11014 5488 11494
rect 5644 11098 5672 11852
rect 5908 11834 5960 11840
rect 5724 11756 5776 11762
rect 6012 11744 6040 13330
rect 6288 13190 6316 13398
rect 6276 13184 6328 13190
rect 6276 13126 6328 13132
rect 6288 12850 6316 13126
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 6092 12096 6144 12102
rect 6092 12038 6144 12044
rect 6104 11830 6132 12038
rect 6092 11824 6144 11830
rect 6092 11766 6144 11772
rect 5776 11716 6040 11744
rect 5724 11698 5776 11704
rect 6000 11144 6052 11150
rect 5644 11070 5764 11098
rect 6000 11086 6052 11092
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 5398 10908 5706 10917
rect 5398 10906 5404 10908
rect 5460 10906 5484 10908
rect 5540 10906 5564 10908
rect 5620 10906 5644 10908
rect 5700 10906 5706 10908
rect 5460 10854 5462 10906
rect 5642 10854 5644 10906
rect 5398 10852 5404 10854
rect 5460 10852 5484 10854
rect 5540 10852 5564 10854
rect 5620 10852 5644 10854
rect 5700 10852 5706 10854
rect 5398 10843 5706 10852
rect 5736 10742 5764 11070
rect 5724 10736 5776 10742
rect 5724 10678 5776 10684
rect 6012 10656 6040 11086
rect 6092 10668 6144 10674
rect 6012 10628 6092 10656
rect 5264 10464 5316 10470
rect 5184 10424 5264 10452
rect 5264 10406 5316 10412
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 5080 8560 5132 8566
rect 5080 8502 5132 8508
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4816 5710 4844 6054
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4816 4282 4844 5646
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 3752 3896 4016 3924
rect 3700 3878 3752 3884
rect 3712 3738 3740 3878
rect 3700 3732 3752 3738
rect 3700 3674 3752 3680
rect 3568 3488 3648 3516
rect 3516 3470 3568 3476
rect 3148 3392 3200 3398
rect 3068 3352 3148 3380
rect 2964 2508 3016 2514
rect 2964 2450 3016 2456
rect 3068 2446 3096 3352
rect 3148 3334 3200 3340
rect 3332 3392 3384 3398
rect 3332 3334 3384 3340
rect 3344 3058 3372 3334
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 3712 2961 3740 3674
rect 3790 3632 3846 3641
rect 3790 3567 3846 3576
rect 3804 3534 3832 3567
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 4068 3052 4120 3058
rect 4172 3040 4200 4014
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 4120 3012 4200 3040
rect 4068 2994 4120 3000
rect 3698 2952 3754 2961
rect 3698 2887 3754 2896
rect 4160 2916 4212 2922
rect 4160 2858 4212 2864
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 3976 2848 4028 2854
rect 3976 2790 4028 2796
rect 3174 2748 3482 2757
rect 3174 2746 3180 2748
rect 3236 2746 3260 2748
rect 3316 2746 3340 2748
rect 3396 2746 3420 2748
rect 3476 2746 3482 2748
rect 3236 2694 3238 2746
rect 3418 2694 3420 2746
rect 3174 2692 3180 2694
rect 3236 2692 3260 2694
rect 3316 2692 3340 2694
rect 3396 2692 3420 2694
rect 3476 2692 3482 2694
rect 3174 2683 3482 2692
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 2870 1184 2926 1193
rect 2870 1119 2926 1128
rect 3252 800 3280 2246
rect 3528 2009 3556 2790
rect 3700 2304 3752 2310
rect 3700 2246 3752 2252
rect 3514 2000 3570 2009
rect 3514 1935 3570 1944
rect 3712 800 3740 2246
rect 938 0 994 800
rect 1398 0 1454 800
rect 1858 0 1914 800
rect 2318 0 2374 800
rect 2778 0 2834 800
rect 3238 0 3294 800
rect 3698 0 3754 800
rect 3988 377 4016 2790
rect 4172 2446 4200 2858
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 4264 2378 4292 3334
rect 5000 3058 5028 7482
rect 5092 7002 5120 8502
rect 5276 8498 5304 10406
rect 6012 10062 6040 10628
rect 6092 10610 6144 10616
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 5908 9920 5960 9926
rect 5908 9862 5960 9868
rect 5398 9820 5706 9829
rect 5398 9818 5404 9820
rect 5460 9818 5484 9820
rect 5540 9818 5564 9820
rect 5620 9818 5644 9820
rect 5700 9818 5706 9820
rect 5460 9766 5462 9818
rect 5642 9766 5644 9818
rect 5398 9764 5404 9766
rect 5460 9764 5484 9766
rect 5540 9764 5564 9766
rect 5620 9764 5644 9766
rect 5700 9764 5706 9766
rect 5398 9755 5706 9764
rect 5724 8900 5776 8906
rect 5724 8842 5776 8848
rect 5398 8732 5706 8741
rect 5398 8730 5404 8732
rect 5460 8730 5484 8732
rect 5540 8730 5564 8732
rect 5620 8730 5644 8732
rect 5700 8730 5706 8732
rect 5460 8678 5462 8730
rect 5642 8678 5644 8730
rect 5398 8676 5404 8678
rect 5460 8676 5484 8678
rect 5540 8676 5564 8678
rect 5620 8676 5644 8678
rect 5700 8676 5706 8678
rect 5398 8667 5706 8676
rect 5736 8566 5764 8842
rect 5724 8560 5776 8566
rect 5724 8502 5776 8508
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 5398 7644 5706 7653
rect 5398 7642 5404 7644
rect 5460 7642 5484 7644
rect 5540 7642 5564 7644
rect 5620 7642 5644 7644
rect 5700 7642 5706 7644
rect 5460 7590 5462 7642
rect 5642 7590 5644 7642
rect 5398 7588 5404 7590
rect 5460 7588 5484 7590
rect 5540 7588 5564 7590
rect 5620 7588 5644 7590
rect 5700 7588 5706 7590
rect 5398 7579 5706 7588
rect 5828 7410 5856 8298
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 4988 3052 5040 3058
rect 4988 2994 5040 3000
rect 4988 2848 5040 2854
rect 4988 2790 5040 2796
rect 5000 2446 5028 2790
rect 5184 2650 5212 7346
rect 5398 6556 5706 6565
rect 5398 6554 5404 6556
rect 5460 6554 5484 6556
rect 5540 6554 5564 6556
rect 5620 6554 5644 6556
rect 5700 6554 5706 6556
rect 5460 6502 5462 6554
rect 5642 6502 5644 6554
rect 5398 6500 5404 6502
rect 5460 6500 5484 6502
rect 5540 6500 5564 6502
rect 5620 6500 5644 6502
rect 5700 6500 5706 6502
rect 5398 6491 5706 6500
rect 5828 6390 5856 7346
rect 5920 6390 5948 9862
rect 6012 9518 6040 9998
rect 6000 9512 6052 9518
rect 6000 9454 6052 9460
rect 6012 8974 6040 9454
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 6000 8560 6052 8566
rect 6000 8502 6052 8508
rect 6012 7750 6040 8502
rect 6104 8401 6132 9114
rect 6090 8392 6146 8401
rect 6090 8327 6146 8336
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 5816 6384 5868 6390
rect 5816 6326 5868 6332
rect 5908 6384 5960 6390
rect 5908 6326 5960 6332
rect 5632 6316 5684 6322
rect 5684 6276 5764 6304
rect 5632 6258 5684 6264
rect 5398 5468 5706 5477
rect 5398 5466 5404 5468
rect 5460 5466 5484 5468
rect 5540 5466 5564 5468
rect 5620 5466 5644 5468
rect 5700 5466 5706 5468
rect 5460 5414 5462 5466
rect 5642 5414 5644 5466
rect 5398 5412 5404 5414
rect 5460 5412 5484 5414
rect 5540 5412 5564 5414
rect 5620 5412 5644 5414
rect 5700 5412 5706 5414
rect 5398 5403 5706 5412
rect 5736 5370 5764 6276
rect 5816 5840 5868 5846
rect 5816 5782 5868 5788
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 5828 5234 5856 5782
rect 5920 5778 5948 6326
rect 6012 5817 6040 7686
rect 6104 6866 6132 8327
rect 6276 7880 6328 7886
rect 6196 7840 6276 7868
rect 6196 7410 6224 7840
rect 6276 7822 6328 7828
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 6092 6724 6144 6730
rect 6092 6666 6144 6672
rect 6104 5914 6132 6666
rect 6196 6322 6224 7346
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 5998 5808 6054 5817
rect 5908 5772 5960 5778
rect 5998 5743 6054 5752
rect 5908 5714 5960 5720
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5920 5098 5948 5714
rect 5908 5092 5960 5098
rect 5908 5034 5960 5040
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 5398 4380 5706 4389
rect 5398 4378 5404 4380
rect 5460 4378 5484 4380
rect 5540 4378 5564 4380
rect 5620 4378 5644 4380
rect 5700 4378 5706 4380
rect 5460 4326 5462 4378
rect 5642 4326 5644 4378
rect 5398 4324 5404 4326
rect 5460 4324 5484 4326
rect 5540 4324 5564 4326
rect 5620 4324 5644 4326
rect 5700 4324 5706 4326
rect 5398 4315 5706 4324
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5552 4078 5580 4218
rect 5828 4214 5856 4966
rect 6104 4690 6132 5850
rect 6092 4684 6144 4690
rect 6092 4626 6144 4632
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6104 4282 6132 4422
rect 6092 4276 6144 4282
rect 6092 4218 6144 4224
rect 5816 4208 5868 4214
rect 5816 4150 5868 4156
rect 6196 4078 6224 5850
rect 6274 5672 6330 5681
rect 6274 5607 6276 5616
rect 6328 5607 6330 5616
rect 6276 5578 6328 5584
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 5816 3392 5868 3398
rect 5816 3334 5868 3340
rect 5398 3292 5706 3301
rect 5398 3290 5404 3292
rect 5460 3290 5484 3292
rect 5540 3290 5564 3292
rect 5620 3290 5644 3292
rect 5700 3290 5706 3292
rect 5460 3238 5462 3290
rect 5642 3238 5644 3290
rect 5398 3236 5404 3238
rect 5460 3236 5484 3238
rect 5540 3236 5564 3238
rect 5620 3236 5644 3238
rect 5700 3236 5706 3238
rect 5398 3227 5706 3236
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 5552 2514 5580 2790
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 5080 2440 5132 2446
rect 5080 2382 5132 2388
rect 4252 2372 4304 2378
rect 4252 2314 4304 2320
rect 5092 2310 5120 2382
rect 5828 2378 5856 3334
rect 6380 2650 6408 13738
rect 6656 13326 6684 14010
rect 6734 13832 6790 13841
rect 6734 13767 6736 13776
rect 6788 13767 6790 13776
rect 6736 13738 6788 13744
rect 6840 13734 6868 14486
rect 7024 13938 7052 14758
rect 7392 14618 7420 16400
rect 7472 14952 7524 14958
rect 7472 14894 7524 14900
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7392 14414 7420 14554
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 7208 13326 7236 13466
rect 7484 13444 7512 14894
rect 7622 14716 7930 14725
rect 7622 14714 7628 14716
rect 7684 14714 7708 14716
rect 7764 14714 7788 14716
rect 7844 14714 7868 14716
rect 7924 14714 7930 14716
rect 7684 14662 7686 14714
rect 7866 14662 7868 14714
rect 7622 14660 7628 14662
rect 7684 14660 7708 14662
rect 7764 14660 7788 14662
rect 7844 14660 7868 14662
rect 7924 14660 7930 14662
rect 7622 14651 7930 14660
rect 7838 13968 7894 13977
rect 7838 13903 7894 13912
rect 7852 13802 7880 13903
rect 7840 13796 7892 13802
rect 7840 13738 7892 13744
rect 7622 13628 7930 13637
rect 7622 13626 7628 13628
rect 7684 13626 7708 13628
rect 7764 13626 7788 13628
rect 7844 13626 7868 13628
rect 7924 13626 7930 13628
rect 7684 13574 7686 13626
rect 7866 13574 7868 13626
rect 7622 13572 7628 13574
rect 7684 13572 7708 13574
rect 7764 13572 7788 13574
rect 7844 13572 7868 13574
rect 7924 13572 7930 13574
rect 7622 13563 7930 13572
rect 7484 13416 7604 13444
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 6920 13252 6972 13258
rect 6920 13194 6972 13200
rect 6932 12918 6960 13194
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 7208 12986 7236 13126
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 7012 12912 7064 12918
rect 7012 12854 7064 12860
rect 6736 12708 6788 12714
rect 6736 12650 6788 12656
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 6458 12064 6514 12073
rect 6458 11999 6514 12008
rect 6472 11830 6500 11999
rect 6460 11824 6512 11830
rect 6460 11766 6512 11772
rect 6472 4146 6500 11766
rect 6564 10198 6592 12242
rect 6656 11830 6684 12582
rect 6748 12084 6776 12650
rect 7024 12434 7052 12854
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 7196 12436 7248 12442
rect 7024 12406 7144 12434
rect 7116 12238 7144 12406
rect 7196 12378 7248 12384
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 7208 12186 7236 12378
rect 7392 12322 7420 12718
rect 7576 12628 7604 13416
rect 7748 13388 7800 13394
rect 7748 13330 7800 13336
rect 7760 12782 7788 13330
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7484 12600 7604 12628
rect 7484 12442 7512 12600
rect 7622 12540 7930 12549
rect 7622 12538 7628 12540
rect 7684 12538 7708 12540
rect 7764 12538 7788 12540
rect 7844 12538 7868 12540
rect 7924 12538 7930 12540
rect 7684 12486 7686 12538
rect 7866 12486 7868 12538
rect 7622 12484 7628 12486
rect 7684 12484 7708 12486
rect 7764 12484 7788 12486
rect 7844 12484 7868 12486
rect 7924 12484 7930 12486
rect 7622 12475 7930 12484
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 7392 12294 7512 12322
rect 7380 12232 7432 12238
rect 7012 12096 7064 12102
rect 6748 12056 7012 12084
rect 6644 11824 6696 11830
rect 6644 11766 6696 11772
rect 6552 10192 6604 10198
rect 6552 10134 6604 10140
rect 6564 9654 6592 10134
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6748 9586 6776 12056
rect 7012 12038 7064 12044
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 7024 11354 7052 11698
rect 7116 11626 7144 12174
rect 7208 12158 7328 12186
rect 7380 12174 7432 12180
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7104 11620 7156 11626
rect 7104 11562 7156 11568
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 7012 11212 7064 11218
rect 7012 11154 7064 11160
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6642 7304 6698 7313
rect 6642 7239 6698 7248
rect 6550 6216 6606 6225
rect 6550 6151 6606 6160
rect 6564 5710 6592 6151
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 6656 4622 6684 7239
rect 6932 7206 6960 7686
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6932 5914 6960 7142
rect 7024 6458 7052 11154
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 7116 5794 7144 11562
rect 7208 10742 7236 11630
rect 7300 11082 7328 12158
rect 7392 11762 7420 12174
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7196 10736 7248 10742
rect 7196 10678 7248 10684
rect 7392 9994 7420 11698
rect 7484 11150 7512 12294
rect 7932 12164 7984 12170
rect 7932 12106 7984 12112
rect 7944 11558 7972 12106
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 7622 11452 7930 11461
rect 7622 11450 7628 11452
rect 7684 11450 7708 11452
rect 7764 11450 7788 11452
rect 7844 11450 7868 11452
rect 7924 11450 7930 11452
rect 7684 11398 7686 11450
rect 7866 11398 7868 11450
rect 7622 11396 7628 11398
rect 7684 11396 7708 11398
rect 7764 11396 7788 11398
rect 7844 11396 7868 11398
rect 7924 11396 7930 11398
rect 7622 11387 7930 11396
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7622 10364 7930 10373
rect 7622 10362 7628 10364
rect 7684 10362 7708 10364
rect 7764 10362 7788 10364
rect 7844 10362 7868 10364
rect 7924 10362 7930 10364
rect 7684 10310 7686 10362
rect 7866 10310 7868 10362
rect 7622 10308 7628 10310
rect 7684 10308 7708 10310
rect 7764 10308 7788 10310
rect 7844 10308 7868 10310
rect 7924 10308 7930 10310
rect 7622 10299 7930 10308
rect 7196 9988 7248 9994
rect 7196 9930 7248 9936
rect 7380 9988 7432 9994
rect 7380 9930 7432 9936
rect 7208 9178 7236 9930
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7196 8900 7248 8906
rect 7196 8842 7248 8848
rect 7208 6644 7236 8842
rect 7300 6905 7328 9522
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7392 8974 7420 9454
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7286 6896 7342 6905
rect 7286 6831 7342 6840
rect 7288 6656 7340 6662
rect 7208 6616 7288 6644
rect 7288 6598 7340 6604
rect 6932 5766 7144 5794
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6748 4690 6776 4966
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6656 4282 6684 4558
rect 6644 4276 6696 4282
rect 6644 4218 6696 4224
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 6656 3505 6684 4218
rect 6840 4214 6868 4626
rect 6828 4208 6880 4214
rect 6828 4150 6880 4156
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6748 3534 6776 3878
rect 6736 3528 6788 3534
rect 6642 3496 6698 3505
rect 6736 3470 6788 3476
rect 6642 3431 6698 3440
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6748 3058 6776 3334
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6932 2990 6960 5766
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 7024 4282 7052 5102
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 6550 2680 6606 2689
rect 6368 2644 6420 2650
rect 6550 2615 6606 2624
rect 6368 2586 6420 2592
rect 6564 2446 6592 2615
rect 7024 2446 7052 3334
rect 7116 3058 7144 5510
rect 7300 5234 7328 6598
rect 7484 5386 7512 9862
rect 8036 9586 8064 16400
rect 8680 14618 8708 16400
rect 8760 14952 8812 14958
rect 8760 14894 8812 14900
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8680 14414 8708 14554
rect 8668 14408 8720 14414
rect 8668 14350 8720 14356
rect 8116 14272 8168 14278
rect 8116 14214 8168 14220
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8128 12434 8156 14214
rect 8300 13728 8352 13734
rect 8300 13670 8352 13676
rect 8128 12406 8248 12434
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 8128 11286 8156 12038
rect 8116 11280 8168 11286
rect 8116 11222 8168 11228
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8128 10742 8156 11086
rect 8116 10736 8168 10742
rect 8116 10678 8168 10684
rect 8128 10198 8156 10678
rect 8116 10192 8168 10198
rect 8116 10134 8168 10140
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 8128 9518 8156 9998
rect 8116 9512 8168 9518
rect 8116 9454 8168 9460
rect 7622 9276 7930 9285
rect 7622 9274 7628 9276
rect 7684 9274 7708 9276
rect 7764 9274 7788 9276
rect 7844 9274 7868 9276
rect 7924 9274 7930 9276
rect 7684 9222 7686 9274
rect 7866 9222 7868 9274
rect 7622 9220 7628 9222
rect 7684 9220 7708 9222
rect 7764 9220 7788 9222
rect 7844 9220 7868 9222
rect 7924 9220 7930 9222
rect 7622 9211 7930 9220
rect 7748 8900 7800 8906
rect 7748 8842 7800 8848
rect 7760 8498 7788 8842
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7622 8188 7930 8197
rect 7622 8186 7628 8188
rect 7684 8186 7708 8188
rect 7764 8186 7788 8188
rect 7844 8186 7868 8188
rect 7924 8186 7930 8188
rect 7684 8134 7686 8186
rect 7866 8134 7868 8186
rect 7622 8132 7628 8134
rect 7684 8132 7708 8134
rect 7764 8132 7788 8134
rect 7844 8132 7868 8134
rect 7924 8132 7930 8134
rect 7622 8123 7930 8132
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 7622 7100 7930 7109
rect 7622 7098 7628 7100
rect 7684 7098 7708 7100
rect 7764 7098 7788 7100
rect 7844 7098 7868 7100
rect 7924 7098 7930 7100
rect 7684 7046 7686 7098
rect 7866 7046 7868 7098
rect 7622 7044 7628 7046
rect 7684 7044 7708 7046
rect 7764 7044 7788 7046
rect 7844 7044 7868 7046
rect 7924 7044 7930 7046
rect 7622 7035 7930 7044
rect 8036 6118 8064 7414
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 7622 6012 7930 6021
rect 7622 6010 7628 6012
rect 7684 6010 7708 6012
rect 7764 6010 7788 6012
rect 7844 6010 7868 6012
rect 7924 6010 7930 6012
rect 7684 5958 7686 6010
rect 7866 5958 7868 6010
rect 7622 5956 7628 5958
rect 7684 5956 7708 5958
rect 7764 5956 7788 5958
rect 7844 5956 7868 5958
rect 7924 5956 7930 5958
rect 7622 5947 7930 5956
rect 7392 5358 7512 5386
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7196 5160 7248 5166
rect 7392 5114 7420 5358
rect 7472 5296 7524 5302
rect 7472 5238 7524 5244
rect 7196 5102 7248 5108
rect 7208 4826 7236 5102
rect 7300 5086 7420 5114
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 7300 2938 7328 5086
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7392 3602 7420 4966
rect 7484 4622 7512 5238
rect 7622 4924 7930 4933
rect 7622 4922 7628 4924
rect 7684 4922 7708 4924
rect 7764 4922 7788 4924
rect 7844 4922 7868 4924
rect 7924 4922 7930 4924
rect 7684 4870 7686 4922
rect 7866 4870 7868 4922
rect 7622 4868 7628 4870
rect 7684 4868 7708 4870
rect 7764 4868 7788 4870
rect 7844 4868 7868 4870
rect 7924 4868 7930 4870
rect 7622 4859 7930 4868
rect 8036 4826 8064 6054
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 7472 4616 7524 4622
rect 7470 4584 7472 4593
rect 7524 4584 7526 4593
rect 7470 4519 7526 4528
rect 7484 4078 7512 4519
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 7622 3836 7930 3845
rect 7622 3834 7628 3836
rect 7684 3834 7708 3836
rect 7764 3834 7788 3836
rect 7844 3834 7868 3836
rect 7924 3834 7930 3836
rect 7684 3782 7686 3834
rect 7866 3782 7868 3834
rect 7622 3780 7628 3782
rect 7684 3780 7708 3782
rect 7764 3780 7788 3782
rect 7844 3780 7868 3782
rect 7924 3780 7930 3782
rect 7622 3771 7930 3780
rect 8128 3670 8156 6394
rect 8220 5710 8248 12406
rect 8312 9926 8340 13670
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8404 11898 8432 13126
rect 8482 12336 8538 12345
rect 8482 12271 8538 12280
rect 8496 11898 8524 12271
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8392 11620 8444 11626
rect 8392 11562 8444 11568
rect 8404 10470 8432 11562
rect 8496 11150 8524 11834
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8496 10282 8524 11086
rect 8404 10254 8524 10282
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8312 7410 8340 7890
rect 8404 7449 8432 10254
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 8496 8294 8524 9522
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8390 7440 8446 7449
rect 8300 7404 8352 7410
rect 8390 7375 8446 7384
rect 8300 7346 8352 7352
rect 8312 6780 8340 7346
rect 8496 7342 8524 7686
rect 8484 7336 8536 7342
rect 8484 7278 8536 7284
rect 8392 6792 8444 6798
rect 8312 6752 8392 6780
rect 8392 6734 8444 6740
rect 8300 5840 8352 5846
rect 8300 5782 8352 5788
rect 8312 5710 8340 5782
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8220 5234 8248 5646
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 8312 4622 8340 5646
rect 8496 5030 8524 7278
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8312 4146 8340 4558
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8206 4040 8262 4049
rect 8206 3975 8262 3984
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 7380 3596 7432 3602
rect 7380 3538 7432 3544
rect 7840 3392 7892 3398
rect 7840 3334 7892 3340
rect 7852 3126 7880 3334
rect 7840 3120 7892 3126
rect 7840 3062 7892 3068
rect 8220 2990 8248 3975
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8496 3602 8524 3878
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8588 3466 8616 11290
rect 8680 3602 8708 14214
rect 8772 14074 8800 14894
rect 9324 14618 9352 16400
rect 9968 14618 9996 16400
rect 10612 14618 10640 16400
rect 11256 14618 11284 16400
rect 11336 14884 11388 14890
rect 11336 14826 11388 14832
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 10600 14612 10652 14618
rect 10600 14554 10652 14560
rect 11244 14612 11296 14618
rect 11244 14554 11296 14560
rect 9324 14414 9352 14554
rect 9968 14414 9996 14554
rect 10612 14414 10640 14554
rect 11060 14544 11112 14550
rect 11060 14486 11112 14492
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 10600 14408 10652 14414
rect 10600 14350 10652 14356
rect 9036 14272 9088 14278
rect 9036 14214 9088 14220
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 8760 14068 8812 14074
rect 8760 14010 8812 14016
rect 8772 13841 8800 14010
rect 8758 13832 8814 13841
rect 8758 13767 8814 13776
rect 8850 12336 8906 12345
rect 8850 12271 8906 12280
rect 8864 12073 8892 12271
rect 8850 12064 8906 12073
rect 8850 11999 8906 12008
rect 8852 11620 8904 11626
rect 8852 11562 8904 11568
rect 8864 11286 8892 11562
rect 8852 11280 8904 11286
rect 8852 11222 8904 11228
rect 8760 11076 8812 11082
rect 8760 11018 8812 11024
rect 8772 9178 8800 11018
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 8956 8974 8984 9318
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 8956 8634 8984 8910
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 8864 3942 8892 6054
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 8956 4214 8984 4966
rect 8944 4208 8996 4214
rect 8944 4150 8996 4156
rect 8852 3936 8904 3942
rect 8852 3878 8904 3884
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 8956 3534 8984 4150
rect 9048 4128 9076 14214
rect 9846 14172 10154 14181
rect 9846 14170 9852 14172
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 10148 14170 10154 14172
rect 9908 14118 9910 14170
rect 10090 14118 10092 14170
rect 9846 14116 9852 14118
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 10148 14116 10154 14118
rect 9846 14107 10154 14116
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 9140 12442 9168 12786
rect 9128 12436 9180 12442
rect 9128 12378 9180 12384
rect 9416 11694 9444 13330
rect 9508 12889 9536 13806
rect 9680 13796 9732 13802
rect 9680 13738 9732 13744
rect 9692 13190 9720 13738
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 9876 13433 9904 13670
rect 9862 13424 9918 13433
rect 9862 13359 9918 13368
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9846 13084 10154 13093
rect 9846 13082 9852 13084
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 10148 13082 10154 13084
rect 9908 13030 9910 13082
rect 10090 13030 10092 13082
rect 9846 13028 9852 13030
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 10148 13028 10154 13030
rect 9846 13019 10154 13028
rect 9494 12880 9550 12889
rect 9494 12815 9550 12824
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9140 11150 9168 11494
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9232 10810 9260 11154
rect 9220 10804 9272 10810
rect 9220 10746 9272 10752
rect 9232 8634 9260 10746
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 9220 7812 9272 7818
rect 9220 7754 9272 7760
rect 9232 7546 9260 7754
rect 9220 7540 9272 7546
rect 9220 7482 9272 7488
rect 9220 7268 9272 7274
rect 9220 7210 9272 7216
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 9140 5642 9168 6054
rect 9128 5636 9180 5642
rect 9128 5578 9180 5584
rect 9232 5030 9260 7210
rect 9404 5092 9456 5098
rect 9404 5034 9456 5040
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 9128 4140 9180 4146
rect 9048 4100 9128 4128
rect 9128 4082 9180 4088
rect 9416 3738 9444 5034
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 8576 3460 8628 3466
rect 8576 3402 8628 3408
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 9220 3392 9272 3398
rect 9220 3334 9272 3340
rect 8208 2984 8260 2990
rect 7300 2910 7420 2938
rect 8208 2926 8260 2932
rect 7392 2854 7420 2910
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 7288 2848 7340 2854
rect 7288 2790 7340 2796
rect 7380 2848 7432 2854
rect 7380 2790 7432 2796
rect 7116 2446 7144 2790
rect 7300 2514 7328 2790
rect 7622 2748 7930 2757
rect 7622 2746 7628 2748
rect 7684 2746 7708 2748
rect 7764 2746 7788 2748
rect 7844 2746 7868 2748
rect 7924 2746 7930 2748
rect 7684 2694 7686 2746
rect 7866 2694 7868 2746
rect 7622 2692 7628 2694
rect 7684 2692 7708 2694
rect 7764 2692 7788 2694
rect 7844 2692 7868 2694
rect 7924 2692 7930 2694
rect 7622 2683 7930 2692
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 8680 2446 8708 3334
rect 9232 2446 9260 3334
rect 9508 2990 9536 12815
rect 10232 12776 10284 12782
rect 10232 12718 10284 12724
rect 10244 12306 10272 12718
rect 10416 12368 10468 12374
rect 10416 12310 10468 12316
rect 10232 12300 10284 12306
rect 10232 12242 10284 12248
rect 9846 11996 10154 12005
rect 9846 11994 9852 11996
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 10148 11994 10154 11996
rect 9908 11942 9910 11994
rect 10090 11942 10092 11994
rect 9846 11940 9852 11942
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 10148 11940 10154 11942
rect 9846 11931 10154 11940
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9692 10962 9720 11834
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9784 11218 9812 11698
rect 10244 11694 10272 12242
rect 10048 11688 10100 11694
rect 10048 11630 10100 11636
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9876 11286 9904 11494
rect 9864 11280 9916 11286
rect 10060 11257 10088 11630
rect 9864 11222 9916 11228
rect 10046 11248 10102 11257
rect 9772 11212 9824 11218
rect 10046 11183 10102 11192
rect 9772 11154 9824 11160
rect 9784 11121 9812 11154
rect 9770 11112 9826 11121
rect 9770 11047 9826 11056
rect 9692 10934 9812 10962
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9692 10062 9720 10542
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9600 6730 9628 7142
rect 9588 6724 9640 6730
rect 9588 6666 9640 6672
rect 9784 6202 9812 10934
rect 9846 10908 10154 10917
rect 9846 10906 9852 10908
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 10148 10906 10154 10908
rect 9908 10854 9910 10906
rect 10090 10854 10092 10906
rect 9846 10852 9852 10854
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 10148 10852 10154 10854
rect 9846 10843 10154 10852
rect 10244 9994 10272 11630
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 10336 10742 10364 10950
rect 10324 10736 10376 10742
rect 10324 10678 10376 10684
rect 10232 9988 10284 9994
rect 10232 9930 10284 9936
rect 9846 9820 10154 9829
rect 9846 9818 9852 9820
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 10148 9818 10154 9820
rect 9908 9766 9910 9818
rect 10090 9766 10092 9818
rect 9846 9764 9852 9766
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 10148 9764 10154 9766
rect 9846 9755 10154 9764
rect 10244 9178 10272 9930
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 9846 8732 10154 8741
rect 9846 8730 9852 8732
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 10148 8730 10154 8732
rect 9908 8678 9910 8730
rect 10090 8678 10092 8730
rect 9846 8676 9852 8678
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 10148 8676 10154 8678
rect 9846 8667 10154 8676
rect 10324 8424 10376 8430
rect 10324 8366 10376 8372
rect 10336 7750 10364 8366
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 9846 7644 10154 7653
rect 9846 7642 9852 7644
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 10148 7642 10154 7644
rect 9908 7590 9910 7642
rect 10090 7590 10092 7642
rect 9846 7588 9852 7590
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 10148 7588 10154 7590
rect 9846 7579 10154 7588
rect 10232 6724 10284 6730
rect 10232 6666 10284 6672
rect 9846 6556 10154 6565
rect 9846 6554 9852 6556
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 10148 6554 10154 6556
rect 9908 6502 9910 6554
rect 10090 6502 10092 6554
rect 9846 6500 9852 6502
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 10148 6500 10154 6502
rect 9846 6491 10154 6500
rect 10244 6322 10272 6666
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 9784 6174 10272 6202
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9692 5234 9720 5510
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9692 4486 9720 5170
rect 9784 4690 9812 5714
rect 9846 5468 10154 5477
rect 9846 5466 9852 5468
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 10148 5466 10154 5468
rect 9908 5414 9910 5466
rect 10090 5414 10092 5466
rect 9846 5412 9852 5414
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 10148 5412 10154 5414
rect 9846 5403 10154 5412
rect 10046 4856 10102 4865
rect 10046 4791 10102 4800
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9600 4078 9628 4422
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9600 3534 9628 4014
rect 9784 3534 9812 4626
rect 10060 4622 10088 4791
rect 10138 4720 10194 4729
rect 10138 4655 10194 4664
rect 10048 4616 10100 4622
rect 10048 4558 10100 4564
rect 10152 4554 10180 4655
rect 10140 4548 10192 4554
rect 10140 4490 10192 4496
rect 9846 4380 10154 4389
rect 9846 4378 9852 4380
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 10148 4378 10154 4380
rect 9908 4326 9910 4378
rect 10090 4326 10092 4378
rect 9846 4324 9852 4326
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 10148 4324 10154 4326
rect 9846 4315 10154 4324
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 10060 3534 10088 3674
rect 10244 3641 10272 6174
rect 10336 5914 10364 7686
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10428 4978 10456 12310
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10612 10266 10640 10406
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10508 8288 10560 8294
rect 10508 8230 10560 8236
rect 10520 7478 10548 8230
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10508 7472 10560 7478
rect 10508 7414 10560 7420
rect 10612 7410 10640 7822
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10520 5914 10548 6190
rect 10508 5908 10560 5914
rect 10508 5850 10560 5856
rect 10336 4950 10456 4978
rect 10336 3942 10364 4950
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10324 3664 10376 3670
rect 10230 3632 10286 3641
rect 10324 3606 10376 3612
rect 10230 3567 10286 3576
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 9600 3194 9628 3470
rect 9680 3392 9732 3398
rect 9864 3392 9916 3398
rect 9680 3334 9732 3340
rect 9784 3352 9864 3380
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9692 3126 9720 3334
rect 9680 3120 9732 3126
rect 9680 3062 9732 3068
rect 9496 2984 9548 2990
rect 9496 2926 9548 2932
rect 9784 2446 9812 3352
rect 9864 3334 9916 3340
rect 10232 3392 10284 3398
rect 10232 3334 10284 3340
rect 9846 3292 10154 3301
rect 9846 3290 9852 3292
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 10148 3290 10154 3292
rect 9908 3238 9910 3290
rect 10090 3238 10092 3290
rect 9846 3236 9852 3238
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 10148 3236 10154 3238
rect 9846 3227 10154 3236
rect 10244 2446 10272 3334
rect 10336 3097 10364 3606
rect 10322 3088 10378 3097
rect 10322 3023 10378 3032
rect 10428 2774 10456 4762
rect 10704 4078 10732 14214
rect 10968 11892 11020 11898
rect 10968 11834 11020 11840
rect 10874 11248 10930 11257
rect 10874 11183 10930 11192
rect 10888 10538 10916 11183
rect 10980 11150 11008 11834
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10876 10532 10928 10538
rect 10876 10474 10928 10480
rect 11072 8378 11100 14486
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 11164 13297 11192 14010
rect 11348 14006 11376 14826
rect 11992 14414 12020 16510
rect 12530 16400 12586 17200
rect 13174 16400 13230 17200
rect 13818 16400 13874 17200
rect 14462 16538 14518 17200
rect 14200 16510 14518 16538
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12070 14716 12378 14725
rect 12070 14714 12076 14716
rect 12132 14714 12156 14716
rect 12212 14714 12236 14716
rect 12292 14714 12316 14716
rect 12372 14714 12378 14716
rect 12132 14662 12134 14714
rect 12314 14662 12316 14714
rect 12070 14660 12076 14662
rect 12132 14660 12156 14662
rect 12212 14660 12236 14662
rect 12292 14660 12316 14662
rect 12372 14660 12378 14662
rect 12070 14651 12378 14660
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 11428 14272 11480 14278
rect 11428 14214 11480 14220
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 11336 14000 11388 14006
rect 11336 13942 11388 13948
rect 11150 13288 11206 13297
rect 11150 13223 11206 13232
rect 11152 13184 11204 13190
rect 11336 13184 11388 13190
rect 11204 13144 11284 13172
rect 11152 13126 11204 13132
rect 11256 12238 11284 13144
rect 11336 13126 11388 13132
rect 11348 12986 11376 13126
rect 11336 12980 11388 12986
rect 11336 12922 11388 12928
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 11244 11144 11296 11150
rect 11242 11112 11244 11121
rect 11296 11112 11298 11121
rect 11242 11047 11298 11056
rect 11244 10464 11296 10470
rect 11348 10452 11376 12242
rect 11296 10424 11376 10452
rect 11244 10406 11296 10412
rect 11256 8566 11284 10406
rect 11244 8560 11296 8566
rect 11244 8502 11296 8508
rect 10784 8356 10836 8362
rect 11072 8350 11284 8378
rect 10784 8298 10836 8304
rect 10796 7886 10824 8298
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10888 6186 10916 6598
rect 10876 6180 10928 6186
rect 10876 6122 10928 6128
rect 10888 5914 10916 6122
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10876 5296 10928 5302
rect 10876 5238 10928 5244
rect 10888 4690 10916 5238
rect 10980 4826 11008 6598
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 10876 4480 10928 4486
rect 10876 4422 10928 4428
rect 10796 4214 10824 4422
rect 10784 4208 10836 4214
rect 10784 4150 10836 4156
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 10796 3534 10824 4150
rect 10888 4049 10916 4422
rect 10874 4040 10930 4049
rect 10874 3975 10930 3984
rect 11072 3602 11100 5510
rect 11164 5166 11192 5646
rect 11256 5234 11284 8350
rect 11336 6724 11388 6730
rect 11336 6666 11388 6672
rect 11348 6458 11376 6666
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11336 6180 11388 6186
rect 11336 6122 11388 6128
rect 11348 5778 11376 6122
rect 11336 5772 11388 5778
rect 11336 5714 11388 5720
rect 11336 5636 11388 5642
rect 11336 5578 11388 5584
rect 11244 5228 11296 5234
rect 11244 5170 11296 5176
rect 11152 5160 11204 5166
rect 11152 5102 11204 5108
rect 11060 3596 11112 3602
rect 11060 3538 11112 3544
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 11164 3482 11192 5102
rect 11348 3534 11376 5578
rect 11440 4690 11468 14214
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11532 10062 11560 11086
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 11624 10674 11652 10746
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11532 8430 11560 8910
rect 11520 8424 11572 8430
rect 11520 8366 11572 8372
rect 11532 7954 11560 8366
rect 11612 8084 11664 8090
rect 11612 8026 11664 8032
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11532 7342 11560 7890
rect 11624 7857 11652 8026
rect 11610 7848 11666 7857
rect 11610 7783 11666 7792
rect 11520 7336 11572 7342
rect 11520 7278 11572 7284
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 11532 6254 11560 6598
rect 11624 6390 11652 7142
rect 11612 6384 11664 6390
rect 11612 6326 11664 6332
rect 11520 6248 11572 6254
rect 11520 6190 11572 6196
rect 11716 5778 11744 14010
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 11428 4684 11480 4690
rect 11428 4626 11480 4632
rect 11808 4146 11836 14214
rect 12452 14074 12480 14758
rect 12544 14618 12572 16400
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12544 14414 12572 14554
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12636 14006 12664 14758
rect 13188 14618 13216 16400
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 12900 14476 12952 14482
rect 12900 14418 12952 14424
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12624 14000 12676 14006
rect 12624 13942 12676 13948
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 11900 13705 11928 13806
rect 11886 13696 11942 13705
rect 11886 13631 11942 13640
rect 11900 13190 11928 13631
rect 12070 13628 12378 13637
rect 12070 13626 12076 13628
rect 12132 13626 12156 13628
rect 12212 13626 12236 13628
rect 12292 13626 12316 13628
rect 12372 13626 12378 13628
rect 12132 13574 12134 13626
rect 12314 13574 12316 13626
rect 12070 13572 12076 13574
rect 12132 13572 12156 13574
rect 12212 13572 12236 13574
rect 12292 13572 12316 13574
rect 12372 13572 12378 13574
rect 12070 13563 12378 13572
rect 12348 13524 12400 13530
rect 12348 13466 12400 13472
rect 12360 13410 12388 13466
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 12176 13382 12388 13410
rect 12440 13388 12492 13394
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11992 12288 12020 13330
rect 12176 12782 12204 13382
rect 12440 13330 12492 13336
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 12360 12850 12388 13262
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12452 12782 12480 13330
rect 12624 13184 12676 13190
rect 12624 13126 12676 13132
rect 12636 12986 12664 13126
rect 12624 12980 12676 12986
rect 12624 12922 12676 12928
rect 12164 12776 12216 12782
rect 12164 12718 12216 12724
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12070 12540 12378 12549
rect 12070 12538 12076 12540
rect 12132 12538 12156 12540
rect 12212 12538 12236 12540
rect 12292 12538 12316 12540
rect 12372 12538 12378 12540
rect 12132 12486 12134 12538
rect 12314 12486 12316 12538
rect 12070 12484 12076 12486
rect 12132 12484 12156 12486
rect 12212 12484 12236 12486
rect 12292 12484 12316 12486
rect 12372 12484 12378 12486
rect 12070 12475 12378 12484
rect 12452 12306 12480 12582
rect 12728 12434 12756 14214
rect 12912 13938 12940 14418
rect 13188 14414 13216 14554
rect 13266 14512 13322 14521
rect 13266 14447 13322 14456
rect 13176 14408 13228 14414
rect 13176 14350 13228 14356
rect 13280 14074 13308 14447
rect 13360 14340 13412 14346
rect 13360 14282 13412 14288
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 12900 13932 12952 13938
rect 12900 13874 12952 13880
rect 13372 13734 13400 14282
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 13004 12442 13032 12786
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 13176 12708 13228 12714
rect 13176 12650 13228 12656
rect 12544 12406 12756 12434
rect 12808 12436 12860 12442
rect 12348 12300 12400 12306
rect 11992 12260 12348 12288
rect 11992 10810 12020 12260
rect 12348 12242 12400 12248
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 12070 11452 12378 11461
rect 12070 11450 12076 11452
rect 12132 11450 12156 11452
rect 12212 11450 12236 11452
rect 12292 11450 12316 11452
rect 12372 11450 12378 11452
rect 12132 11398 12134 11450
rect 12314 11398 12316 11450
rect 12070 11396 12076 11398
rect 12132 11396 12156 11398
rect 12212 11396 12236 11398
rect 12292 11396 12316 11398
rect 12372 11396 12378 11398
rect 12070 11387 12378 11396
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 12070 10364 12378 10373
rect 12070 10362 12076 10364
rect 12132 10362 12156 10364
rect 12212 10362 12236 10364
rect 12292 10362 12316 10364
rect 12372 10362 12378 10364
rect 12132 10310 12134 10362
rect 12314 10310 12316 10362
rect 12070 10308 12076 10310
rect 12132 10308 12156 10310
rect 12212 10308 12236 10310
rect 12292 10308 12316 10310
rect 12372 10308 12378 10310
rect 12070 10299 12378 10308
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11900 7410 11928 9318
rect 11992 8974 12020 9998
rect 12070 9276 12378 9285
rect 12070 9274 12076 9276
rect 12132 9274 12156 9276
rect 12212 9274 12236 9276
rect 12292 9274 12316 9276
rect 12372 9274 12378 9276
rect 12132 9222 12134 9274
rect 12314 9222 12316 9274
rect 12070 9220 12076 9222
rect 12132 9220 12156 9222
rect 12212 9220 12236 9222
rect 12292 9220 12316 9222
rect 12372 9220 12378 9222
rect 12070 9211 12378 9220
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 12070 8188 12378 8197
rect 12070 8186 12076 8188
rect 12132 8186 12156 8188
rect 12212 8186 12236 8188
rect 12292 8186 12316 8188
rect 12372 8186 12378 8188
rect 12132 8134 12134 8186
rect 12314 8134 12316 8186
rect 12070 8132 12076 8134
rect 12132 8132 12156 8134
rect 12212 8132 12236 8134
rect 12292 8132 12316 8134
rect 12372 8132 12378 8134
rect 12070 8123 12378 8132
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 12084 7478 12112 7686
rect 12072 7472 12124 7478
rect 12072 7414 12124 7420
rect 11888 7404 11940 7410
rect 11888 7346 11940 7352
rect 11980 7336 12032 7342
rect 11980 7278 12032 7284
rect 11992 7002 12020 7278
rect 12360 7188 12388 8026
rect 12360 7160 12480 7188
rect 12070 7100 12378 7109
rect 12070 7098 12076 7100
rect 12132 7098 12156 7100
rect 12212 7098 12236 7100
rect 12292 7098 12316 7100
rect 12372 7098 12378 7100
rect 12132 7046 12134 7098
rect 12314 7046 12316 7098
rect 12070 7044 12076 7046
rect 12132 7044 12156 7046
rect 12212 7044 12236 7046
rect 12292 7044 12316 7046
rect 12372 7044 12378 7046
rect 12070 7035 12378 7044
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 12452 6914 12480 7160
rect 12360 6886 12480 6914
rect 12360 6390 12388 6886
rect 12348 6384 12400 6390
rect 12348 6326 12400 6332
rect 12360 6202 12388 6326
rect 12360 6174 12480 6202
rect 12070 6012 12378 6021
rect 12070 6010 12076 6012
rect 12132 6010 12156 6012
rect 12212 6010 12236 6012
rect 12292 6010 12316 6012
rect 12372 6010 12378 6012
rect 12132 5958 12134 6010
rect 12314 5958 12316 6010
rect 12070 5956 12076 5958
rect 12132 5956 12156 5958
rect 12212 5956 12236 5958
rect 12292 5956 12316 5958
rect 12372 5956 12378 5958
rect 12070 5947 12378 5956
rect 12452 5778 12480 6174
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12164 5636 12216 5642
rect 12164 5578 12216 5584
rect 12176 5302 12204 5578
rect 12164 5296 12216 5302
rect 12164 5238 12216 5244
rect 12164 5160 12216 5166
rect 12162 5128 12164 5137
rect 12216 5128 12218 5137
rect 12162 5063 12218 5072
rect 12070 4924 12378 4933
rect 12070 4922 12076 4924
rect 12132 4922 12156 4924
rect 12212 4922 12236 4924
rect 12292 4922 12316 4924
rect 12372 4922 12378 4924
rect 12132 4870 12134 4922
rect 12314 4870 12316 4922
rect 12070 4868 12076 4870
rect 12132 4868 12156 4870
rect 12212 4868 12236 4870
rect 12292 4868 12316 4870
rect 12372 4868 12378 4870
rect 11886 4856 11942 4865
rect 12070 4859 12378 4868
rect 11886 4791 11942 4800
rect 11900 4758 11928 4791
rect 11888 4752 11940 4758
rect 11888 4694 11940 4700
rect 12544 4690 12572 12406
rect 12808 12378 12860 12384
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 12714 12336 12770 12345
rect 12714 12271 12770 12280
rect 12728 11762 12756 12271
rect 12820 12170 12848 12378
rect 12808 12164 12860 12170
rect 12808 12106 12860 12112
rect 13188 12102 13216 12650
rect 13372 12306 13400 12718
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 12624 11688 12676 11694
rect 13188 11665 13216 12038
rect 13280 11898 13308 12038
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13266 11792 13322 11801
rect 13266 11727 13268 11736
rect 13320 11727 13322 11736
rect 13268 11698 13320 11704
rect 12624 11630 12676 11636
rect 13174 11656 13230 11665
rect 12636 10674 12664 11630
rect 13084 11620 13136 11626
rect 13174 11591 13230 11600
rect 13084 11562 13136 11568
rect 13096 11014 13124 11562
rect 13188 11558 13216 11591
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 13084 11008 13136 11014
rect 13084 10950 13136 10956
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12636 9178 12664 10610
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12912 10062 12940 10542
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 13096 9994 13124 10950
rect 13372 10742 13400 12242
rect 13360 10736 13412 10742
rect 13360 10678 13412 10684
rect 13084 9988 13136 9994
rect 13084 9930 13136 9936
rect 13268 9512 13320 9518
rect 13268 9454 13320 9460
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 13280 8974 13308 9454
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 12808 8900 12860 8906
rect 12808 8842 12860 8848
rect 12992 8900 13044 8906
rect 12992 8842 13044 8848
rect 13452 8900 13504 8906
rect 13452 8842 13504 8848
rect 12714 4856 12770 4865
rect 12714 4791 12716 4800
rect 12768 4791 12770 4800
rect 12716 4762 12768 4768
rect 12820 4690 12848 8842
rect 13004 8498 13032 8842
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 13268 7812 13320 7818
rect 13268 7754 13320 7760
rect 13084 7472 13136 7478
rect 13084 7414 13136 7420
rect 12900 6724 12952 6730
rect 12900 6666 12952 6672
rect 12992 6724 13044 6730
rect 12992 6666 13044 6672
rect 12912 5166 12940 6666
rect 13004 5914 13032 6666
rect 13096 6202 13124 7414
rect 13280 6458 13308 7754
rect 13464 7750 13492 8842
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13268 6452 13320 6458
rect 13268 6394 13320 6400
rect 13464 6254 13492 7686
rect 13452 6248 13504 6254
rect 13096 6174 13216 6202
rect 13452 6190 13504 6196
rect 13084 6112 13136 6118
rect 13084 6054 13136 6060
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 12900 5160 12952 5166
rect 12900 5102 12952 5108
rect 12532 4684 12584 4690
rect 12532 4626 12584 4632
rect 12808 4684 12860 4690
rect 12808 4626 12860 4632
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 12624 4072 12676 4078
rect 13096 4026 13124 6054
rect 13188 5914 13216 6174
rect 13176 5908 13228 5914
rect 13176 5850 13228 5856
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 12624 4014 12676 4020
rect 12070 3836 12378 3845
rect 12070 3834 12076 3836
rect 12132 3834 12156 3836
rect 12212 3834 12236 3836
rect 12292 3834 12316 3836
rect 12372 3834 12378 3836
rect 12132 3782 12134 3834
rect 12314 3782 12316 3834
rect 12070 3780 12076 3782
rect 12132 3780 12156 3782
rect 12212 3780 12236 3782
rect 12292 3780 12316 3782
rect 12372 3780 12378 3782
rect 12070 3771 12378 3780
rect 12636 3738 12664 4014
rect 12912 3998 13124 4026
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 12532 3664 12584 3670
rect 12532 3606 12584 3612
rect 11336 3528 11388 3534
rect 11164 3454 11284 3482
rect 11336 3470 11388 3476
rect 11702 3496 11758 3505
rect 10692 3392 10744 3398
rect 10692 3334 10744 3340
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 10336 2746 10456 2774
rect 10336 2582 10364 2746
rect 10324 2576 10376 2582
rect 10324 2518 10376 2524
rect 10704 2446 10732 3334
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10888 2854 10916 3130
rect 10876 2848 10928 2854
rect 10876 2790 10928 2796
rect 10980 2650 11008 3334
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 6000 2440 6052 2446
rect 6000 2382 6052 2388
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 11072 2428 11100 2790
rect 11164 2582 11192 3334
rect 11256 2774 11284 3454
rect 11520 3460 11572 3466
rect 11702 3431 11758 3440
rect 11520 3402 11572 3408
rect 11428 2984 11480 2990
rect 11428 2926 11480 2932
rect 11256 2746 11376 2774
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 11244 2440 11296 2446
rect 11072 2400 11244 2428
rect 5816 2372 5868 2378
rect 5816 2314 5868 2320
rect 4160 2304 4212 2310
rect 4160 2246 4212 2252
rect 4620 2304 4672 2310
rect 4620 2246 4672 2252
rect 5080 2304 5132 2310
rect 5080 2246 5132 2252
rect 5724 2304 5776 2310
rect 5724 2246 5776 2252
rect 4172 800 4200 2246
rect 4632 800 4660 2246
rect 5092 800 5120 2246
rect 5398 2204 5706 2213
rect 5398 2202 5404 2204
rect 5460 2202 5484 2204
rect 5540 2202 5564 2204
rect 5620 2202 5644 2204
rect 5700 2202 5706 2204
rect 5460 2150 5462 2202
rect 5642 2150 5644 2202
rect 5398 2148 5404 2150
rect 5460 2148 5484 2150
rect 5540 2148 5564 2150
rect 5620 2148 5644 2150
rect 5700 2148 5706 2150
rect 5398 2139 5706 2148
rect 5736 1170 5764 2246
rect 5552 1142 5764 1170
rect 5552 800 5580 1142
rect 6012 800 6040 2382
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 7380 2304 7432 2310
rect 7380 2246 7432 2252
rect 7840 2304 7892 2310
rect 7840 2246 7892 2252
rect 8300 2304 8352 2310
rect 8300 2246 8352 2252
rect 8760 2304 8812 2310
rect 8760 2246 8812 2252
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 10232 2304 10284 2310
rect 10232 2246 10284 2252
rect 10600 2304 10652 2310
rect 10600 2246 10652 2252
rect 6472 800 6500 2246
rect 6932 800 6960 2246
rect 7392 800 7420 2246
rect 7852 800 7880 2246
rect 8312 800 8340 2246
rect 8772 800 8800 2246
rect 9232 800 9260 2246
rect 9692 800 9720 2246
rect 9846 2204 10154 2213
rect 9846 2202 9852 2204
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 10148 2202 10154 2204
rect 9908 2150 9910 2202
rect 10090 2150 10092 2202
rect 9846 2148 9852 2150
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 10148 2148 10154 2150
rect 9846 2139 10154 2148
rect 10244 1170 10272 2246
rect 10152 1142 10272 1170
rect 10152 800 10180 1142
rect 10612 800 10640 2246
rect 11072 800 11100 2400
rect 11244 2382 11296 2388
rect 11348 2378 11376 2746
rect 11440 2582 11468 2926
rect 11428 2576 11480 2582
rect 11428 2518 11480 2524
rect 11336 2372 11388 2378
rect 11336 2314 11388 2320
rect 11532 800 11560 3402
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11624 3058 11652 3334
rect 11716 3194 11744 3431
rect 12440 3392 12492 3398
rect 12440 3334 12492 3340
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 12070 2748 12378 2757
rect 12070 2746 12076 2748
rect 12132 2746 12156 2748
rect 12212 2746 12236 2748
rect 12292 2746 12316 2748
rect 12372 2746 12378 2748
rect 12132 2694 12134 2746
rect 12314 2694 12316 2746
rect 12070 2692 12076 2694
rect 12132 2692 12156 2694
rect 12212 2692 12236 2694
rect 12292 2692 12316 2694
rect 12372 2692 12378 2694
rect 12070 2683 12378 2692
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 11992 2378 12020 2586
rect 11980 2372 12032 2378
rect 11980 2314 12032 2320
rect 12256 2372 12308 2378
rect 12256 2314 12308 2320
rect 11992 870 12112 898
rect 11992 800 12020 870
rect 3974 368 4030 377
rect 3974 303 4030 312
rect 4158 0 4214 800
rect 4618 0 4674 800
rect 5078 0 5134 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 6918 0 6974 800
rect 7378 0 7434 800
rect 7838 0 7894 800
rect 8298 0 8354 800
rect 8758 0 8814 800
rect 9218 0 9274 800
rect 9678 0 9734 800
rect 10138 0 10194 800
rect 10598 0 10654 800
rect 11058 0 11114 800
rect 11518 0 11574 800
rect 11978 0 12034 800
rect 12084 762 12112 870
rect 12268 762 12296 2314
rect 12452 800 12480 3334
rect 12544 2514 12572 3606
rect 12636 3466 12664 3674
rect 12820 3534 12848 3878
rect 12808 3528 12860 3534
rect 12808 3470 12860 3476
rect 12624 3460 12676 3466
rect 12624 3402 12676 3408
rect 12912 3346 12940 3998
rect 13084 3936 13136 3942
rect 13084 3878 13136 3884
rect 12820 3318 12940 3346
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 12820 2922 12848 3318
rect 12900 3188 12952 3194
rect 12900 3130 12952 3136
rect 12808 2916 12860 2922
rect 12808 2858 12860 2864
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 12912 800 12940 3130
rect 13004 2922 13032 3334
rect 12992 2916 13044 2922
rect 12992 2858 13044 2864
rect 13096 2394 13124 3878
rect 13188 3738 13216 4014
rect 13280 3942 13308 4082
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 13176 2984 13228 2990
rect 13176 2926 13228 2932
rect 13004 2378 13124 2394
rect 12992 2372 13124 2378
rect 13044 2366 13124 2372
rect 12992 2314 13044 2320
rect 13188 2310 13216 2926
rect 13280 2530 13308 3878
rect 13372 3534 13400 4558
rect 13452 4004 13504 4010
rect 13452 3946 13504 3952
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13464 3058 13492 3946
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 13360 2984 13412 2990
rect 13360 2926 13412 2932
rect 13372 2650 13400 2926
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 13280 2502 13400 2530
rect 13556 2514 13584 14758
rect 13832 14414 13860 16400
rect 14200 14482 14228 16510
rect 14462 16400 14518 16510
rect 15106 16400 15162 17200
rect 15474 16552 15530 16561
rect 15474 16487 15530 16496
rect 14924 15020 14976 15026
rect 14924 14962 14976 14968
rect 14188 14476 14240 14482
rect 14188 14418 14240 14424
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13636 11892 13688 11898
rect 13636 11834 13688 11840
rect 13648 11082 13676 11834
rect 13636 11076 13688 11082
rect 13636 11018 13688 11024
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13648 7274 13676 7346
rect 13636 7268 13688 7274
rect 13636 7210 13688 7216
rect 13740 4690 13768 14214
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13832 13190 13860 13466
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 14094 11520 14150 11529
rect 14094 11455 14150 11464
rect 14108 9450 14136 11455
rect 14096 9444 14148 9450
rect 14096 9386 14148 9392
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13832 5370 13860 6054
rect 13924 5794 13952 8910
rect 14200 7834 14228 14418
rect 14294 14172 14602 14181
rect 14294 14170 14300 14172
rect 14356 14170 14380 14172
rect 14436 14170 14460 14172
rect 14516 14170 14540 14172
rect 14596 14170 14602 14172
rect 14356 14118 14358 14170
rect 14538 14118 14540 14170
rect 14294 14116 14300 14118
rect 14356 14116 14380 14118
rect 14436 14116 14460 14118
rect 14516 14116 14540 14118
rect 14596 14116 14602 14118
rect 14294 14107 14602 14116
rect 14936 14074 14964 14962
rect 14924 14068 14976 14074
rect 14924 14010 14976 14016
rect 15120 13954 15148 16400
rect 15292 14544 15344 14550
rect 15292 14486 15344 14492
rect 15028 13938 15148 13954
rect 15016 13932 15148 13938
rect 15068 13926 15148 13932
rect 15016 13874 15068 13880
rect 14294 13084 14602 13093
rect 14294 13082 14300 13084
rect 14356 13082 14380 13084
rect 14436 13082 14460 13084
rect 14516 13082 14540 13084
rect 14596 13082 14602 13084
rect 14356 13030 14358 13082
rect 14538 13030 14540 13082
rect 14294 13028 14300 13030
rect 14356 13028 14380 13030
rect 14436 13028 14460 13030
rect 14516 13028 14540 13030
rect 14596 13028 14602 13030
rect 14294 13019 14602 13028
rect 14464 12776 14516 12782
rect 14464 12718 14516 12724
rect 14476 12434 14504 12718
rect 15120 12434 15148 13926
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 15212 12850 15240 13126
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 14476 12406 14688 12434
rect 14660 12306 14688 12406
rect 14844 12406 15148 12434
rect 14648 12300 14700 12306
rect 14648 12242 14700 12248
rect 14294 11996 14602 12005
rect 14294 11994 14300 11996
rect 14356 11994 14380 11996
rect 14436 11994 14460 11996
rect 14516 11994 14540 11996
rect 14596 11994 14602 11996
rect 14356 11942 14358 11994
rect 14538 11942 14540 11994
rect 14294 11940 14300 11942
rect 14356 11940 14380 11942
rect 14436 11940 14460 11942
rect 14516 11940 14540 11942
rect 14596 11940 14602 11942
rect 14294 11931 14602 11940
rect 14556 11756 14608 11762
rect 14556 11698 14608 11704
rect 14568 11558 14596 11698
rect 14660 11694 14688 12242
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14556 11552 14608 11558
rect 14554 11520 14556 11529
rect 14608 11520 14610 11529
rect 14554 11455 14610 11464
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 14648 11076 14700 11082
rect 14648 11018 14700 11024
rect 14294 10908 14602 10917
rect 14294 10906 14300 10908
rect 14356 10906 14380 10908
rect 14436 10906 14460 10908
rect 14516 10906 14540 10908
rect 14596 10906 14602 10908
rect 14356 10854 14358 10906
rect 14538 10854 14540 10906
rect 14294 10852 14300 10854
rect 14356 10852 14380 10854
rect 14436 10852 14460 10854
rect 14516 10852 14540 10854
rect 14596 10852 14602 10854
rect 14294 10843 14602 10852
rect 14660 10810 14688 11018
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 14462 10704 14518 10713
rect 14462 10639 14464 10648
rect 14516 10639 14518 10648
rect 14464 10610 14516 10616
rect 14752 10266 14780 11154
rect 14740 10260 14792 10266
rect 14740 10202 14792 10208
rect 14294 9820 14602 9829
rect 14294 9818 14300 9820
rect 14356 9818 14380 9820
rect 14436 9818 14460 9820
rect 14516 9818 14540 9820
rect 14596 9818 14602 9820
rect 14356 9766 14358 9818
rect 14538 9766 14540 9818
rect 14294 9764 14300 9766
rect 14356 9764 14380 9766
rect 14436 9764 14460 9766
rect 14516 9764 14540 9766
rect 14596 9764 14602 9766
rect 14294 9755 14602 9764
rect 14740 9172 14792 9178
rect 14740 9114 14792 9120
rect 14752 8974 14780 9114
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14294 8732 14602 8741
rect 14294 8730 14300 8732
rect 14356 8730 14380 8732
rect 14436 8730 14460 8732
rect 14516 8730 14540 8732
rect 14596 8730 14602 8732
rect 14356 8678 14358 8730
rect 14538 8678 14540 8730
rect 14294 8676 14300 8678
rect 14356 8676 14380 8678
rect 14436 8676 14460 8678
rect 14516 8676 14540 8678
rect 14596 8676 14602 8678
rect 14294 8667 14602 8676
rect 14660 8537 14688 8774
rect 14646 8528 14702 8537
rect 14646 8463 14702 8472
rect 14200 7806 14780 7834
rect 14294 7644 14602 7653
rect 14294 7642 14300 7644
rect 14356 7642 14380 7644
rect 14436 7642 14460 7644
rect 14516 7642 14540 7644
rect 14596 7642 14602 7644
rect 14356 7590 14358 7642
rect 14538 7590 14540 7642
rect 14294 7588 14300 7590
rect 14356 7588 14380 7590
rect 14436 7588 14460 7590
rect 14516 7588 14540 7590
rect 14596 7588 14602 7590
rect 14294 7579 14602 7588
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14108 5817 14136 6598
rect 14294 6556 14602 6565
rect 14294 6554 14300 6556
rect 14356 6554 14380 6556
rect 14436 6554 14460 6556
rect 14516 6554 14540 6556
rect 14596 6554 14602 6556
rect 14356 6502 14358 6554
rect 14538 6502 14540 6554
rect 14294 6500 14300 6502
rect 14356 6500 14380 6502
rect 14436 6500 14460 6502
rect 14516 6500 14540 6502
rect 14596 6500 14602 6502
rect 14294 6491 14602 6500
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14094 5808 14150 5817
rect 13924 5766 14044 5794
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13728 4684 13780 4690
rect 13728 4626 13780 4632
rect 13832 4622 13860 5306
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13832 3942 13860 4082
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13648 3670 13676 3878
rect 13636 3664 13688 3670
rect 13636 3606 13688 3612
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13648 3126 13676 3334
rect 13740 3194 13768 3470
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13636 3120 13688 3126
rect 13636 3062 13688 3068
rect 13176 2304 13228 2310
rect 13176 2246 13228 2252
rect 13372 800 13400 2502
rect 13544 2508 13596 2514
rect 13544 2450 13596 2456
rect 13832 800 13860 3878
rect 13924 3738 13952 5646
rect 14016 5234 14044 5766
rect 14094 5743 14150 5752
rect 14004 5228 14056 5234
rect 14004 5170 14056 5176
rect 14004 5092 14056 5098
rect 14004 5034 14056 5040
rect 14016 4758 14044 5034
rect 14004 4752 14056 4758
rect 14004 4694 14056 4700
rect 14108 4604 14136 5743
rect 14200 5710 14228 5850
rect 14188 5704 14240 5710
rect 14188 5646 14240 5652
rect 14556 5636 14608 5642
rect 14608 5596 14688 5624
rect 14556 5578 14608 5584
rect 14294 5468 14602 5477
rect 14294 5466 14300 5468
rect 14356 5466 14380 5468
rect 14436 5466 14460 5468
rect 14516 5466 14540 5468
rect 14596 5466 14602 5468
rect 14356 5414 14358 5466
rect 14538 5414 14540 5466
rect 14294 5412 14300 5414
rect 14356 5412 14380 5414
rect 14436 5412 14460 5414
rect 14516 5412 14540 5414
rect 14596 5412 14602 5414
rect 14294 5403 14602 5412
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 14292 4865 14320 5170
rect 14278 4856 14334 4865
rect 14278 4791 14334 4800
rect 14188 4752 14240 4758
rect 14188 4694 14240 4700
rect 14016 4576 14136 4604
rect 14016 4185 14044 4576
rect 14096 4480 14148 4486
rect 14096 4422 14148 4428
rect 14002 4176 14058 4185
rect 14002 4111 14058 4120
rect 14004 3936 14056 3942
rect 14004 3878 14056 3884
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 14016 3534 14044 3878
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 14108 1986 14136 4422
rect 14200 2514 14228 4694
rect 14292 4554 14320 4791
rect 14660 4622 14688 5596
rect 14648 4616 14700 4622
rect 14648 4558 14700 4564
rect 14280 4548 14332 4554
rect 14280 4490 14332 4496
rect 14294 4380 14602 4389
rect 14294 4378 14300 4380
rect 14356 4378 14380 4380
rect 14436 4378 14460 4380
rect 14516 4378 14540 4380
rect 14596 4378 14602 4380
rect 14356 4326 14358 4378
rect 14538 4326 14540 4378
rect 14294 4324 14300 4326
rect 14356 4324 14380 4326
rect 14436 4324 14460 4326
rect 14516 4324 14540 4326
rect 14596 4324 14602 4326
rect 14294 4315 14602 4324
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 14476 3602 14504 4082
rect 14646 4040 14702 4049
rect 14646 3975 14702 3984
rect 14660 3942 14688 3975
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14752 3754 14780 7806
rect 14660 3726 14780 3754
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 14294 3292 14602 3301
rect 14294 3290 14300 3292
rect 14356 3290 14380 3292
rect 14436 3290 14460 3292
rect 14516 3290 14540 3292
rect 14596 3290 14602 3292
rect 14356 3238 14358 3290
rect 14538 3238 14540 3290
rect 14294 3236 14300 3238
rect 14356 3236 14380 3238
rect 14436 3236 14460 3238
rect 14516 3236 14540 3238
rect 14596 3236 14602 3238
rect 14294 3227 14602 3236
rect 14372 3120 14424 3126
rect 14370 3088 14372 3097
rect 14424 3088 14426 3097
rect 14370 3023 14426 3032
rect 14660 2990 14688 3726
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 14648 2984 14700 2990
rect 14648 2926 14700 2932
rect 14188 2508 14240 2514
rect 14188 2450 14240 2456
rect 14294 2204 14602 2213
rect 14294 2202 14300 2204
rect 14356 2202 14380 2204
rect 14436 2202 14460 2204
rect 14516 2202 14540 2204
rect 14596 2202 14602 2204
rect 14356 2150 14358 2202
rect 14538 2150 14540 2202
rect 14294 2148 14300 2150
rect 14356 2148 14380 2150
rect 14436 2148 14460 2150
rect 14516 2148 14540 2150
rect 14596 2148 14602 2150
rect 14294 2139 14602 2148
rect 14108 1958 14320 1986
rect 14292 800 14320 1958
rect 14752 800 14780 3130
rect 14844 2582 14872 12406
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 15212 11830 15240 12174
rect 15200 11824 15252 11830
rect 15200 11766 15252 11772
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 14924 11008 14976 11014
rect 14924 10950 14976 10956
rect 14936 7410 14964 10950
rect 15028 9654 15056 11494
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15108 11076 15160 11082
rect 15108 11018 15160 11024
rect 15120 10606 15148 11018
rect 15212 10742 15240 11086
rect 15200 10736 15252 10742
rect 15200 10678 15252 10684
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 15016 9648 15068 9654
rect 15016 9590 15068 9596
rect 15028 8634 15056 9590
rect 15304 8922 15332 14486
rect 15488 14414 15516 16487
rect 15750 16400 15806 17200
rect 16394 16400 16450 17200
rect 17038 16538 17094 17200
rect 17682 16538 17738 17200
rect 17038 16510 17356 16538
rect 17038 16400 17094 16510
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 15396 12209 15424 14214
rect 15764 13938 15792 16400
rect 16302 16144 16358 16153
rect 16302 16079 16358 16088
rect 16210 14920 16266 14929
rect 16210 14855 16266 14864
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 15844 14000 15896 14006
rect 15844 13942 15896 13948
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15764 12434 15792 13874
rect 15856 12714 15884 13942
rect 15844 12708 15896 12714
rect 15844 12650 15896 12656
rect 15672 12406 15792 12434
rect 15382 12200 15438 12209
rect 15382 12135 15438 12144
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15396 11218 15424 11494
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15488 11218 15516 11290
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 15580 11150 15608 11494
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15396 9178 15424 9318
rect 15384 9172 15436 9178
rect 15384 9114 15436 9120
rect 15304 8894 15608 8922
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 15028 7954 15056 8570
rect 15016 7948 15068 7954
rect 15016 7890 15068 7896
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 15028 6934 15056 7890
rect 15016 6928 15068 6934
rect 15016 6870 15068 6876
rect 15120 6866 15148 8774
rect 15384 8288 15436 8294
rect 15384 8230 15436 8236
rect 15396 7954 15424 8230
rect 15384 7948 15436 7954
rect 15384 7890 15436 7896
rect 15488 7886 15516 8774
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15384 7744 15436 7750
rect 15384 7686 15436 7692
rect 15396 7546 15424 7686
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 15200 7336 15252 7342
rect 15200 7278 15252 7284
rect 15108 6860 15160 6866
rect 15108 6802 15160 6808
rect 15014 6760 15070 6769
rect 15014 6695 15070 6704
rect 15028 5302 15056 6695
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 15120 5914 15148 6258
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 15212 5794 15240 7278
rect 15304 7002 15332 7346
rect 15292 6996 15344 7002
rect 15292 6938 15344 6944
rect 15384 6792 15436 6798
rect 15384 6734 15436 6740
rect 15396 6254 15424 6734
rect 15384 6248 15436 6254
rect 15384 6190 15436 6196
rect 15476 6248 15528 6254
rect 15476 6190 15528 6196
rect 15488 5914 15516 6190
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 15120 5766 15240 5794
rect 15016 5296 15068 5302
rect 14922 5264 14978 5273
rect 15016 5238 15068 5244
rect 14922 5199 14924 5208
rect 14976 5199 14978 5208
rect 14924 5170 14976 5176
rect 15014 5128 15070 5137
rect 15014 5063 15070 5072
rect 15028 4690 15056 5063
rect 15120 4729 15148 5766
rect 15292 5636 15344 5642
rect 15292 5578 15344 5584
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 15212 5370 15240 5510
rect 15304 5370 15332 5578
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 15474 5264 15530 5273
rect 15474 5199 15476 5208
rect 15528 5199 15530 5208
rect 15476 5170 15528 5176
rect 15106 4720 15162 4729
rect 15016 4684 15068 4690
rect 15106 4655 15162 4664
rect 15016 4626 15068 4632
rect 14924 4616 14976 4622
rect 14924 4558 14976 4564
rect 14936 3058 14964 4558
rect 15580 3466 15608 8894
rect 15672 4078 15700 12406
rect 15752 11348 15804 11354
rect 15752 11290 15804 11296
rect 15764 7342 15792 11290
rect 15752 7336 15804 7342
rect 15752 7278 15804 7284
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15764 6390 15792 6598
rect 15752 6384 15804 6390
rect 15752 6326 15804 6332
rect 15752 6248 15804 6254
rect 15752 6190 15804 6196
rect 15764 5778 15792 6190
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15752 5296 15804 5302
rect 15752 5238 15804 5244
rect 15764 4690 15792 5238
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 15660 4072 15712 4078
rect 15660 4014 15712 4020
rect 15856 3602 15884 12650
rect 16040 12102 16068 14350
rect 16224 13938 16252 14855
rect 16316 14414 16344 16079
rect 16408 14958 16436 16400
rect 16854 15736 16910 15745
rect 16854 15671 16910 15680
rect 16396 14952 16448 14958
rect 16396 14894 16448 14900
rect 16518 14716 16826 14725
rect 16518 14714 16524 14716
rect 16580 14714 16604 14716
rect 16660 14714 16684 14716
rect 16740 14714 16764 14716
rect 16820 14714 16826 14716
rect 16580 14662 16582 14714
rect 16762 14662 16764 14714
rect 16518 14660 16524 14662
rect 16580 14660 16604 14662
rect 16660 14660 16684 14662
rect 16740 14660 16764 14662
rect 16820 14660 16826 14662
rect 16518 14651 16826 14660
rect 16762 14512 16818 14521
rect 16762 14447 16764 14456
rect 16816 14447 16818 14456
rect 16764 14418 16816 14424
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 16868 14226 16896 15671
rect 17130 15328 17186 15337
rect 17130 15263 17186 15272
rect 16948 14408 17000 14414
rect 16948 14350 17000 14356
rect 16776 14198 16896 14226
rect 16486 14104 16542 14113
rect 16486 14039 16542 14048
rect 16500 13938 16528 14039
rect 16212 13932 16264 13938
rect 16212 13874 16264 13880
rect 16488 13932 16540 13938
rect 16488 13874 16540 13880
rect 16776 13870 16804 14198
rect 16854 14104 16910 14113
rect 16854 14039 16910 14048
rect 16764 13864 16816 13870
rect 16764 13806 16816 13812
rect 16120 13796 16172 13802
rect 16120 13738 16172 13744
rect 16132 13394 16160 13738
rect 16776 13734 16804 13806
rect 16304 13728 16356 13734
rect 16304 13670 16356 13676
rect 16764 13728 16816 13734
rect 16764 13670 16816 13676
rect 16120 13388 16172 13394
rect 16120 13330 16172 13336
rect 16316 12889 16344 13670
rect 16518 13628 16826 13637
rect 16518 13626 16524 13628
rect 16580 13626 16604 13628
rect 16660 13626 16684 13628
rect 16740 13626 16764 13628
rect 16820 13626 16826 13628
rect 16580 13574 16582 13626
rect 16762 13574 16764 13626
rect 16518 13572 16524 13574
rect 16580 13572 16604 13574
rect 16660 13572 16684 13574
rect 16740 13572 16764 13574
rect 16820 13572 16826 13574
rect 16518 13563 16826 13572
rect 16868 13530 16896 14039
rect 16856 13524 16908 13530
rect 16856 13466 16908 13472
rect 16960 13394 16988 14350
rect 17040 13728 17092 13734
rect 17040 13670 17092 13676
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 17052 13274 17080 13670
rect 16580 13252 16632 13258
rect 16580 13194 16632 13200
rect 16960 13246 17080 13274
rect 17144 13258 17172 15263
rect 17224 14408 17276 14414
rect 17224 14350 17276 14356
rect 17132 13252 17184 13258
rect 16302 12880 16358 12889
rect 16212 12844 16264 12850
rect 16592 12850 16620 13194
rect 16960 12918 16988 13246
rect 17132 13194 17184 13200
rect 17040 13184 17092 13190
rect 17040 13126 17092 13132
rect 16948 12912 17000 12918
rect 16948 12854 17000 12860
rect 16302 12815 16358 12824
rect 16580 12844 16632 12850
rect 16212 12786 16264 12792
rect 16580 12786 16632 12792
rect 15936 12096 15988 12102
rect 15936 12038 15988 12044
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 15948 11830 15976 12038
rect 15936 11824 15988 11830
rect 15936 11766 15988 11772
rect 16040 11694 16068 12038
rect 16028 11688 16080 11694
rect 16028 11630 16080 11636
rect 16040 9926 16068 11630
rect 16224 10130 16252 12786
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16518 12540 16826 12549
rect 16518 12538 16524 12540
rect 16580 12538 16604 12540
rect 16660 12538 16684 12540
rect 16740 12538 16764 12540
rect 16820 12538 16826 12540
rect 16580 12486 16582 12538
rect 16762 12486 16764 12538
rect 16518 12484 16524 12486
rect 16580 12484 16604 12486
rect 16660 12484 16684 12486
rect 16740 12484 16764 12486
rect 16820 12484 16826 12486
rect 16518 12475 16826 12484
rect 16868 12434 16896 12582
rect 16868 12406 16988 12434
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16518 11452 16826 11461
rect 16518 11450 16524 11452
rect 16580 11450 16604 11452
rect 16660 11450 16684 11452
rect 16740 11450 16764 11452
rect 16820 11450 16826 11452
rect 16580 11398 16582 11450
rect 16762 11398 16764 11450
rect 16518 11396 16524 11398
rect 16580 11396 16604 11398
rect 16660 11396 16684 11398
rect 16740 11396 16764 11398
rect 16820 11396 16826 11398
rect 16518 11387 16826 11396
rect 16868 11150 16896 11494
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 16396 11076 16448 11082
rect 16396 11018 16448 11024
rect 16408 10266 16436 11018
rect 16854 10704 16910 10713
rect 16854 10639 16910 10648
rect 16518 10364 16826 10373
rect 16518 10362 16524 10364
rect 16580 10362 16604 10364
rect 16660 10362 16684 10364
rect 16740 10362 16764 10364
rect 16820 10362 16826 10364
rect 16580 10310 16582 10362
rect 16762 10310 16764 10362
rect 16518 10308 16524 10310
rect 16580 10308 16604 10310
rect 16660 10308 16684 10310
rect 16740 10308 16764 10310
rect 16820 10308 16826 10310
rect 16518 10299 16826 10308
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 16028 9920 16080 9926
rect 16028 9862 16080 9868
rect 16868 9466 16896 10639
rect 16960 10062 16988 12406
rect 17052 11286 17080 13126
rect 17144 12918 17172 13194
rect 17132 12912 17184 12918
rect 17132 12854 17184 12860
rect 17236 12434 17264 14350
rect 17328 13297 17356 16510
rect 17682 16510 17908 16538
rect 17682 16400 17738 16510
rect 17684 14408 17736 14414
rect 17684 14350 17736 14356
rect 17696 13705 17724 14350
rect 17776 13864 17828 13870
rect 17776 13806 17828 13812
rect 17682 13696 17738 13705
rect 17682 13631 17738 13640
rect 17696 13462 17724 13631
rect 17684 13456 17736 13462
rect 17684 13398 17736 13404
rect 17684 13320 17736 13326
rect 17314 13288 17370 13297
rect 17788 13297 17816 13806
rect 17684 13262 17736 13268
rect 17774 13288 17830 13297
rect 17314 13223 17370 13232
rect 17592 13252 17644 13258
rect 17592 13194 17644 13200
rect 17408 13184 17460 13190
rect 17408 13126 17460 13132
rect 17236 12406 17356 12434
rect 17224 12368 17276 12374
rect 17224 12310 17276 12316
rect 17236 11830 17264 12310
rect 17224 11824 17276 11830
rect 17224 11766 17276 11772
rect 17328 11778 17356 12406
rect 17420 11937 17448 13126
rect 17604 12918 17632 13194
rect 17592 12912 17644 12918
rect 17590 12880 17592 12889
rect 17644 12880 17646 12889
rect 17500 12844 17552 12850
rect 17590 12815 17646 12824
rect 17500 12786 17552 12792
rect 17406 11928 17462 11937
rect 17406 11863 17462 11872
rect 17130 11656 17186 11665
rect 17130 11591 17186 11600
rect 17040 11280 17092 11286
rect 17040 11222 17092 11228
rect 17144 11150 17172 11591
rect 17132 11144 17184 11150
rect 17038 11112 17094 11121
rect 17132 11086 17184 11092
rect 17038 11047 17094 11056
rect 17052 10810 17080 11047
rect 17040 10804 17092 10810
rect 17040 10746 17092 10752
rect 17132 10600 17184 10606
rect 17132 10542 17184 10548
rect 17144 10266 17172 10542
rect 17236 10266 17264 11766
rect 17328 11750 17448 11778
rect 17316 11688 17368 11694
rect 17316 11630 17368 11636
rect 17328 10606 17356 11630
rect 17316 10600 17368 10606
rect 17316 10542 17368 10548
rect 17132 10260 17184 10266
rect 17132 10202 17184 10208
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 17328 10130 17356 10542
rect 17420 10418 17448 11750
rect 17512 11150 17540 12786
rect 17696 12481 17724 13262
rect 17774 13223 17830 13232
rect 17788 12986 17816 13223
rect 17776 12980 17828 12986
rect 17776 12922 17828 12928
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 17682 12472 17738 12481
rect 17682 12407 17738 12416
rect 17592 12096 17644 12102
rect 17592 12038 17644 12044
rect 17684 12096 17736 12102
rect 17788 12073 17816 12718
rect 17880 12345 17908 16510
rect 18326 16400 18382 17200
rect 18970 16400 19026 17200
rect 19614 16400 19670 17200
rect 18340 14822 18368 16400
rect 18984 14890 19012 16400
rect 18972 14884 19024 14890
rect 18972 14826 19024 14832
rect 18328 14816 18380 14822
rect 18328 14758 18380 14764
rect 17960 14408 18012 14414
rect 17960 14350 18012 14356
rect 17972 12442 18000 14350
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 17960 12436 18012 12442
rect 17960 12378 18012 12384
rect 17866 12336 17922 12345
rect 17866 12271 17922 12280
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 17684 12038 17736 12044
rect 17774 12064 17830 12073
rect 17604 11762 17632 12038
rect 17592 11756 17644 11762
rect 17592 11698 17644 11704
rect 17696 11694 17724 12038
rect 17774 11999 17830 12008
rect 17774 11928 17830 11937
rect 17774 11863 17830 11872
rect 17684 11688 17736 11694
rect 17684 11630 17736 11636
rect 17592 11280 17644 11286
rect 17696 11257 17724 11630
rect 17592 11222 17644 11228
rect 17682 11248 17738 11257
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17420 10390 17540 10418
rect 17408 10260 17460 10266
rect 17408 10202 17460 10208
rect 17420 10130 17448 10202
rect 17040 10124 17092 10130
rect 17040 10066 17092 10072
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 17408 10124 17460 10130
rect 17408 10066 17460 10072
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 16960 9722 16988 9998
rect 16948 9716 17000 9722
rect 16948 9658 17000 9664
rect 16868 9438 16988 9466
rect 16518 9276 16826 9285
rect 16518 9274 16524 9276
rect 16580 9274 16604 9276
rect 16660 9274 16684 9276
rect 16740 9274 16764 9276
rect 16820 9274 16826 9276
rect 16580 9222 16582 9274
rect 16762 9222 16764 9274
rect 16518 9220 16524 9222
rect 16580 9220 16604 9222
rect 16660 9220 16684 9222
rect 16740 9220 16764 9222
rect 16820 9220 16826 9222
rect 16518 9211 16826 9220
rect 16028 9036 16080 9042
rect 16028 8978 16080 8984
rect 16040 8566 16068 8978
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16028 8560 16080 8566
rect 16028 8502 16080 8508
rect 15936 8492 15988 8498
rect 15936 8434 15988 8440
rect 15948 6186 15976 8434
rect 16040 8430 16068 8502
rect 16028 8424 16080 8430
rect 16028 8366 16080 8372
rect 16028 7812 16080 7818
rect 16028 7754 16080 7760
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 15948 5778 15976 6122
rect 16040 5778 16068 7754
rect 16212 7268 16264 7274
rect 16212 7210 16264 7216
rect 16224 6866 16252 7210
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 16212 6384 16264 6390
rect 16212 6326 16264 6332
rect 15936 5772 15988 5778
rect 15936 5714 15988 5720
rect 16028 5772 16080 5778
rect 16028 5714 16080 5720
rect 15948 5234 15976 5714
rect 16040 5352 16068 5714
rect 16224 5710 16252 6326
rect 16316 5778 16344 8910
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 16592 8634 16620 8774
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16518 8188 16826 8197
rect 16518 8186 16524 8188
rect 16580 8186 16604 8188
rect 16660 8186 16684 8188
rect 16740 8186 16764 8188
rect 16820 8186 16826 8188
rect 16580 8134 16582 8186
rect 16762 8134 16764 8186
rect 16518 8132 16524 8134
rect 16580 8132 16604 8134
rect 16660 8132 16684 8134
rect 16740 8132 16764 8134
rect 16820 8132 16826 8134
rect 16518 8123 16826 8132
rect 16394 7848 16450 7857
rect 16394 7783 16450 7792
rect 16408 7546 16436 7783
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16518 7100 16826 7109
rect 16518 7098 16524 7100
rect 16580 7098 16604 7100
rect 16660 7098 16684 7100
rect 16740 7098 16764 7100
rect 16820 7098 16826 7100
rect 16580 7046 16582 7098
rect 16762 7046 16764 7098
rect 16518 7044 16524 7046
rect 16580 7044 16604 7046
rect 16660 7044 16684 7046
rect 16740 7044 16764 7046
rect 16820 7044 16826 7046
rect 16518 7035 16826 7044
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16592 6254 16620 6802
rect 16868 6474 16896 8774
rect 16960 8090 16988 9438
rect 17052 8498 17080 10066
rect 17512 10010 17540 10390
rect 17132 9988 17184 9994
rect 17132 9930 17184 9936
rect 17236 9982 17540 10010
rect 17144 9654 17172 9930
rect 17132 9648 17184 9654
rect 17132 9590 17184 9596
rect 17132 8900 17184 8906
rect 17132 8842 17184 8848
rect 17040 8492 17092 8498
rect 17040 8434 17092 8440
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 16960 7886 16988 8026
rect 16948 7880 17000 7886
rect 16948 7822 17000 7828
rect 17144 7698 17172 8842
rect 16776 6446 16896 6474
rect 16960 7670 17172 7698
rect 16960 6458 16988 7670
rect 17236 7426 17264 9982
rect 17500 9920 17552 9926
rect 17500 9862 17552 9868
rect 17408 9512 17460 9518
rect 17314 9480 17370 9489
rect 17408 9454 17460 9460
rect 17314 9415 17370 9424
rect 17328 9178 17356 9415
rect 17420 9217 17448 9454
rect 17406 9208 17462 9217
rect 17316 9172 17368 9178
rect 17406 9143 17462 9152
rect 17316 9114 17368 9120
rect 17328 8974 17356 9114
rect 17316 8968 17368 8974
rect 17316 8910 17368 8916
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17316 8084 17368 8090
rect 17316 8026 17368 8032
rect 17328 7750 17356 8026
rect 17316 7744 17368 7750
rect 17316 7686 17368 7692
rect 17052 7398 17264 7426
rect 17328 7410 17356 7686
rect 17316 7404 17368 7410
rect 16948 6452 17000 6458
rect 16776 6254 16804 6446
rect 16948 6394 17000 6400
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 16764 6248 16816 6254
rect 16764 6190 16816 6196
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16408 5914 16436 6054
rect 16518 6012 16826 6021
rect 16518 6010 16524 6012
rect 16580 6010 16604 6012
rect 16660 6010 16684 6012
rect 16740 6010 16764 6012
rect 16820 6010 16826 6012
rect 16580 5958 16582 6010
rect 16762 5958 16764 6010
rect 16518 5956 16524 5958
rect 16580 5956 16604 5958
rect 16660 5956 16684 5958
rect 16740 5956 16764 5958
rect 16820 5956 16826 5958
rect 16518 5947 16826 5956
rect 16396 5908 16448 5914
rect 16396 5850 16448 5856
rect 16672 5840 16724 5846
rect 16672 5782 16724 5788
rect 16304 5772 16356 5778
rect 16304 5714 16356 5720
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 16684 5522 16712 5782
rect 16500 5494 16712 5522
rect 16500 5370 16528 5494
rect 16868 5370 16896 6258
rect 16948 6248 17000 6254
rect 16946 6216 16948 6225
rect 17000 6216 17002 6225
rect 16946 6151 17002 6160
rect 16948 6112 17000 6118
rect 16948 6054 17000 6060
rect 16960 5642 16988 6054
rect 17052 5846 17080 7398
rect 17316 7346 17368 7352
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 17236 6866 17264 7278
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 17328 6458 17356 6734
rect 17224 6452 17276 6458
rect 17224 6394 17276 6400
rect 17316 6452 17368 6458
rect 17316 6394 17368 6400
rect 17040 5840 17092 5846
rect 17040 5782 17092 5788
rect 17040 5704 17092 5710
rect 17040 5646 17092 5652
rect 16948 5636 17000 5642
rect 16948 5578 17000 5584
rect 17052 5370 17080 5646
rect 16488 5364 16540 5370
rect 16040 5324 16252 5352
rect 15936 5228 15988 5234
rect 15936 5170 15988 5176
rect 16040 5166 16068 5324
rect 16118 5264 16174 5273
rect 16118 5199 16174 5208
rect 16028 5160 16080 5166
rect 16028 5102 16080 5108
rect 16132 4486 16160 5199
rect 16224 5098 16252 5324
rect 16488 5306 16540 5312
rect 16856 5364 16908 5370
rect 16856 5306 16908 5312
rect 17040 5364 17092 5370
rect 17040 5306 17092 5312
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 17132 5160 17184 5166
rect 17236 5148 17264 6394
rect 17314 5808 17370 5817
rect 17314 5743 17316 5752
rect 17368 5743 17370 5752
rect 17316 5714 17368 5720
rect 17184 5120 17264 5148
rect 17132 5102 17184 5108
rect 16212 5092 16264 5098
rect 16212 5034 16264 5040
rect 16304 5024 16356 5030
rect 16304 4966 16356 4972
rect 16212 4752 16264 4758
rect 16212 4694 16264 4700
rect 16120 4480 16172 4486
rect 16120 4422 16172 4428
rect 15844 3596 15896 3602
rect 15844 3538 15896 3544
rect 15568 3460 15620 3466
rect 15568 3402 15620 3408
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 16132 2961 16160 4422
rect 16118 2952 16174 2961
rect 16118 2887 16174 2896
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 15660 2848 15712 2854
rect 15660 2790 15712 2796
rect 16120 2848 16172 2854
rect 16120 2790 16172 2796
rect 14832 2576 14884 2582
rect 14832 2518 14884 2524
rect 15212 2514 15240 2790
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 15200 2304 15252 2310
rect 15200 2246 15252 2252
rect 15212 800 15240 2246
rect 15672 800 15700 2790
rect 16132 2446 16160 2790
rect 16224 2446 16252 4694
rect 16316 3466 16344 4966
rect 16518 4924 16826 4933
rect 16518 4922 16524 4924
rect 16580 4922 16604 4924
rect 16660 4922 16684 4924
rect 16740 4922 16764 4924
rect 16820 4922 16826 4924
rect 16580 4870 16582 4922
rect 16762 4870 16764 4922
rect 16518 4868 16524 4870
rect 16580 4868 16604 4870
rect 16660 4868 16684 4870
rect 16740 4868 16764 4870
rect 16820 4868 16826 4870
rect 16518 4859 16826 4868
rect 16396 4684 16448 4690
rect 16396 4626 16448 4632
rect 16408 4486 16436 4626
rect 16764 4616 16816 4622
rect 16868 4604 16896 5102
rect 16816 4576 16896 4604
rect 16764 4558 16816 4564
rect 16396 4480 16448 4486
rect 16396 4422 16448 4428
rect 16856 4480 16908 4486
rect 16856 4422 16908 4428
rect 17224 4480 17276 4486
rect 17224 4422 17276 4428
rect 17316 4480 17368 4486
rect 17316 4422 17368 4428
rect 16408 4282 16436 4422
rect 16396 4276 16448 4282
rect 16396 4218 16448 4224
rect 16396 4004 16448 4010
rect 16396 3946 16448 3952
rect 16408 3738 16436 3946
rect 16518 3836 16826 3845
rect 16518 3834 16524 3836
rect 16580 3834 16604 3836
rect 16660 3834 16684 3836
rect 16740 3834 16764 3836
rect 16820 3834 16826 3836
rect 16580 3782 16582 3834
rect 16762 3782 16764 3834
rect 16518 3780 16524 3782
rect 16580 3780 16604 3782
rect 16660 3780 16684 3782
rect 16740 3780 16764 3782
rect 16820 3780 16826 3782
rect 16518 3771 16826 3780
rect 16396 3732 16448 3738
rect 16396 3674 16448 3680
rect 16304 3460 16356 3466
rect 16304 3402 16356 3408
rect 16868 3058 16896 4422
rect 16960 4146 17080 4162
rect 16960 4140 17092 4146
rect 16960 4134 17040 4140
rect 16960 3670 16988 4134
rect 17040 4082 17092 4088
rect 17040 4004 17092 4010
rect 17040 3946 17092 3952
rect 16948 3664 17000 3670
rect 16948 3606 17000 3612
rect 16948 3528 17000 3534
rect 16948 3470 17000 3476
rect 16960 3194 16988 3470
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 16304 2916 16356 2922
rect 16304 2858 16356 2864
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 16212 2440 16264 2446
rect 16212 2382 16264 2388
rect 16316 1057 16344 2858
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 16518 2748 16826 2757
rect 16518 2746 16524 2748
rect 16580 2746 16604 2748
rect 16660 2746 16684 2748
rect 16740 2746 16764 2748
rect 16820 2746 16826 2748
rect 16580 2694 16582 2746
rect 16762 2694 16764 2746
rect 16518 2692 16524 2694
rect 16580 2692 16604 2694
rect 16660 2692 16684 2694
rect 16740 2692 16764 2694
rect 16820 2692 16826 2694
rect 16518 2683 16826 2692
rect 16580 2576 16632 2582
rect 16580 2518 16632 2524
rect 16396 2304 16448 2310
rect 16396 2246 16448 2252
rect 16302 1048 16358 1057
rect 16302 983 16358 992
rect 16132 870 16252 898
rect 16132 800 16160 870
rect 12084 734 12296 762
rect 12438 0 12494 800
rect 12898 0 12954 800
rect 13358 0 13414 800
rect 13818 0 13874 800
rect 14278 0 14334 800
rect 14738 0 14794 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 16224 762 16252 870
rect 16408 762 16436 2246
rect 16592 800 16620 2518
rect 16960 1465 16988 2790
rect 17052 2446 17080 3946
rect 17132 3936 17184 3942
rect 17132 3878 17184 3884
rect 17144 2446 17172 3878
rect 17236 3126 17264 4422
rect 17224 3120 17276 3126
rect 17224 3062 17276 3068
rect 17328 2990 17356 4422
rect 17420 3058 17448 8570
rect 17512 3534 17540 9862
rect 17604 8401 17632 11222
rect 17682 11183 17738 11192
rect 17684 11144 17736 11150
rect 17684 11086 17736 11092
rect 17696 10849 17724 11086
rect 17682 10840 17738 10849
rect 17682 10775 17738 10784
rect 17788 10656 17816 11863
rect 17880 11665 17908 12174
rect 17972 11801 18000 12174
rect 17958 11792 18014 11801
rect 17958 11727 18014 11736
rect 17866 11656 17922 11665
rect 17866 11591 17922 11600
rect 18064 11393 18092 13262
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 18156 11898 18184 12378
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 18050 11384 18106 11393
rect 18050 11319 18106 11328
rect 17960 11144 18012 11150
rect 17960 11086 18012 11092
rect 17972 10810 18000 11086
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 17960 10804 18012 10810
rect 17960 10746 18012 10752
rect 17788 10628 17908 10656
rect 17684 10600 17736 10606
rect 17684 10542 17736 10548
rect 17696 10441 17724 10542
rect 17682 10432 17738 10441
rect 17682 10367 17738 10376
rect 17880 10282 17908 10628
rect 17696 10254 17908 10282
rect 17590 8392 17646 8401
rect 17590 8327 17646 8336
rect 17604 7970 17632 8327
rect 17696 8090 17724 10254
rect 18064 10112 18092 10950
rect 17788 10084 18092 10112
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17604 7942 17724 7970
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17604 7449 17632 7822
rect 17696 7562 17724 7942
rect 17788 7886 17816 10084
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 17880 8498 17908 9318
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17866 8392 17922 8401
rect 17866 8327 17922 8336
rect 17776 7880 17828 7886
rect 17776 7822 17828 7828
rect 17696 7534 17816 7562
rect 17684 7472 17736 7478
rect 17590 7440 17646 7449
rect 17684 7414 17736 7420
rect 17590 7375 17592 7384
rect 17644 7375 17646 7384
rect 17592 7346 17644 7352
rect 17696 7002 17724 7414
rect 17788 7002 17816 7534
rect 17684 6996 17736 7002
rect 17684 6938 17736 6944
rect 17776 6996 17828 7002
rect 17776 6938 17828 6944
rect 17880 6882 17908 8327
rect 17696 6854 17908 6882
rect 17592 6316 17644 6322
rect 17592 6258 17644 6264
rect 17604 5234 17632 6258
rect 17592 5228 17644 5234
rect 17592 5170 17644 5176
rect 17592 4140 17644 4146
rect 17592 4082 17644 4088
rect 17604 3641 17632 4082
rect 17696 4026 17724 6854
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 17880 5914 17908 6734
rect 17972 6202 18000 9862
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 18064 8974 18092 9522
rect 18248 9518 18276 12718
rect 19628 12714 19656 16400
rect 19616 12708 19668 12714
rect 19616 12650 19668 12656
rect 18696 12368 18748 12374
rect 18696 12310 18748 12316
rect 18420 11756 18472 11762
rect 18420 11698 18472 11704
rect 18328 10600 18380 10606
rect 18328 10542 18380 10548
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 18144 9104 18196 9110
rect 18144 9046 18196 9052
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 18052 8356 18104 8362
rect 18052 8298 18104 8304
rect 18064 7993 18092 8298
rect 18050 7984 18106 7993
rect 18050 7919 18106 7928
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 18064 6361 18092 6598
rect 18050 6352 18106 6361
rect 18156 6322 18184 9046
rect 18248 8498 18276 9318
rect 18340 9058 18368 10542
rect 18432 10266 18460 11698
rect 18604 11076 18656 11082
rect 18604 11018 18656 11024
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18418 10024 18474 10033
rect 18418 9959 18420 9968
rect 18472 9959 18474 9968
rect 18420 9930 18472 9936
rect 18510 9616 18566 9625
rect 18420 9580 18472 9586
rect 18510 9551 18566 9560
rect 18420 9522 18472 9528
rect 18432 9217 18460 9522
rect 18418 9208 18474 9217
rect 18418 9143 18474 9152
rect 18340 9030 18460 9058
rect 18328 8968 18380 8974
rect 18328 8910 18380 8916
rect 18340 8809 18368 8910
rect 18326 8800 18382 8809
rect 18326 8735 18382 8744
rect 18432 8514 18460 9030
rect 18524 8974 18552 9551
rect 18512 8968 18564 8974
rect 18512 8910 18564 8916
rect 18236 8492 18288 8498
rect 18432 8486 18552 8514
rect 18236 8434 18288 8440
rect 18418 8392 18474 8401
rect 18418 8327 18420 8336
rect 18472 8327 18474 8336
rect 18420 8298 18472 8304
rect 18328 8016 18380 8022
rect 18328 7958 18380 7964
rect 18236 7200 18288 7206
rect 18236 7142 18288 7148
rect 18248 6798 18276 7142
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18050 6287 18106 6296
rect 18144 6316 18196 6322
rect 18144 6258 18196 6264
rect 17972 6174 18276 6202
rect 17960 6112 18012 6118
rect 17960 6054 18012 6060
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 17972 4570 18000 6054
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 18064 4729 18092 4966
rect 18144 4752 18196 4758
rect 18050 4720 18106 4729
rect 18144 4694 18196 4700
rect 18050 4655 18106 4664
rect 17788 4542 18000 4570
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 17788 4146 17816 4542
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 17696 3998 17816 4026
rect 17684 3936 17736 3942
rect 17684 3878 17736 3884
rect 17590 3632 17646 3641
rect 17590 3567 17646 3576
rect 17500 3528 17552 3534
rect 17500 3470 17552 3476
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 17316 2984 17368 2990
rect 17316 2926 17368 2932
rect 17040 2440 17092 2446
rect 17040 2382 17092 2388
rect 17132 2440 17184 2446
rect 17132 2382 17184 2388
rect 17040 2304 17092 2310
rect 17040 2246 17092 2252
rect 16946 1456 17002 1465
rect 16946 1391 17002 1400
rect 17052 800 17080 2246
rect 17604 1873 17632 3334
rect 17696 2446 17724 3878
rect 17788 3505 17816 3998
rect 17880 3534 17908 4422
rect 17972 4146 18000 4422
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 18064 3534 18092 4558
rect 17868 3528 17920 3534
rect 17774 3496 17830 3505
rect 17868 3470 17920 3476
rect 18052 3528 18104 3534
rect 18052 3470 18104 3476
rect 17774 3431 17830 3440
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 18064 3097 18092 3334
rect 18050 3088 18106 3097
rect 18050 3023 18106 3032
rect 17868 2848 17920 2854
rect 17868 2790 17920 2796
rect 17684 2440 17736 2446
rect 17684 2382 17736 2388
rect 17776 2304 17828 2310
rect 17880 2281 17908 2790
rect 18156 2446 18184 4694
rect 18248 3058 18276 6174
rect 18340 4622 18368 7958
rect 18420 7744 18472 7750
rect 18420 7686 18472 7692
rect 18432 7585 18460 7686
rect 18418 7576 18474 7585
rect 18418 7511 18474 7520
rect 18420 7200 18472 7206
rect 18418 7168 18420 7177
rect 18472 7168 18474 7177
rect 18418 7103 18474 7112
rect 18418 6760 18474 6769
rect 18418 6695 18474 6704
rect 18432 6662 18460 6695
rect 18420 6656 18472 6662
rect 18420 6598 18472 6604
rect 18420 6112 18472 6118
rect 18420 6054 18472 6060
rect 18432 5953 18460 6054
rect 18418 5944 18474 5953
rect 18418 5879 18474 5888
rect 18420 5568 18472 5574
rect 18418 5536 18420 5545
rect 18472 5536 18474 5545
rect 18418 5471 18474 5480
rect 18418 5128 18474 5137
rect 18418 5063 18420 5072
rect 18472 5063 18474 5072
rect 18420 5034 18472 5040
rect 18328 4616 18380 4622
rect 18524 4593 18552 8486
rect 18616 5234 18644 11018
rect 18604 5228 18656 5234
rect 18604 5170 18656 5176
rect 18328 4558 18380 4564
rect 18510 4584 18566 4593
rect 18510 4519 18566 4528
rect 18420 4480 18472 4486
rect 18420 4422 18472 4428
rect 18432 4321 18460 4422
rect 18418 4312 18474 4321
rect 18418 4247 18474 4256
rect 18420 3936 18472 3942
rect 18418 3904 18420 3913
rect 18472 3904 18474 3913
rect 18418 3839 18474 3848
rect 18512 3664 18564 3670
rect 18512 3606 18564 3612
rect 18418 3496 18474 3505
rect 18418 3431 18474 3440
rect 18432 3398 18460 3431
rect 18420 3392 18472 3398
rect 18420 3334 18472 3340
rect 18236 3052 18288 3058
rect 18236 2994 18288 3000
rect 18328 2916 18380 2922
rect 18328 2858 18380 2864
rect 18144 2440 18196 2446
rect 18144 2382 18196 2388
rect 18052 2304 18104 2310
rect 17776 2246 17828 2252
rect 17866 2272 17922 2281
rect 17590 1864 17646 1873
rect 17590 1799 17646 1808
rect 17512 870 17632 898
rect 17512 800 17540 870
rect 16224 734 16436 762
rect 16578 0 16634 800
rect 17038 0 17094 800
rect 17498 0 17554 800
rect 17604 762 17632 870
rect 17788 762 17816 2246
rect 17866 2207 17922 2216
rect 17972 2264 18052 2292
rect 17972 800 18000 2264
rect 18052 2246 18104 2252
rect 18340 1442 18368 2858
rect 18420 2848 18472 2854
rect 18420 2790 18472 2796
rect 18432 2689 18460 2790
rect 18418 2680 18474 2689
rect 18418 2615 18474 2624
rect 18340 1414 18460 1442
rect 18432 800 18460 1414
rect 17604 734 17816 762
rect 17958 0 18014 800
rect 18418 0 18474 800
rect 18524 649 18552 3606
rect 18708 3534 18736 12310
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 18786 8528 18842 8537
rect 18786 8463 18842 8472
rect 18800 6186 18828 8463
rect 18788 6180 18840 6186
rect 18788 6122 18840 6128
rect 18892 5273 18920 11630
rect 18878 5264 18934 5273
rect 18878 5199 18934 5208
rect 18880 4004 18932 4010
rect 18880 3946 18932 3952
rect 18696 3528 18748 3534
rect 18696 3470 18748 3476
rect 18892 800 18920 3946
rect 18510 640 18566 649
rect 18510 575 18566 584
rect 18878 0 18934 800
<< via2 >>
rect 1950 14356 1952 14376
rect 1952 14356 2004 14376
rect 2004 14356 2006 14376
rect 1950 14320 2006 14356
rect 2226 13776 2282 13832
rect 3790 16632 3846 16688
rect 2778 15816 2834 15872
rect 3054 15000 3110 15056
rect 2962 14592 3018 14648
rect 3180 14714 3236 14716
rect 3260 14714 3316 14716
rect 3340 14714 3396 14716
rect 3420 14714 3476 14716
rect 3180 14662 3226 14714
rect 3226 14662 3236 14714
rect 3260 14662 3290 14714
rect 3290 14662 3302 14714
rect 3302 14662 3316 14714
rect 3340 14662 3354 14714
rect 3354 14662 3366 14714
rect 3366 14662 3396 14714
rect 3420 14662 3430 14714
rect 3430 14662 3476 14714
rect 3180 14660 3236 14662
rect 3260 14660 3316 14662
rect 3340 14660 3396 14662
rect 3420 14660 3476 14662
rect 4066 16224 4122 16280
rect 3606 14456 3662 14512
rect 2962 14184 3018 14240
rect 2042 13368 2098 13424
rect 2778 12960 2834 13016
rect 2778 12824 2834 12880
rect 3180 13626 3236 13628
rect 3260 13626 3316 13628
rect 3340 13626 3396 13628
rect 3420 13626 3476 13628
rect 3180 13574 3226 13626
rect 3226 13574 3236 13626
rect 3260 13574 3290 13626
rect 3290 13574 3302 13626
rect 3302 13574 3316 13626
rect 3340 13574 3354 13626
rect 3354 13574 3366 13626
rect 3366 13574 3396 13626
rect 3420 13574 3430 13626
rect 3430 13574 3476 13626
rect 3180 13572 3236 13574
rect 3260 13572 3316 13574
rect 3340 13572 3396 13574
rect 3420 13572 3476 13574
rect 4158 15408 4214 15464
rect 3514 13368 3570 13424
rect 1490 10104 1546 10160
rect 1490 9580 1546 9616
rect 1490 9560 1492 9580
rect 1492 9560 1544 9580
rect 1544 9560 1546 9580
rect 1490 9288 1546 9344
rect 1490 8472 1546 8528
rect 1490 8084 1546 8120
rect 1490 8064 1492 8084
rect 1492 8064 1544 8084
rect 1544 8064 1546 8084
rect 1490 7248 1546 7304
rect 1582 6840 1638 6896
rect 1582 6704 1638 6760
rect 1950 11212 2006 11248
rect 1950 11192 1952 11212
rect 1952 11192 2004 11212
rect 2004 11192 2006 11212
rect 2870 12688 2926 12744
rect 2226 12552 2282 12608
rect 2410 12164 2466 12200
rect 2410 12144 2412 12164
rect 2412 12144 2464 12164
rect 2464 12144 2466 12164
rect 2226 11328 2282 11384
rect 2226 10920 2282 10976
rect 2134 10648 2190 10704
rect 2226 10548 2228 10568
rect 2228 10548 2280 10568
rect 2280 10548 2282 10568
rect 2226 10512 2282 10548
rect 1950 8900 2006 8936
rect 1950 8880 1952 8900
rect 1952 8880 2004 8900
rect 2004 8880 2006 8900
rect 1858 7692 1860 7712
rect 1860 7692 1912 7712
rect 1912 7692 1914 7712
rect 1858 7656 1914 7692
rect 1490 6024 1546 6080
rect 1674 5772 1730 5808
rect 1674 5752 1676 5772
rect 1676 5752 1728 5772
rect 1728 5752 1730 5772
rect 2778 11736 2834 11792
rect 2502 11600 2558 11656
rect 2318 8472 2374 8528
rect 2134 6840 2190 6896
rect 1950 5616 2006 5672
rect 1490 4820 1546 4856
rect 1490 4800 1492 4820
rect 1492 4800 1544 4820
rect 1544 4800 1546 4820
rect 1858 4428 1860 4448
rect 1860 4428 1912 4448
rect 1912 4428 1914 4448
rect 1858 4392 1914 4428
rect 1490 4004 1546 4040
rect 1490 3984 1492 4004
rect 1492 3984 1544 4004
rect 1544 3984 1546 4004
rect 1858 3576 1914 3632
rect 1490 3168 1546 3224
rect 1490 2760 1546 2816
rect 2410 5344 2466 5400
rect 3514 12724 3516 12744
rect 3516 12724 3568 12744
rect 3568 12724 3570 12744
rect 3514 12688 3570 12724
rect 3180 12538 3236 12540
rect 3260 12538 3316 12540
rect 3340 12538 3396 12540
rect 3420 12538 3476 12540
rect 3180 12486 3226 12538
rect 3226 12486 3236 12538
rect 3260 12486 3290 12538
rect 3290 12486 3302 12538
rect 3302 12486 3316 12538
rect 3340 12486 3354 12538
rect 3354 12486 3366 12538
rect 3366 12486 3396 12538
rect 3420 12486 3430 12538
rect 3430 12486 3476 12538
rect 3180 12484 3236 12486
rect 3260 12484 3316 12486
rect 3340 12484 3396 12486
rect 3420 12484 3476 12486
rect 3146 12164 3202 12200
rect 3146 12144 3148 12164
rect 3148 12144 3200 12164
rect 3200 12144 3202 12164
rect 3790 12960 3846 13016
rect 3698 12280 3754 12336
rect 3180 11450 3236 11452
rect 3260 11450 3316 11452
rect 3340 11450 3396 11452
rect 3420 11450 3476 11452
rect 3180 11398 3226 11450
rect 3226 11398 3236 11450
rect 3260 11398 3290 11450
rect 3290 11398 3302 11450
rect 3302 11398 3316 11450
rect 3340 11398 3354 11450
rect 3354 11398 3366 11450
rect 3366 11398 3396 11450
rect 3420 11398 3430 11450
rect 3430 11398 3476 11450
rect 3180 11396 3236 11398
rect 3260 11396 3316 11398
rect 3340 11396 3396 11398
rect 3420 11396 3476 11398
rect 3606 11600 3662 11656
rect 4066 13268 4068 13288
rect 4068 13268 4120 13288
rect 4120 13268 4122 13288
rect 4066 13232 4122 13268
rect 2686 9596 2688 9616
rect 2688 9596 2740 9616
rect 2740 9596 2742 9616
rect 2686 9560 2742 9596
rect 3180 10362 3236 10364
rect 3260 10362 3316 10364
rect 3340 10362 3396 10364
rect 3420 10362 3476 10364
rect 3180 10310 3226 10362
rect 3226 10310 3236 10362
rect 3260 10310 3290 10362
rect 3290 10310 3302 10362
rect 3302 10310 3316 10362
rect 3340 10310 3354 10362
rect 3354 10310 3366 10362
rect 3366 10310 3396 10362
rect 3420 10310 3430 10362
rect 3430 10310 3476 10362
rect 3180 10308 3236 10310
rect 3260 10308 3316 10310
rect 3340 10308 3396 10310
rect 3420 10308 3476 10310
rect 3238 9696 3294 9752
rect 3180 9274 3236 9276
rect 3260 9274 3316 9276
rect 3340 9274 3396 9276
rect 3420 9274 3476 9276
rect 3180 9222 3226 9274
rect 3226 9222 3236 9274
rect 3260 9222 3290 9274
rect 3290 9222 3302 9274
rect 3302 9222 3316 9274
rect 3340 9222 3354 9274
rect 3354 9222 3366 9274
rect 3366 9222 3396 9274
rect 3420 9222 3430 9274
rect 3430 9222 3476 9274
rect 3180 9220 3236 9222
rect 3260 9220 3316 9222
rect 3340 9220 3396 9222
rect 3420 9220 3476 9222
rect 2870 8608 2926 8664
rect 2962 8336 3018 8392
rect 3180 8186 3236 8188
rect 3260 8186 3316 8188
rect 3340 8186 3396 8188
rect 3420 8186 3476 8188
rect 3180 8134 3226 8186
rect 3226 8134 3236 8186
rect 3260 8134 3290 8186
rect 3290 8134 3302 8186
rect 3302 8134 3316 8186
rect 3340 8134 3354 8186
rect 3354 8134 3366 8186
rect 3366 8134 3396 8186
rect 3420 8134 3430 8186
rect 3430 8134 3476 8186
rect 3180 8132 3236 8134
rect 3260 8132 3316 8134
rect 3340 8132 3396 8134
rect 3420 8132 3476 8134
rect 3180 7098 3236 7100
rect 3260 7098 3316 7100
rect 3340 7098 3396 7100
rect 3420 7098 3476 7100
rect 3180 7046 3226 7098
rect 3226 7046 3236 7098
rect 3260 7046 3290 7098
rect 3290 7046 3302 7098
rect 3302 7046 3316 7098
rect 3340 7046 3354 7098
rect 3354 7046 3366 7098
rect 3366 7046 3396 7098
rect 3420 7046 3430 7098
rect 3430 7046 3476 7098
rect 3180 7044 3236 7046
rect 3260 7044 3316 7046
rect 3340 7044 3396 7046
rect 3420 7044 3476 7046
rect 3330 6568 3386 6624
rect 3146 6296 3202 6352
rect 2410 5228 2466 5264
rect 2410 5208 2412 5228
rect 2412 5208 2464 5228
rect 2464 5208 2466 5228
rect 2318 4564 2320 4584
rect 2320 4564 2372 4584
rect 2372 4564 2374 4584
rect 2318 4528 2374 4564
rect 3180 6010 3236 6012
rect 3260 6010 3316 6012
rect 3340 6010 3396 6012
rect 3420 6010 3476 6012
rect 3180 5958 3226 6010
rect 3226 5958 3236 6010
rect 3260 5958 3290 6010
rect 3290 5958 3302 6010
rect 3302 5958 3316 6010
rect 3340 5958 3354 6010
rect 3354 5958 3366 6010
rect 3366 5958 3396 6010
rect 3420 5958 3430 6010
rect 3430 5958 3476 6010
rect 3180 5956 3236 5958
rect 3260 5956 3316 5958
rect 3340 5956 3396 5958
rect 3420 5956 3476 5958
rect 3238 5480 3294 5536
rect 3514 5208 3570 5264
rect 3180 4922 3236 4924
rect 3260 4922 3316 4924
rect 3340 4922 3396 4924
rect 3420 4922 3476 4924
rect 3180 4870 3226 4922
rect 3226 4870 3236 4922
rect 3260 4870 3290 4922
rect 3290 4870 3302 4922
rect 3302 4870 3316 4922
rect 3340 4870 3354 4922
rect 3354 4870 3366 4922
rect 3366 4870 3396 4922
rect 3420 4870 3430 4922
rect 3430 4870 3476 4922
rect 3180 4868 3236 4870
rect 3260 4868 3316 4870
rect 3340 4868 3396 4870
rect 3420 4868 3476 4870
rect 2778 4004 2834 4040
rect 2778 3984 2780 4004
rect 2780 3984 2832 4004
rect 2832 3984 2834 4004
rect 1858 2352 1914 2408
rect 2226 856 2282 912
rect 2686 1536 2742 1592
rect 3180 3834 3236 3836
rect 3260 3834 3316 3836
rect 3340 3834 3396 3836
rect 3420 3834 3476 3836
rect 3180 3782 3226 3834
rect 3226 3782 3236 3834
rect 3260 3782 3290 3834
rect 3290 3782 3302 3834
rect 3302 3782 3316 3834
rect 3340 3782 3354 3834
rect 3354 3782 3366 3834
rect 3366 3782 3396 3834
rect 3420 3782 3430 3834
rect 3430 3782 3476 3834
rect 3180 3780 3236 3782
rect 3260 3780 3316 3782
rect 3340 3780 3396 3782
rect 3420 3780 3476 3782
rect 3790 6704 3846 6760
rect 5404 14170 5460 14172
rect 5484 14170 5540 14172
rect 5564 14170 5620 14172
rect 5644 14170 5700 14172
rect 5404 14118 5450 14170
rect 5450 14118 5460 14170
rect 5484 14118 5514 14170
rect 5514 14118 5526 14170
rect 5526 14118 5540 14170
rect 5564 14118 5578 14170
rect 5578 14118 5590 14170
rect 5590 14118 5620 14170
rect 5644 14118 5654 14170
rect 5654 14118 5700 14170
rect 5404 14116 5460 14118
rect 5484 14116 5540 14118
rect 5564 14116 5620 14118
rect 5644 14116 5700 14118
rect 5538 13932 5594 13968
rect 5538 13912 5540 13932
rect 5540 13912 5592 13932
rect 5592 13912 5594 13932
rect 5998 13640 6054 13696
rect 5404 13082 5460 13084
rect 5484 13082 5540 13084
rect 5564 13082 5620 13084
rect 5644 13082 5700 13084
rect 5404 13030 5450 13082
rect 5450 13030 5460 13082
rect 5484 13030 5514 13082
rect 5514 13030 5526 13082
rect 5526 13030 5540 13082
rect 5564 13030 5578 13082
rect 5578 13030 5590 13082
rect 5590 13030 5620 13082
rect 5644 13030 5654 13082
rect 5654 13030 5700 13082
rect 5404 13028 5460 13030
rect 5484 13028 5540 13030
rect 5564 13028 5620 13030
rect 5644 13028 5700 13030
rect 4250 8336 4306 8392
rect 4066 6568 4122 6624
rect 3974 6432 4030 6488
rect 4158 6296 4214 6352
rect 3790 4664 3846 4720
rect 3882 3984 3938 4040
rect 4526 5616 4582 5672
rect 4250 4564 4252 4584
rect 4252 4564 4304 4584
rect 4304 4564 4306 4584
rect 4250 4528 4306 4564
rect 4066 4120 4122 4176
rect 5354 12860 5356 12880
rect 5356 12860 5408 12880
rect 5408 12860 5410 12880
rect 5354 12824 5410 12860
rect 4986 9424 5042 9480
rect 5404 11994 5460 11996
rect 5484 11994 5540 11996
rect 5564 11994 5620 11996
rect 5644 11994 5700 11996
rect 5404 11942 5450 11994
rect 5450 11942 5460 11994
rect 5484 11942 5514 11994
rect 5514 11942 5526 11994
rect 5526 11942 5540 11994
rect 5564 11942 5578 11994
rect 5578 11942 5590 11994
rect 5590 11942 5620 11994
rect 5644 11942 5654 11994
rect 5654 11942 5700 11994
rect 5404 11940 5460 11942
rect 5484 11940 5540 11942
rect 5564 11940 5620 11942
rect 5644 11940 5700 11942
rect 5404 10906 5460 10908
rect 5484 10906 5540 10908
rect 5564 10906 5620 10908
rect 5644 10906 5700 10908
rect 5404 10854 5450 10906
rect 5450 10854 5460 10906
rect 5484 10854 5514 10906
rect 5514 10854 5526 10906
rect 5526 10854 5540 10906
rect 5564 10854 5578 10906
rect 5578 10854 5590 10906
rect 5590 10854 5620 10906
rect 5644 10854 5654 10906
rect 5654 10854 5700 10906
rect 5404 10852 5460 10854
rect 5484 10852 5540 10854
rect 5564 10852 5620 10854
rect 5644 10852 5700 10854
rect 3790 3576 3846 3632
rect 3698 2896 3754 2952
rect 3180 2746 3236 2748
rect 3260 2746 3316 2748
rect 3340 2746 3396 2748
rect 3420 2746 3476 2748
rect 3180 2694 3226 2746
rect 3226 2694 3236 2746
rect 3260 2694 3290 2746
rect 3290 2694 3302 2746
rect 3302 2694 3316 2746
rect 3340 2694 3354 2746
rect 3354 2694 3366 2746
rect 3366 2694 3396 2746
rect 3420 2694 3430 2746
rect 3430 2694 3476 2746
rect 3180 2692 3236 2694
rect 3260 2692 3316 2694
rect 3340 2692 3396 2694
rect 3420 2692 3476 2694
rect 2870 1128 2926 1184
rect 3514 1944 3570 2000
rect 5404 9818 5460 9820
rect 5484 9818 5540 9820
rect 5564 9818 5620 9820
rect 5644 9818 5700 9820
rect 5404 9766 5450 9818
rect 5450 9766 5460 9818
rect 5484 9766 5514 9818
rect 5514 9766 5526 9818
rect 5526 9766 5540 9818
rect 5564 9766 5578 9818
rect 5578 9766 5590 9818
rect 5590 9766 5620 9818
rect 5644 9766 5654 9818
rect 5654 9766 5700 9818
rect 5404 9764 5460 9766
rect 5484 9764 5540 9766
rect 5564 9764 5620 9766
rect 5644 9764 5700 9766
rect 5404 8730 5460 8732
rect 5484 8730 5540 8732
rect 5564 8730 5620 8732
rect 5644 8730 5700 8732
rect 5404 8678 5450 8730
rect 5450 8678 5460 8730
rect 5484 8678 5514 8730
rect 5514 8678 5526 8730
rect 5526 8678 5540 8730
rect 5564 8678 5578 8730
rect 5578 8678 5590 8730
rect 5590 8678 5620 8730
rect 5644 8678 5654 8730
rect 5654 8678 5700 8730
rect 5404 8676 5460 8678
rect 5484 8676 5540 8678
rect 5564 8676 5620 8678
rect 5644 8676 5700 8678
rect 5404 7642 5460 7644
rect 5484 7642 5540 7644
rect 5564 7642 5620 7644
rect 5644 7642 5700 7644
rect 5404 7590 5450 7642
rect 5450 7590 5460 7642
rect 5484 7590 5514 7642
rect 5514 7590 5526 7642
rect 5526 7590 5540 7642
rect 5564 7590 5578 7642
rect 5578 7590 5590 7642
rect 5590 7590 5620 7642
rect 5644 7590 5654 7642
rect 5654 7590 5700 7642
rect 5404 7588 5460 7590
rect 5484 7588 5540 7590
rect 5564 7588 5620 7590
rect 5644 7588 5700 7590
rect 5404 6554 5460 6556
rect 5484 6554 5540 6556
rect 5564 6554 5620 6556
rect 5644 6554 5700 6556
rect 5404 6502 5450 6554
rect 5450 6502 5460 6554
rect 5484 6502 5514 6554
rect 5514 6502 5526 6554
rect 5526 6502 5540 6554
rect 5564 6502 5578 6554
rect 5578 6502 5590 6554
rect 5590 6502 5620 6554
rect 5644 6502 5654 6554
rect 5654 6502 5700 6554
rect 5404 6500 5460 6502
rect 5484 6500 5540 6502
rect 5564 6500 5620 6502
rect 5644 6500 5700 6502
rect 6090 8336 6146 8392
rect 5404 5466 5460 5468
rect 5484 5466 5540 5468
rect 5564 5466 5620 5468
rect 5644 5466 5700 5468
rect 5404 5414 5450 5466
rect 5450 5414 5460 5466
rect 5484 5414 5514 5466
rect 5514 5414 5526 5466
rect 5526 5414 5540 5466
rect 5564 5414 5578 5466
rect 5578 5414 5590 5466
rect 5590 5414 5620 5466
rect 5644 5414 5654 5466
rect 5654 5414 5700 5466
rect 5404 5412 5460 5414
rect 5484 5412 5540 5414
rect 5564 5412 5620 5414
rect 5644 5412 5700 5414
rect 5998 5752 6054 5808
rect 5404 4378 5460 4380
rect 5484 4378 5540 4380
rect 5564 4378 5620 4380
rect 5644 4378 5700 4380
rect 5404 4326 5450 4378
rect 5450 4326 5460 4378
rect 5484 4326 5514 4378
rect 5514 4326 5526 4378
rect 5526 4326 5540 4378
rect 5564 4326 5578 4378
rect 5578 4326 5590 4378
rect 5590 4326 5620 4378
rect 5644 4326 5654 4378
rect 5654 4326 5700 4378
rect 5404 4324 5460 4326
rect 5484 4324 5540 4326
rect 5564 4324 5620 4326
rect 5644 4324 5700 4326
rect 6274 5636 6330 5672
rect 6274 5616 6276 5636
rect 6276 5616 6328 5636
rect 6328 5616 6330 5636
rect 5404 3290 5460 3292
rect 5484 3290 5540 3292
rect 5564 3290 5620 3292
rect 5644 3290 5700 3292
rect 5404 3238 5450 3290
rect 5450 3238 5460 3290
rect 5484 3238 5514 3290
rect 5514 3238 5526 3290
rect 5526 3238 5540 3290
rect 5564 3238 5578 3290
rect 5578 3238 5590 3290
rect 5590 3238 5620 3290
rect 5644 3238 5654 3290
rect 5654 3238 5700 3290
rect 5404 3236 5460 3238
rect 5484 3236 5540 3238
rect 5564 3236 5620 3238
rect 5644 3236 5700 3238
rect 6734 13796 6790 13832
rect 6734 13776 6736 13796
rect 6736 13776 6788 13796
rect 6788 13776 6790 13796
rect 7628 14714 7684 14716
rect 7708 14714 7764 14716
rect 7788 14714 7844 14716
rect 7868 14714 7924 14716
rect 7628 14662 7674 14714
rect 7674 14662 7684 14714
rect 7708 14662 7738 14714
rect 7738 14662 7750 14714
rect 7750 14662 7764 14714
rect 7788 14662 7802 14714
rect 7802 14662 7814 14714
rect 7814 14662 7844 14714
rect 7868 14662 7878 14714
rect 7878 14662 7924 14714
rect 7628 14660 7684 14662
rect 7708 14660 7764 14662
rect 7788 14660 7844 14662
rect 7868 14660 7924 14662
rect 7838 13912 7894 13968
rect 7628 13626 7684 13628
rect 7708 13626 7764 13628
rect 7788 13626 7844 13628
rect 7868 13626 7924 13628
rect 7628 13574 7674 13626
rect 7674 13574 7684 13626
rect 7708 13574 7738 13626
rect 7738 13574 7750 13626
rect 7750 13574 7764 13626
rect 7788 13574 7802 13626
rect 7802 13574 7814 13626
rect 7814 13574 7844 13626
rect 7868 13574 7878 13626
rect 7878 13574 7924 13626
rect 7628 13572 7684 13574
rect 7708 13572 7764 13574
rect 7788 13572 7844 13574
rect 7868 13572 7924 13574
rect 6458 12008 6514 12064
rect 7628 12538 7684 12540
rect 7708 12538 7764 12540
rect 7788 12538 7844 12540
rect 7868 12538 7924 12540
rect 7628 12486 7674 12538
rect 7674 12486 7684 12538
rect 7708 12486 7738 12538
rect 7738 12486 7750 12538
rect 7750 12486 7764 12538
rect 7788 12486 7802 12538
rect 7802 12486 7814 12538
rect 7814 12486 7844 12538
rect 7868 12486 7878 12538
rect 7878 12486 7924 12538
rect 7628 12484 7684 12486
rect 7708 12484 7764 12486
rect 7788 12484 7844 12486
rect 7868 12484 7924 12486
rect 6642 7248 6698 7304
rect 6550 6160 6606 6216
rect 7628 11450 7684 11452
rect 7708 11450 7764 11452
rect 7788 11450 7844 11452
rect 7868 11450 7924 11452
rect 7628 11398 7674 11450
rect 7674 11398 7684 11450
rect 7708 11398 7738 11450
rect 7738 11398 7750 11450
rect 7750 11398 7764 11450
rect 7788 11398 7802 11450
rect 7802 11398 7814 11450
rect 7814 11398 7844 11450
rect 7868 11398 7878 11450
rect 7878 11398 7924 11450
rect 7628 11396 7684 11398
rect 7708 11396 7764 11398
rect 7788 11396 7844 11398
rect 7868 11396 7924 11398
rect 7628 10362 7684 10364
rect 7708 10362 7764 10364
rect 7788 10362 7844 10364
rect 7868 10362 7924 10364
rect 7628 10310 7674 10362
rect 7674 10310 7684 10362
rect 7708 10310 7738 10362
rect 7738 10310 7750 10362
rect 7750 10310 7764 10362
rect 7788 10310 7802 10362
rect 7802 10310 7814 10362
rect 7814 10310 7844 10362
rect 7868 10310 7878 10362
rect 7878 10310 7924 10362
rect 7628 10308 7684 10310
rect 7708 10308 7764 10310
rect 7788 10308 7844 10310
rect 7868 10308 7924 10310
rect 7286 6840 7342 6896
rect 6642 3440 6698 3496
rect 6550 2624 6606 2680
rect 7628 9274 7684 9276
rect 7708 9274 7764 9276
rect 7788 9274 7844 9276
rect 7868 9274 7924 9276
rect 7628 9222 7674 9274
rect 7674 9222 7684 9274
rect 7708 9222 7738 9274
rect 7738 9222 7750 9274
rect 7750 9222 7764 9274
rect 7788 9222 7802 9274
rect 7802 9222 7814 9274
rect 7814 9222 7844 9274
rect 7868 9222 7878 9274
rect 7878 9222 7924 9274
rect 7628 9220 7684 9222
rect 7708 9220 7764 9222
rect 7788 9220 7844 9222
rect 7868 9220 7924 9222
rect 7628 8186 7684 8188
rect 7708 8186 7764 8188
rect 7788 8186 7844 8188
rect 7868 8186 7924 8188
rect 7628 8134 7674 8186
rect 7674 8134 7684 8186
rect 7708 8134 7738 8186
rect 7738 8134 7750 8186
rect 7750 8134 7764 8186
rect 7788 8134 7802 8186
rect 7802 8134 7814 8186
rect 7814 8134 7844 8186
rect 7868 8134 7878 8186
rect 7878 8134 7924 8186
rect 7628 8132 7684 8134
rect 7708 8132 7764 8134
rect 7788 8132 7844 8134
rect 7868 8132 7924 8134
rect 7628 7098 7684 7100
rect 7708 7098 7764 7100
rect 7788 7098 7844 7100
rect 7868 7098 7924 7100
rect 7628 7046 7674 7098
rect 7674 7046 7684 7098
rect 7708 7046 7738 7098
rect 7738 7046 7750 7098
rect 7750 7046 7764 7098
rect 7788 7046 7802 7098
rect 7802 7046 7814 7098
rect 7814 7046 7844 7098
rect 7868 7046 7878 7098
rect 7878 7046 7924 7098
rect 7628 7044 7684 7046
rect 7708 7044 7764 7046
rect 7788 7044 7844 7046
rect 7868 7044 7924 7046
rect 7628 6010 7684 6012
rect 7708 6010 7764 6012
rect 7788 6010 7844 6012
rect 7868 6010 7924 6012
rect 7628 5958 7674 6010
rect 7674 5958 7684 6010
rect 7708 5958 7738 6010
rect 7738 5958 7750 6010
rect 7750 5958 7764 6010
rect 7788 5958 7802 6010
rect 7802 5958 7814 6010
rect 7814 5958 7844 6010
rect 7868 5958 7878 6010
rect 7878 5958 7924 6010
rect 7628 5956 7684 5958
rect 7708 5956 7764 5958
rect 7788 5956 7844 5958
rect 7868 5956 7924 5958
rect 7628 4922 7684 4924
rect 7708 4922 7764 4924
rect 7788 4922 7844 4924
rect 7868 4922 7924 4924
rect 7628 4870 7674 4922
rect 7674 4870 7684 4922
rect 7708 4870 7738 4922
rect 7738 4870 7750 4922
rect 7750 4870 7764 4922
rect 7788 4870 7802 4922
rect 7802 4870 7814 4922
rect 7814 4870 7844 4922
rect 7868 4870 7878 4922
rect 7878 4870 7924 4922
rect 7628 4868 7684 4870
rect 7708 4868 7764 4870
rect 7788 4868 7844 4870
rect 7868 4868 7924 4870
rect 7470 4564 7472 4584
rect 7472 4564 7524 4584
rect 7524 4564 7526 4584
rect 7470 4528 7526 4564
rect 7628 3834 7684 3836
rect 7708 3834 7764 3836
rect 7788 3834 7844 3836
rect 7868 3834 7924 3836
rect 7628 3782 7674 3834
rect 7674 3782 7684 3834
rect 7708 3782 7738 3834
rect 7738 3782 7750 3834
rect 7750 3782 7764 3834
rect 7788 3782 7802 3834
rect 7802 3782 7814 3834
rect 7814 3782 7844 3834
rect 7868 3782 7878 3834
rect 7878 3782 7924 3834
rect 7628 3780 7684 3782
rect 7708 3780 7764 3782
rect 7788 3780 7844 3782
rect 7868 3780 7924 3782
rect 8482 12280 8538 12336
rect 8390 7384 8446 7440
rect 8206 3984 8262 4040
rect 8758 13776 8814 13832
rect 8850 12280 8906 12336
rect 8850 12008 8906 12064
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9898 14170
rect 9898 14118 9908 14170
rect 9932 14118 9962 14170
rect 9962 14118 9974 14170
rect 9974 14118 9988 14170
rect 10012 14118 10026 14170
rect 10026 14118 10038 14170
rect 10038 14118 10068 14170
rect 10092 14118 10102 14170
rect 10102 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 9862 13368 9918 13424
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9898 13082
rect 9898 13030 9908 13082
rect 9932 13030 9962 13082
rect 9962 13030 9974 13082
rect 9974 13030 9988 13082
rect 10012 13030 10026 13082
rect 10026 13030 10038 13082
rect 10038 13030 10068 13082
rect 10092 13030 10102 13082
rect 10102 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 9494 12824 9550 12880
rect 7628 2746 7684 2748
rect 7708 2746 7764 2748
rect 7788 2746 7844 2748
rect 7868 2746 7924 2748
rect 7628 2694 7674 2746
rect 7674 2694 7684 2746
rect 7708 2694 7738 2746
rect 7738 2694 7750 2746
rect 7750 2694 7764 2746
rect 7788 2694 7802 2746
rect 7802 2694 7814 2746
rect 7814 2694 7844 2746
rect 7868 2694 7878 2746
rect 7878 2694 7924 2746
rect 7628 2692 7684 2694
rect 7708 2692 7764 2694
rect 7788 2692 7844 2694
rect 7868 2692 7924 2694
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9898 11994
rect 9898 11942 9908 11994
rect 9932 11942 9962 11994
rect 9962 11942 9974 11994
rect 9974 11942 9988 11994
rect 10012 11942 10026 11994
rect 10026 11942 10038 11994
rect 10038 11942 10068 11994
rect 10092 11942 10102 11994
rect 10102 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 10046 11192 10102 11248
rect 9770 11056 9826 11112
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9898 10906
rect 9898 10854 9908 10906
rect 9932 10854 9962 10906
rect 9962 10854 9974 10906
rect 9974 10854 9988 10906
rect 10012 10854 10026 10906
rect 10026 10854 10038 10906
rect 10038 10854 10068 10906
rect 10092 10854 10102 10906
rect 10102 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9898 9818
rect 9898 9766 9908 9818
rect 9932 9766 9962 9818
rect 9962 9766 9974 9818
rect 9974 9766 9988 9818
rect 10012 9766 10026 9818
rect 10026 9766 10038 9818
rect 10038 9766 10068 9818
rect 10092 9766 10102 9818
rect 10102 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9898 8730
rect 9898 8678 9908 8730
rect 9932 8678 9962 8730
rect 9962 8678 9974 8730
rect 9974 8678 9988 8730
rect 10012 8678 10026 8730
rect 10026 8678 10038 8730
rect 10038 8678 10068 8730
rect 10092 8678 10102 8730
rect 10102 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9898 7642
rect 9898 7590 9908 7642
rect 9932 7590 9962 7642
rect 9962 7590 9974 7642
rect 9974 7590 9988 7642
rect 10012 7590 10026 7642
rect 10026 7590 10038 7642
rect 10038 7590 10068 7642
rect 10092 7590 10102 7642
rect 10102 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9898 6554
rect 9898 6502 9908 6554
rect 9932 6502 9962 6554
rect 9962 6502 9974 6554
rect 9974 6502 9988 6554
rect 10012 6502 10026 6554
rect 10026 6502 10038 6554
rect 10038 6502 10068 6554
rect 10092 6502 10102 6554
rect 10102 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9898 5466
rect 9898 5414 9908 5466
rect 9932 5414 9962 5466
rect 9962 5414 9974 5466
rect 9974 5414 9988 5466
rect 10012 5414 10026 5466
rect 10026 5414 10038 5466
rect 10038 5414 10068 5466
rect 10092 5414 10102 5466
rect 10102 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 10046 4800 10102 4856
rect 10138 4664 10194 4720
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9898 4378
rect 9898 4326 9908 4378
rect 9932 4326 9962 4378
rect 9962 4326 9974 4378
rect 9974 4326 9988 4378
rect 10012 4326 10026 4378
rect 10026 4326 10038 4378
rect 10038 4326 10068 4378
rect 10092 4326 10102 4378
rect 10102 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 10230 3576 10286 3632
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9898 3290
rect 9898 3238 9908 3290
rect 9932 3238 9962 3290
rect 9962 3238 9974 3290
rect 9974 3238 9988 3290
rect 10012 3238 10026 3290
rect 10026 3238 10038 3290
rect 10038 3238 10068 3290
rect 10092 3238 10102 3290
rect 10102 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 10322 3032 10378 3088
rect 10874 11192 10930 11248
rect 12076 14714 12132 14716
rect 12156 14714 12212 14716
rect 12236 14714 12292 14716
rect 12316 14714 12372 14716
rect 12076 14662 12122 14714
rect 12122 14662 12132 14714
rect 12156 14662 12186 14714
rect 12186 14662 12198 14714
rect 12198 14662 12212 14714
rect 12236 14662 12250 14714
rect 12250 14662 12262 14714
rect 12262 14662 12292 14714
rect 12316 14662 12326 14714
rect 12326 14662 12372 14714
rect 12076 14660 12132 14662
rect 12156 14660 12212 14662
rect 12236 14660 12292 14662
rect 12316 14660 12372 14662
rect 11150 13232 11206 13288
rect 11242 11092 11244 11112
rect 11244 11092 11296 11112
rect 11296 11092 11298 11112
rect 11242 11056 11298 11092
rect 10874 3984 10930 4040
rect 11610 7792 11666 7848
rect 11886 13640 11942 13696
rect 12076 13626 12132 13628
rect 12156 13626 12212 13628
rect 12236 13626 12292 13628
rect 12316 13626 12372 13628
rect 12076 13574 12122 13626
rect 12122 13574 12132 13626
rect 12156 13574 12186 13626
rect 12186 13574 12198 13626
rect 12198 13574 12212 13626
rect 12236 13574 12250 13626
rect 12250 13574 12262 13626
rect 12262 13574 12292 13626
rect 12316 13574 12326 13626
rect 12326 13574 12372 13626
rect 12076 13572 12132 13574
rect 12156 13572 12212 13574
rect 12236 13572 12292 13574
rect 12316 13572 12372 13574
rect 12076 12538 12132 12540
rect 12156 12538 12212 12540
rect 12236 12538 12292 12540
rect 12316 12538 12372 12540
rect 12076 12486 12122 12538
rect 12122 12486 12132 12538
rect 12156 12486 12186 12538
rect 12186 12486 12198 12538
rect 12198 12486 12212 12538
rect 12236 12486 12250 12538
rect 12250 12486 12262 12538
rect 12262 12486 12292 12538
rect 12316 12486 12326 12538
rect 12326 12486 12372 12538
rect 12076 12484 12132 12486
rect 12156 12484 12212 12486
rect 12236 12484 12292 12486
rect 12316 12484 12372 12486
rect 13266 14456 13322 14512
rect 12076 11450 12132 11452
rect 12156 11450 12212 11452
rect 12236 11450 12292 11452
rect 12316 11450 12372 11452
rect 12076 11398 12122 11450
rect 12122 11398 12132 11450
rect 12156 11398 12186 11450
rect 12186 11398 12198 11450
rect 12198 11398 12212 11450
rect 12236 11398 12250 11450
rect 12250 11398 12262 11450
rect 12262 11398 12292 11450
rect 12316 11398 12326 11450
rect 12326 11398 12372 11450
rect 12076 11396 12132 11398
rect 12156 11396 12212 11398
rect 12236 11396 12292 11398
rect 12316 11396 12372 11398
rect 12076 10362 12132 10364
rect 12156 10362 12212 10364
rect 12236 10362 12292 10364
rect 12316 10362 12372 10364
rect 12076 10310 12122 10362
rect 12122 10310 12132 10362
rect 12156 10310 12186 10362
rect 12186 10310 12198 10362
rect 12198 10310 12212 10362
rect 12236 10310 12250 10362
rect 12250 10310 12262 10362
rect 12262 10310 12292 10362
rect 12316 10310 12326 10362
rect 12326 10310 12372 10362
rect 12076 10308 12132 10310
rect 12156 10308 12212 10310
rect 12236 10308 12292 10310
rect 12316 10308 12372 10310
rect 12076 9274 12132 9276
rect 12156 9274 12212 9276
rect 12236 9274 12292 9276
rect 12316 9274 12372 9276
rect 12076 9222 12122 9274
rect 12122 9222 12132 9274
rect 12156 9222 12186 9274
rect 12186 9222 12198 9274
rect 12198 9222 12212 9274
rect 12236 9222 12250 9274
rect 12250 9222 12262 9274
rect 12262 9222 12292 9274
rect 12316 9222 12326 9274
rect 12326 9222 12372 9274
rect 12076 9220 12132 9222
rect 12156 9220 12212 9222
rect 12236 9220 12292 9222
rect 12316 9220 12372 9222
rect 12076 8186 12132 8188
rect 12156 8186 12212 8188
rect 12236 8186 12292 8188
rect 12316 8186 12372 8188
rect 12076 8134 12122 8186
rect 12122 8134 12132 8186
rect 12156 8134 12186 8186
rect 12186 8134 12198 8186
rect 12198 8134 12212 8186
rect 12236 8134 12250 8186
rect 12250 8134 12262 8186
rect 12262 8134 12292 8186
rect 12316 8134 12326 8186
rect 12326 8134 12372 8186
rect 12076 8132 12132 8134
rect 12156 8132 12212 8134
rect 12236 8132 12292 8134
rect 12316 8132 12372 8134
rect 12076 7098 12132 7100
rect 12156 7098 12212 7100
rect 12236 7098 12292 7100
rect 12316 7098 12372 7100
rect 12076 7046 12122 7098
rect 12122 7046 12132 7098
rect 12156 7046 12186 7098
rect 12186 7046 12198 7098
rect 12198 7046 12212 7098
rect 12236 7046 12250 7098
rect 12250 7046 12262 7098
rect 12262 7046 12292 7098
rect 12316 7046 12326 7098
rect 12326 7046 12372 7098
rect 12076 7044 12132 7046
rect 12156 7044 12212 7046
rect 12236 7044 12292 7046
rect 12316 7044 12372 7046
rect 12076 6010 12132 6012
rect 12156 6010 12212 6012
rect 12236 6010 12292 6012
rect 12316 6010 12372 6012
rect 12076 5958 12122 6010
rect 12122 5958 12132 6010
rect 12156 5958 12186 6010
rect 12186 5958 12198 6010
rect 12198 5958 12212 6010
rect 12236 5958 12250 6010
rect 12250 5958 12262 6010
rect 12262 5958 12292 6010
rect 12316 5958 12326 6010
rect 12326 5958 12372 6010
rect 12076 5956 12132 5958
rect 12156 5956 12212 5958
rect 12236 5956 12292 5958
rect 12316 5956 12372 5958
rect 12162 5108 12164 5128
rect 12164 5108 12216 5128
rect 12216 5108 12218 5128
rect 12162 5072 12218 5108
rect 12076 4922 12132 4924
rect 12156 4922 12212 4924
rect 12236 4922 12292 4924
rect 12316 4922 12372 4924
rect 12076 4870 12122 4922
rect 12122 4870 12132 4922
rect 12156 4870 12186 4922
rect 12186 4870 12198 4922
rect 12198 4870 12212 4922
rect 12236 4870 12250 4922
rect 12250 4870 12262 4922
rect 12262 4870 12292 4922
rect 12316 4870 12326 4922
rect 12326 4870 12372 4922
rect 12076 4868 12132 4870
rect 12156 4868 12212 4870
rect 12236 4868 12292 4870
rect 12316 4868 12372 4870
rect 11886 4800 11942 4856
rect 12714 12280 12770 12336
rect 13266 11756 13322 11792
rect 13266 11736 13268 11756
rect 13268 11736 13320 11756
rect 13320 11736 13322 11756
rect 13174 11600 13230 11656
rect 12714 4820 12770 4856
rect 12714 4800 12716 4820
rect 12716 4800 12768 4820
rect 12768 4800 12770 4820
rect 12076 3834 12132 3836
rect 12156 3834 12212 3836
rect 12236 3834 12292 3836
rect 12316 3834 12372 3836
rect 12076 3782 12122 3834
rect 12122 3782 12132 3834
rect 12156 3782 12186 3834
rect 12186 3782 12198 3834
rect 12198 3782 12212 3834
rect 12236 3782 12250 3834
rect 12250 3782 12262 3834
rect 12262 3782 12292 3834
rect 12316 3782 12326 3834
rect 12326 3782 12372 3834
rect 12076 3780 12132 3782
rect 12156 3780 12212 3782
rect 12236 3780 12292 3782
rect 12316 3780 12372 3782
rect 11702 3440 11758 3496
rect 5404 2202 5460 2204
rect 5484 2202 5540 2204
rect 5564 2202 5620 2204
rect 5644 2202 5700 2204
rect 5404 2150 5450 2202
rect 5450 2150 5460 2202
rect 5484 2150 5514 2202
rect 5514 2150 5526 2202
rect 5526 2150 5540 2202
rect 5564 2150 5578 2202
rect 5578 2150 5590 2202
rect 5590 2150 5620 2202
rect 5644 2150 5654 2202
rect 5654 2150 5700 2202
rect 5404 2148 5460 2150
rect 5484 2148 5540 2150
rect 5564 2148 5620 2150
rect 5644 2148 5700 2150
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9898 2202
rect 9898 2150 9908 2202
rect 9932 2150 9962 2202
rect 9962 2150 9974 2202
rect 9974 2150 9988 2202
rect 10012 2150 10026 2202
rect 10026 2150 10038 2202
rect 10038 2150 10068 2202
rect 10092 2150 10102 2202
rect 10102 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 12076 2746 12132 2748
rect 12156 2746 12212 2748
rect 12236 2746 12292 2748
rect 12316 2746 12372 2748
rect 12076 2694 12122 2746
rect 12122 2694 12132 2746
rect 12156 2694 12186 2746
rect 12186 2694 12198 2746
rect 12198 2694 12212 2746
rect 12236 2694 12250 2746
rect 12250 2694 12262 2746
rect 12262 2694 12292 2746
rect 12316 2694 12326 2746
rect 12326 2694 12372 2746
rect 12076 2692 12132 2694
rect 12156 2692 12212 2694
rect 12236 2692 12292 2694
rect 12316 2692 12372 2694
rect 3974 312 4030 368
rect 15474 16496 15530 16552
rect 14094 11464 14150 11520
rect 14300 14170 14356 14172
rect 14380 14170 14436 14172
rect 14460 14170 14516 14172
rect 14540 14170 14596 14172
rect 14300 14118 14346 14170
rect 14346 14118 14356 14170
rect 14380 14118 14410 14170
rect 14410 14118 14422 14170
rect 14422 14118 14436 14170
rect 14460 14118 14474 14170
rect 14474 14118 14486 14170
rect 14486 14118 14516 14170
rect 14540 14118 14550 14170
rect 14550 14118 14596 14170
rect 14300 14116 14356 14118
rect 14380 14116 14436 14118
rect 14460 14116 14516 14118
rect 14540 14116 14596 14118
rect 14300 13082 14356 13084
rect 14380 13082 14436 13084
rect 14460 13082 14516 13084
rect 14540 13082 14596 13084
rect 14300 13030 14346 13082
rect 14346 13030 14356 13082
rect 14380 13030 14410 13082
rect 14410 13030 14422 13082
rect 14422 13030 14436 13082
rect 14460 13030 14474 13082
rect 14474 13030 14486 13082
rect 14486 13030 14516 13082
rect 14540 13030 14550 13082
rect 14550 13030 14596 13082
rect 14300 13028 14356 13030
rect 14380 13028 14436 13030
rect 14460 13028 14516 13030
rect 14540 13028 14596 13030
rect 14300 11994 14356 11996
rect 14380 11994 14436 11996
rect 14460 11994 14516 11996
rect 14540 11994 14596 11996
rect 14300 11942 14346 11994
rect 14346 11942 14356 11994
rect 14380 11942 14410 11994
rect 14410 11942 14422 11994
rect 14422 11942 14436 11994
rect 14460 11942 14474 11994
rect 14474 11942 14486 11994
rect 14486 11942 14516 11994
rect 14540 11942 14550 11994
rect 14550 11942 14596 11994
rect 14300 11940 14356 11942
rect 14380 11940 14436 11942
rect 14460 11940 14516 11942
rect 14540 11940 14596 11942
rect 14554 11500 14556 11520
rect 14556 11500 14608 11520
rect 14608 11500 14610 11520
rect 14554 11464 14610 11500
rect 14300 10906 14356 10908
rect 14380 10906 14436 10908
rect 14460 10906 14516 10908
rect 14540 10906 14596 10908
rect 14300 10854 14346 10906
rect 14346 10854 14356 10906
rect 14380 10854 14410 10906
rect 14410 10854 14422 10906
rect 14422 10854 14436 10906
rect 14460 10854 14474 10906
rect 14474 10854 14486 10906
rect 14486 10854 14516 10906
rect 14540 10854 14550 10906
rect 14550 10854 14596 10906
rect 14300 10852 14356 10854
rect 14380 10852 14436 10854
rect 14460 10852 14516 10854
rect 14540 10852 14596 10854
rect 14462 10668 14518 10704
rect 14462 10648 14464 10668
rect 14464 10648 14516 10668
rect 14516 10648 14518 10668
rect 14300 9818 14356 9820
rect 14380 9818 14436 9820
rect 14460 9818 14516 9820
rect 14540 9818 14596 9820
rect 14300 9766 14346 9818
rect 14346 9766 14356 9818
rect 14380 9766 14410 9818
rect 14410 9766 14422 9818
rect 14422 9766 14436 9818
rect 14460 9766 14474 9818
rect 14474 9766 14486 9818
rect 14486 9766 14516 9818
rect 14540 9766 14550 9818
rect 14550 9766 14596 9818
rect 14300 9764 14356 9766
rect 14380 9764 14436 9766
rect 14460 9764 14516 9766
rect 14540 9764 14596 9766
rect 14300 8730 14356 8732
rect 14380 8730 14436 8732
rect 14460 8730 14516 8732
rect 14540 8730 14596 8732
rect 14300 8678 14346 8730
rect 14346 8678 14356 8730
rect 14380 8678 14410 8730
rect 14410 8678 14422 8730
rect 14422 8678 14436 8730
rect 14460 8678 14474 8730
rect 14474 8678 14486 8730
rect 14486 8678 14516 8730
rect 14540 8678 14550 8730
rect 14550 8678 14596 8730
rect 14300 8676 14356 8678
rect 14380 8676 14436 8678
rect 14460 8676 14516 8678
rect 14540 8676 14596 8678
rect 14646 8472 14702 8528
rect 14300 7642 14356 7644
rect 14380 7642 14436 7644
rect 14460 7642 14516 7644
rect 14540 7642 14596 7644
rect 14300 7590 14346 7642
rect 14346 7590 14356 7642
rect 14380 7590 14410 7642
rect 14410 7590 14422 7642
rect 14422 7590 14436 7642
rect 14460 7590 14474 7642
rect 14474 7590 14486 7642
rect 14486 7590 14516 7642
rect 14540 7590 14550 7642
rect 14550 7590 14596 7642
rect 14300 7588 14356 7590
rect 14380 7588 14436 7590
rect 14460 7588 14516 7590
rect 14540 7588 14596 7590
rect 14300 6554 14356 6556
rect 14380 6554 14436 6556
rect 14460 6554 14516 6556
rect 14540 6554 14596 6556
rect 14300 6502 14346 6554
rect 14346 6502 14356 6554
rect 14380 6502 14410 6554
rect 14410 6502 14422 6554
rect 14422 6502 14436 6554
rect 14460 6502 14474 6554
rect 14474 6502 14486 6554
rect 14486 6502 14516 6554
rect 14540 6502 14550 6554
rect 14550 6502 14596 6554
rect 14300 6500 14356 6502
rect 14380 6500 14436 6502
rect 14460 6500 14516 6502
rect 14540 6500 14596 6502
rect 14094 5752 14150 5808
rect 14300 5466 14356 5468
rect 14380 5466 14436 5468
rect 14460 5466 14516 5468
rect 14540 5466 14596 5468
rect 14300 5414 14346 5466
rect 14346 5414 14356 5466
rect 14380 5414 14410 5466
rect 14410 5414 14422 5466
rect 14422 5414 14436 5466
rect 14460 5414 14474 5466
rect 14474 5414 14486 5466
rect 14486 5414 14516 5466
rect 14540 5414 14550 5466
rect 14550 5414 14596 5466
rect 14300 5412 14356 5414
rect 14380 5412 14436 5414
rect 14460 5412 14516 5414
rect 14540 5412 14596 5414
rect 14278 4800 14334 4856
rect 14002 4120 14058 4176
rect 14300 4378 14356 4380
rect 14380 4378 14436 4380
rect 14460 4378 14516 4380
rect 14540 4378 14596 4380
rect 14300 4326 14346 4378
rect 14346 4326 14356 4378
rect 14380 4326 14410 4378
rect 14410 4326 14422 4378
rect 14422 4326 14436 4378
rect 14460 4326 14474 4378
rect 14474 4326 14486 4378
rect 14486 4326 14516 4378
rect 14540 4326 14550 4378
rect 14550 4326 14596 4378
rect 14300 4324 14356 4326
rect 14380 4324 14436 4326
rect 14460 4324 14516 4326
rect 14540 4324 14596 4326
rect 14646 3984 14702 4040
rect 14300 3290 14356 3292
rect 14380 3290 14436 3292
rect 14460 3290 14516 3292
rect 14540 3290 14596 3292
rect 14300 3238 14346 3290
rect 14346 3238 14356 3290
rect 14380 3238 14410 3290
rect 14410 3238 14422 3290
rect 14422 3238 14436 3290
rect 14460 3238 14474 3290
rect 14474 3238 14486 3290
rect 14486 3238 14516 3290
rect 14540 3238 14550 3290
rect 14550 3238 14596 3290
rect 14300 3236 14356 3238
rect 14380 3236 14436 3238
rect 14460 3236 14516 3238
rect 14540 3236 14596 3238
rect 14370 3068 14372 3088
rect 14372 3068 14424 3088
rect 14424 3068 14426 3088
rect 14370 3032 14426 3068
rect 14300 2202 14356 2204
rect 14380 2202 14436 2204
rect 14460 2202 14516 2204
rect 14540 2202 14596 2204
rect 14300 2150 14346 2202
rect 14346 2150 14356 2202
rect 14380 2150 14410 2202
rect 14410 2150 14422 2202
rect 14422 2150 14436 2202
rect 14460 2150 14474 2202
rect 14474 2150 14486 2202
rect 14486 2150 14516 2202
rect 14540 2150 14550 2202
rect 14550 2150 14596 2202
rect 14300 2148 14356 2150
rect 14380 2148 14436 2150
rect 14460 2148 14516 2150
rect 14540 2148 14596 2150
rect 16302 16088 16358 16144
rect 16210 14864 16266 14920
rect 15382 12144 15438 12200
rect 15014 6704 15070 6760
rect 14922 5228 14978 5264
rect 14922 5208 14924 5228
rect 14924 5208 14976 5228
rect 14976 5208 14978 5228
rect 15014 5072 15070 5128
rect 15474 5228 15530 5264
rect 15474 5208 15476 5228
rect 15476 5208 15528 5228
rect 15528 5208 15530 5228
rect 15106 4664 15162 4720
rect 16854 15680 16910 15736
rect 16524 14714 16580 14716
rect 16604 14714 16660 14716
rect 16684 14714 16740 14716
rect 16764 14714 16820 14716
rect 16524 14662 16570 14714
rect 16570 14662 16580 14714
rect 16604 14662 16634 14714
rect 16634 14662 16646 14714
rect 16646 14662 16660 14714
rect 16684 14662 16698 14714
rect 16698 14662 16710 14714
rect 16710 14662 16740 14714
rect 16764 14662 16774 14714
rect 16774 14662 16820 14714
rect 16524 14660 16580 14662
rect 16604 14660 16660 14662
rect 16684 14660 16740 14662
rect 16764 14660 16820 14662
rect 16762 14476 16818 14512
rect 16762 14456 16764 14476
rect 16764 14456 16816 14476
rect 16816 14456 16818 14476
rect 17130 15272 17186 15328
rect 16486 14048 16542 14104
rect 16854 14048 16910 14104
rect 16524 13626 16580 13628
rect 16604 13626 16660 13628
rect 16684 13626 16740 13628
rect 16764 13626 16820 13628
rect 16524 13574 16570 13626
rect 16570 13574 16580 13626
rect 16604 13574 16634 13626
rect 16634 13574 16646 13626
rect 16646 13574 16660 13626
rect 16684 13574 16698 13626
rect 16698 13574 16710 13626
rect 16710 13574 16740 13626
rect 16764 13574 16774 13626
rect 16774 13574 16820 13626
rect 16524 13572 16580 13574
rect 16604 13572 16660 13574
rect 16684 13572 16740 13574
rect 16764 13572 16820 13574
rect 16302 12824 16358 12880
rect 16524 12538 16580 12540
rect 16604 12538 16660 12540
rect 16684 12538 16740 12540
rect 16764 12538 16820 12540
rect 16524 12486 16570 12538
rect 16570 12486 16580 12538
rect 16604 12486 16634 12538
rect 16634 12486 16646 12538
rect 16646 12486 16660 12538
rect 16684 12486 16698 12538
rect 16698 12486 16710 12538
rect 16710 12486 16740 12538
rect 16764 12486 16774 12538
rect 16774 12486 16820 12538
rect 16524 12484 16580 12486
rect 16604 12484 16660 12486
rect 16684 12484 16740 12486
rect 16764 12484 16820 12486
rect 16524 11450 16580 11452
rect 16604 11450 16660 11452
rect 16684 11450 16740 11452
rect 16764 11450 16820 11452
rect 16524 11398 16570 11450
rect 16570 11398 16580 11450
rect 16604 11398 16634 11450
rect 16634 11398 16646 11450
rect 16646 11398 16660 11450
rect 16684 11398 16698 11450
rect 16698 11398 16710 11450
rect 16710 11398 16740 11450
rect 16764 11398 16774 11450
rect 16774 11398 16820 11450
rect 16524 11396 16580 11398
rect 16604 11396 16660 11398
rect 16684 11396 16740 11398
rect 16764 11396 16820 11398
rect 16854 10648 16910 10704
rect 16524 10362 16580 10364
rect 16604 10362 16660 10364
rect 16684 10362 16740 10364
rect 16764 10362 16820 10364
rect 16524 10310 16570 10362
rect 16570 10310 16580 10362
rect 16604 10310 16634 10362
rect 16634 10310 16646 10362
rect 16646 10310 16660 10362
rect 16684 10310 16698 10362
rect 16698 10310 16710 10362
rect 16710 10310 16740 10362
rect 16764 10310 16774 10362
rect 16774 10310 16820 10362
rect 16524 10308 16580 10310
rect 16604 10308 16660 10310
rect 16684 10308 16740 10310
rect 16764 10308 16820 10310
rect 17682 13640 17738 13696
rect 17314 13232 17370 13288
rect 17590 12860 17592 12880
rect 17592 12860 17644 12880
rect 17644 12860 17646 12880
rect 17590 12824 17646 12860
rect 17406 11872 17462 11928
rect 17130 11600 17186 11656
rect 17038 11056 17094 11112
rect 17774 13232 17830 13288
rect 17682 12416 17738 12472
rect 17866 12280 17922 12336
rect 17774 12008 17830 12064
rect 17774 11872 17830 11928
rect 16524 9274 16580 9276
rect 16604 9274 16660 9276
rect 16684 9274 16740 9276
rect 16764 9274 16820 9276
rect 16524 9222 16570 9274
rect 16570 9222 16580 9274
rect 16604 9222 16634 9274
rect 16634 9222 16646 9274
rect 16646 9222 16660 9274
rect 16684 9222 16698 9274
rect 16698 9222 16710 9274
rect 16710 9222 16740 9274
rect 16764 9222 16774 9274
rect 16774 9222 16820 9274
rect 16524 9220 16580 9222
rect 16604 9220 16660 9222
rect 16684 9220 16740 9222
rect 16764 9220 16820 9222
rect 16524 8186 16580 8188
rect 16604 8186 16660 8188
rect 16684 8186 16740 8188
rect 16764 8186 16820 8188
rect 16524 8134 16570 8186
rect 16570 8134 16580 8186
rect 16604 8134 16634 8186
rect 16634 8134 16646 8186
rect 16646 8134 16660 8186
rect 16684 8134 16698 8186
rect 16698 8134 16710 8186
rect 16710 8134 16740 8186
rect 16764 8134 16774 8186
rect 16774 8134 16820 8186
rect 16524 8132 16580 8134
rect 16604 8132 16660 8134
rect 16684 8132 16740 8134
rect 16764 8132 16820 8134
rect 16394 7792 16450 7848
rect 16524 7098 16580 7100
rect 16604 7098 16660 7100
rect 16684 7098 16740 7100
rect 16764 7098 16820 7100
rect 16524 7046 16570 7098
rect 16570 7046 16580 7098
rect 16604 7046 16634 7098
rect 16634 7046 16646 7098
rect 16646 7046 16660 7098
rect 16684 7046 16698 7098
rect 16698 7046 16710 7098
rect 16710 7046 16740 7098
rect 16764 7046 16774 7098
rect 16774 7046 16820 7098
rect 16524 7044 16580 7046
rect 16604 7044 16660 7046
rect 16684 7044 16740 7046
rect 16764 7044 16820 7046
rect 17314 9424 17370 9480
rect 17406 9152 17462 9208
rect 16524 6010 16580 6012
rect 16604 6010 16660 6012
rect 16684 6010 16740 6012
rect 16764 6010 16820 6012
rect 16524 5958 16570 6010
rect 16570 5958 16580 6010
rect 16604 5958 16634 6010
rect 16634 5958 16646 6010
rect 16646 5958 16660 6010
rect 16684 5958 16698 6010
rect 16698 5958 16710 6010
rect 16710 5958 16740 6010
rect 16764 5958 16774 6010
rect 16774 5958 16820 6010
rect 16524 5956 16580 5958
rect 16604 5956 16660 5958
rect 16684 5956 16740 5958
rect 16764 5956 16820 5958
rect 16946 6196 16948 6216
rect 16948 6196 17000 6216
rect 17000 6196 17002 6216
rect 16946 6160 17002 6196
rect 16118 5208 16174 5264
rect 17314 5772 17370 5808
rect 17314 5752 17316 5772
rect 17316 5752 17368 5772
rect 17368 5752 17370 5772
rect 16118 2896 16174 2952
rect 16524 4922 16580 4924
rect 16604 4922 16660 4924
rect 16684 4922 16740 4924
rect 16764 4922 16820 4924
rect 16524 4870 16570 4922
rect 16570 4870 16580 4922
rect 16604 4870 16634 4922
rect 16634 4870 16646 4922
rect 16646 4870 16660 4922
rect 16684 4870 16698 4922
rect 16698 4870 16710 4922
rect 16710 4870 16740 4922
rect 16764 4870 16774 4922
rect 16774 4870 16820 4922
rect 16524 4868 16580 4870
rect 16604 4868 16660 4870
rect 16684 4868 16740 4870
rect 16764 4868 16820 4870
rect 16524 3834 16580 3836
rect 16604 3834 16660 3836
rect 16684 3834 16740 3836
rect 16764 3834 16820 3836
rect 16524 3782 16570 3834
rect 16570 3782 16580 3834
rect 16604 3782 16634 3834
rect 16634 3782 16646 3834
rect 16646 3782 16660 3834
rect 16684 3782 16698 3834
rect 16698 3782 16710 3834
rect 16710 3782 16740 3834
rect 16764 3782 16774 3834
rect 16774 3782 16820 3834
rect 16524 3780 16580 3782
rect 16604 3780 16660 3782
rect 16684 3780 16740 3782
rect 16764 3780 16820 3782
rect 16524 2746 16580 2748
rect 16604 2746 16660 2748
rect 16684 2746 16740 2748
rect 16764 2746 16820 2748
rect 16524 2694 16570 2746
rect 16570 2694 16580 2746
rect 16604 2694 16634 2746
rect 16634 2694 16646 2746
rect 16646 2694 16660 2746
rect 16684 2694 16698 2746
rect 16698 2694 16710 2746
rect 16710 2694 16740 2746
rect 16764 2694 16774 2746
rect 16774 2694 16820 2746
rect 16524 2692 16580 2694
rect 16604 2692 16660 2694
rect 16684 2692 16740 2694
rect 16764 2692 16820 2694
rect 16302 992 16358 1048
rect 17682 11192 17738 11248
rect 17682 10784 17738 10840
rect 17958 11736 18014 11792
rect 17866 11600 17922 11656
rect 18050 11328 18106 11384
rect 17682 10376 17738 10432
rect 17590 8336 17646 8392
rect 17866 8336 17922 8392
rect 17590 7404 17646 7440
rect 17590 7384 17592 7404
rect 17592 7384 17644 7404
rect 17644 7384 17646 7404
rect 18050 7928 18106 7984
rect 18050 6296 18106 6352
rect 18418 9988 18474 10024
rect 18418 9968 18420 9988
rect 18420 9968 18472 9988
rect 18472 9968 18474 9988
rect 18510 9560 18566 9616
rect 18418 9152 18474 9208
rect 18326 8744 18382 8800
rect 18418 8356 18474 8392
rect 18418 8336 18420 8356
rect 18420 8336 18472 8356
rect 18472 8336 18474 8356
rect 18050 4664 18106 4720
rect 17590 3576 17646 3632
rect 16946 1400 17002 1456
rect 17774 3440 17830 3496
rect 18050 3032 18106 3088
rect 18418 7520 18474 7576
rect 18418 7148 18420 7168
rect 18420 7148 18472 7168
rect 18472 7148 18474 7168
rect 18418 7112 18474 7148
rect 18418 6704 18474 6760
rect 18418 5888 18474 5944
rect 18418 5516 18420 5536
rect 18420 5516 18472 5536
rect 18472 5516 18474 5536
rect 18418 5480 18474 5516
rect 18418 5092 18474 5128
rect 18418 5072 18420 5092
rect 18420 5072 18472 5092
rect 18472 5072 18474 5092
rect 18510 4528 18566 4584
rect 18418 4256 18474 4312
rect 18418 3884 18420 3904
rect 18420 3884 18472 3904
rect 18472 3884 18474 3904
rect 18418 3848 18474 3884
rect 18418 3440 18474 3496
rect 17590 1808 17646 1864
rect 17866 2216 17922 2272
rect 18418 2624 18474 2680
rect 18786 8472 18842 8528
rect 18878 5208 18934 5264
rect 18510 584 18566 640
<< metal3 >>
rect 0 16690 800 16720
rect 3785 16690 3851 16693
rect 0 16688 3851 16690
rect 0 16632 3790 16688
rect 3846 16632 3851 16688
rect 0 16630 3851 16632
rect 0 16600 800 16630
rect 3785 16627 3851 16630
rect 15469 16554 15535 16557
rect 19200 16554 20000 16584
rect 15469 16552 20000 16554
rect 15469 16496 15474 16552
rect 15530 16496 20000 16552
rect 15469 16494 20000 16496
rect 15469 16491 15535 16494
rect 19200 16464 20000 16494
rect 0 16282 800 16312
rect 4061 16282 4127 16285
rect 0 16280 4127 16282
rect 0 16224 4066 16280
rect 4122 16224 4127 16280
rect 0 16222 4127 16224
rect 0 16192 800 16222
rect 4061 16219 4127 16222
rect 16297 16146 16363 16149
rect 19200 16146 20000 16176
rect 16297 16144 20000 16146
rect 16297 16088 16302 16144
rect 16358 16088 20000 16144
rect 16297 16086 20000 16088
rect 16297 16083 16363 16086
rect 19200 16056 20000 16086
rect 0 15874 800 15904
rect 2773 15874 2839 15877
rect 0 15872 2839 15874
rect 0 15816 2778 15872
rect 2834 15816 2839 15872
rect 0 15814 2839 15816
rect 0 15784 800 15814
rect 2773 15811 2839 15814
rect 16849 15738 16915 15741
rect 19200 15738 20000 15768
rect 16849 15736 20000 15738
rect 16849 15680 16854 15736
rect 16910 15680 20000 15736
rect 16849 15678 20000 15680
rect 16849 15675 16915 15678
rect 19200 15648 20000 15678
rect 0 15466 800 15496
rect 4153 15466 4219 15469
rect 0 15464 4219 15466
rect 0 15408 4158 15464
rect 4214 15408 4219 15464
rect 0 15406 4219 15408
rect 0 15376 800 15406
rect 4153 15403 4219 15406
rect 17125 15330 17191 15333
rect 19200 15330 20000 15360
rect 17125 15328 20000 15330
rect 17125 15272 17130 15328
rect 17186 15272 20000 15328
rect 17125 15270 20000 15272
rect 17125 15267 17191 15270
rect 19200 15240 20000 15270
rect 0 15058 800 15088
rect 3049 15058 3115 15061
rect 0 15056 3115 15058
rect 0 15000 3054 15056
rect 3110 15000 3115 15056
rect 0 14998 3115 15000
rect 0 14968 800 14998
rect 3049 14995 3115 14998
rect 16205 14922 16271 14925
rect 19200 14922 20000 14952
rect 16205 14920 20000 14922
rect 16205 14864 16210 14920
rect 16266 14864 20000 14920
rect 16205 14862 20000 14864
rect 16205 14859 16271 14862
rect 19200 14832 20000 14862
rect 3170 14720 3486 14721
rect 0 14650 800 14680
rect 3170 14656 3176 14720
rect 3240 14656 3256 14720
rect 3320 14656 3336 14720
rect 3400 14656 3416 14720
rect 3480 14656 3486 14720
rect 3170 14655 3486 14656
rect 7618 14720 7934 14721
rect 7618 14656 7624 14720
rect 7688 14656 7704 14720
rect 7768 14656 7784 14720
rect 7848 14656 7864 14720
rect 7928 14656 7934 14720
rect 7618 14655 7934 14656
rect 12066 14720 12382 14721
rect 12066 14656 12072 14720
rect 12136 14656 12152 14720
rect 12216 14656 12232 14720
rect 12296 14656 12312 14720
rect 12376 14656 12382 14720
rect 12066 14655 12382 14656
rect 16514 14720 16830 14721
rect 16514 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16760 14720
rect 16824 14656 16830 14720
rect 16514 14655 16830 14656
rect 2957 14650 3023 14653
rect 0 14648 3023 14650
rect 0 14592 2962 14648
rect 3018 14592 3023 14648
rect 0 14590 3023 14592
rect 0 14560 800 14590
rect 2957 14587 3023 14590
rect 3601 14514 3667 14517
rect 13261 14514 13327 14517
rect 3601 14512 13327 14514
rect 3601 14456 3606 14512
rect 3662 14456 13266 14512
rect 13322 14456 13327 14512
rect 3601 14454 13327 14456
rect 3601 14451 3667 14454
rect 13261 14451 13327 14454
rect 16757 14514 16823 14517
rect 19200 14514 20000 14544
rect 16757 14512 20000 14514
rect 16757 14456 16762 14512
rect 16818 14456 20000 14512
rect 16757 14454 20000 14456
rect 16757 14451 16823 14454
rect 19200 14424 20000 14454
rect 1945 14378 2011 14381
rect 2998 14378 3004 14380
rect 1945 14376 3004 14378
rect 1945 14320 1950 14376
rect 2006 14320 3004 14376
rect 1945 14318 3004 14320
rect 1945 14315 2011 14318
rect 2998 14316 3004 14318
rect 3068 14316 3074 14380
rect 0 14242 800 14272
rect 2957 14242 3023 14245
rect 0 14240 3023 14242
rect 0 14184 2962 14240
rect 3018 14184 3023 14240
rect 0 14182 3023 14184
rect 0 14152 800 14182
rect 2957 14179 3023 14182
rect 5394 14176 5710 14177
rect 5394 14112 5400 14176
rect 5464 14112 5480 14176
rect 5544 14112 5560 14176
rect 5624 14112 5640 14176
rect 5704 14112 5710 14176
rect 5394 14111 5710 14112
rect 9842 14176 10158 14177
rect 9842 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10158 14176
rect 9842 14111 10158 14112
rect 14290 14176 14606 14177
rect 14290 14112 14296 14176
rect 14360 14112 14376 14176
rect 14440 14112 14456 14176
rect 14520 14112 14536 14176
rect 14600 14112 14606 14176
rect 14290 14111 14606 14112
rect 16481 14106 16547 14109
rect 16849 14106 16915 14109
rect 19200 14106 20000 14136
rect 16481 14104 20000 14106
rect 16481 14048 16486 14104
rect 16542 14048 16854 14104
rect 16910 14048 20000 14104
rect 16481 14046 20000 14048
rect 16481 14043 16547 14046
rect 16849 14043 16915 14046
rect 19200 14016 20000 14046
rect 5533 13970 5599 13973
rect 7833 13970 7899 13973
rect 5533 13968 7899 13970
rect 5533 13912 5538 13968
rect 5594 13912 7838 13968
rect 7894 13912 7899 13968
rect 5533 13910 7899 13912
rect 5533 13907 5599 13910
rect 7833 13907 7899 13910
rect 0 13834 800 13864
rect 2221 13834 2287 13837
rect 6729 13836 6795 13837
rect 8753 13836 8819 13837
rect 6678 13834 6684 13836
rect 0 13832 2287 13834
rect 0 13776 2226 13832
rect 2282 13776 2287 13832
rect 0 13774 2287 13776
rect 6638 13774 6684 13834
rect 6748 13832 6795 13836
rect 8702 13834 8708 13836
rect 6790 13776 6795 13832
rect 0 13744 800 13774
rect 2221 13771 2287 13774
rect 6678 13772 6684 13774
rect 6748 13772 6795 13776
rect 6729 13771 6795 13772
rect 7422 13774 8218 13834
rect 8662 13774 8708 13834
rect 8772 13832 8819 13836
rect 8814 13776 8819 13832
rect 5993 13698 6059 13701
rect 7422 13698 7482 13774
rect 5993 13696 7482 13698
rect 5993 13640 5998 13696
rect 6054 13640 7482 13696
rect 5993 13638 7482 13640
rect 8158 13698 8218 13774
rect 8702 13772 8708 13774
rect 8772 13772 8819 13776
rect 8753 13771 8819 13772
rect 11881 13698 11947 13701
rect 8158 13696 11947 13698
rect 8158 13640 11886 13696
rect 11942 13640 11947 13696
rect 8158 13638 11947 13640
rect 5993 13635 6059 13638
rect 11881 13635 11947 13638
rect 17677 13698 17743 13701
rect 19200 13698 20000 13728
rect 17677 13696 20000 13698
rect 17677 13640 17682 13696
rect 17738 13640 20000 13696
rect 17677 13638 20000 13640
rect 17677 13635 17743 13638
rect 3170 13632 3486 13633
rect 3170 13568 3176 13632
rect 3240 13568 3256 13632
rect 3320 13568 3336 13632
rect 3400 13568 3416 13632
rect 3480 13568 3486 13632
rect 3170 13567 3486 13568
rect 7618 13632 7934 13633
rect 7618 13568 7624 13632
rect 7688 13568 7704 13632
rect 7768 13568 7784 13632
rect 7848 13568 7864 13632
rect 7928 13568 7934 13632
rect 7618 13567 7934 13568
rect 12066 13632 12382 13633
rect 12066 13568 12072 13632
rect 12136 13568 12152 13632
rect 12216 13568 12232 13632
rect 12296 13568 12312 13632
rect 12376 13568 12382 13632
rect 12066 13567 12382 13568
rect 16514 13632 16830 13633
rect 16514 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16760 13632
rect 16824 13568 16830 13632
rect 19200 13608 20000 13638
rect 16514 13567 16830 13568
rect 0 13426 800 13456
rect 2037 13426 2103 13429
rect 0 13424 2103 13426
rect 0 13368 2042 13424
rect 2098 13368 2103 13424
rect 0 13366 2103 13368
rect 0 13336 800 13366
rect 2037 13363 2103 13366
rect 3509 13426 3575 13429
rect 9857 13426 9923 13429
rect 3509 13424 9923 13426
rect 3509 13368 3514 13424
rect 3570 13368 9862 13424
rect 9918 13368 9923 13424
rect 3509 13366 9923 13368
rect 3509 13363 3575 13366
rect 9857 13363 9923 13366
rect 4061 13290 4127 13293
rect 11145 13290 11211 13293
rect 17309 13290 17375 13293
rect 4061 13288 11211 13290
rect 4061 13232 4066 13288
rect 4122 13232 11150 13288
rect 11206 13232 11211 13288
rect 4061 13230 11211 13232
rect 4061 13227 4127 13230
rect 11145 13227 11211 13230
rect 12390 13288 17375 13290
rect 12390 13232 17314 13288
rect 17370 13232 17375 13288
rect 12390 13230 17375 13232
rect 5394 13088 5710 13089
rect 0 13018 800 13048
rect 5394 13024 5400 13088
rect 5464 13024 5480 13088
rect 5544 13024 5560 13088
rect 5624 13024 5640 13088
rect 5704 13024 5710 13088
rect 5394 13023 5710 13024
rect 9842 13088 10158 13089
rect 9842 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10158 13088
rect 9842 13023 10158 13024
rect 2773 13018 2839 13021
rect 3785 13018 3851 13021
rect 12390 13018 12450 13230
rect 17309 13227 17375 13230
rect 17769 13290 17835 13293
rect 19200 13290 20000 13320
rect 17769 13288 20000 13290
rect 17769 13232 17774 13288
rect 17830 13232 20000 13288
rect 17769 13230 20000 13232
rect 17769 13227 17835 13230
rect 19200 13200 20000 13230
rect 14290 13088 14606 13089
rect 14290 13024 14296 13088
rect 14360 13024 14376 13088
rect 14440 13024 14456 13088
rect 14520 13024 14536 13088
rect 14600 13024 14606 13088
rect 14290 13023 14606 13024
rect 0 13016 3851 13018
rect 0 12960 2778 13016
rect 2834 12960 3790 13016
rect 3846 12960 3851 13016
rect 0 12958 3851 12960
rect 0 12928 800 12958
rect 2773 12955 2839 12958
rect 3785 12955 3851 12958
rect 10366 12958 12450 13018
rect 2773 12882 2839 12885
rect 5349 12882 5415 12885
rect 2773 12880 5415 12882
rect 2773 12824 2778 12880
rect 2834 12824 5354 12880
rect 5410 12824 5415 12880
rect 2773 12822 5415 12824
rect 2773 12819 2839 12822
rect 5349 12819 5415 12822
rect 9489 12882 9555 12885
rect 10366 12882 10426 12958
rect 16297 12882 16363 12885
rect 9489 12880 10426 12882
rect 9489 12824 9494 12880
rect 9550 12824 10426 12880
rect 9489 12822 10426 12824
rect 12390 12880 16363 12882
rect 12390 12824 16302 12880
rect 16358 12824 16363 12880
rect 12390 12822 16363 12824
rect 9489 12819 9555 12822
rect 2865 12746 2931 12749
rect 3509 12746 3575 12749
rect 12390 12746 12450 12822
rect 16297 12819 16363 12822
rect 17585 12882 17651 12885
rect 19200 12882 20000 12912
rect 17585 12880 20000 12882
rect 17585 12824 17590 12880
rect 17646 12824 20000 12880
rect 17585 12822 20000 12824
rect 17585 12819 17651 12822
rect 19200 12792 20000 12822
rect 2865 12744 12450 12746
rect 2865 12688 2870 12744
rect 2926 12688 3514 12744
rect 3570 12688 12450 12744
rect 2865 12686 12450 12688
rect 2865 12683 2931 12686
rect 3509 12683 3575 12686
rect 0 12610 800 12640
rect 2221 12610 2287 12613
rect 0 12608 2287 12610
rect 0 12552 2226 12608
rect 2282 12552 2287 12608
rect 0 12550 2287 12552
rect 0 12520 800 12550
rect 2221 12547 2287 12550
rect 3170 12544 3486 12545
rect 3170 12480 3176 12544
rect 3240 12480 3256 12544
rect 3320 12480 3336 12544
rect 3400 12480 3416 12544
rect 3480 12480 3486 12544
rect 3170 12479 3486 12480
rect 7618 12544 7934 12545
rect 7618 12480 7624 12544
rect 7688 12480 7704 12544
rect 7768 12480 7784 12544
rect 7848 12480 7864 12544
rect 7928 12480 7934 12544
rect 7618 12479 7934 12480
rect 12066 12544 12382 12545
rect 12066 12480 12072 12544
rect 12136 12480 12152 12544
rect 12216 12480 12232 12544
rect 12296 12480 12312 12544
rect 12376 12480 12382 12544
rect 12066 12479 12382 12480
rect 16514 12544 16830 12545
rect 16514 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16760 12544
rect 16824 12480 16830 12544
rect 16514 12479 16830 12480
rect 17677 12474 17743 12477
rect 19200 12474 20000 12504
rect 17677 12472 20000 12474
rect 17677 12416 17682 12472
rect 17738 12416 20000 12472
rect 17677 12414 20000 12416
rect 17677 12411 17743 12414
rect 19200 12384 20000 12414
rect 3693 12338 3759 12341
rect 8477 12338 8543 12341
rect 3693 12336 8543 12338
rect 3693 12280 3698 12336
rect 3754 12280 8482 12336
rect 8538 12280 8543 12336
rect 3693 12278 8543 12280
rect 3693 12275 3759 12278
rect 8477 12275 8543 12278
rect 8845 12338 8911 12341
rect 12709 12338 12775 12341
rect 8845 12336 12775 12338
rect 8845 12280 8850 12336
rect 8906 12280 12714 12336
rect 12770 12280 12775 12336
rect 8845 12278 12775 12280
rect 8845 12275 8911 12278
rect 12709 12275 12775 12278
rect 17861 12340 17927 12341
rect 17861 12336 17908 12340
rect 17972 12338 17978 12340
rect 17861 12280 17866 12336
rect 17861 12276 17908 12280
rect 17972 12278 18018 12338
rect 17972 12276 17978 12278
rect 17861 12275 17927 12276
rect 0 12202 800 12232
rect 2405 12202 2471 12205
rect 0 12200 2471 12202
rect 0 12144 2410 12200
rect 2466 12144 2471 12200
rect 0 12142 2471 12144
rect 0 12112 800 12142
rect 2405 12139 2471 12142
rect 3141 12202 3207 12205
rect 15377 12202 15443 12205
rect 3141 12200 15443 12202
rect 3141 12144 3146 12200
rect 3202 12144 15382 12200
rect 15438 12144 15443 12200
rect 3141 12142 15443 12144
rect 3141 12139 3207 12142
rect 15377 12139 15443 12142
rect 6453 12066 6519 12069
rect 8845 12066 8911 12069
rect 6453 12064 8911 12066
rect 6453 12008 6458 12064
rect 6514 12008 8850 12064
rect 8906 12008 8911 12064
rect 6453 12006 8911 12008
rect 6453 12003 6519 12006
rect 8845 12003 8911 12006
rect 17769 12066 17835 12069
rect 19200 12066 20000 12096
rect 17769 12064 20000 12066
rect 17769 12008 17774 12064
rect 17830 12008 20000 12064
rect 17769 12006 20000 12008
rect 17769 12003 17835 12006
rect 5394 12000 5710 12001
rect 5394 11936 5400 12000
rect 5464 11936 5480 12000
rect 5544 11936 5560 12000
rect 5624 11936 5640 12000
rect 5704 11936 5710 12000
rect 5394 11935 5710 11936
rect 9842 12000 10158 12001
rect 9842 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10158 12000
rect 9842 11935 10158 11936
rect 14290 12000 14606 12001
rect 14290 11936 14296 12000
rect 14360 11936 14376 12000
rect 14440 11936 14456 12000
rect 14520 11936 14536 12000
rect 14600 11936 14606 12000
rect 19200 11976 20000 12006
rect 14290 11935 14606 11936
rect 17401 11930 17467 11933
rect 17769 11930 17835 11933
rect 17401 11928 17835 11930
rect 17401 11872 17406 11928
rect 17462 11872 17774 11928
rect 17830 11872 17835 11928
rect 17401 11870 17835 11872
rect 17401 11867 17467 11870
rect 17769 11867 17835 11870
rect 0 11794 800 11824
rect 2773 11794 2839 11797
rect 0 11792 2839 11794
rect 0 11736 2778 11792
rect 2834 11736 2839 11792
rect 0 11734 2839 11736
rect 0 11704 800 11734
rect 2773 11731 2839 11734
rect 13261 11794 13327 11797
rect 17953 11794 18019 11797
rect 13261 11792 18019 11794
rect 13261 11736 13266 11792
rect 13322 11736 17958 11792
rect 18014 11736 18019 11792
rect 13261 11734 18019 11736
rect 13261 11731 13327 11734
rect 17953 11731 18019 11734
rect 2497 11658 2563 11661
rect 2998 11658 3004 11660
rect 2497 11656 3004 11658
rect 2497 11600 2502 11656
rect 2558 11600 3004 11656
rect 2497 11598 3004 11600
rect 2497 11595 2563 11598
rect 2998 11596 3004 11598
rect 3068 11596 3074 11660
rect 3601 11658 3667 11661
rect 13169 11658 13235 11661
rect 17125 11658 17191 11661
rect 3601 11656 13002 11658
rect 3601 11600 3606 11656
rect 3662 11600 13002 11656
rect 3601 11598 13002 11600
rect 3601 11595 3667 11598
rect 12942 11522 13002 11598
rect 13169 11656 17191 11658
rect 13169 11600 13174 11656
rect 13230 11600 17130 11656
rect 17186 11600 17191 11656
rect 13169 11598 17191 11600
rect 13169 11595 13235 11598
rect 17125 11595 17191 11598
rect 17861 11658 17927 11661
rect 19200 11658 20000 11688
rect 17861 11656 20000 11658
rect 17861 11600 17866 11656
rect 17922 11600 20000 11656
rect 17861 11598 20000 11600
rect 17861 11595 17927 11598
rect 19200 11568 20000 11598
rect 14089 11522 14155 11525
rect 14549 11522 14615 11525
rect 12942 11520 14615 11522
rect 12942 11464 14094 11520
rect 14150 11464 14554 11520
rect 14610 11464 14615 11520
rect 12942 11462 14615 11464
rect 14089 11459 14155 11462
rect 14549 11459 14615 11462
rect 3170 11456 3486 11457
rect 0 11386 800 11416
rect 3170 11392 3176 11456
rect 3240 11392 3256 11456
rect 3320 11392 3336 11456
rect 3400 11392 3416 11456
rect 3480 11392 3486 11456
rect 3170 11391 3486 11392
rect 7618 11456 7934 11457
rect 7618 11392 7624 11456
rect 7688 11392 7704 11456
rect 7768 11392 7784 11456
rect 7848 11392 7864 11456
rect 7928 11392 7934 11456
rect 7618 11391 7934 11392
rect 12066 11456 12382 11457
rect 12066 11392 12072 11456
rect 12136 11392 12152 11456
rect 12216 11392 12232 11456
rect 12296 11392 12312 11456
rect 12376 11392 12382 11456
rect 12066 11391 12382 11392
rect 16514 11456 16830 11457
rect 16514 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16760 11456
rect 16824 11392 16830 11456
rect 16514 11391 16830 11392
rect 2221 11386 2287 11389
rect 18045 11386 18111 11389
rect 0 11384 2287 11386
rect 0 11328 2226 11384
rect 2282 11328 2287 11384
rect 0 11326 2287 11328
rect 0 11296 800 11326
rect 2221 11323 2287 11326
rect 16990 11384 18111 11386
rect 16990 11328 18050 11384
rect 18106 11328 18111 11384
rect 16990 11326 18111 11328
rect 1945 11250 2011 11253
rect 10041 11250 10107 11253
rect 10869 11250 10935 11253
rect 16990 11250 17050 11326
rect 18045 11323 18111 11326
rect 1945 11248 10935 11250
rect 1945 11192 1950 11248
rect 2006 11192 10046 11248
rect 10102 11192 10874 11248
rect 10930 11192 10935 11248
rect 1945 11190 10935 11192
rect 1945 11187 2011 11190
rect 10041 11187 10107 11190
rect 10869 11187 10935 11190
rect 11102 11190 17050 11250
rect 17677 11250 17743 11253
rect 19200 11250 20000 11280
rect 17677 11248 20000 11250
rect 17677 11192 17682 11248
rect 17738 11192 20000 11248
rect 17677 11190 20000 11192
rect 9622 11052 9628 11116
rect 9692 11114 9698 11116
rect 9765 11114 9831 11117
rect 11102 11114 11162 11190
rect 17677 11187 17743 11190
rect 19200 11160 20000 11190
rect 9692 11112 11162 11114
rect 9692 11056 9770 11112
rect 9826 11056 11162 11112
rect 9692 11054 11162 11056
rect 11237 11114 11303 11117
rect 17033 11114 17099 11117
rect 11237 11112 17099 11114
rect 11237 11056 11242 11112
rect 11298 11056 17038 11112
rect 17094 11056 17099 11112
rect 11237 11054 17099 11056
rect 9692 11052 9698 11054
rect 9765 11051 9831 11054
rect 11237 11051 11303 11054
rect 17033 11051 17099 11054
rect 0 10978 800 11008
rect 2221 10978 2287 10981
rect 0 10976 2287 10978
rect 0 10920 2226 10976
rect 2282 10920 2287 10976
rect 0 10918 2287 10920
rect 0 10888 800 10918
rect 2221 10915 2287 10918
rect 5394 10912 5710 10913
rect 5394 10848 5400 10912
rect 5464 10848 5480 10912
rect 5544 10848 5560 10912
rect 5624 10848 5640 10912
rect 5704 10848 5710 10912
rect 5394 10847 5710 10848
rect 9842 10912 10158 10913
rect 9842 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10158 10912
rect 9842 10847 10158 10848
rect 14290 10912 14606 10913
rect 14290 10848 14296 10912
rect 14360 10848 14376 10912
rect 14440 10848 14456 10912
rect 14520 10848 14536 10912
rect 14600 10848 14606 10912
rect 14290 10847 14606 10848
rect 17677 10842 17743 10845
rect 19200 10842 20000 10872
rect 17677 10840 20000 10842
rect 17677 10784 17682 10840
rect 17738 10784 20000 10840
rect 17677 10782 20000 10784
rect 17677 10779 17743 10782
rect 19200 10752 20000 10782
rect 2129 10706 2195 10709
rect 14457 10706 14523 10709
rect 16849 10706 16915 10709
rect 2129 10704 16915 10706
rect 2129 10648 2134 10704
rect 2190 10648 14462 10704
rect 14518 10648 16854 10704
rect 16910 10648 16915 10704
rect 2129 10646 16915 10648
rect 2129 10643 2195 10646
rect 14457 10643 14523 10646
rect 16849 10643 16915 10646
rect 0 10570 800 10600
rect 2221 10570 2287 10573
rect 0 10568 2287 10570
rect 0 10512 2226 10568
rect 2282 10512 2287 10568
rect 0 10510 2287 10512
rect 0 10480 800 10510
rect 2221 10507 2287 10510
rect 17677 10434 17743 10437
rect 19200 10434 20000 10464
rect 17677 10432 20000 10434
rect 17677 10376 17682 10432
rect 17738 10376 20000 10432
rect 17677 10374 20000 10376
rect 17677 10371 17743 10374
rect 3170 10368 3486 10369
rect 3170 10304 3176 10368
rect 3240 10304 3256 10368
rect 3320 10304 3336 10368
rect 3400 10304 3416 10368
rect 3480 10304 3486 10368
rect 3170 10303 3486 10304
rect 7618 10368 7934 10369
rect 7618 10304 7624 10368
rect 7688 10304 7704 10368
rect 7768 10304 7784 10368
rect 7848 10304 7864 10368
rect 7928 10304 7934 10368
rect 7618 10303 7934 10304
rect 12066 10368 12382 10369
rect 12066 10304 12072 10368
rect 12136 10304 12152 10368
rect 12216 10304 12232 10368
rect 12296 10304 12312 10368
rect 12376 10304 12382 10368
rect 12066 10303 12382 10304
rect 16514 10368 16830 10369
rect 16514 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16760 10368
rect 16824 10304 16830 10368
rect 19200 10344 20000 10374
rect 16514 10303 16830 10304
rect 0 10162 800 10192
rect 1485 10162 1551 10165
rect 0 10160 1551 10162
rect 0 10104 1490 10160
rect 1546 10104 1551 10160
rect 0 10102 1551 10104
rect 0 10072 800 10102
rect 1485 10099 1551 10102
rect 18413 10026 18479 10029
rect 19200 10026 20000 10056
rect 18413 10024 20000 10026
rect 18413 9968 18418 10024
rect 18474 9968 20000 10024
rect 18413 9966 20000 9968
rect 18413 9963 18479 9966
rect 19200 9936 20000 9966
rect 5394 9824 5710 9825
rect 0 9754 800 9784
rect 5394 9760 5400 9824
rect 5464 9760 5480 9824
rect 5544 9760 5560 9824
rect 5624 9760 5640 9824
rect 5704 9760 5710 9824
rect 5394 9759 5710 9760
rect 9842 9824 10158 9825
rect 9842 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10158 9824
rect 9842 9759 10158 9760
rect 14290 9824 14606 9825
rect 14290 9760 14296 9824
rect 14360 9760 14376 9824
rect 14440 9760 14456 9824
rect 14520 9760 14536 9824
rect 14600 9760 14606 9824
rect 14290 9759 14606 9760
rect 3233 9754 3299 9757
rect 0 9752 3299 9754
rect 0 9696 3238 9752
rect 3294 9696 3299 9752
rect 0 9694 3299 9696
rect 0 9664 800 9694
rect 3233 9691 3299 9694
rect 1485 9618 1551 9621
rect 2681 9618 2747 9621
rect 1485 9616 2747 9618
rect 1485 9560 1490 9616
rect 1546 9560 2686 9616
rect 2742 9560 2747 9616
rect 1485 9558 2747 9560
rect 1485 9555 1551 9558
rect 2681 9555 2747 9558
rect 18505 9618 18571 9621
rect 19200 9618 20000 9648
rect 18505 9616 20000 9618
rect 18505 9560 18510 9616
rect 18566 9560 20000 9616
rect 18505 9558 20000 9560
rect 18505 9555 18571 9558
rect 19200 9528 20000 9558
rect 4981 9482 5047 9485
rect 17309 9482 17375 9485
rect 4981 9480 17375 9482
rect 4981 9424 4986 9480
rect 5042 9424 17314 9480
rect 17370 9424 17375 9480
rect 4981 9422 17375 9424
rect 4981 9419 5047 9422
rect 17309 9419 17375 9422
rect 0 9346 800 9376
rect 1485 9346 1551 9349
rect 0 9344 1551 9346
rect 0 9288 1490 9344
rect 1546 9288 1551 9344
rect 0 9286 1551 9288
rect 0 9256 800 9286
rect 1485 9283 1551 9286
rect 3170 9280 3486 9281
rect 3170 9216 3176 9280
rect 3240 9216 3256 9280
rect 3320 9216 3336 9280
rect 3400 9216 3416 9280
rect 3480 9216 3486 9280
rect 3170 9215 3486 9216
rect 7618 9280 7934 9281
rect 7618 9216 7624 9280
rect 7688 9216 7704 9280
rect 7768 9216 7784 9280
rect 7848 9216 7864 9280
rect 7928 9216 7934 9280
rect 7618 9215 7934 9216
rect 12066 9280 12382 9281
rect 12066 9216 12072 9280
rect 12136 9216 12152 9280
rect 12216 9216 12232 9280
rect 12296 9216 12312 9280
rect 12376 9216 12382 9280
rect 12066 9215 12382 9216
rect 16514 9280 16830 9281
rect 16514 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16760 9280
rect 16824 9216 16830 9280
rect 16514 9215 16830 9216
rect 17401 9210 17467 9213
rect 18413 9210 18479 9213
rect 19200 9210 20000 9240
rect 17401 9208 20000 9210
rect 17401 9152 17406 9208
rect 17462 9152 18418 9208
rect 18474 9152 20000 9208
rect 17401 9150 20000 9152
rect 17401 9147 17467 9150
rect 18413 9147 18479 9150
rect 19200 9120 20000 9150
rect 0 8938 800 8968
rect 1945 8938 2011 8941
rect 0 8936 2011 8938
rect 0 8880 1950 8936
rect 2006 8880 2011 8936
rect 0 8878 2011 8880
rect 0 8848 800 8878
rect 1945 8875 2011 8878
rect 18321 8802 18387 8805
rect 19200 8802 20000 8832
rect 18321 8800 20000 8802
rect 18321 8744 18326 8800
rect 18382 8744 20000 8800
rect 18321 8742 20000 8744
rect 18321 8739 18387 8742
rect 5394 8736 5710 8737
rect 5394 8672 5400 8736
rect 5464 8672 5480 8736
rect 5544 8672 5560 8736
rect 5624 8672 5640 8736
rect 5704 8672 5710 8736
rect 5394 8671 5710 8672
rect 9842 8736 10158 8737
rect 9842 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10158 8736
rect 9842 8671 10158 8672
rect 14290 8736 14606 8737
rect 14290 8672 14296 8736
rect 14360 8672 14376 8736
rect 14440 8672 14456 8736
rect 14520 8672 14536 8736
rect 14600 8672 14606 8736
rect 19200 8712 20000 8742
rect 14290 8671 14606 8672
rect 2865 8664 2931 8669
rect 2865 8608 2870 8664
rect 2926 8608 2931 8664
rect 2865 8603 2931 8608
rect 0 8530 800 8560
rect 1485 8530 1551 8533
rect 0 8528 1551 8530
rect 0 8472 1490 8528
rect 1546 8472 1551 8528
rect 0 8470 1551 8472
rect 0 8440 800 8470
rect 1485 8467 1551 8470
rect 2313 8530 2379 8533
rect 2868 8530 2928 8603
rect 2313 8528 2928 8530
rect 2313 8472 2318 8528
rect 2374 8472 2928 8528
rect 2313 8470 2928 8472
rect 14641 8530 14707 8533
rect 18781 8530 18847 8533
rect 14641 8528 18847 8530
rect 14641 8472 14646 8528
rect 14702 8472 18786 8528
rect 18842 8472 18847 8528
rect 14641 8470 18847 8472
rect 2313 8467 2379 8470
rect 14641 8467 14707 8470
rect 18781 8467 18847 8470
rect 2957 8394 3023 8397
rect 4245 8394 4311 8397
rect 2957 8392 4311 8394
rect 2957 8336 2962 8392
rect 3018 8336 4250 8392
rect 4306 8336 4311 8392
rect 2957 8334 4311 8336
rect 2957 8331 3023 8334
rect 4245 8331 4311 8334
rect 6085 8394 6151 8397
rect 17585 8394 17651 8397
rect 17861 8396 17927 8397
rect 17861 8394 17908 8396
rect 6085 8392 17651 8394
rect 6085 8336 6090 8392
rect 6146 8336 17590 8392
rect 17646 8336 17651 8392
rect 6085 8334 17651 8336
rect 17816 8392 17908 8394
rect 17816 8336 17866 8392
rect 17816 8334 17908 8336
rect 6085 8331 6151 8334
rect 17585 8331 17651 8334
rect 17861 8332 17908 8334
rect 17972 8332 17978 8396
rect 18413 8394 18479 8397
rect 19200 8394 20000 8424
rect 18413 8392 20000 8394
rect 18413 8336 18418 8392
rect 18474 8336 20000 8392
rect 18413 8334 20000 8336
rect 17861 8331 17927 8332
rect 18413 8331 18479 8334
rect 19200 8304 20000 8334
rect 3170 8192 3486 8193
rect 0 8122 800 8152
rect 3170 8128 3176 8192
rect 3240 8128 3256 8192
rect 3320 8128 3336 8192
rect 3400 8128 3416 8192
rect 3480 8128 3486 8192
rect 3170 8127 3486 8128
rect 7618 8192 7934 8193
rect 7618 8128 7624 8192
rect 7688 8128 7704 8192
rect 7768 8128 7784 8192
rect 7848 8128 7864 8192
rect 7928 8128 7934 8192
rect 7618 8127 7934 8128
rect 12066 8192 12382 8193
rect 12066 8128 12072 8192
rect 12136 8128 12152 8192
rect 12216 8128 12232 8192
rect 12296 8128 12312 8192
rect 12376 8128 12382 8192
rect 12066 8127 12382 8128
rect 16514 8192 16830 8193
rect 16514 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16760 8192
rect 16824 8128 16830 8192
rect 16514 8127 16830 8128
rect 1485 8122 1551 8125
rect 0 8120 1551 8122
rect 0 8064 1490 8120
rect 1546 8064 1551 8120
rect 0 8062 1551 8064
rect 0 8032 800 8062
rect 1485 8059 1551 8062
rect 18045 7986 18111 7989
rect 19200 7986 20000 8016
rect 18045 7984 20000 7986
rect 18045 7928 18050 7984
rect 18106 7928 20000 7984
rect 18045 7926 20000 7928
rect 18045 7923 18111 7926
rect 19200 7896 20000 7926
rect 11605 7850 11671 7853
rect 16389 7850 16455 7853
rect 11605 7848 16455 7850
rect 11605 7792 11610 7848
rect 11666 7792 16394 7848
rect 16450 7792 16455 7848
rect 11605 7790 16455 7792
rect 11605 7787 11671 7790
rect 16389 7787 16455 7790
rect 0 7714 800 7744
rect 1853 7714 1919 7717
rect 0 7712 1919 7714
rect 0 7656 1858 7712
rect 1914 7656 1919 7712
rect 0 7654 1919 7656
rect 0 7624 800 7654
rect 1853 7651 1919 7654
rect 5394 7648 5710 7649
rect 5394 7584 5400 7648
rect 5464 7584 5480 7648
rect 5544 7584 5560 7648
rect 5624 7584 5640 7648
rect 5704 7584 5710 7648
rect 5394 7583 5710 7584
rect 9842 7648 10158 7649
rect 9842 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10158 7648
rect 9842 7583 10158 7584
rect 14290 7648 14606 7649
rect 14290 7584 14296 7648
rect 14360 7584 14376 7648
rect 14440 7584 14456 7648
rect 14520 7584 14536 7648
rect 14600 7584 14606 7648
rect 14290 7583 14606 7584
rect 18413 7578 18479 7581
rect 19200 7578 20000 7608
rect 18413 7576 20000 7578
rect 18413 7520 18418 7576
rect 18474 7520 20000 7576
rect 18413 7518 20000 7520
rect 18413 7515 18479 7518
rect 19200 7488 20000 7518
rect 8385 7442 8451 7445
rect 17585 7442 17651 7445
rect 8385 7440 17651 7442
rect 8385 7384 8390 7440
rect 8446 7384 17590 7440
rect 17646 7384 17651 7440
rect 8385 7382 17651 7384
rect 8385 7379 8451 7382
rect 17585 7379 17651 7382
rect 0 7306 800 7336
rect 1485 7306 1551 7309
rect 0 7304 1551 7306
rect 0 7248 1490 7304
rect 1546 7248 1551 7304
rect 0 7246 1551 7248
rect 0 7216 800 7246
rect 1485 7243 1551 7246
rect 2998 7244 3004 7308
rect 3068 7306 3074 7308
rect 6637 7306 6703 7309
rect 3068 7304 6703 7306
rect 3068 7248 6642 7304
rect 6698 7248 6703 7304
rect 3068 7246 6703 7248
rect 3068 7244 3074 7246
rect 6637 7243 6703 7246
rect 18413 7170 18479 7173
rect 19200 7170 20000 7200
rect 18413 7168 20000 7170
rect 18413 7112 18418 7168
rect 18474 7112 20000 7168
rect 18413 7110 20000 7112
rect 18413 7107 18479 7110
rect 3170 7104 3486 7105
rect 3170 7040 3176 7104
rect 3240 7040 3256 7104
rect 3320 7040 3336 7104
rect 3400 7040 3416 7104
rect 3480 7040 3486 7104
rect 3170 7039 3486 7040
rect 7618 7104 7934 7105
rect 7618 7040 7624 7104
rect 7688 7040 7704 7104
rect 7768 7040 7784 7104
rect 7848 7040 7864 7104
rect 7928 7040 7934 7104
rect 7618 7039 7934 7040
rect 12066 7104 12382 7105
rect 12066 7040 12072 7104
rect 12136 7040 12152 7104
rect 12216 7040 12232 7104
rect 12296 7040 12312 7104
rect 12376 7040 12382 7104
rect 12066 7039 12382 7040
rect 16514 7104 16830 7105
rect 16514 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16760 7104
rect 16824 7040 16830 7104
rect 19200 7080 20000 7110
rect 16514 7039 16830 7040
rect 0 6898 800 6928
rect 1577 6898 1643 6901
rect 0 6896 1643 6898
rect 0 6840 1582 6896
rect 1638 6840 1643 6896
rect 0 6838 1643 6840
rect 0 6808 800 6838
rect 1577 6835 1643 6838
rect 2129 6898 2195 6901
rect 7281 6898 7347 6901
rect 2129 6896 7347 6898
rect 2129 6840 2134 6896
rect 2190 6840 7286 6896
rect 7342 6840 7347 6896
rect 2129 6838 7347 6840
rect 2129 6835 2195 6838
rect 7281 6835 7347 6838
rect 1577 6762 1643 6765
rect 3785 6762 3851 6765
rect 15009 6762 15075 6765
rect 1577 6760 3851 6762
rect 1577 6704 1582 6760
rect 1638 6704 3790 6760
rect 3846 6704 3851 6760
rect 1577 6702 3851 6704
rect 1577 6699 1643 6702
rect 3785 6699 3851 6702
rect 4294 6760 15075 6762
rect 4294 6704 15014 6760
rect 15070 6704 15075 6760
rect 4294 6702 15075 6704
rect 3325 6626 3391 6629
rect 4061 6626 4127 6629
rect 4294 6626 4354 6702
rect 15009 6699 15075 6702
rect 18413 6762 18479 6765
rect 19200 6762 20000 6792
rect 18413 6760 20000 6762
rect 18413 6704 18418 6760
rect 18474 6704 20000 6760
rect 18413 6702 20000 6704
rect 18413 6699 18479 6702
rect 19200 6672 20000 6702
rect 3325 6624 4354 6626
rect 3325 6568 3330 6624
rect 3386 6568 4066 6624
rect 4122 6568 4354 6624
rect 3325 6566 4354 6568
rect 3325 6563 3391 6566
rect 4061 6563 4127 6566
rect 5394 6560 5710 6561
rect 0 6490 800 6520
rect 5394 6496 5400 6560
rect 5464 6496 5480 6560
rect 5544 6496 5560 6560
rect 5624 6496 5640 6560
rect 5704 6496 5710 6560
rect 5394 6495 5710 6496
rect 9842 6560 10158 6561
rect 9842 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10158 6560
rect 9842 6495 10158 6496
rect 14290 6560 14606 6561
rect 14290 6496 14296 6560
rect 14360 6496 14376 6560
rect 14440 6496 14456 6560
rect 14520 6496 14536 6560
rect 14600 6496 14606 6560
rect 14290 6495 14606 6496
rect 3969 6490 4035 6493
rect 0 6488 4035 6490
rect 0 6432 3974 6488
rect 4030 6432 4035 6488
rect 0 6430 4035 6432
rect 0 6400 800 6430
rect 3969 6427 4035 6430
rect 3141 6354 3207 6357
rect 4153 6354 4219 6357
rect 3141 6352 4219 6354
rect 3141 6296 3146 6352
rect 3202 6296 4158 6352
rect 4214 6296 4219 6352
rect 3141 6294 4219 6296
rect 3141 6291 3207 6294
rect 4153 6291 4219 6294
rect 18045 6354 18111 6357
rect 19200 6354 20000 6384
rect 18045 6352 20000 6354
rect 18045 6296 18050 6352
rect 18106 6296 20000 6352
rect 18045 6294 20000 6296
rect 18045 6291 18111 6294
rect 19200 6264 20000 6294
rect 6545 6218 6611 6221
rect 16941 6218 17007 6221
rect 6545 6216 17007 6218
rect 6545 6160 6550 6216
rect 6606 6160 16946 6216
rect 17002 6160 17007 6216
rect 6545 6158 17007 6160
rect 6545 6155 6611 6158
rect 16941 6155 17007 6158
rect 0 6082 800 6112
rect 1485 6082 1551 6085
rect 0 6080 1551 6082
rect 0 6024 1490 6080
rect 1546 6024 1551 6080
rect 0 6022 1551 6024
rect 0 5992 800 6022
rect 1485 6019 1551 6022
rect 3170 6016 3486 6017
rect 3170 5952 3176 6016
rect 3240 5952 3256 6016
rect 3320 5952 3336 6016
rect 3400 5952 3416 6016
rect 3480 5952 3486 6016
rect 3170 5951 3486 5952
rect 7618 6016 7934 6017
rect 7618 5952 7624 6016
rect 7688 5952 7704 6016
rect 7768 5952 7784 6016
rect 7848 5952 7864 6016
rect 7928 5952 7934 6016
rect 7618 5951 7934 5952
rect 12066 6016 12382 6017
rect 12066 5952 12072 6016
rect 12136 5952 12152 6016
rect 12216 5952 12232 6016
rect 12296 5952 12312 6016
rect 12376 5952 12382 6016
rect 12066 5951 12382 5952
rect 16514 6016 16830 6017
rect 16514 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16760 6016
rect 16824 5952 16830 6016
rect 16514 5951 16830 5952
rect 18413 5946 18479 5949
rect 19200 5946 20000 5976
rect 18413 5944 20000 5946
rect 18413 5888 18418 5944
rect 18474 5888 20000 5944
rect 18413 5886 20000 5888
rect 18413 5883 18479 5886
rect 19200 5856 20000 5886
rect 1669 5810 1735 5813
rect 5993 5810 6059 5813
rect 1669 5808 6059 5810
rect 1669 5752 1674 5808
rect 1730 5752 5998 5808
rect 6054 5752 6059 5808
rect 1669 5750 6059 5752
rect 1669 5747 1735 5750
rect 5993 5747 6059 5750
rect 14089 5810 14155 5813
rect 17309 5810 17375 5813
rect 14089 5808 17375 5810
rect 14089 5752 14094 5808
rect 14150 5752 17314 5808
rect 17370 5752 17375 5808
rect 14089 5750 17375 5752
rect 14089 5747 14155 5750
rect 17309 5747 17375 5750
rect 0 5674 800 5704
rect 1945 5674 2011 5677
rect 0 5672 2011 5674
rect 0 5616 1950 5672
rect 2006 5616 2011 5672
rect 0 5614 2011 5616
rect 0 5584 800 5614
rect 1945 5611 2011 5614
rect 4521 5674 4587 5677
rect 6269 5674 6335 5677
rect 4521 5672 6335 5674
rect 4521 5616 4526 5672
rect 4582 5616 6274 5672
rect 6330 5616 6335 5672
rect 4521 5614 6335 5616
rect 4521 5611 4587 5614
rect 6269 5611 6335 5614
rect 2814 5476 2820 5540
rect 2884 5538 2890 5540
rect 3233 5538 3299 5541
rect 2884 5536 3299 5538
rect 2884 5480 3238 5536
rect 3294 5480 3299 5536
rect 2884 5478 3299 5480
rect 2884 5476 2890 5478
rect 3233 5475 3299 5478
rect 18413 5538 18479 5541
rect 19200 5538 20000 5568
rect 18413 5536 20000 5538
rect 18413 5480 18418 5536
rect 18474 5480 20000 5536
rect 18413 5478 20000 5480
rect 18413 5475 18479 5478
rect 5394 5472 5710 5473
rect 5394 5408 5400 5472
rect 5464 5408 5480 5472
rect 5544 5408 5560 5472
rect 5624 5408 5640 5472
rect 5704 5408 5710 5472
rect 5394 5407 5710 5408
rect 9842 5472 10158 5473
rect 9842 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10158 5472
rect 9842 5407 10158 5408
rect 14290 5472 14606 5473
rect 14290 5408 14296 5472
rect 14360 5408 14376 5472
rect 14440 5408 14456 5472
rect 14520 5408 14536 5472
rect 14600 5408 14606 5472
rect 19200 5448 20000 5478
rect 14290 5407 14606 5408
rect 2405 5402 2471 5405
rect 1166 5400 2471 5402
rect 1166 5344 2410 5400
rect 2466 5344 2471 5400
rect 1166 5342 2471 5344
rect 0 5266 800 5296
rect 1166 5266 1226 5342
rect 2405 5339 2471 5342
rect 0 5206 1226 5266
rect 2405 5266 2471 5269
rect 3509 5266 3575 5269
rect 14917 5266 14983 5269
rect 2405 5264 14983 5266
rect 2405 5208 2410 5264
rect 2466 5208 3514 5264
rect 3570 5208 14922 5264
rect 14978 5208 14983 5264
rect 2405 5206 14983 5208
rect 0 5176 800 5206
rect 2405 5203 2471 5206
rect 3509 5203 3575 5206
rect 14917 5203 14983 5206
rect 15469 5266 15535 5269
rect 16113 5266 16179 5269
rect 18873 5266 18939 5269
rect 15469 5264 18939 5266
rect 15469 5208 15474 5264
rect 15530 5208 16118 5264
rect 16174 5208 18878 5264
rect 18934 5208 18939 5264
rect 15469 5206 18939 5208
rect 15469 5203 15535 5206
rect 16113 5203 16179 5206
rect 18873 5203 18939 5206
rect 12157 5130 12223 5133
rect 15009 5130 15075 5133
rect 12157 5128 15075 5130
rect 12157 5072 12162 5128
rect 12218 5072 15014 5128
rect 15070 5072 15075 5128
rect 12157 5070 15075 5072
rect 12157 5067 12223 5070
rect 15009 5067 15075 5070
rect 18413 5130 18479 5133
rect 19200 5130 20000 5160
rect 18413 5128 20000 5130
rect 18413 5072 18418 5128
rect 18474 5072 20000 5128
rect 18413 5070 20000 5072
rect 18413 5067 18479 5070
rect 19200 5040 20000 5070
rect 3170 4928 3486 4929
rect 0 4858 800 4888
rect 3170 4864 3176 4928
rect 3240 4864 3256 4928
rect 3320 4864 3336 4928
rect 3400 4864 3416 4928
rect 3480 4864 3486 4928
rect 3170 4863 3486 4864
rect 7618 4928 7934 4929
rect 7618 4864 7624 4928
rect 7688 4864 7704 4928
rect 7768 4864 7784 4928
rect 7848 4864 7864 4928
rect 7928 4864 7934 4928
rect 7618 4863 7934 4864
rect 12066 4928 12382 4929
rect 12066 4864 12072 4928
rect 12136 4864 12152 4928
rect 12216 4864 12232 4928
rect 12296 4864 12312 4928
rect 12376 4864 12382 4928
rect 12066 4863 12382 4864
rect 16514 4928 16830 4929
rect 16514 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16760 4928
rect 16824 4864 16830 4928
rect 16514 4863 16830 4864
rect 1485 4858 1551 4861
rect 0 4856 1551 4858
rect 0 4800 1490 4856
rect 1546 4800 1551 4856
rect 0 4798 1551 4800
rect 0 4768 800 4798
rect 1485 4795 1551 4798
rect 10041 4858 10107 4861
rect 11881 4858 11947 4861
rect 10041 4856 11947 4858
rect 10041 4800 10046 4856
rect 10102 4800 11886 4856
rect 11942 4800 11947 4856
rect 10041 4798 11947 4800
rect 10041 4795 10107 4798
rect 11881 4795 11947 4798
rect 12709 4858 12775 4861
rect 14273 4858 14339 4861
rect 12709 4856 14339 4858
rect 12709 4800 12714 4856
rect 12770 4800 14278 4856
rect 14334 4800 14339 4856
rect 12709 4798 14339 4800
rect 12709 4795 12775 4798
rect 14273 4795 14339 4798
rect 3785 4722 3851 4725
rect 9622 4722 9628 4724
rect 3785 4720 9628 4722
rect 3785 4664 3790 4720
rect 3846 4664 9628 4720
rect 3785 4662 9628 4664
rect 3785 4659 3851 4662
rect 9622 4660 9628 4662
rect 9692 4660 9698 4724
rect 10133 4722 10199 4725
rect 15101 4722 15167 4725
rect 10133 4720 15167 4722
rect 10133 4664 10138 4720
rect 10194 4664 15106 4720
rect 15162 4664 15167 4720
rect 10133 4662 15167 4664
rect 10133 4659 10199 4662
rect 15101 4659 15167 4662
rect 18045 4722 18111 4725
rect 19200 4722 20000 4752
rect 18045 4720 20000 4722
rect 18045 4664 18050 4720
rect 18106 4664 20000 4720
rect 18045 4662 20000 4664
rect 18045 4659 18111 4662
rect 19200 4632 20000 4662
rect 2313 4586 2379 4589
rect 4245 4586 4311 4589
rect 2313 4584 4311 4586
rect 2313 4528 2318 4584
rect 2374 4528 4250 4584
rect 4306 4528 4311 4584
rect 2313 4526 4311 4528
rect 2313 4523 2379 4526
rect 4245 4523 4311 4526
rect 7465 4586 7531 4589
rect 18505 4586 18571 4589
rect 7465 4584 18571 4586
rect 7465 4528 7470 4584
rect 7526 4528 18510 4584
rect 18566 4528 18571 4584
rect 7465 4526 18571 4528
rect 7465 4523 7531 4526
rect 18505 4523 18571 4526
rect 0 4450 800 4480
rect 1853 4450 1919 4453
rect 0 4448 1919 4450
rect 0 4392 1858 4448
rect 1914 4392 1919 4448
rect 0 4390 1919 4392
rect 0 4360 800 4390
rect 1853 4387 1919 4390
rect 5394 4384 5710 4385
rect 5394 4320 5400 4384
rect 5464 4320 5480 4384
rect 5544 4320 5560 4384
rect 5624 4320 5640 4384
rect 5704 4320 5710 4384
rect 5394 4319 5710 4320
rect 9842 4384 10158 4385
rect 9842 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10158 4384
rect 9842 4319 10158 4320
rect 14290 4384 14606 4385
rect 14290 4320 14296 4384
rect 14360 4320 14376 4384
rect 14440 4320 14456 4384
rect 14520 4320 14536 4384
rect 14600 4320 14606 4384
rect 14290 4319 14606 4320
rect 18413 4314 18479 4317
rect 19200 4314 20000 4344
rect 18413 4312 20000 4314
rect 18413 4256 18418 4312
rect 18474 4256 20000 4312
rect 18413 4254 20000 4256
rect 18413 4251 18479 4254
rect 19200 4224 20000 4254
rect 4061 4178 4127 4181
rect 13997 4178 14063 4181
rect 4061 4176 14063 4178
rect 4061 4120 4066 4176
rect 4122 4120 14002 4176
rect 14058 4120 14063 4176
rect 4061 4118 14063 4120
rect 4061 4115 4127 4118
rect 13997 4115 14063 4118
rect 0 4042 800 4072
rect 1485 4042 1551 4045
rect 0 4040 1551 4042
rect 0 3984 1490 4040
rect 1546 3984 1551 4040
rect 0 3982 1551 3984
rect 0 3952 800 3982
rect 1485 3979 1551 3982
rect 2773 4042 2839 4045
rect 3877 4042 3943 4045
rect 2773 4040 3943 4042
rect 2773 3984 2778 4040
rect 2834 3984 3882 4040
rect 3938 3984 3943 4040
rect 2773 3982 3943 3984
rect 2773 3979 2839 3982
rect 3877 3979 3943 3982
rect 8201 4042 8267 4045
rect 8702 4042 8708 4044
rect 8201 4040 8708 4042
rect 8201 3984 8206 4040
rect 8262 3984 8708 4040
rect 8201 3982 8708 3984
rect 8201 3979 8267 3982
rect 8702 3980 8708 3982
rect 8772 3980 8778 4044
rect 10869 4042 10935 4045
rect 14641 4042 14707 4045
rect 10869 4040 14707 4042
rect 10869 3984 10874 4040
rect 10930 3984 14646 4040
rect 14702 3984 14707 4040
rect 10869 3982 14707 3984
rect 10869 3979 10935 3982
rect 14641 3979 14707 3982
rect 18413 3906 18479 3909
rect 19200 3906 20000 3936
rect 18413 3904 20000 3906
rect 18413 3848 18418 3904
rect 18474 3848 20000 3904
rect 18413 3846 20000 3848
rect 18413 3843 18479 3846
rect 3170 3840 3486 3841
rect 3170 3776 3176 3840
rect 3240 3776 3256 3840
rect 3320 3776 3336 3840
rect 3400 3776 3416 3840
rect 3480 3776 3486 3840
rect 3170 3775 3486 3776
rect 7618 3840 7934 3841
rect 7618 3776 7624 3840
rect 7688 3776 7704 3840
rect 7768 3776 7784 3840
rect 7848 3776 7864 3840
rect 7928 3776 7934 3840
rect 7618 3775 7934 3776
rect 12066 3840 12382 3841
rect 12066 3776 12072 3840
rect 12136 3776 12152 3840
rect 12216 3776 12232 3840
rect 12296 3776 12312 3840
rect 12376 3776 12382 3840
rect 12066 3775 12382 3776
rect 16514 3840 16830 3841
rect 16514 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16760 3840
rect 16824 3776 16830 3840
rect 19200 3816 20000 3846
rect 16514 3775 16830 3776
rect 0 3634 800 3664
rect 1853 3634 1919 3637
rect 0 3632 1919 3634
rect 0 3576 1858 3632
rect 1914 3576 1919 3632
rect 0 3574 1919 3576
rect 0 3544 800 3574
rect 1853 3571 1919 3574
rect 3785 3634 3851 3637
rect 10225 3634 10291 3637
rect 17585 3634 17651 3637
rect 3785 3632 10291 3634
rect 3785 3576 3790 3632
rect 3846 3576 10230 3632
rect 10286 3576 10291 3632
rect 3785 3574 10291 3576
rect 3785 3571 3851 3574
rect 10225 3571 10291 3574
rect 10366 3632 17651 3634
rect 10366 3576 17590 3632
rect 17646 3576 17651 3632
rect 10366 3574 17651 3576
rect 6637 3498 6703 3501
rect 10366 3498 10426 3574
rect 17585 3571 17651 3574
rect 6637 3496 10426 3498
rect 6637 3440 6642 3496
rect 6698 3440 10426 3496
rect 6637 3438 10426 3440
rect 11697 3498 11763 3501
rect 17769 3498 17835 3501
rect 11697 3496 17835 3498
rect 11697 3440 11702 3496
rect 11758 3440 17774 3496
rect 17830 3440 17835 3496
rect 11697 3438 17835 3440
rect 6637 3435 6703 3438
rect 11697 3435 11763 3438
rect 17769 3435 17835 3438
rect 18413 3498 18479 3501
rect 19200 3498 20000 3528
rect 18413 3496 20000 3498
rect 18413 3440 18418 3496
rect 18474 3440 20000 3496
rect 18413 3438 20000 3440
rect 18413 3435 18479 3438
rect 19200 3408 20000 3438
rect 5394 3296 5710 3297
rect 0 3226 800 3256
rect 5394 3232 5400 3296
rect 5464 3232 5480 3296
rect 5544 3232 5560 3296
rect 5624 3232 5640 3296
rect 5704 3232 5710 3296
rect 5394 3231 5710 3232
rect 9842 3296 10158 3297
rect 9842 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10158 3296
rect 9842 3231 10158 3232
rect 14290 3296 14606 3297
rect 14290 3232 14296 3296
rect 14360 3232 14376 3296
rect 14440 3232 14456 3296
rect 14520 3232 14536 3296
rect 14600 3232 14606 3296
rect 14290 3231 14606 3232
rect 1485 3226 1551 3229
rect 0 3224 1551 3226
rect 0 3168 1490 3224
rect 1546 3168 1551 3224
rect 0 3166 1551 3168
rect 0 3136 800 3166
rect 1485 3163 1551 3166
rect 10317 3090 10383 3093
rect 14365 3090 14431 3093
rect 10317 3088 14431 3090
rect 10317 3032 10322 3088
rect 10378 3032 14370 3088
rect 14426 3032 14431 3088
rect 10317 3030 14431 3032
rect 10317 3027 10383 3030
rect 14365 3027 14431 3030
rect 18045 3090 18111 3093
rect 19200 3090 20000 3120
rect 18045 3088 20000 3090
rect 18045 3032 18050 3088
rect 18106 3032 20000 3088
rect 18045 3030 20000 3032
rect 18045 3027 18111 3030
rect 19200 3000 20000 3030
rect 3693 2954 3759 2957
rect 16113 2954 16179 2957
rect 3693 2952 16179 2954
rect 3693 2896 3698 2952
rect 3754 2896 16118 2952
rect 16174 2896 16179 2952
rect 3693 2894 16179 2896
rect 3693 2891 3759 2894
rect 16113 2891 16179 2894
rect 0 2818 800 2848
rect 1485 2818 1551 2821
rect 0 2816 1551 2818
rect 0 2760 1490 2816
rect 1546 2760 1551 2816
rect 0 2758 1551 2760
rect 0 2728 800 2758
rect 1485 2755 1551 2758
rect 3170 2752 3486 2753
rect 3170 2688 3176 2752
rect 3240 2688 3256 2752
rect 3320 2688 3336 2752
rect 3400 2688 3416 2752
rect 3480 2688 3486 2752
rect 3170 2687 3486 2688
rect 7618 2752 7934 2753
rect 7618 2688 7624 2752
rect 7688 2688 7704 2752
rect 7768 2688 7784 2752
rect 7848 2688 7864 2752
rect 7928 2688 7934 2752
rect 7618 2687 7934 2688
rect 12066 2752 12382 2753
rect 12066 2688 12072 2752
rect 12136 2688 12152 2752
rect 12216 2688 12232 2752
rect 12296 2688 12312 2752
rect 12376 2688 12382 2752
rect 12066 2687 12382 2688
rect 16514 2752 16830 2753
rect 16514 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16760 2752
rect 16824 2688 16830 2752
rect 16514 2687 16830 2688
rect 6545 2682 6611 2685
rect 6678 2682 6684 2684
rect 6545 2680 6684 2682
rect 6545 2624 6550 2680
rect 6606 2624 6684 2680
rect 6545 2622 6684 2624
rect 6545 2619 6611 2622
rect 6678 2620 6684 2622
rect 6748 2620 6754 2684
rect 18413 2682 18479 2685
rect 19200 2682 20000 2712
rect 18413 2680 20000 2682
rect 18413 2624 18418 2680
rect 18474 2624 20000 2680
rect 18413 2622 20000 2624
rect 18413 2619 18479 2622
rect 19200 2592 20000 2622
rect 0 2410 800 2440
rect 1853 2410 1919 2413
rect 0 2408 1919 2410
rect 0 2352 1858 2408
rect 1914 2352 1919 2408
rect 0 2350 1919 2352
rect 0 2320 800 2350
rect 1853 2347 1919 2350
rect 17861 2274 17927 2277
rect 19200 2274 20000 2304
rect 17861 2272 20000 2274
rect 17861 2216 17866 2272
rect 17922 2216 20000 2272
rect 17861 2214 20000 2216
rect 17861 2211 17927 2214
rect 5394 2208 5710 2209
rect 5394 2144 5400 2208
rect 5464 2144 5480 2208
rect 5544 2144 5560 2208
rect 5624 2144 5640 2208
rect 5704 2144 5710 2208
rect 5394 2143 5710 2144
rect 9842 2208 10158 2209
rect 9842 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10158 2208
rect 9842 2143 10158 2144
rect 14290 2208 14606 2209
rect 14290 2144 14296 2208
rect 14360 2144 14376 2208
rect 14440 2144 14456 2208
rect 14520 2144 14536 2208
rect 14600 2144 14606 2208
rect 19200 2184 20000 2214
rect 14290 2143 14606 2144
rect 0 2002 800 2032
rect 3509 2002 3575 2005
rect 0 2000 3575 2002
rect 0 1944 3514 2000
rect 3570 1944 3575 2000
rect 0 1942 3575 1944
rect 0 1912 800 1942
rect 3509 1939 3575 1942
rect 17585 1866 17651 1869
rect 19200 1866 20000 1896
rect 17585 1864 20000 1866
rect 17585 1808 17590 1864
rect 17646 1808 20000 1864
rect 17585 1806 20000 1808
rect 17585 1803 17651 1806
rect 19200 1776 20000 1806
rect 0 1594 800 1624
rect 2681 1594 2747 1597
rect 0 1592 2747 1594
rect 0 1536 2686 1592
rect 2742 1536 2747 1592
rect 0 1534 2747 1536
rect 0 1504 800 1534
rect 2681 1531 2747 1534
rect 16941 1458 17007 1461
rect 19200 1458 20000 1488
rect 16941 1456 20000 1458
rect 16941 1400 16946 1456
rect 17002 1400 20000 1456
rect 16941 1398 20000 1400
rect 16941 1395 17007 1398
rect 19200 1368 20000 1398
rect 0 1186 800 1216
rect 2865 1186 2931 1189
rect 0 1184 2931 1186
rect 0 1128 2870 1184
rect 2926 1128 2931 1184
rect 0 1126 2931 1128
rect 0 1096 800 1126
rect 2865 1123 2931 1126
rect 16297 1050 16363 1053
rect 19200 1050 20000 1080
rect 16297 1048 20000 1050
rect 16297 992 16302 1048
rect 16358 992 20000 1048
rect 16297 990 20000 992
rect 16297 987 16363 990
rect 19200 960 20000 990
rect 2221 914 2287 917
rect 1166 912 2287 914
rect 1166 856 2226 912
rect 2282 856 2287 912
rect 1166 854 2287 856
rect 0 778 800 808
rect 1166 778 1226 854
rect 2221 851 2287 854
rect 0 718 1226 778
rect 0 688 800 718
rect 18505 642 18571 645
rect 19200 642 20000 672
rect 18505 640 20000 642
rect 18505 584 18510 640
rect 18566 584 20000 640
rect 18505 582 20000 584
rect 18505 579 18571 582
rect 19200 552 20000 582
rect 0 370 800 400
rect 3969 370 4035 373
rect 0 368 4035 370
rect 0 312 3974 368
rect 4030 312 4035 368
rect 0 310 4035 312
rect 0 280 800 310
rect 3969 307 4035 310
<< via3 >>
rect 3176 14716 3240 14720
rect 3176 14660 3180 14716
rect 3180 14660 3236 14716
rect 3236 14660 3240 14716
rect 3176 14656 3240 14660
rect 3256 14716 3320 14720
rect 3256 14660 3260 14716
rect 3260 14660 3316 14716
rect 3316 14660 3320 14716
rect 3256 14656 3320 14660
rect 3336 14716 3400 14720
rect 3336 14660 3340 14716
rect 3340 14660 3396 14716
rect 3396 14660 3400 14716
rect 3336 14656 3400 14660
rect 3416 14716 3480 14720
rect 3416 14660 3420 14716
rect 3420 14660 3476 14716
rect 3476 14660 3480 14716
rect 3416 14656 3480 14660
rect 7624 14716 7688 14720
rect 7624 14660 7628 14716
rect 7628 14660 7684 14716
rect 7684 14660 7688 14716
rect 7624 14656 7688 14660
rect 7704 14716 7768 14720
rect 7704 14660 7708 14716
rect 7708 14660 7764 14716
rect 7764 14660 7768 14716
rect 7704 14656 7768 14660
rect 7784 14716 7848 14720
rect 7784 14660 7788 14716
rect 7788 14660 7844 14716
rect 7844 14660 7848 14716
rect 7784 14656 7848 14660
rect 7864 14716 7928 14720
rect 7864 14660 7868 14716
rect 7868 14660 7924 14716
rect 7924 14660 7928 14716
rect 7864 14656 7928 14660
rect 12072 14716 12136 14720
rect 12072 14660 12076 14716
rect 12076 14660 12132 14716
rect 12132 14660 12136 14716
rect 12072 14656 12136 14660
rect 12152 14716 12216 14720
rect 12152 14660 12156 14716
rect 12156 14660 12212 14716
rect 12212 14660 12216 14716
rect 12152 14656 12216 14660
rect 12232 14716 12296 14720
rect 12232 14660 12236 14716
rect 12236 14660 12292 14716
rect 12292 14660 12296 14716
rect 12232 14656 12296 14660
rect 12312 14716 12376 14720
rect 12312 14660 12316 14716
rect 12316 14660 12372 14716
rect 12372 14660 12376 14716
rect 12312 14656 12376 14660
rect 16520 14716 16584 14720
rect 16520 14660 16524 14716
rect 16524 14660 16580 14716
rect 16580 14660 16584 14716
rect 16520 14656 16584 14660
rect 16600 14716 16664 14720
rect 16600 14660 16604 14716
rect 16604 14660 16660 14716
rect 16660 14660 16664 14716
rect 16600 14656 16664 14660
rect 16680 14716 16744 14720
rect 16680 14660 16684 14716
rect 16684 14660 16740 14716
rect 16740 14660 16744 14716
rect 16680 14656 16744 14660
rect 16760 14716 16824 14720
rect 16760 14660 16764 14716
rect 16764 14660 16820 14716
rect 16820 14660 16824 14716
rect 16760 14656 16824 14660
rect 3004 14316 3068 14380
rect 5400 14172 5464 14176
rect 5400 14116 5404 14172
rect 5404 14116 5460 14172
rect 5460 14116 5464 14172
rect 5400 14112 5464 14116
rect 5480 14172 5544 14176
rect 5480 14116 5484 14172
rect 5484 14116 5540 14172
rect 5540 14116 5544 14172
rect 5480 14112 5544 14116
rect 5560 14172 5624 14176
rect 5560 14116 5564 14172
rect 5564 14116 5620 14172
rect 5620 14116 5624 14172
rect 5560 14112 5624 14116
rect 5640 14172 5704 14176
rect 5640 14116 5644 14172
rect 5644 14116 5700 14172
rect 5700 14116 5704 14172
rect 5640 14112 5704 14116
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 14296 14172 14360 14176
rect 14296 14116 14300 14172
rect 14300 14116 14356 14172
rect 14356 14116 14360 14172
rect 14296 14112 14360 14116
rect 14376 14172 14440 14176
rect 14376 14116 14380 14172
rect 14380 14116 14436 14172
rect 14436 14116 14440 14172
rect 14376 14112 14440 14116
rect 14456 14172 14520 14176
rect 14456 14116 14460 14172
rect 14460 14116 14516 14172
rect 14516 14116 14520 14172
rect 14456 14112 14520 14116
rect 14536 14172 14600 14176
rect 14536 14116 14540 14172
rect 14540 14116 14596 14172
rect 14596 14116 14600 14172
rect 14536 14112 14600 14116
rect 6684 13832 6748 13836
rect 6684 13776 6734 13832
rect 6734 13776 6748 13832
rect 6684 13772 6748 13776
rect 8708 13832 8772 13836
rect 8708 13776 8758 13832
rect 8758 13776 8772 13832
rect 8708 13772 8772 13776
rect 3176 13628 3240 13632
rect 3176 13572 3180 13628
rect 3180 13572 3236 13628
rect 3236 13572 3240 13628
rect 3176 13568 3240 13572
rect 3256 13628 3320 13632
rect 3256 13572 3260 13628
rect 3260 13572 3316 13628
rect 3316 13572 3320 13628
rect 3256 13568 3320 13572
rect 3336 13628 3400 13632
rect 3336 13572 3340 13628
rect 3340 13572 3396 13628
rect 3396 13572 3400 13628
rect 3336 13568 3400 13572
rect 3416 13628 3480 13632
rect 3416 13572 3420 13628
rect 3420 13572 3476 13628
rect 3476 13572 3480 13628
rect 3416 13568 3480 13572
rect 7624 13628 7688 13632
rect 7624 13572 7628 13628
rect 7628 13572 7684 13628
rect 7684 13572 7688 13628
rect 7624 13568 7688 13572
rect 7704 13628 7768 13632
rect 7704 13572 7708 13628
rect 7708 13572 7764 13628
rect 7764 13572 7768 13628
rect 7704 13568 7768 13572
rect 7784 13628 7848 13632
rect 7784 13572 7788 13628
rect 7788 13572 7844 13628
rect 7844 13572 7848 13628
rect 7784 13568 7848 13572
rect 7864 13628 7928 13632
rect 7864 13572 7868 13628
rect 7868 13572 7924 13628
rect 7924 13572 7928 13628
rect 7864 13568 7928 13572
rect 12072 13628 12136 13632
rect 12072 13572 12076 13628
rect 12076 13572 12132 13628
rect 12132 13572 12136 13628
rect 12072 13568 12136 13572
rect 12152 13628 12216 13632
rect 12152 13572 12156 13628
rect 12156 13572 12212 13628
rect 12212 13572 12216 13628
rect 12152 13568 12216 13572
rect 12232 13628 12296 13632
rect 12232 13572 12236 13628
rect 12236 13572 12292 13628
rect 12292 13572 12296 13628
rect 12232 13568 12296 13572
rect 12312 13628 12376 13632
rect 12312 13572 12316 13628
rect 12316 13572 12372 13628
rect 12372 13572 12376 13628
rect 12312 13568 12376 13572
rect 16520 13628 16584 13632
rect 16520 13572 16524 13628
rect 16524 13572 16580 13628
rect 16580 13572 16584 13628
rect 16520 13568 16584 13572
rect 16600 13628 16664 13632
rect 16600 13572 16604 13628
rect 16604 13572 16660 13628
rect 16660 13572 16664 13628
rect 16600 13568 16664 13572
rect 16680 13628 16744 13632
rect 16680 13572 16684 13628
rect 16684 13572 16740 13628
rect 16740 13572 16744 13628
rect 16680 13568 16744 13572
rect 16760 13628 16824 13632
rect 16760 13572 16764 13628
rect 16764 13572 16820 13628
rect 16820 13572 16824 13628
rect 16760 13568 16824 13572
rect 5400 13084 5464 13088
rect 5400 13028 5404 13084
rect 5404 13028 5460 13084
rect 5460 13028 5464 13084
rect 5400 13024 5464 13028
rect 5480 13084 5544 13088
rect 5480 13028 5484 13084
rect 5484 13028 5540 13084
rect 5540 13028 5544 13084
rect 5480 13024 5544 13028
rect 5560 13084 5624 13088
rect 5560 13028 5564 13084
rect 5564 13028 5620 13084
rect 5620 13028 5624 13084
rect 5560 13024 5624 13028
rect 5640 13084 5704 13088
rect 5640 13028 5644 13084
rect 5644 13028 5700 13084
rect 5700 13028 5704 13084
rect 5640 13024 5704 13028
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 14296 13084 14360 13088
rect 14296 13028 14300 13084
rect 14300 13028 14356 13084
rect 14356 13028 14360 13084
rect 14296 13024 14360 13028
rect 14376 13084 14440 13088
rect 14376 13028 14380 13084
rect 14380 13028 14436 13084
rect 14436 13028 14440 13084
rect 14376 13024 14440 13028
rect 14456 13084 14520 13088
rect 14456 13028 14460 13084
rect 14460 13028 14516 13084
rect 14516 13028 14520 13084
rect 14456 13024 14520 13028
rect 14536 13084 14600 13088
rect 14536 13028 14540 13084
rect 14540 13028 14596 13084
rect 14596 13028 14600 13084
rect 14536 13024 14600 13028
rect 3176 12540 3240 12544
rect 3176 12484 3180 12540
rect 3180 12484 3236 12540
rect 3236 12484 3240 12540
rect 3176 12480 3240 12484
rect 3256 12540 3320 12544
rect 3256 12484 3260 12540
rect 3260 12484 3316 12540
rect 3316 12484 3320 12540
rect 3256 12480 3320 12484
rect 3336 12540 3400 12544
rect 3336 12484 3340 12540
rect 3340 12484 3396 12540
rect 3396 12484 3400 12540
rect 3336 12480 3400 12484
rect 3416 12540 3480 12544
rect 3416 12484 3420 12540
rect 3420 12484 3476 12540
rect 3476 12484 3480 12540
rect 3416 12480 3480 12484
rect 7624 12540 7688 12544
rect 7624 12484 7628 12540
rect 7628 12484 7684 12540
rect 7684 12484 7688 12540
rect 7624 12480 7688 12484
rect 7704 12540 7768 12544
rect 7704 12484 7708 12540
rect 7708 12484 7764 12540
rect 7764 12484 7768 12540
rect 7704 12480 7768 12484
rect 7784 12540 7848 12544
rect 7784 12484 7788 12540
rect 7788 12484 7844 12540
rect 7844 12484 7848 12540
rect 7784 12480 7848 12484
rect 7864 12540 7928 12544
rect 7864 12484 7868 12540
rect 7868 12484 7924 12540
rect 7924 12484 7928 12540
rect 7864 12480 7928 12484
rect 12072 12540 12136 12544
rect 12072 12484 12076 12540
rect 12076 12484 12132 12540
rect 12132 12484 12136 12540
rect 12072 12480 12136 12484
rect 12152 12540 12216 12544
rect 12152 12484 12156 12540
rect 12156 12484 12212 12540
rect 12212 12484 12216 12540
rect 12152 12480 12216 12484
rect 12232 12540 12296 12544
rect 12232 12484 12236 12540
rect 12236 12484 12292 12540
rect 12292 12484 12296 12540
rect 12232 12480 12296 12484
rect 12312 12540 12376 12544
rect 12312 12484 12316 12540
rect 12316 12484 12372 12540
rect 12372 12484 12376 12540
rect 12312 12480 12376 12484
rect 16520 12540 16584 12544
rect 16520 12484 16524 12540
rect 16524 12484 16580 12540
rect 16580 12484 16584 12540
rect 16520 12480 16584 12484
rect 16600 12540 16664 12544
rect 16600 12484 16604 12540
rect 16604 12484 16660 12540
rect 16660 12484 16664 12540
rect 16600 12480 16664 12484
rect 16680 12540 16744 12544
rect 16680 12484 16684 12540
rect 16684 12484 16740 12540
rect 16740 12484 16744 12540
rect 16680 12480 16744 12484
rect 16760 12540 16824 12544
rect 16760 12484 16764 12540
rect 16764 12484 16820 12540
rect 16820 12484 16824 12540
rect 16760 12480 16824 12484
rect 17908 12336 17972 12340
rect 17908 12280 17922 12336
rect 17922 12280 17972 12336
rect 17908 12276 17972 12280
rect 5400 11996 5464 12000
rect 5400 11940 5404 11996
rect 5404 11940 5460 11996
rect 5460 11940 5464 11996
rect 5400 11936 5464 11940
rect 5480 11996 5544 12000
rect 5480 11940 5484 11996
rect 5484 11940 5540 11996
rect 5540 11940 5544 11996
rect 5480 11936 5544 11940
rect 5560 11996 5624 12000
rect 5560 11940 5564 11996
rect 5564 11940 5620 11996
rect 5620 11940 5624 11996
rect 5560 11936 5624 11940
rect 5640 11996 5704 12000
rect 5640 11940 5644 11996
rect 5644 11940 5700 11996
rect 5700 11940 5704 11996
rect 5640 11936 5704 11940
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 14296 11996 14360 12000
rect 14296 11940 14300 11996
rect 14300 11940 14356 11996
rect 14356 11940 14360 11996
rect 14296 11936 14360 11940
rect 14376 11996 14440 12000
rect 14376 11940 14380 11996
rect 14380 11940 14436 11996
rect 14436 11940 14440 11996
rect 14376 11936 14440 11940
rect 14456 11996 14520 12000
rect 14456 11940 14460 11996
rect 14460 11940 14516 11996
rect 14516 11940 14520 11996
rect 14456 11936 14520 11940
rect 14536 11996 14600 12000
rect 14536 11940 14540 11996
rect 14540 11940 14596 11996
rect 14596 11940 14600 11996
rect 14536 11936 14600 11940
rect 3004 11596 3068 11660
rect 3176 11452 3240 11456
rect 3176 11396 3180 11452
rect 3180 11396 3236 11452
rect 3236 11396 3240 11452
rect 3176 11392 3240 11396
rect 3256 11452 3320 11456
rect 3256 11396 3260 11452
rect 3260 11396 3316 11452
rect 3316 11396 3320 11452
rect 3256 11392 3320 11396
rect 3336 11452 3400 11456
rect 3336 11396 3340 11452
rect 3340 11396 3396 11452
rect 3396 11396 3400 11452
rect 3336 11392 3400 11396
rect 3416 11452 3480 11456
rect 3416 11396 3420 11452
rect 3420 11396 3476 11452
rect 3476 11396 3480 11452
rect 3416 11392 3480 11396
rect 7624 11452 7688 11456
rect 7624 11396 7628 11452
rect 7628 11396 7684 11452
rect 7684 11396 7688 11452
rect 7624 11392 7688 11396
rect 7704 11452 7768 11456
rect 7704 11396 7708 11452
rect 7708 11396 7764 11452
rect 7764 11396 7768 11452
rect 7704 11392 7768 11396
rect 7784 11452 7848 11456
rect 7784 11396 7788 11452
rect 7788 11396 7844 11452
rect 7844 11396 7848 11452
rect 7784 11392 7848 11396
rect 7864 11452 7928 11456
rect 7864 11396 7868 11452
rect 7868 11396 7924 11452
rect 7924 11396 7928 11452
rect 7864 11392 7928 11396
rect 12072 11452 12136 11456
rect 12072 11396 12076 11452
rect 12076 11396 12132 11452
rect 12132 11396 12136 11452
rect 12072 11392 12136 11396
rect 12152 11452 12216 11456
rect 12152 11396 12156 11452
rect 12156 11396 12212 11452
rect 12212 11396 12216 11452
rect 12152 11392 12216 11396
rect 12232 11452 12296 11456
rect 12232 11396 12236 11452
rect 12236 11396 12292 11452
rect 12292 11396 12296 11452
rect 12232 11392 12296 11396
rect 12312 11452 12376 11456
rect 12312 11396 12316 11452
rect 12316 11396 12372 11452
rect 12372 11396 12376 11452
rect 12312 11392 12376 11396
rect 16520 11452 16584 11456
rect 16520 11396 16524 11452
rect 16524 11396 16580 11452
rect 16580 11396 16584 11452
rect 16520 11392 16584 11396
rect 16600 11452 16664 11456
rect 16600 11396 16604 11452
rect 16604 11396 16660 11452
rect 16660 11396 16664 11452
rect 16600 11392 16664 11396
rect 16680 11452 16744 11456
rect 16680 11396 16684 11452
rect 16684 11396 16740 11452
rect 16740 11396 16744 11452
rect 16680 11392 16744 11396
rect 16760 11452 16824 11456
rect 16760 11396 16764 11452
rect 16764 11396 16820 11452
rect 16820 11396 16824 11452
rect 16760 11392 16824 11396
rect 9628 11052 9692 11116
rect 5400 10908 5464 10912
rect 5400 10852 5404 10908
rect 5404 10852 5460 10908
rect 5460 10852 5464 10908
rect 5400 10848 5464 10852
rect 5480 10908 5544 10912
rect 5480 10852 5484 10908
rect 5484 10852 5540 10908
rect 5540 10852 5544 10908
rect 5480 10848 5544 10852
rect 5560 10908 5624 10912
rect 5560 10852 5564 10908
rect 5564 10852 5620 10908
rect 5620 10852 5624 10908
rect 5560 10848 5624 10852
rect 5640 10908 5704 10912
rect 5640 10852 5644 10908
rect 5644 10852 5700 10908
rect 5700 10852 5704 10908
rect 5640 10848 5704 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 14296 10908 14360 10912
rect 14296 10852 14300 10908
rect 14300 10852 14356 10908
rect 14356 10852 14360 10908
rect 14296 10848 14360 10852
rect 14376 10908 14440 10912
rect 14376 10852 14380 10908
rect 14380 10852 14436 10908
rect 14436 10852 14440 10908
rect 14376 10848 14440 10852
rect 14456 10908 14520 10912
rect 14456 10852 14460 10908
rect 14460 10852 14516 10908
rect 14516 10852 14520 10908
rect 14456 10848 14520 10852
rect 14536 10908 14600 10912
rect 14536 10852 14540 10908
rect 14540 10852 14596 10908
rect 14596 10852 14600 10908
rect 14536 10848 14600 10852
rect 3176 10364 3240 10368
rect 3176 10308 3180 10364
rect 3180 10308 3236 10364
rect 3236 10308 3240 10364
rect 3176 10304 3240 10308
rect 3256 10364 3320 10368
rect 3256 10308 3260 10364
rect 3260 10308 3316 10364
rect 3316 10308 3320 10364
rect 3256 10304 3320 10308
rect 3336 10364 3400 10368
rect 3336 10308 3340 10364
rect 3340 10308 3396 10364
rect 3396 10308 3400 10364
rect 3336 10304 3400 10308
rect 3416 10364 3480 10368
rect 3416 10308 3420 10364
rect 3420 10308 3476 10364
rect 3476 10308 3480 10364
rect 3416 10304 3480 10308
rect 7624 10364 7688 10368
rect 7624 10308 7628 10364
rect 7628 10308 7684 10364
rect 7684 10308 7688 10364
rect 7624 10304 7688 10308
rect 7704 10364 7768 10368
rect 7704 10308 7708 10364
rect 7708 10308 7764 10364
rect 7764 10308 7768 10364
rect 7704 10304 7768 10308
rect 7784 10364 7848 10368
rect 7784 10308 7788 10364
rect 7788 10308 7844 10364
rect 7844 10308 7848 10364
rect 7784 10304 7848 10308
rect 7864 10364 7928 10368
rect 7864 10308 7868 10364
rect 7868 10308 7924 10364
rect 7924 10308 7928 10364
rect 7864 10304 7928 10308
rect 12072 10364 12136 10368
rect 12072 10308 12076 10364
rect 12076 10308 12132 10364
rect 12132 10308 12136 10364
rect 12072 10304 12136 10308
rect 12152 10364 12216 10368
rect 12152 10308 12156 10364
rect 12156 10308 12212 10364
rect 12212 10308 12216 10364
rect 12152 10304 12216 10308
rect 12232 10364 12296 10368
rect 12232 10308 12236 10364
rect 12236 10308 12292 10364
rect 12292 10308 12296 10364
rect 12232 10304 12296 10308
rect 12312 10364 12376 10368
rect 12312 10308 12316 10364
rect 12316 10308 12372 10364
rect 12372 10308 12376 10364
rect 12312 10304 12376 10308
rect 16520 10364 16584 10368
rect 16520 10308 16524 10364
rect 16524 10308 16580 10364
rect 16580 10308 16584 10364
rect 16520 10304 16584 10308
rect 16600 10364 16664 10368
rect 16600 10308 16604 10364
rect 16604 10308 16660 10364
rect 16660 10308 16664 10364
rect 16600 10304 16664 10308
rect 16680 10364 16744 10368
rect 16680 10308 16684 10364
rect 16684 10308 16740 10364
rect 16740 10308 16744 10364
rect 16680 10304 16744 10308
rect 16760 10364 16824 10368
rect 16760 10308 16764 10364
rect 16764 10308 16820 10364
rect 16820 10308 16824 10364
rect 16760 10304 16824 10308
rect 5400 9820 5464 9824
rect 5400 9764 5404 9820
rect 5404 9764 5460 9820
rect 5460 9764 5464 9820
rect 5400 9760 5464 9764
rect 5480 9820 5544 9824
rect 5480 9764 5484 9820
rect 5484 9764 5540 9820
rect 5540 9764 5544 9820
rect 5480 9760 5544 9764
rect 5560 9820 5624 9824
rect 5560 9764 5564 9820
rect 5564 9764 5620 9820
rect 5620 9764 5624 9820
rect 5560 9760 5624 9764
rect 5640 9820 5704 9824
rect 5640 9764 5644 9820
rect 5644 9764 5700 9820
rect 5700 9764 5704 9820
rect 5640 9760 5704 9764
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 14296 9820 14360 9824
rect 14296 9764 14300 9820
rect 14300 9764 14356 9820
rect 14356 9764 14360 9820
rect 14296 9760 14360 9764
rect 14376 9820 14440 9824
rect 14376 9764 14380 9820
rect 14380 9764 14436 9820
rect 14436 9764 14440 9820
rect 14376 9760 14440 9764
rect 14456 9820 14520 9824
rect 14456 9764 14460 9820
rect 14460 9764 14516 9820
rect 14516 9764 14520 9820
rect 14456 9760 14520 9764
rect 14536 9820 14600 9824
rect 14536 9764 14540 9820
rect 14540 9764 14596 9820
rect 14596 9764 14600 9820
rect 14536 9760 14600 9764
rect 3176 9276 3240 9280
rect 3176 9220 3180 9276
rect 3180 9220 3236 9276
rect 3236 9220 3240 9276
rect 3176 9216 3240 9220
rect 3256 9276 3320 9280
rect 3256 9220 3260 9276
rect 3260 9220 3316 9276
rect 3316 9220 3320 9276
rect 3256 9216 3320 9220
rect 3336 9276 3400 9280
rect 3336 9220 3340 9276
rect 3340 9220 3396 9276
rect 3396 9220 3400 9276
rect 3336 9216 3400 9220
rect 3416 9276 3480 9280
rect 3416 9220 3420 9276
rect 3420 9220 3476 9276
rect 3476 9220 3480 9276
rect 3416 9216 3480 9220
rect 7624 9276 7688 9280
rect 7624 9220 7628 9276
rect 7628 9220 7684 9276
rect 7684 9220 7688 9276
rect 7624 9216 7688 9220
rect 7704 9276 7768 9280
rect 7704 9220 7708 9276
rect 7708 9220 7764 9276
rect 7764 9220 7768 9276
rect 7704 9216 7768 9220
rect 7784 9276 7848 9280
rect 7784 9220 7788 9276
rect 7788 9220 7844 9276
rect 7844 9220 7848 9276
rect 7784 9216 7848 9220
rect 7864 9276 7928 9280
rect 7864 9220 7868 9276
rect 7868 9220 7924 9276
rect 7924 9220 7928 9276
rect 7864 9216 7928 9220
rect 12072 9276 12136 9280
rect 12072 9220 12076 9276
rect 12076 9220 12132 9276
rect 12132 9220 12136 9276
rect 12072 9216 12136 9220
rect 12152 9276 12216 9280
rect 12152 9220 12156 9276
rect 12156 9220 12212 9276
rect 12212 9220 12216 9276
rect 12152 9216 12216 9220
rect 12232 9276 12296 9280
rect 12232 9220 12236 9276
rect 12236 9220 12292 9276
rect 12292 9220 12296 9276
rect 12232 9216 12296 9220
rect 12312 9276 12376 9280
rect 12312 9220 12316 9276
rect 12316 9220 12372 9276
rect 12372 9220 12376 9276
rect 12312 9216 12376 9220
rect 16520 9276 16584 9280
rect 16520 9220 16524 9276
rect 16524 9220 16580 9276
rect 16580 9220 16584 9276
rect 16520 9216 16584 9220
rect 16600 9276 16664 9280
rect 16600 9220 16604 9276
rect 16604 9220 16660 9276
rect 16660 9220 16664 9276
rect 16600 9216 16664 9220
rect 16680 9276 16744 9280
rect 16680 9220 16684 9276
rect 16684 9220 16740 9276
rect 16740 9220 16744 9276
rect 16680 9216 16744 9220
rect 16760 9276 16824 9280
rect 16760 9220 16764 9276
rect 16764 9220 16820 9276
rect 16820 9220 16824 9276
rect 16760 9216 16824 9220
rect 5400 8732 5464 8736
rect 5400 8676 5404 8732
rect 5404 8676 5460 8732
rect 5460 8676 5464 8732
rect 5400 8672 5464 8676
rect 5480 8732 5544 8736
rect 5480 8676 5484 8732
rect 5484 8676 5540 8732
rect 5540 8676 5544 8732
rect 5480 8672 5544 8676
rect 5560 8732 5624 8736
rect 5560 8676 5564 8732
rect 5564 8676 5620 8732
rect 5620 8676 5624 8732
rect 5560 8672 5624 8676
rect 5640 8732 5704 8736
rect 5640 8676 5644 8732
rect 5644 8676 5700 8732
rect 5700 8676 5704 8732
rect 5640 8672 5704 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 14296 8732 14360 8736
rect 14296 8676 14300 8732
rect 14300 8676 14356 8732
rect 14356 8676 14360 8732
rect 14296 8672 14360 8676
rect 14376 8732 14440 8736
rect 14376 8676 14380 8732
rect 14380 8676 14436 8732
rect 14436 8676 14440 8732
rect 14376 8672 14440 8676
rect 14456 8732 14520 8736
rect 14456 8676 14460 8732
rect 14460 8676 14516 8732
rect 14516 8676 14520 8732
rect 14456 8672 14520 8676
rect 14536 8732 14600 8736
rect 14536 8676 14540 8732
rect 14540 8676 14596 8732
rect 14596 8676 14600 8732
rect 14536 8672 14600 8676
rect 17908 8392 17972 8396
rect 17908 8336 17922 8392
rect 17922 8336 17972 8392
rect 17908 8332 17972 8336
rect 3176 8188 3240 8192
rect 3176 8132 3180 8188
rect 3180 8132 3236 8188
rect 3236 8132 3240 8188
rect 3176 8128 3240 8132
rect 3256 8188 3320 8192
rect 3256 8132 3260 8188
rect 3260 8132 3316 8188
rect 3316 8132 3320 8188
rect 3256 8128 3320 8132
rect 3336 8188 3400 8192
rect 3336 8132 3340 8188
rect 3340 8132 3396 8188
rect 3396 8132 3400 8188
rect 3336 8128 3400 8132
rect 3416 8188 3480 8192
rect 3416 8132 3420 8188
rect 3420 8132 3476 8188
rect 3476 8132 3480 8188
rect 3416 8128 3480 8132
rect 7624 8188 7688 8192
rect 7624 8132 7628 8188
rect 7628 8132 7684 8188
rect 7684 8132 7688 8188
rect 7624 8128 7688 8132
rect 7704 8188 7768 8192
rect 7704 8132 7708 8188
rect 7708 8132 7764 8188
rect 7764 8132 7768 8188
rect 7704 8128 7768 8132
rect 7784 8188 7848 8192
rect 7784 8132 7788 8188
rect 7788 8132 7844 8188
rect 7844 8132 7848 8188
rect 7784 8128 7848 8132
rect 7864 8188 7928 8192
rect 7864 8132 7868 8188
rect 7868 8132 7924 8188
rect 7924 8132 7928 8188
rect 7864 8128 7928 8132
rect 12072 8188 12136 8192
rect 12072 8132 12076 8188
rect 12076 8132 12132 8188
rect 12132 8132 12136 8188
rect 12072 8128 12136 8132
rect 12152 8188 12216 8192
rect 12152 8132 12156 8188
rect 12156 8132 12212 8188
rect 12212 8132 12216 8188
rect 12152 8128 12216 8132
rect 12232 8188 12296 8192
rect 12232 8132 12236 8188
rect 12236 8132 12292 8188
rect 12292 8132 12296 8188
rect 12232 8128 12296 8132
rect 12312 8188 12376 8192
rect 12312 8132 12316 8188
rect 12316 8132 12372 8188
rect 12372 8132 12376 8188
rect 12312 8128 12376 8132
rect 16520 8188 16584 8192
rect 16520 8132 16524 8188
rect 16524 8132 16580 8188
rect 16580 8132 16584 8188
rect 16520 8128 16584 8132
rect 16600 8188 16664 8192
rect 16600 8132 16604 8188
rect 16604 8132 16660 8188
rect 16660 8132 16664 8188
rect 16600 8128 16664 8132
rect 16680 8188 16744 8192
rect 16680 8132 16684 8188
rect 16684 8132 16740 8188
rect 16740 8132 16744 8188
rect 16680 8128 16744 8132
rect 16760 8188 16824 8192
rect 16760 8132 16764 8188
rect 16764 8132 16820 8188
rect 16820 8132 16824 8188
rect 16760 8128 16824 8132
rect 5400 7644 5464 7648
rect 5400 7588 5404 7644
rect 5404 7588 5460 7644
rect 5460 7588 5464 7644
rect 5400 7584 5464 7588
rect 5480 7644 5544 7648
rect 5480 7588 5484 7644
rect 5484 7588 5540 7644
rect 5540 7588 5544 7644
rect 5480 7584 5544 7588
rect 5560 7644 5624 7648
rect 5560 7588 5564 7644
rect 5564 7588 5620 7644
rect 5620 7588 5624 7644
rect 5560 7584 5624 7588
rect 5640 7644 5704 7648
rect 5640 7588 5644 7644
rect 5644 7588 5700 7644
rect 5700 7588 5704 7644
rect 5640 7584 5704 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 14296 7644 14360 7648
rect 14296 7588 14300 7644
rect 14300 7588 14356 7644
rect 14356 7588 14360 7644
rect 14296 7584 14360 7588
rect 14376 7644 14440 7648
rect 14376 7588 14380 7644
rect 14380 7588 14436 7644
rect 14436 7588 14440 7644
rect 14376 7584 14440 7588
rect 14456 7644 14520 7648
rect 14456 7588 14460 7644
rect 14460 7588 14516 7644
rect 14516 7588 14520 7644
rect 14456 7584 14520 7588
rect 14536 7644 14600 7648
rect 14536 7588 14540 7644
rect 14540 7588 14596 7644
rect 14596 7588 14600 7644
rect 14536 7584 14600 7588
rect 3004 7244 3068 7308
rect 3176 7100 3240 7104
rect 3176 7044 3180 7100
rect 3180 7044 3236 7100
rect 3236 7044 3240 7100
rect 3176 7040 3240 7044
rect 3256 7100 3320 7104
rect 3256 7044 3260 7100
rect 3260 7044 3316 7100
rect 3316 7044 3320 7100
rect 3256 7040 3320 7044
rect 3336 7100 3400 7104
rect 3336 7044 3340 7100
rect 3340 7044 3396 7100
rect 3396 7044 3400 7100
rect 3336 7040 3400 7044
rect 3416 7100 3480 7104
rect 3416 7044 3420 7100
rect 3420 7044 3476 7100
rect 3476 7044 3480 7100
rect 3416 7040 3480 7044
rect 7624 7100 7688 7104
rect 7624 7044 7628 7100
rect 7628 7044 7684 7100
rect 7684 7044 7688 7100
rect 7624 7040 7688 7044
rect 7704 7100 7768 7104
rect 7704 7044 7708 7100
rect 7708 7044 7764 7100
rect 7764 7044 7768 7100
rect 7704 7040 7768 7044
rect 7784 7100 7848 7104
rect 7784 7044 7788 7100
rect 7788 7044 7844 7100
rect 7844 7044 7848 7100
rect 7784 7040 7848 7044
rect 7864 7100 7928 7104
rect 7864 7044 7868 7100
rect 7868 7044 7924 7100
rect 7924 7044 7928 7100
rect 7864 7040 7928 7044
rect 12072 7100 12136 7104
rect 12072 7044 12076 7100
rect 12076 7044 12132 7100
rect 12132 7044 12136 7100
rect 12072 7040 12136 7044
rect 12152 7100 12216 7104
rect 12152 7044 12156 7100
rect 12156 7044 12212 7100
rect 12212 7044 12216 7100
rect 12152 7040 12216 7044
rect 12232 7100 12296 7104
rect 12232 7044 12236 7100
rect 12236 7044 12292 7100
rect 12292 7044 12296 7100
rect 12232 7040 12296 7044
rect 12312 7100 12376 7104
rect 12312 7044 12316 7100
rect 12316 7044 12372 7100
rect 12372 7044 12376 7100
rect 12312 7040 12376 7044
rect 16520 7100 16584 7104
rect 16520 7044 16524 7100
rect 16524 7044 16580 7100
rect 16580 7044 16584 7100
rect 16520 7040 16584 7044
rect 16600 7100 16664 7104
rect 16600 7044 16604 7100
rect 16604 7044 16660 7100
rect 16660 7044 16664 7100
rect 16600 7040 16664 7044
rect 16680 7100 16744 7104
rect 16680 7044 16684 7100
rect 16684 7044 16740 7100
rect 16740 7044 16744 7100
rect 16680 7040 16744 7044
rect 16760 7100 16824 7104
rect 16760 7044 16764 7100
rect 16764 7044 16820 7100
rect 16820 7044 16824 7100
rect 16760 7040 16824 7044
rect 5400 6556 5464 6560
rect 5400 6500 5404 6556
rect 5404 6500 5460 6556
rect 5460 6500 5464 6556
rect 5400 6496 5464 6500
rect 5480 6556 5544 6560
rect 5480 6500 5484 6556
rect 5484 6500 5540 6556
rect 5540 6500 5544 6556
rect 5480 6496 5544 6500
rect 5560 6556 5624 6560
rect 5560 6500 5564 6556
rect 5564 6500 5620 6556
rect 5620 6500 5624 6556
rect 5560 6496 5624 6500
rect 5640 6556 5704 6560
rect 5640 6500 5644 6556
rect 5644 6500 5700 6556
rect 5700 6500 5704 6556
rect 5640 6496 5704 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 14296 6556 14360 6560
rect 14296 6500 14300 6556
rect 14300 6500 14356 6556
rect 14356 6500 14360 6556
rect 14296 6496 14360 6500
rect 14376 6556 14440 6560
rect 14376 6500 14380 6556
rect 14380 6500 14436 6556
rect 14436 6500 14440 6556
rect 14376 6496 14440 6500
rect 14456 6556 14520 6560
rect 14456 6500 14460 6556
rect 14460 6500 14516 6556
rect 14516 6500 14520 6556
rect 14456 6496 14520 6500
rect 14536 6556 14600 6560
rect 14536 6500 14540 6556
rect 14540 6500 14596 6556
rect 14596 6500 14600 6556
rect 14536 6496 14600 6500
rect 3176 6012 3240 6016
rect 3176 5956 3180 6012
rect 3180 5956 3236 6012
rect 3236 5956 3240 6012
rect 3176 5952 3240 5956
rect 3256 6012 3320 6016
rect 3256 5956 3260 6012
rect 3260 5956 3316 6012
rect 3316 5956 3320 6012
rect 3256 5952 3320 5956
rect 3336 6012 3400 6016
rect 3336 5956 3340 6012
rect 3340 5956 3396 6012
rect 3396 5956 3400 6012
rect 3336 5952 3400 5956
rect 3416 6012 3480 6016
rect 3416 5956 3420 6012
rect 3420 5956 3476 6012
rect 3476 5956 3480 6012
rect 3416 5952 3480 5956
rect 7624 6012 7688 6016
rect 7624 5956 7628 6012
rect 7628 5956 7684 6012
rect 7684 5956 7688 6012
rect 7624 5952 7688 5956
rect 7704 6012 7768 6016
rect 7704 5956 7708 6012
rect 7708 5956 7764 6012
rect 7764 5956 7768 6012
rect 7704 5952 7768 5956
rect 7784 6012 7848 6016
rect 7784 5956 7788 6012
rect 7788 5956 7844 6012
rect 7844 5956 7848 6012
rect 7784 5952 7848 5956
rect 7864 6012 7928 6016
rect 7864 5956 7868 6012
rect 7868 5956 7924 6012
rect 7924 5956 7928 6012
rect 7864 5952 7928 5956
rect 12072 6012 12136 6016
rect 12072 5956 12076 6012
rect 12076 5956 12132 6012
rect 12132 5956 12136 6012
rect 12072 5952 12136 5956
rect 12152 6012 12216 6016
rect 12152 5956 12156 6012
rect 12156 5956 12212 6012
rect 12212 5956 12216 6012
rect 12152 5952 12216 5956
rect 12232 6012 12296 6016
rect 12232 5956 12236 6012
rect 12236 5956 12292 6012
rect 12292 5956 12296 6012
rect 12232 5952 12296 5956
rect 12312 6012 12376 6016
rect 12312 5956 12316 6012
rect 12316 5956 12372 6012
rect 12372 5956 12376 6012
rect 12312 5952 12376 5956
rect 16520 6012 16584 6016
rect 16520 5956 16524 6012
rect 16524 5956 16580 6012
rect 16580 5956 16584 6012
rect 16520 5952 16584 5956
rect 16600 6012 16664 6016
rect 16600 5956 16604 6012
rect 16604 5956 16660 6012
rect 16660 5956 16664 6012
rect 16600 5952 16664 5956
rect 16680 6012 16744 6016
rect 16680 5956 16684 6012
rect 16684 5956 16740 6012
rect 16740 5956 16744 6012
rect 16680 5952 16744 5956
rect 16760 6012 16824 6016
rect 16760 5956 16764 6012
rect 16764 5956 16820 6012
rect 16820 5956 16824 6012
rect 16760 5952 16824 5956
rect 2820 5476 2884 5540
rect 5400 5468 5464 5472
rect 5400 5412 5404 5468
rect 5404 5412 5460 5468
rect 5460 5412 5464 5468
rect 5400 5408 5464 5412
rect 5480 5468 5544 5472
rect 5480 5412 5484 5468
rect 5484 5412 5540 5468
rect 5540 5412 5544 5468
rect 5480 5408 5544 5412
rect 5560 5468 5624 5472
rect 5560 5412 5564 5468
rect 5564 5412 5620 5468
rect 5620 5412 5624 5468
rect 5560 5408 5624 5412
rect 5640 5468 5704 5472
rect 5640 5412 5644 5468
rect 5644 5412 5700 5468
rect 5700 5412 5704 5468
rect 5640 5408 5704 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 14296 5468 14360 5472
rect 14296 5412 14300 5468
rect 14300 5412 14356 5468
rect 14356 5412 14360 5468
rect 14296 5408 14360 5412
rect 14376 5468 14440 5472
rect 14376 5412 14380 5468
rect 14380 5412 14436 5468
rect 14436 5412 14440 5468
rect 14376 5408 14440 5412
rect 14456 5468 14520 5472
rect 14456 5412 14460 5468
rect 14460 5412 14516 5468
rect 14516 5412 14520 5468
rect 14456 5408 14520 5412
rect 14536 5468 14600 5472
rect 14536 5412 14540 5468
rect 14540 5412 14596 5468
rect 14596 5412 14600 5468
rect 14536 5408 14600 5412
rect 3176 4924 3240 4928
rect 3176 4868 3180 4924
rect 3180 4868 3236 4924
rect 3236 4868 3240 4924
rect 3176 4864 3240 4868
rect 3256 4924 3320 4928
rect 3256 4868 3260 4924
rect 3260 4868 3316 4924
rect 3316 4868 3320 4924
rect 3256 4864 3320 4868
rect 3336 4924 3400 4928
rect 3336 4868 3340 4924
rect 3340 4868 3396 4924
rect 3396 4868 3400 4924
rect 3336 4864 3400 4868
rect 3416 4924 3480 4928
rect 3416 4868 3420 4924
rect 3420 4868 3476 4924
rect 3476 4868 3480 4924
rect 3416 4864 3480 4868
rect 7624 4924 7688 4928
rect 7624 4868 7628 4924
rect 7628 4868 7684 4924
rect 7684 4868 7688 4924
rect 7624 4864 7688 4868
rect 7704 4924 7768 4928
rect 7704 4868 7708 4924
rect 7708 4868 7764 4924
rect 7764 4868 7768 4924
rect 7704 4864 7768 4868
rect 7784 4924 7848 4928
rect 7784 4868 7788 4924
rect 7788 4868 7844 4924
rect 7844 4868 7848 4924
rect 7784 4864 7848 4868
rect 7864 4924 7928 4928
rect 7864 4868 7868 4924
rect 7868 4868 7924 4924
rect 7924 4868 7928 4924
rect 7864 4864 7928 4868
rect 12072 4924 12136 4928
rect 12072 4868 12076 4924
rect 12076 4868 12132 4924
rect 12132 4868 12136 4924
rect 12072 4864 12136 4868
rect 12152 4924 12216 4928
rect 12152 4868 12156 4924
rect 12156 4868 12212 4924
rect 12212 4868 12216 4924
rect 12152 4864 12216 4868
rect 12232 4924 12296 4928
rect 12232 4868 12236 4924
rect 12236 4868 12292 4924
rect 12292 4868 12296 4924
rect 12232 4864 12296 4868
rect 12312 4924 12376 4928
rect 12312 4868 12316 4924
rect 12316 4868 12372 4924
rect 12372 4868 12376 4924
rect 12312 4864 12376 4868
rect 16520 4924 16584 4928
rect 16520 4868 16524 4924
rect 16524 4868 16580 4924
rect 16580 4868 16584 4924
rect 16520 4864 16584 4868
rect 16600 4924 16664 4928
rect 16600 4868 16604 4924
rect 16604 4868 16660 4924
rect 16660 4868 16664 4924
rect 16600 4864 16664 4868
rect 16680 4924 16744 4928
rect 16680 4868 16684 4924
rect 16684 4868 16740 4924
rect 16740 4868 16744 4924
rect 16680 4864 16744 4868
rect 16760 4924 16824 4928
rect 16760 4868 16764 4924
rect 16764 4868 16820 4924
rect 16820 4868 16824 4924
rect 16760 4864 16824 4868
rect 9628 4660 9692 4724
rect 5400 4380 5464 4384
rect 5400 4324 5404 4380
rect 5404 4324 5460 4380
rect 5460 4324 5464 4380
rect 5400 4320 5464 4324
rect 5480 4380 5544 4384
rect 5480 4324 5484 4380
rect 5484 4324 5540 4380
rect 5540 4324 5544 4380
rect 5480 4320 5544 4324
rect 5560 4380 5624 4384
rect 5560 4324 5564 4380
rect 5564 4324 5620 4380
rect 5620 4324 5624 4380
rect 5560 4320 5624 4324
rect 5640 4380 5704 4384
rect 5640 4324 5644 4380
rect 5644 4324 5700 4380
rect 5700 4324 5704 4380
rect 5640 4320 5704 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 14296 4380 14360 4384
rect 14296 4324 14300 4380
rect 14300 4324 14356 4380
rect 14356 4324 14360 4380
rect 14296 4320 14360 4324
rect 14376 4380 14440 4384
rect 14376 4324 14380 4380
rect 14380 4324 14436 4380
rect 14436 4324 14440 4380
rect 14376 4320 14440 4324
rect 14456 4380 14520 4384
rect 14456 4324 14460 4380
rect 14460 4324 14516 4380
rect 14516 4324 14520 4380
rect 14456 4320 14520 4324
rect 14536 4380 14600 4384
rect 14536 4324 14540 4380
rect 14540 4324 14596 4380
rect 14596 4324 14600 4380
rect 14536 4320 14600 4324
rect 8708 3980 8772 4044
rect 3176 3836 3240 3840
rect 3176 3780 3180 3836
rect 3180 3780 3236 3836
rect 3236 3780 3240 3836
rect 3176 3776 3240 3780
rect 3256 3836 3320 3840
rect 3256 3780 3260 3836
rect 3260 3780 3316 3836
rect 3316 3780 3320 3836
rect 3256 3776 3320 3780
rect 3336 3836 3400 3840
rect 3336 3780 3340 3836
rect 3340 3780 3396 3836
rect 3396 3780 3400 3836
rect 3336 3776 3400 3780
rect 3416 3836 3480 3840
rect 3416 3780 3420 3836
rect 3420 3780 3476 3836
rect 3476 3780 3480 3836
rect 3416 3776 3480 3780
rect 7624 3836 7688 3840
rect 7624 3780 7628 3836
rect 7628 3780 7684 3836
rect 7684 3780 7688 3836
rect 7624 3776 7688 3780
rect 7704 3836 7768 3840
rect 7704 3780 7708 3836
rect 7708 3780 7764 3836
rect 7764 3780 7768 3836
rect 7704 3776 7768 3780
rect 7784 3836 7848 3840
rect 7784 3780 7788 3836
rect 7788 3780 7844 3836
rect 7844 3780 7848 3836
rect 7784 3776 7848 3780
rect 7864 3836 7928 3840
rect 7864 3780 7868 3836
rect 7868 3780 7924 3836
rect 7924 3780 7928 3836
rect 7864 3776 7928 3780
rect 12072 3836 12136 3840
rect 12072 3780 12076 3836
rect 12076 3780 12132 3836
rect 12132 3780 12136 3836
rect 12072 3776 12136 3780
rect 12152 3836 12216 3840
rect 12152 3780 12156 3836
rect 12156 3780 12212 3836
rect 12212 3780 12216 3836
rect 12152 3776 12216 3780
rect 12232 3836 12296 3840
rect 12232 3780 12236 3836
rect 12236 3780 12292 3836
rect 12292 3780 12296 3836
rect 12232 3776 12296 3780
rect 12312 3836 12376 3840
rect 12312 3780 12316 3836
rect 12316 3780 12372 3836
rect 12372 3780 12376 3836
rect 12312 3776 12376 3780
rect 16520 3836 16584 3840
rect 16520 3780 16524 3836
rect 16524 3780 16580 3836
rect 16580 3780 16584 3836
rect 16520 3776 16584 3780
rect 16600 3836 16664 3840
rect 16600 3780 16604 3836
rect 16604 3780 16660 3836
rect 16660 3780 16664 3836
rect 16600 3776 16664 3780
rect 16680 3836 16744 3840
rect 16680 3780 16684 3836
rect 16684 3780 16740 3836
rect 16740 3780 16744 3836
rect 16680 3776 16744 3780
rect 16760 3836 16824 3840
rect 16760 3780 16764 3836
rect 16764 3780 16820 3836
rect 16820 3780 16824 3836
rect 16760 3776 16824 3780
rect 5400 3292 5464 3296
rect 5400 3236 5404 3292
rect 5404 3236 5460 3292
rect 5460 3236 5464 3292
rect 5400 3232 5464 3236
rect 5480 3292 5544 3296
rect 5480 3236 5484 3292
rect 5484 3236 5540 3292
rect 5540 3236 5544 3292
rect 5480 3232 5544 3236
rect 5560 3292 5624 3296
rect 5560 3236 5564 3292
rect 5564 3236 5620 3292
rect 5620 3236 5624 3292
rect 5560 3232 5624 3236
rect 5640 3292 5704 3296
rect 5640 3236 5644 3292
rect 5644 3236 5700 3292
rect 5700 3236 5704 3292
rect 5640 3232 5704 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 14296 3292 14360 3296
rect 14296 3236 14300 3292
rect 14300 3236 14356 3292
rect 14356 3236 14360 3292
rect 14296 3232 14360 3236
rect 14376 3292 14440 3296
rect 14376 3236 14380 3292
rect 14380 3236 14436 3292
rect 14436 3236 14440 3292
rect 14376 3232 14440 3236
rect 14456 3292 14520 3296
rect 14456 3236 14460 3292
rect 14460 3236 14516 3292
rect 14516 3236 14520 3292
rect 14456 3232 14520 3236
rect 14536 3292 14600 3296
rect 14536 3236 14540 3292
rect 14540 3236 14596 3292
rect 14596 3236 14600 3292
rect 14536 3232 14600 3236
rect 3176 2748 3240 2752
rect 3176 2692 3180 2748
rect 3180 2692 3236 2748
rect 3236 2692 3240 2748
rect 3176 2688 3240 2692
rect 3256 2748 3320 2752
rect 3256 2692 3260 2748
rect 3260 2692 3316 2748
rect 3316 2692 3320 2748
rect 3256 2688 3320 2692
rect 3336 2748 3400 2752
rect 3336 2692 3340 2748
rect 3340 2692 3396 2748
rect 3396 2692 3400 2748
rect 3336 2688 3400 2692
rect 3416 2748 3480 2752
rect 3416 2692 3420 2748
rect 3420 2692 3476 2748
rect 3476 2692 3480 2748
rect 3416 2688 3480 2692
rect 7624 2748 7688 2752
rect 7624 2692 7628 2748
rect 7628 2692 7684 2748
rect 7684 2692 7688 2748
rect 7624 2688 7688 2692
rect 7704 2748 7768 2752
rect 7704 2692 7708 2748
rect 7708 2692 7764 2748
rect 7764 2692 7768 2748
rect 7704 2688 7768 2692
rect 7784 2748 7848 2752
rect 7784 2692 7788 2748
rect 7788 2692 7844 2748
rect 7844 2692 7848 2748
rect 7784 2688 7848 2692
rect 7864 2748 7928 2752
rect 7864 2692 7868 2748
rect 7868 2692 7924 2748
rect 7924 2692 7928 2748
rect 7864 2688 7928 2692
rect 12072 2748 12136 2752
rect 12072 2692 12076 2748
rect 12076 2692 12132 2748
rect 12132 2692 12136 2748
rect 12072 2688 12136 2692
rect 12152 2748 12216 2752
rect 12152 2692 12156 2748
rect 12156 2692 12212 2748
rect 12212 2692 12216 2748
rect 12152 2688 12216 2692
rect 12232 2748 12296 2752
rect 12232 2692 12236 2748
rect 12236 2692 12292 2748
rect 12292 2692 12296 2748
rect 12232 2688 12296 2692
rect 12312 2748 12376 2752
rect 12312 2692 12316 2748
rect 12316 2692 12372 2748
rect 12372 2692 12376 2748
rect 12312 2688 12376 2692
rect 16520 2748 16584 2752
rect 16520 2692 16524 2748
rect 16524 2692 16580 2748
rect 16580 2692 16584 2748
rect 16520 2688 16584 2692
rect 16600 2748 16664 2752
rect 16600 2692 16604 2748
rect 16604 2692 16660 2748
rect 16660 2692 16664 2748
rect 16600 2688 16664 2692
rect 16680 2748 16744 2752
rect 16680 2692 16684 2748
rect 16684 2692 16740 2748
rect 16740 2692 16744 2748
rect 16680 2688 16744 2692
rect 16760 2748 16824 2752
rect 16760 2692 16764 2748
rect 16764 2692 16820 2748
rect 16820 2692 16824 2748
rect 16760 2688 16824 2692
rect 6684 2620 6748 2684
rect 5400 2204 5464 2208
rect 5400 2148 5404 2204
rect 5404 2148 5460 2204
rect 5460 2148 5464 2204
rect 5400 2144 5464 2148
rect 5480 2204 5544 2208
rect 5480 2148 5484 2204
rect 5484 2148 5540 2204
rect 5540 2148 5544 2204
rect 5480 2144 5544 2148
rect 5560 2204 5624 2208
rect 5560 2148 5564 2204
rect 5564 2148 5620 2204
rect 5620 2148 5624 2204
rect 5560 2144 5624 2148
rect 5640 2204 5704 2208
rect 5640 2148 5644 2204
rect 5644 2148 5700 2204
rect 5700 2148 5704 2204
rect 5640 2144 5704 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 14296 2204 14360 2208
rect 14296 2148 14300 2204
rect 14300 2148 14356 2204
rect 14356 2148 14360 2204
rect 14296 2144 14360 2148
rect 14376 2204 14440 2208
rect 14376 2148 14380 2204
rect 14380 2148 14436 2204
rect 14436 2148 14440 2204
rect 14376 2144 14440 2148
rect 14456 2204 14520 2208
rect 14456 2148 14460 2204
rect 14460 2148 14516 2204
rect 14516 2148 14520 2204
rect 14456 2144 14520 2148
rect 14536 2204 14600 2208
rect 14536 2148 14540 2204
rect 14540 2148 14596 2204
rect 14596 2148 14600 2204
rect 14536 2144 14600 2148
<< metal4 >>
rect 3168 14720 3488 14736
rect 3168 14656 3176 14720
rect 3240 14656 3256 14720
rect 3320 14656 3336 14720
rect 3400 14656 3416 14720
rect 3480 14656 3488 14720
rect 3003 14380 3069 14381
rect 3003 14316 3004 14380
rect 3068 14316 3069 14380
rect 3003 14315 3069 14316
rect 3006 12450 3066 14315
rect 2822 12390 3066 12450
rect 3168 13632 3488 14656
rect 3168 13568 3176 13632
rect 3240 13568 3256 13632
rect 3320 13568 3336 13632
rect 3400 13568 3416 13632
rect 3480 13568 3488 13632
rect 3168 12544 3488 13568
rect 3168 12480 3176 12544
rect 3240 12480 3256 12544
rect 3320 12480 3336 12544
rect 3400 12480 3416 12544
rect 3480 12480 3488 12544
rect 2822 5541 2882 12390
rect 3003 11660 3069 11661
rect 3003 11596 3004 11660
rect 3068 11596 3069 11660
rect 3003 11595 3069 11596
rect 3006 7309 3066 11595
rect 3168 11456 3488 12480
rect 3168 11392 3176 11456
rect 3240 11392 3256 11456
rect 3320 11392 3336 11456
rect 3400 11392 3416 11456
rect 3480 11392 3488 11456
rect 3168 10368 3488 11392
rect 3168 10304 3176 10368
rect 3240 10304 3256 10368
rect 3320 10304 3336 10368
rect 3400 10304 3416 10368
rect 3480 10304 3488 10368
rect 3168 9280 3488 10304
rect 3168 9216 3176 9280
rect 3240 9216 3256 9280
rect 3320 9216 3336 9280
rect 3400 9216 3416 9280
rect 3480 9216 3488 9280
rect 3168 8192 3488 9216
rect 3168 8128 3176 8192
rect 3240 8128 3256 8192
rect 3320 8128 3336 8192
rect 3400 8128 3416 8192
rect 3480 8128 3488 8192
rect 3003 7308 3069 7309
rect 3003 7244 3004 7308
rect 3068 7244 3069 7308
rect 3003 7243 3069 7244
rect 3168 7104 3488 8128
rect 3168 7040 3176 7104
rect 3240 7040 3256 7104
rect 3320 7040 3336 7104
rect 3400 7040 3416 7104
rect 3480 7040 3488 7104
rect 3168 6016 3488 7040
rect 3168 5952 3176 6016
rect 3240 5952 3256 6016
rect 3320 5952 3336 6016
rect 3400 5952 3416 6016
rect 3480 5952 3488 6016
rect 2819 5540 2885 5541
rect 2819 5476 2820 5540
rect 2884 5476 2885 5540
rect 2819 5475 2885 5476
rect 3168 4928 3488 5952
rect 3168 4864 3176 4928
rect 3240 4864 3256 4928
rect 3320 4864 3336 4928
rect 3400 4864 3416 4928
rect 3480 4864 3488 4928
rect 3168 3840 3488 4864
rect 3168 3776 3176 3840
rect 3240 3776 3256 3840
rect 3320 3776 3336 3840
rect 3400 3776 3416 3840
rect 3480 3776 3488 3840
rect 3168 2752 3488 3776
rect 3168 2688 3176 2752
rect 3240 2688 3256 2752
rect 3320 2688 3336 2752
rect 3400 2688 3416 2752
rect 3480 2688 3488 2752
rect 3168 2128 3488 2688
rect 5392 14176 5712 14736
rect 5392 14112 5400 14176
rect 5464 14112 5480 14176
rect 5544 14112 5560 14176
rect 5624 14112 5640 14176
rect 5704 14112 5712 14176
rect 5392 13088 5712 14112
rect 7616 14720 7936 14736
rect 7616 14656 7624 14720
rect 7688 14656 7704 14720
rect 7768 14656 7784 14720
rect 7848 14656 7864 14720
rect 7928 14656 7936 14720
rect 6683 13836 6749 13837
rect 6683 13772 6684 13836
rect 6748 13772 6749 13836
rect 6683 13771 6749 13772
rect 5392 13024 5400 13088
rect 5464 13024 5480 13088
rect 5544 13024 5560 13088
rect 5624 13024 5640 13088
rect 5704 13024 5712 13088
rect 5392 12000 5712 13024
rect 5392 11936 5400 12000
rect 5464 11936 5480 12000
rect 5544 11936 5560 12000
rect 5624 11936 5640 12000
rect 5704 11936 5712 12000
rect 5392 10912 5712 11936
rect 5392 10848 5400 10912
rect 5464 10848 5480 10912
rect 5544 10848 5560 10912
rect 5624 10848 5640 10912
rect 5704 10848 5712 10912
rect 5392 9824 5712 10848
rect 5392 9760 5400 9824
rect 5464 9760 5480 9824
rect 5544 9760 5560 9824
rect 5624 9760 5640 9824
rect 5704 9760 5712 9824
rect 5392 8736 5712 9760
rect 5392 8672 5400 8736
rect 5464 8672 5480 8736
rect 5544 8672 5560 8736
rect 5624 8672 5640 8736
rect 5704 8672 5712 8736
rect 5392 7648 5712 8672
rect 5392 7584 5400 7648
rect 5464 7584 5480 7648
rect 5544 7584 5560 7648
rect 5624 7584 5640 7648
rect 5704 7584 5712 7648
rect 5392 6560 5712 7584
rect 5392 6496 5400 6560
rect 5464 6496 5480 6560
rect 5544 6496 5560 6560
rect 5624 6496 5640 6560
rect 5704 6496 5712 6560
rect 5392 5472 5712 6496
rect 5392 5408 5400 5472
rect 5464 5408 5480 5472
rect 5544 5408 5560 5472
rect 5624 5408 5640 5472
rect 5704 5408 5712 5472
rect 5392 4384 5712 5408
rect 5392 4320 5400 4384
rect 5464 4320 5480 4384
rect 5544 4320 5560 4384
rect 5624 4320 5640 4384
rect 5704 4320 5712 4384
rect 5392 3296 5712 4320
rect 5392 3232 5400 3296
rect 5464 3232 5480 3296
rect 5544 3232 5560 3296
rect 5624 3232 5640 3296
rect 5704 3232 5712 3296
rect 5392 2208 5712 3232
rect 6686 2685 6746 13771
rect 7616 13632 7936 14656
rect 9840 14176 10160 14736
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 8707 13836 8773 13837
rect 8707 13772 8708 13836
rect 8772 13772 8773 13836
rect 8707 13771 8773 13772
rect 7616 13568 7624 13632
rect 7688 13568 7704 13632
rect 7768 13568 7784 13632
rect 7848 13568 7864 13632
rect 7928 13568 7936 13632
rect 7616 12544 7936 13568
rect 7616 12480 7624 12544
rect 7688 12480 7704 12544
rect 7768 12480 7784 12544
rect 7848 12480 7864 12544
rect 7928 12480 7936 12544
rect 7616 11456 7936 12480
rect 7616 11392 7624 11456
rect 7688 11392 7704 11456
rect 7768 11392 7784 11456
rect 7848 11392 7864 11456
rect 7928 11392 7936 11456
rect 7616 10368 7936 11392
rect 7616 10304 7624 10368
rect 7688 10304 7704 10368
rect 7768 10304 7784 10368
rect 7848 10304 7864 10368
rect 7928 10304 7936 10368
rect 7616 9280 7936 10304
rect 7616 9216 7624 9280
rect 7688 9216 7704 9280
rect 7768 9216 7784 9280
rect 7848 9216 7864 9280
rect 7928 9216 7936 9280
rect 7616 8192 7936 9216
rect 7616 8128 7624 8192
rect 7688 8128 7704 8192
rect 7768 8128 7784 8192
rect 7848 8128 7864 8192
rect 7928 8128 7936 8192
rect 7616 7104 7936 8128
rect 7616 7040 7624 7104
rect 7688 7040 7704 7104
rect 7768 7040 7784 7104
rect 7848 7040 7864 7104
rect 7928 7040 7936 7104
rect 7616 6016 7936 7040
rect 7616 5952 7624 6016
rect 7688 5952 7704 6016
rect 7768 5952 7784 6016
rect 7848 5952 7864 6016
rect 7928 5952 7936 6016
rect 7616 4928 7936 5952
rect 7616 4864 7624 4928
rect 7688 4864 7704 4928
rect 7768 4864 7784 4928
rect 7848 4864 7864 4928
rect 7928 4864 7936 4928
rect 7616 3840 7936 4864
rect 8710 4045 8770 13771
rect 9840 13088 10160 14112
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 12000 10160 13024
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9627 11116 9693 11117
rect 9627 11052 9628 11116
rect 9692 11052 9693 11116
rect 9627 11051 9693 11052
rect 9630 4725 9690 11051
rect 9840 10912 10160 11936
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 9824 10160 10848
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 8736 10160 9760
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 6560 10160 7584
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 5472 10160 6496
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9627 4724 9693 4725
rect 9627 4660 9628 4724
rect 9692 4660 9693 4724
rect 9627 4659 9693 4660
rect 9840 4384 10160 5408
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 8707 4044 8773 4045
rect 8707 3980 8708 4044
rect 8772 3980 8773 4044
rect 8707 3979 8773 3980
rect 7616 3776 7624 3840
rect 7688 3776 7704 3840
rect 7768 3776 7784 3840
rect 7848 3776 7864 3840
rect 7928 3776 7936 3840
rect 7616 2752 7936 3776
rect 7616 2688 7624 2752
rect 7688 2688 7704 2752
rect 7768 2688 7784 2752
rect 7848 2688 7864 2752
rect 7928 2688 7936 2752
rect 6683 2684 6749 2685
rect 6683 2620 6684 2684
rect 6748 2620 6749 2684
rect 6683 2619 6749 2620
rect 5392 2144 5400 2208
rect 5464 2144 5480 2208
rect 5544 2144 5560 2208
rect 5624 2144 5640 2208
rect 5704 2144 5712 2208
rect 5392 2128 5712 2144
rect 7616 2128 7936 2688
rect 9840 3296 10160 4320
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 2208 10160 3232
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 12064 14720 12384 14736
rect 12064 14656 12072 14720
rect 12136 14656 12152 14720
rect 12216 14656 12232 14720
rect 12296 14656 12312 14720
rect 12376 14656 12384 14720
rect 12064 13632 12384 14656
rect 12064 13568 12072 13632
rect 12136 13568 12152 13632
rect 12216 13568 12232 13632
rect 12296 13568 12312 13632
rect 12376 13568 12384 13632
rect 12064 12544 12384 13568
rect 12064 12480 12072 12544
rect 12136 12480 12152 12544
rect 12216 12480 12232 12544
rect 12296 12480 12312 12544
rect 12376 12480 12384 12544
rect 12064 11456 12384 12480
rect 12064 11392 12072 11456
rect 12136 11392 12152 11456
rect 12216 11392 12232 11456
rect 12296 11392 12312 11456
rect 12376 11392 12384 11456
rect 12064 10368 12384 11392
rect 12064 10304 12072 10368
rect 12136 10304 12152 10368
rect 12216 10304 12232 10368
rect 12296 10304 12312 10368
rect 12376 10304 12384 10368
rect 12064 9280 12384 10304
rect 12064 9216 12072 9280
rect 12136 9216 12152 9280
rect 12216 9216 12232 9280
rect 12296 9216 12312 9280
rect 12376 9216 12384 9280
rect 12064 8192 12384 9216
rect 12064 8128 12072 8192
rect 12136 8128 12152 8192
rect 12216 8128 12232 8192
rect 12296 8128 12312 8192
rect 12376 8128 12384 8192
rect 12064 7104 12384 8128
rect 12064 7040 12072 7104
rect 12136 7040 12152 7104
rect 12216 7040 12232 7104
rect 12296 7040 12312 7104
rect 12376 7040 12384 7104
rect 12064 6016 12384 7040
rect 12064 5952 12072 6016
rect 12136 5952 12152 6016
rect 12216 5952 12232 6016
rect 12296 5952 12312 6016
rect 12376 5952 12384 6016
rect 12064 4928 12384 5952
rect 12064 4864 12072 4928
rect 12136 4864 12152 4928
rect 12216 4864 12232 4928
rect 12296 4864 12312 4928
rect 12376 4864 12384 4928
rect 12064 3840 12384 4864
rect 12064 3776 12072 3840
rect 12136 3776 12152 3840
rect 12216 3776 12232 3840
rect 12296 3776 12312 3840
rect 12376 3776 12384 3840
rect 12064 2752 12384 3776
rect 12064 2688 12072 2752
rect 12136 2688 12152 2752
rect 12216 2688 12232 2752
rect 12296 2688 12312 2752
rect 12376 2688 12384 2752
rect 12064 2128 12384 2688
rect 14288 14176 14608 14736
rect 14288 14112 14296 14176
rect 14360 14112 14376 14176
rect 14440 14112 14456 14176
rect 14520 14112 14536 14176
rect 14600 14112 14608 14176
rect 14288 13088 14608 14112
rect 14288 13024 14296 13088
rect 14360 13024 14376 13088
rect 14440 13024 14456 13088
rect 14520 13024 14536 13088
rect 14600 13024 14608 13088
rect 14288 12000 14608 13024
rect 14288 11936 14296 12000
rect 14360 11936 14376 12000
rect 14440 11936 14456 12000
rect 14520 11936 14536 12000
rect 14600 11936 14608 12000
rect 14288 10912 14608 11936
rect 14288 10848 14296 10912
rect 14360 10848 14376 10912
rect 14440 10848 14456 10912
rect 14520 10848 14536 10912
rect 14600 10848 14608 10912
rect 14288 9824 14608 10848
rect 14288 9760 14296 9824
rect 14360 9760 14376 9824
rect 14440 9760 14456 9824
rect 14520 9760 14536 9824
rect 14600 9760 14608 9824
rect 14288 8736 14608 9760
rect 14288 8672 14296 8736
rect 14360 8672 14376 8736
rect 14440 8672 14456 8736
rect 14520 8672 14536 8736
rect 14600 8672 14608 8736
rect 14288 7648 14608 8672
rect 14288 7584 14296 7648
rect 14360 7584 14376 7648
rect 14440 7584 14456 7648
rect 14520 7584 14536 7648
rect 14600 7584 14608 7648
rect 14288 6560 14608 7584
rect 14288 6496 14296 6560
rect 14360 6496 14376 6560
rect 14440 6496 14456 6560
rect 14520 6496 14536 6560
rect 14600 6496 14608 6560
rect 14288 5472 14608 6496
rect 14288 5408 14296 5472
rect 14360 5408 14376 5472
rect 14440 5408 14456 5472
rect 14520 5408 14536 5472
rect 14600 5408 14608 5472
rect 14288 4384 14608 5408
rect 14288 4320 14296 4384
rect 14360 4320 14376 4384
rect 14440 4320 14456 4384
rect 14520 4320 14536 4384
rect 14600 4320 14608 4384
rect 14288 3296 14608 4320
rect 14288 3232 14296 3296
rect 14360 3232 14376 3296
rect 14440 3232 14456 3296
rect 14520 3232 14536 3296
rect 14600 3232 14608 3296
rect 14288 2208 14608 3232
rect 14288 2144 14296 2208
rect 14360 2144 14376 2208
rect 14440 2144 14456 2208
rect 14520 2144 14536 2208
rect 14600 2144 14608 2208
rect 14288 2128 14608 2144
rect 16512 14720 16832 14736
rect 16512 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16760 14720
rect 16824 14656 16832 14720
rect 16512 13632 16832 14656
rect 16512 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16760 13632
rect 16824 13568 16832 13632
rect 16512 12544 16832 13568
rect 16512 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16760 12544
rect 16824 12480 16832 12544
rect 16512 11456 16832 12480
rect 17907 12340 17973 12341
rect 17907 12276 17908 12340
rect 17972 12276 17973 12340
rect 17907 12275 17973 12276
rect 16512 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16760 11456
rect 16824 11392 16832 11456
rect 16512 10368 16832 11392
rect 16512 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16760 10368
rect 16824 10304 16832 10368
rect 16512 9280 16832 10304
rect 16512 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16760 9280
rect 16824 9216 16832 9280
rect 16512 8192 16832 9216
rect 17910 8397 17970 12275
rect 17907 8396 17973 8397
rect 17907 8332 17908 8396
rect 17972 8332 17973 8396
rect 17907 8331 17973 8332
rect 16512 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16760 8192
rect 16824 8128 16832 8192
rect 16512 7104 16832 8128
rect 16512 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16760 7104
rect 16824 7040 16832 7104
rect 16512 6016 16832 7040
rect 16512 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16760 6016
rect 16824 5952 16832 6016
rect 16512 4928 16832 5952
rect 16512 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16760 4928
rect 16824 4864 16832 4928
rect 16512 3840 16832 4864
rect 16512 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16760 3840
rect 16824 3776 16832 3840
rect 16512 2752 16832 3776
rect 16512 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16760 2752
rect 16824 2688 16832 2752
rect 16512 2128 16832 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__18__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3956 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__19__A
timestamp 1649977179
transform -1 0 3588 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__20__A
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__21__A
timestamp 1649977179
transform -1 0 3772 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__22__A
timestamp 1649977179
transform -1 0 3956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__23__A
timestamp 1649977179
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__24__A
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__25__A
timestamp 1649977179
transform 1 0 4140 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__27__A
timestamp 1649977179
transform -1 0 3496 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__29__A
timestamp 1649977179
transform -1 0 3404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__31__A
timestamp 1649977179
transform 1 0 5888 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__33__A
timestamp 1649977179
transform -1 0 2208 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1649977179
transform -1 0 17572 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1649977179
transform 1 0 16376 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1649977179
transform 1 0 15916 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1649977179
transform -1 0 18124 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1649977179
transform 1 0 16836 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1649977179
transform -1 0 17940 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1649977179
transform 1 0 16928 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1649977179
transform 1 0 17296 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1649977179
transform 1 0 17204 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1649977179
transform -1 0 17848 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1649977179
transform -1 0 17388 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1649977179
transform -1 0 17940 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1649977179
transform 1 0 13892 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1649977179
transform 1 0 8372 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1649977179
transform 1 0 7544 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__80__A
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__81__A
timestamp 1649977179
transform 1 0 10120 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__85__A
timestamp 1649977179
transform -1 0 5244 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 7452 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 6532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 6808 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 5612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 3680 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 5980 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 6992 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 7176 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 4232 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 6808 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 5980 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 6164 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 5060 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 5796 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 4784 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 3680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 3680 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 4140 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 3956 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 3956 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 3956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 5428 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 2852 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 5796 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 17296 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 17664 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 16928 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 16376 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 16744 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 15180 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 16008 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 17480 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 17112 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 16928 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 15364 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 17020 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 17112 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 17204 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 16560 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 16100 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 17204 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 17020 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 17296 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 16560 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 11408 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 11592 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 13248 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 12512 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 14352 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 13432 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 13892 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 13984 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 12420 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 12604 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 13248 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 14536 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 9384 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1649977179
transform -1 0 10028 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1649977179
transform -1 0 10672 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1649977179
transform -1 0 11960 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 1932 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 2392 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 2944 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 3128 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 3956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 3312 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10396 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 10672 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 9660 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 10396 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 7544 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 3864 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 2668 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 4140 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 3404 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 4232 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 4048 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7728 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6716 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 8740 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 7544 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 4232 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 4600 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 7360 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 6532 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 13616 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 14168 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 17388 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 16376 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 17388 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 16744 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 17480 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 14444 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 8556 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 9752 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 16100 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 15732 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 14168 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 17756 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 17756 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14720 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 13892 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 15088 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 13984 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 13156 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 14168 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 14444 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 14536 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 16560 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 8556 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_W_FTB01_A
timestamp 1649977179
transform -1 0 1932 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2300 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18
timestamp 1649977179
transform 1 0 2760 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23
timestamp 1649977179
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33
timestamp 1649977179
transform 1 0 4140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38
timestamp 1649977179
transform 1 0 4600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43
timestamp 1649977179
transform 1 0 5060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63
timestamp 1649977179
transform 1 0 6900 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68
timestamp 1649977179
transform 1 0 7360 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73
timestamp 1649977179
transform 1 0 7820 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78
timestamp 1649977179
transform 1 0 8280 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1649977179
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93
timestamp 1649977179
transform 1 0 9660 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98
timestamp 1649977179
transform 1 0 10120 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103
timestamp 1649977179
transform 1 0 10580 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1649977179
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1649977179
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_189
timestamp 1649977179
transform 1 0 18492 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_34 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_45
timestamp 1649977179
transform 1 0 5244 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_49 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_158
timestamp 1649977179
transform 1 0 15640 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_33 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_45
timestamp 1649977179
transform 1 0 5244 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_49 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5612 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_57
timestamp 1649977179
transform 1 0 6348 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_65 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_69
timestamp 1649977179
transform 1 0 7452 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_73
timestamp 1649977179
transform 1 0 7820 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_88
timestamp 1649977179
transform 1 0 9200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_104
timestamp 1649977179
transform 1 0 10672 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_117
timestamp 1649977179
transform 1 0 11868 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_173
timestamp 1649977179
transform 1 0 17020 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_31
timestamp 1649977179
transform 1 0 3956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_43
timestamp 1649977179
transform 1 0 5060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_59
timestamp 1649977179
transform 1 0 6532 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_71
timestamp 1649977179
transform 1 0 7636 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_79
timestamp 1649977179
transform 1 0 8372 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_95
timestamp 1649977179
transform 1 0 9844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_106
timestamp 1649977179
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1649977179
transform 1 0 12236 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_178
timestamp 1649977179
transform 1 0 17480 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_35
timestamp 1649977179
transform 1 0 4324 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_70
timestamp 1649977179
transform 1 0 7544 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_114
timestamp 1649977179
transform 1 0 11592 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_128
timestamp 1649977179
transform 1 0 12880 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_136
timestamp 1649977179
transform 1 0 13616 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_147
timestamp 1649977179
transform 1 0 14628 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_44
timestamp 1649977179
transform 1 0 5152 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_83
timestamp 1649977179
transform 1 0 8740 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_92
timestamp 1649977179
transform 1 0 9568 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_104
timestamp 1649977179
transform 1 0 10672 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_124
timestamp 1649977179
transform 1 0 12512 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_178
timestamp 1649977179
transform 1 0 17480 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_32
timestamp 1649977179
transform 1 0 4048 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_36
timestamp 1649977179
transform 1 0 4416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_64
timestamp 1649977179
transform 1 0 6992 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_71
timestamp 1649977179
transform 1 0 7636 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_75
timestamp 1649977179
transform 1 0 8004 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_79
timestamp 1649977179
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_94
timestamp 1649977179
transform 1 0 9752 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_98
timestamp 1649977179
transform 1 0 10120 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_185
timestamp 1649977179
transform 1 0 18124 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_75
timestamp 1649977179
transform 1 0 8004 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_100
timestamp 1649977179
transform 1 0 10304 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_133
timestamp 1649977179
transform 1 0 13340 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_162
timestamp 1649977179
transform 1 0 16008 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_185
timestamp 1649977179
transform 1 0 18124 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_54
timestamp 1649977179
transform 1 0 6072 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_62
timestamp 1649977179
transform 1 0 6808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_81
timestamp 1649977179
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_105
timestamp 1649977179
transform 1 0 10764 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_156
timestamp 1649977179
transform 1 0 15456 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1649977179
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_77
timestamp 1649977179
transform 1 0 8188 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_135
timestamp 1649977179
transform 1 0 13524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_159
timestamp 1649977179
transform 1 0 15732 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_165
timestamp 1649977179
transform 1 0 16284 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_178
timestamp 1649977179
transform 1 0 17480 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_185
timestamp 1649977179
transform 1 0 18124 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1649977179
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_79
timestamp 1649977179
transform 1 0 8372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_101
timestamp 1649977179
transform 1 0 10396 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_118
timestamp 1649977179
transform 1 0 11960 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1649977179
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_158
timestamp 1649977179
transform 1 0 15640 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_170
timestamp 1649977179
transform 1 0 16744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_176
timestamp 1649977179
transform 1 0 17296 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_181
timestamp 1649977179
transform 1 0 17756 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_185
timestamp 1649977179
transform 1 0 18124 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_33
timestamp 1649977179
transform 1 0 4140 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_73
timestamp 1649977179
transform 1 0 7820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_85
timestamp 1649977179
transform 1 0 8924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1649977179
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_145
timestamp 1649977179
transform 1 0 14444 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_153
timestamp 1649977179
transform 1 0 15180 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1649977179
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_14
timestamp 1649977179
transform 1 0 2392 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_63
timestamp 1649977179
transform 1 0 6900 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_67
timestamp 1649977179
transform 1 0 7268 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_114
timestamp 1649977179
transform 1 0 11592 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_134
timestamp 1649977179
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_155
timestamp 1649977179
transform 1 0 15364 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_171
timestamp 1649977179
transform 1 0 16836 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_183
timestamp 1649977179
transform 1 0 17940 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_28
timestamp 1649977179
transform 1 0 3680 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1649977179
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_65
timestamp 1649977179
transform 1 0 7084 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_97
timestamp 1649977179
transform 1 0 10028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1649977179
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_133
timestamp 1649977179
transform 1 0 13340 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_145
timestamp 1649977179
transform 1 0 14444 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_157
timestamp 1649977179
transform 1 0 15548 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 1649977179
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_185
timestamp 1649977179
transform 1 0 18124 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_19
timestamp 1649977179
transform 1 0 2852 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_33
timestamp 1649977179
transform 1 0 4140 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_75
timestamp 1649977179
transform 1 0 8004 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_102
timestamp 1649977179
transform 1 0 10488 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_110
timestamp 1649977179
transform 1 0 11224 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_128
timestamp 1649977179
transform 1 0 12880 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_185
timestamp 1649977179
transform 1 0 18124 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_13
timestamp 1649977179
transform 1 0 2300 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_36
timestamp 1649977179
transform 1 0 4416 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_61
timestamp 1649977179
transform 1 0 6716 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_94
timestamp 1649977179
transform 1 0 9752 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_156
timestamp 1649977179
transform 1 0 15456 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_164
timestamp 1649977179
transform 1 0 16192 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_31
timestamp 1649977179
transform 1 0 3956 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_69
timestamp 1649977179
transform 1 0 7452 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_96
timestamp 1649977179
transform 1 0 9936 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_108
timestamp 1649977179
transform 1 0 11040 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_114
timestamp 1649977179
transform 1 0 11592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_131
timestamp 1649977179
transform 1 0 13156 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_159
timestamp 1649977179
transform 1 0 15732 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_19
timestamp 1649977179
transform 1 0 2852 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_40
timestamp 1649977179
transform 1 0 4784 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_46
timestamp 1649977179
transform 1 0 5336 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_59
timestamp 1649977179
transform 1 0 6532 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_103
timestamp 1649977179
transform 1 0 10580 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1649977179
transform 1 0 12236 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_133
timestamp 1649977179
transform 1 0 13340 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_145
timestamp 1649977179
transform 1 0 14444 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_179
timestamp 1649977179
transform 1 0 17572 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_47
timestamp 1649977179
transform 1 0 5428 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_104
timestamp 1649977179
transform 1 0 10672 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_115
timestamp 1649977179
transform 1 0 11684 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_136
timestamp 1649977179
transform 1 0 13616 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_155
timestamp 1649977179
transform 1 0 15364 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_163
timestamp 1649977179
transform 1 0 16100 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_170
timestamp 1649977179
transform 1 0 16744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1649977179
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_63
timestamp 1649977179
transform 1 0 6900 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_75
timestamp 1649977179
transform 1 0 8004 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_103
timestamp 1649977179
transform 1 0 10580 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1649977179
transform 1 0 12420 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_127
timestamp 1649977179
transform 1 0 12788 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_150
timestamp 1649977179
transform 1 0 14904 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_162
timestamp 1649977179
transform 1 0 16008 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_43
timestamp 1649977179
transform 1 0 5060 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_71
timestamp 1649977179
transform 1 0 7636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_100
timestamp 1649977179
transform 1 0 10304 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_106
timestamp 1649977179
transform 1 0 10856 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_128
timestamp 1649977179
transform 1 0 12880 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_136
timestamp 1649977179
transform 1 0 13616 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_161
timestamp 1649977179
transform 1 0 15916 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_33
timestamp 1649977179
transform 1 0 4140 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_40
timestamp 1649977179
transform 1 0 4784 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_66
timestamp 1649977179
transform 1 0 7176 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_72
timestamp 1649977179
transform 1 0 7728 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_83
timestamp 1649977179
transform 1 0 8740 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_100
timestamp 1649977179
transform 1 0 10304 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_115
timestamp 1649977179
transform 1 0 11684 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_123
timestamp 1649977179
transform 1 0 12420 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_127
timestamp 1649977179
transform 1 0 12788 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_131
timestamp 1649977179
transform 1 0 13156 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_135
timestamp 1649977179
transform 1 0 13524 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_141
timestamp 1649977179
transform 1 0 14076 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_153
timestamp 1649977179
transform 1 0 15180 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_159
timestamp 1649977179
transform 1 0 15732 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_23
timestamp 1649977179
transform 1 0 3220 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_55
timestamp 1649977179
transform 1 0 6164 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_66
timestamp 1649977179
transform 1 0 7176 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_72
timestamp 1649977179
transform 1 0 7728 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_80
timestamp 1649977179
transform 1 0 8464 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1649977179
transform 1 0 9660 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_100
timestamp 1649977179
transform 1 0 10304 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_107
timestamp 1649977179
transform 1 0 10948 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_111
timestamp 1649977179
transform 1 0 11316 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_128
timestamp 1649977179
transform 1 0 12880 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_135
timestamp 1649977179
transform 1 0 13524 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_146
timestamp 1649977179
transform 1 0 14536 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_150
timestamp 1649977179
transform 1 0 14904 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_169
timestamp 1649977179
transform 1 0 16652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 6256 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 16560 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _18_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3128 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _19_
timestamp 1649977179
transform 1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _20_
timestamp 1649977179
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _21_
timestamp 1649977179
transform 1 0 2392 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _22_
timestamp 1649977179
transform 1 0 2116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 1649977179
transform 1 0 3220 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _24_
timestamp 1649977179
transform 1 0 2944 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _25_
timestamp 1649977179
transform 1 0 2116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _26_
timestamp 1649977179
transform 1 0 2576 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _27_
timestamp 1649977179
transform 1 0 1748 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _28_
timestamp 1649977179
transform 1 0 2300 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _29_
timestamp 1649977179
transform -1 0 2392 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _30_
timestamp 1649977179
transform 1 0 4324 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _31_
timestamp 1649977179
transform 1 0 4140 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _32_
timestamp 1649977179
transform 1 0 3220 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _33_
timestamp 1649977179
transform 1 0 1748 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _34_
timestamp 1649977179
transform 1 0 2300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1649977179
transform -1 0 16376 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _36_
timestamp 1649977179
transform 1 0 17572 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _37_
timestamp 1649977179
transform -1 0 16836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp 1649977179
transform 1 0 17572 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1649977179
transform -1 0 17112 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1649977179
transform -1 0 18124 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp 1649977179
transform -1 0 17940 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1649977179
transform -1 0 17664 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _43_
timestamp 1649977179
transform -1 0 17848 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _44_
timestamp 1649977179
transform -1 0 17296 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _45_
timestamp 1649977179
transform -1 0 17848 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _46_
timestamp 1649977179
transform -1 0 17388 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _47_
timestamp 1649977179
transform -1 0 17848 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1649977179
transform -1 0 17756 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1649977179
transform 1 0 17848 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1649977179
transform -1 0 17848 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1649977179
transform -1 0 18124 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1649977179
transform -1 0 17664 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1649977179
transform -1 0 17848 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1649977179
transform -1 0 18124 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1649977179
transform -1 0 7084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1649977179
transform -1 0 7084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1649977179
transform -1 0 7360 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1649977179
transform 1 0 9292 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1649977179
transform 1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1649977179
transform 1 0 10120 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1649977179
transform -1 0 10672 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 1649977179
transform 1 0 16100 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1649977179
transform -1 0 13064 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1649977179
transform -1 0 15732 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1649977179
transform -1 0 16928 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1649977179
transform -1 0 17204 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1649977179
transform -1 0 17480 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1649977179
transform -1 0 17664 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1649977179
transform -1 0 17388 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1649977179
transform 1 0 17940 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp 1649977179
transform 1 0 13248 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp 1649977179
transform 1 0 12512 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _75_
timestamp 1649977179
transform 1 0 13616 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _76_
timestamp 1649977179
transform 1 0 14904 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _77_
timestamp 1649977179
transform 1 0 8096 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _78_
timestamp 1649977179
transform 1 0 7820 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _79_
timestamp 1649977179
transform 1 0 7268 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _80_
timestamp 1649977179
transform 1 0 11040 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _81_
timestamp 1649977179
transform 1 0 9844 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _82_
timestamp 1649977179
transform -1 0 6624 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _83_
timestamp 1649977179
transform -1 0 6256 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _84_
timestamp 1649977179
transform 1 0 2668 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _85_
timestamp 1649977179
transform 1 0 4508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _86_
timestamp 1649977179
transform 1 0 2392 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10672 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1649977179
transform 1 0 6164 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1649977179
transform -1 0 11224 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1649977179
transform -1 0 11408 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1649977179
transform 1 0 8464 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1649977179
transform -1 0 8832 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1649977179
transform 1 0 11316 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 7728 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 6256 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform 1 0 6348 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform 1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 2392 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2300 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1649977179
transform -1 0 2300 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1649977179
transform -1 0 2300 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1649977179
transform -1 0 3220 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1649977179
transform -1 0 3220 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1649977179
transform -1 0 3220 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1649977179
transform -1 0 4692 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 1649977179
transform -1 0 3220 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1649977179
transform -1 0 4140 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1649977179
transform 1 0 4692 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input16 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 3496 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1649977179
transform -1 0 2300 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1649977179
transform -1 0 2300 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1649977179
transform -1 0 2300 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1649977179
transform -1 0 2300 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1649977179
transform 1 0 2300 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1649977179
transform -1 0 2300 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform 1 0 18032 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1649977179
transform -1 0 17664 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1649977179
transform 1 0 17664 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1649977179
transform 1 0 17664 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input30
timestamp 1649977179
transform 1 0 16744 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform 1 0 16008 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1649977179
transform -1 0 17296 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1649977179
transform 1 0 16744 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1649977179
transform -1 0 16560 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform 1 0 15364 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1649977179
transform -1 0 18584 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform 1 0 18308 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1649977179
transform -1 0 18584 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1649977179
transform 1 0 17664 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1649977179
transform 1 0 17664 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input41
timestamp 1649977179
transform 1 0 17664 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1649977179
transform 1 0 17664 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43
timestamp 1649977179
transform 1 0 17664 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp 1649977179
transform 1 0 17664 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1649977179
transform 1 0 11592 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1649977179
transform 1 0 12512 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1649977179
transform -1 0 13892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1649977179
transform -1 0 13708 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1649977179
transform 1 0 13892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1649977179
transform 1 0 14352 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1649977179
transform 1 0 16744 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1649977179
transform -1 0 12236 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1649977179
transform 1 0 12604 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1649977179
transform -1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1649977179
transform -1 0 14352 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1649977179
transform 1 0 9384 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1649977179
transform -1 0 10304 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1649977179
transform 1 0 10672 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1649977179
transform 1 0 11500 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7544 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 9292 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 9108 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 8740 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10304 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1649977179
transform 1 0 9568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1649977179
transform -1 0 11224 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1649977179
transform 1 0 8280 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 9108 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6532 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1649977179
transform 1 0 11040 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1649977179
transform -1 0 13432 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1649977179
transform -1 0 7636 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8188 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1649977179
transform 1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1649977179
transform 1 0 11776 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1649977179
transform 1 0 8188 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 10120 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6900 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1649977179
transform 1 0 12236 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1649977179
transform -1 0 13984 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform -1 0 11592 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1649977179
transform 1 0 13064 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1649977179
transform -1 0 9568 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 12328 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10672 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1649977179
transform 1 0 13432 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1649977179
transform 1 0 10764 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 12144 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9292 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1649977179
transform -1 0 15640 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1649977179
transform 1 0 14168 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1649977179
transform 1 0 10212 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 14720 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13892 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1649977179
transform 1 0 14352 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1649977179
transform -1 0 16560 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1649977179
transform 1 0 10304 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 16008 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12420 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 4508 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4416 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11592 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10488 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 9752 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 6256 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 7820 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5980 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 5428 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4508 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 5428 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8004 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 5888 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 5980 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4508 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 6256 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4508 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 8556 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7360 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11684 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12880 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6808 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9016 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 10488 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11868 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 12052 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13432 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12972 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 12972 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 9844 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12972 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13340 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 12052 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3036 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1649977179
transform -1 0 3588 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 1932 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3128 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2208 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2300 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_0.mux_l2_in_3__149 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2116 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1649977179
transform 1 0 2208 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1649977179
transform 1 0 1472 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9568 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9660 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 9568 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8740 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7728 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1649977179
transform 1 0 6808 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_1.mux_l2_in_3__150
timestamp 1649977179
transform -1 0 6716 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6624 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1649977179
transform 1 0 5152 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4784 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3680 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_1_
timestamp 1649977179
transform 1 0 3404 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_2_
timestamp 1649977179
transform 1 0 3036 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2208 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 2576 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2392 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1649977179
transform 1 0 3220 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_2.mux_l2_in_3__151
timestamp 1649977179
transform -1 0 3220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1649977179
transform -1 0 2208 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1649977179
transform 1 0 2024 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1649977179
transform -1 0 2300 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6900 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7728 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1649977179
transform 1 0 5428 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6072 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4416 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1649977179
transform 1 0 3496 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_3.mux_l2_in_3__152
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1649977179
transform -1 0 3680 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3956 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1649977179
transform 1 0 2944 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1649977179
transform -1 0 3404 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3128 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6164 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1649977179
transform -1 0 6164 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6532 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 6164 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6256 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1649977179
transform 1 0 13616 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_4.mux_l2_in_3__153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14444 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 6256 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1649977179
transform 1 0 12788 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1649977179
transform 1 0 7360 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 5336 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16560 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 16744 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16100 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14628 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1649977179
transform 1 0 8740 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_5.mux_l2_in_3__154
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 9200 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1649977179
transform -1 0 8740 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1649977179
transform 1 0 15456 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_1_
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_2_
timestamp 1649977179
transform 1 0 15272 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15180 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1649977179
transform -1 0 15180 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_6.mux_l2_in_3__155
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1649977179
transform 1 0 16560 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14352 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1649977179
transform 1 0 15732 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1649977179
transform 1 0 13524 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 5336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1649977179
transform 1 0 13892 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1649977179
transform -1 0 13156 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1649977179
transform 1 0 13064 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12788 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1649977179
transform 1 0 11776 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_7.mux_l2_in_3__156
timestamp 1649977179
transform 1 0 12604 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1649977179
transform 1 0 11592 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1649977179
transform 1 0 11960 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1649977179
transform 1 0 10948 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1649977179
transform 1 0 10856 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 6532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 15364 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1649977179
transform 1 0 15456 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1649977179
transform -1 0 15180 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1649977179
transform -1 0 15640 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1649977179
transform -1 0 15456 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1649977179
transform -1 0 15548 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_8.mux_l2_in_3__157
timestamp 1649977179
transform -1 0 15364 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 15548 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14904 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1649977179
transform 1 0 14904 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1649977179
transform 1 0 14076 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 4784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output63 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform 1 0 6808 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform 1 0 2576 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform -1 0 3680 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform -1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform -1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform -1 0 5060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform -1 0 2576 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform -1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform -1 0 2760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform -1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform -1 0 5980 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform -1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform -1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform -1 0 2668 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform 1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform -1 0 2116 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform -1 0 1748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform -1 0 2116 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform -1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform -1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform -1 0 3312 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform 1 0 3312 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform -1 0 2116 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform -1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform -1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform -1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform -1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform -1 0 2116 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform 1 0 17112 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform 1 0 17848 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform 1 0 18216 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform 1 0 18216 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform 1 0 18216 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform 1 0 17848 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform 1 0 18216 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform 1 0 18216 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1649977179
transform 1 0 18216 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1649977179
transform 1 0 17848 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1649977179
transform 1 0 18216 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1649977179
transform -1 0 17480 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1649977179
transform 1 0 16744 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1649977179
transform 1 0 17480 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1649977179
transform 1 0 17480 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1649977179
transform 1 0 18216 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1649977179
transform 1 0 17848 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1649977179
transform 1 0 18216 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1649977179
transform 1 0 18216 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1649977179
transform 1 0 18216 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1649977179
transform 1 0 6992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1649977179
transform 1 0 7912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1649977179
transform -1 0 8740 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1649977179
transform -1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1649977179
transform -1 0 9660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1649977179
transform -1 0 10120 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1649977179
transform -1 0 10580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1649977179
transform 1 0 10672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1649977179
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1649977179
transform 1 0 15732 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1649977179
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1649977179
transform 1 0 17388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1649977179
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1649977179
transform 1 0 17848 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1649977179
transform 1 0 17848 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output133
timestamp 1649977179
transform 1 0 3956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1649977179
transform -1 0 3680 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1649977179
transform -1 0 4600 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1649977179
transform -1 0 5244 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1649977179
transform -1 0 5980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1649977179
transform -1 0 4876 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1649977179
transform -1 0 5612 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1649977179
transform -1 0 4508 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1649977179
transform -1 0 4140 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1649977179
transform -1 0 3588 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2208 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater143
timestamp 1649977179
transform 1 0 4232 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater144
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater145
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater146
timestamp 1649977179
transform 1 0 3864 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater147
timestamp 1649977179
transform -1 0 9752 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater148
timestamp 1649977179
transform -1 0 8372 0 1 5440
box -38 -48 314 592
<< labels >>
flabel metal2 s 7378 16400 7434 17200 0 FreeSans 224 90 0 0 IO_ISOL_N
port 0 nsew signal input
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 SC_IN_BOT
port 1 nsew signal input
flabel metal2 s 6090 16400 6146 17200 0 FreeSans 224 90 0 0 SC_IN_TOP
port 2 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 SC_OUT_BOT
port 3 nsew signal tristate
flabel metal2 s 6734 16400 6790 17200 0 FreeSans 224 90 0 0 SC_OUT_TOP
port 4 nsew signal tristate
flabel metal4 s 5392 2128 5712 14736 0 FreeSans 1920 90 0 0 VGND
port 5 nsew ground bidirectional
flabel metal4 s 9840 2128 10160 14736 0 FreeSans 1920 90 0 0 VGND
port 5 nsew ground bidirectional
flabel metal4 s 14288 2128 14608 14736 0 FreeSans 1920 90 0 0 VGND
port 5 nsew ground bidirectional
flabel metal4 s 3168 2128 3488 14736 0 FreeSans 1920 90 0 0 VPWR
port 6 nsew power bidirectional
flabel metal4 s 7616 2128 7936 14736 0 FreeSans 1920 90 0 0 VPWR
port 6 nsew power bidirectional
flabel metal4 s 12064 2128 12384 14736 0 FreeSans 1920 90 0 0 VPWR
port 6 nsew power bidirectional
flabel metal4 s 16512 2128 16832 14736 0 FreeSans 1920 90 0 0 VPWR
port 6 nsew power bidirectional
flabel metal2 s 938 0 994 800 0 FreeSans 224 90 0 0 bottom_grid_pin_0_
port 7 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 bottom_grid_pin_10_
port 8 nsew signal tristate
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 bottom_grid_pin_12_
port 9 nsew signal tristate
flabel metal2 s 4158 0 4214 800 0 FreeSans 224 90 0 0 bottom_grid_pin_14_
port 10 nsew signal tristate
flabel metal2 s 4618 0 4674 800 0 FreeSans 224 90 0 0 bottom_grid_pin_16_
port 11 nsew signal tristate
flabel metal2 s 1398 0 1454 800 0 FreeSans 224 90 0 0 bottom_grid_pin_2_
port 12 nsew signal tristate
flabel metal2 s 1858 0 1914 800 0 FreeSans 224 90 0 0 bottom_grid_pin_4_
port 13 nsew signal tristate
flabel metal2 s 2318 0 2374 800 0 FreeSans 224 90 0 0 bottom_grid_pin_6_
port 14 nsew signal tristate
flabel metal2 s 2778 0 2834 800 0 FreeSans 224 90 0 0 bottom_grid_pin_8_
port 15 nsew signal tristate
flabel metal2 s 5078 0 5134 800 0 FreeSans 224 90 0 0 ccff_head
port 16 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 ccff_tail
port 17 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 18 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 19 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 20 nsew signal input
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 21 nsew signal input
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 22 nsew signal input
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 23 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 24 nsew signal input
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 25 nsew signal input
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 26 nsew signal input
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 27 nsew signal input
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 28 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 29 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 30 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 31 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 32 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 33 nsew signal input
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 34 nsew signal input
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 35 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 36 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 37 nsew signal input
flabel metal3 s 0 688 800 808 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 38 nsew signal tristate
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 39 nsew signal tristate
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 40 nsew signal tristate
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 41 nsew signal tristate
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 42 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 43 nsew signal tristate
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 44 nsew signal tristate
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 45 nsew signal tristate
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 46 nsew signal tristate
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 47 nsew signal tristate
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 48 nsew signal tristate
flabel metal3 s 0 1096 800 1216 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 49 nsew signal tristate
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 50 nsew signal tristate
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 51 nsew signal tristate
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 52 nsew signal tristate
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 53 nsew signal tristate
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 54 nsew signal tristate
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 55 nsew signal tristate
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 56 nsew signal tristate
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 57 nsew signal tristate
flabel metal3 s 19200 8712 20000 8832 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 58 nsew signal input
flabel metal3 s 19200 12792 20000 12912 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 59 nsew signal input
flabel metal3 s 19200 13200 20000 13320 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 60 nsew signal input
flabel metal3 s 19200 13608 20000 13728 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 61 nsew signal input
flabel metal3 s 19200 14016 20000 14136 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 62 nsew signal input
flabel metal3 s 19200 14424 20000 14544 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 63 nsew signal input
flabel metal3 s 19200 14832 20000 14952 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 64 nsew signal input
flabel metal3 s 19200 15240 20000 15360 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 65 nsew signal input
flabel metal3 s 19200 15648 20000 15768 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 66 nsew signal input
flabel metal3 s 19200 16056 20000 16176 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 67 nsew signal input
flabel metal3 s 19200 16464 20000 16584 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 68 nsew signal input
flabel metal3 s 19200 9120 20000 9240 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 69 nsew signal input
flabel metal3 s 19200 9528 20000 9648 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 70 nsew signal input
flabel metal3 s 19200 9936 20000 10056 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 71 nsew signal input
flabel metal3 s 19200 10344 20000 10464 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 72 nsew signal input
flabel metal3 s 19200 10752 20000 10872 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 73 nsew signal input
flabel metal3 s 19200 11160 20000 11280 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 74 nsew signal input
flabel metal3 s 19200 11568 20000 11688 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 75 nsew signal input
flabel metal3 s 19200 11976 20000 12096 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 76 nsew signal input
flabel metal3 s 19200 12384 20000 12504 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 77 nsew signal input
flabel metal3 s 19200 552 20000 672 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 78 nsew signal tristate
flabel metal3 s 19200 4632 20000 4752 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 79 nsew signal tristate
flabel metal3 s 19200 5040 20000 5160 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 80 nsew signal tristate
flabel metal3 s 19200 5448 20000 5568 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 81 nsew signal tristate
flabel metal3 s 19200 5856 20000 5976 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 82 nsew signal tristate
flabel metal3 s 19200 6264 20000 6384 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 83 nsew signal tristate
flabel metal3 s 19200 6672 20000 6792 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 84 nsew signal tristate
flabel metal3 s 19200 7080 20000 7200 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 85 nsew signal tristate
flabel metal3 s 19200 7488 20000 7608 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 86 nsew signal tristate
flabel metal3 s 19200 7896 20000 8016 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 87 nsew signal tristate
flabel metal3 s 19200 8304 20000 8424 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 88 nsew signal tristate
flabel metal3 s 19200 960 20000 1080 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 89 nsew signal tristate
flabel metal3 s 19200 1368 20000 1488 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 90 nsew signal tristate
flabel metal3 s 19200 1776 20000 1896 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 91 nsew signal tristate
flabel metal3 s 19200 2184 20000 2304 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 92 nsew signal tristate
flabel metal3 s 19200 2592 20000 2712 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 93 nsew signal tristate
flabel metal3 s 19200 3000 20000 3120 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 94 nsew signal tristate
flabel metal3 s 19200 3408 20000 3528 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 95 nsew signal tristate
flabel metal3 s 19200 3816 20000 3936 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 96 nsew signal tristate
flabel metal3 s 19200 4224 20000 4344 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 97 nsew signal tristate
flabel metal2 s 6918 0 6974 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
port 98 nsew signal tristate
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
port 99 nsew signal tristate
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
port 100 nsew signal tristate
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
port 101 nsew signal tristate
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
port 102 nsew signal tristate
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
port 103 nsew signal tristate
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
port 104 nsew signal tristate
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
port 105 nsew signal tristate
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
port 106 nsew signal tristate
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
port 107 nsew signal input
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
port 108 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
port 109 nsew signal input
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
port 110 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
port 111 nsew signal input
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
port 112 nsew signal input
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
port 113 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
port 114 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
port 115 nsew signal input
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
port 116 nsew signal tristate
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
port 117 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
port 118 nsew signal tristate
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
port 119 nsew signal tristate
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
port 120 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
port 121 nsew signal tristate
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
port 122 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
port 123 nsew signal tristate
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
port 124 nsew signal tristate
flabel metal2 s 8022 16400 8078 17200 0 FreeSans 224 90 0 0 prog_clk_0_N_in
port 125 nsew signal input
flabel metal3 s 0 280 800 400 0 FreeSans 480 0 0 0 prog_clk_0_W_out
port 126 nsew signal tristate
flabel metal2 s 8666 16400 8722 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_0_
port 127 nsew signal input
flabel metal2 s 11886 16400 11942 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_10_
port 128 nsew signal input
flabel metal2 s 19614 16400 19670 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_11_lower
port 129 nsew signal tristate
flabel metal2 s 3514 16400 3570 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_11_upper
port 130 nsew signal tristate
flabel metal2 s 12530 16400 12586 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_12_
port 131 nsew signal input
flabel metal2 s 14462 16400 14518 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_13_lower
port 132 nsew signal tristate
flabel metal2 s 4158 16400 4214 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_13_upper
port 133 nsew signal tristate
flabel metal2 s 13174 16400 13230 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_14_
port 134 nsew signal input
flabel metal2 s 15106 16400 15162 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_15_lower
port 135 nsew signal tristate
flabel metal2 s 4802 16400 4858 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_15_upper
port 136 nsew signal tristate
flabel metal2 s 13818 16400 13874 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_16_
port 137 nsew signal input
flabel metal2 s 15750 16400 15806 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_17_lower
port 138 nsew signal tristate
flabel metal2 s 5446 16400 5502 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_17_upper
port 139 nsew signal tristate
flabel metal2 s 16394 16400 16450 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_1_lower
port 140 nsew signal tristate
flabel metal2 s 294 16400 350 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_1_upper
port 141 nsew signal tristate
flabel metal2 s 9310 16400 9366 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_2_
port 142 nsew signal input
flabel metal2 s 17038 16400 17094 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_3_lower
port 143 nsew signal tristate
flabel metal2 s 938 16400 994 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_3_upper
port 144 nsew signal tristate
flabel metal2 s 9954 16400 10010 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_4_
port 145 nsew signal input
flabel metal2 s 17682 16400 17738 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_5_lower
port 146 nsew signal tristate
flabel metal2 s 1582 16400 1638 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_5_upper
port 147 nsew signal tristate
flabel metal2 s 10598 16400 10654 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_6_
port 148 nsew signal input
flabel metal2 s 18326 16400 18382 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_7_lower
port 149 nsew signal tristate
flabel metal2 s 2226 16400 2282 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_7_upper
port 150 nsew signal tristate
flabel metal2 s 11242 16400 11298 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_8_
port 151 nsew signal input
flabel metal2 s 18970 16400 19026 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_9_lower
port 152 nsew signal tristate
flabel metal2 s 2870 16400 2926 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_9_upper
port 153 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 20000 17200
<< end >>
