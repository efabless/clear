magic
tech sky130A
magscale 1 2
timestamp 1656942944
<< obsli1 >>
rect 1104 2159 16008 17425
<< obsm1 >>
rect 1104 2128 16008 17944
<< metal2 >>
rect 1214 19200 1270 20000
rect 1582 19200 1638 20000
rect 1950 19200 2006 20000
rect 2318 19200 2374 20000
rect 2686 19200 2742 20000
rect 3054 19200 3110 20000
rect 3422 19200 3478 20000
rect 3790 19200 3846 20000
rect 4158 19200 4214 20000
rect 4526 19200 4582 20000
rect 4894 19200 4950 20000
rect 5262 19200 5318 20000
rect 5630 19200 5686 20000
rect 5998 19200 6054 20000
rect 6366 19200 6422 20000
rect 6734 19200 6790 20000
rect 7102 19200 7158 20000
rect 7470 19200 7526 20000
rect 7838 19200 7894 20000
rect 8206 19200 8262 20000
rect 8574 19200 8630 20000
rect 8942 19200 8998 20000
rect 9310 19200 9366 20000
rect 9678 19200 9734 20000
rect 10046 19200 10102 20000
rect 10414 19200 10470 20000
rect 10782 19200 10838 20000
rect 11150 19200 11206 20000
rect 11518 19200 11574 20000
rect 11886 19200 11942 20000
rect 12254 19200 12310 20000
rect 12622 19200 12678 20000
rect 12990 19200 13046 20000
rect 13358 19200 13414 20000
rect 13726 19200 13782 20000
rect 14094 19200 14150 20000
rect 14462 19200 14518 20000
rect 14830 19200 14886 20000
rect 15198 19200 15254 20000
rect 15566 19200 15622 20000
rect 15934 19200 15990 20000
rect 1398 0 1454 800
rect 1766 0 1822 800
rect 2134 0 2190 800
rect 2502 0 2558 800
rect 2870 0 2926 800
rect 3238 0 3294 800
rect 3606 0 3662 800
rect 3974 0 4030 800
rect 4342 0 4398 800
rect 4710 0 4766 800
rect 5078 0 5134 800
rect 5446 0 5502 800
rect 5814 0 5870 800
rect 6182 0 6238 800
rect 6550 0 6606 800
rect 6918 0 6974 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 8022 0 8078 800
rect 8390 0 8446 800
rect 8758 0 8814 800
rect 9126 0 9182 800
rect 9494 0 9550 800
rect 9862 0 9918 800
rect 10230 0 10286 800
rect 10598 0 10654 800
rect 10966 0 11022 800
rect 11334 0 11390 800
rect 11702 0 11758 800
rect 12070 0 12126 800
rect 12438 0 12494 800
rect 12806 0 12862 800
rect 13174 0 13230 800
rect 13542 0 13598 800
rect 13910 0 13966 800
rect 14278 0 14334 800
rect 14646 0 14702 800
rect 15014 0 15070 800
rect 15382 0 15438 800
rect 15750 0 15806 800
<< obsm2 >>
rect 1326 19144 1526 19258
rect 1694 19144 1894 19258
rect 2062 19144 2262 19258
rect 2430 19144 2630 19258
rect 2798 19144 2998 19258
rect 3166 19144 3366 19258
rect 3534 19144 3734 19258
rect 3902 19144 4102 19258
rect 4270 19144 4470 19258
rect 4638 19144 4838 19258
rect 5006 19144 5206 19258
rect 5374 19144 5574 19258
rect 5742 19144 5942 19258
rect 6110 19144 6310 19258
rect 6478 19144 6678 19258
rect 6846 19144 7046 19258
rect 7214 19144 7414 19258
rect 7582 19144 7782 19258
rect 7950 19144 8150 19258
rect 8318 19144 8518 19258
rect 8686 19144 8886 19258
rect 9054 19144 9254 19258
rect 9422 19144 9622 19258
rect 9790 19144 9990 19258
rect 10158 19144 10358 19258
rect 10526 19144 10726 19258
rect 10894 19144 11094 19258
rect 11262 19144 11462 19258
rect 11630 19144 11830 19258
rect 11998 19144 12198 19258
rect 12366 19144 12566 19258
rect 12734 19144 12934 19258
rect 13102 19144 13302 19258
rect 13470 19144 13670 19258
rect 13838 19144 14038 19258
rect 14206 19144 14406 19258
rect 14574 19144 14774 19258
rect 14942 19144 15142 19258
rect 15310 19144 15510 19258
rect 15678 19144 15878 19258
rect 1216 856 15988 19144
rect 1216 734 1342 856
rect 1510 734 1710 856
rect 1878 734 2078 856
rect 2246 734 2446 856
rect 2614 734 2814 856
rect 2982 734 3182 856
rect 3350 734 3550 856
rect 3718 734 3918 856
rect 4086 734 4286 856
rect 4454 734 4654 856
rect 4822 734 5022 856
rect 5190 734 5390 856
rect 5558 734 5758 856
rect 5926 734 6126 856
rect 6294 734 6494 856
rect 6662 734 6862 856
rect 7030 734 7230 856
rect 7398 734 7598 856
rect 7766 734 7966 856
rect 8134 734 8334 856
rect 8502 734 8702 856
rect 8870 734 9070 856
rect 9238 734 9438 856
rect 9606 734 9806 856
rect 9974 734 10174 856
rect 10342 734 10542 856
rect 10710 734 10910 856
rect 11078 734 11278 856
rect 11446 734 11646 856
rect 11814 734 12014 856
rect 12182 734 12382 856
rect 12550 734 12750 856
rect 12918 734 13118 856
rect 13286 734 13486 856
rect 13654 734 13854 856
rect 14022 734 14222 856
rect 14390 734 14590 856
rect 14758 734 14958 856
rect 15126 734 15326 856
rect 15494 734 15694 856
rect 15862 734 15988 856
<< metal3 >>
rect 0 18096 800 18216
rect 16400 17280 17200 17400
rect 0 14832 800 14952
rect 16400 12384 17200 12504
rect 0 11568 800 11688
rect 0 8304 800 8424
rect 16400 7488 17200 7608
rect 0 5040 800 5160
rect 16400 2592 17200 2712
rect 0 1776 800 1896
<< obsm3 >>
rect 880 18016 16400 18189
rect 800 17480 16400 18016
rect 800 17200 16320 17480
rect 800 15032 16400 17200
rect 880 14752 16400 15032
rect 800 12584 16400 14752
rect 800 12304 16320 12584
rect 800 11768 16400 12304
rect 880 11488 16400 11768
rect 800 8504 16400 11488
rect 880 8224 16400 8504
rect 800 7688 16400 8224
rect 800 7408 16320 7688
rect 800 5240 16400 7408
rect 880 4960 16400 5240
rect 800 2792 16400 4960
rect 800 2512 16320 2792
rect 800 1976 16400 2512
rect 880 1803 16400 1976
<< metal4 >>
rect 2818 2128 3138 17456
rect 4692 2128 5012 17456
rect 6566 2128 6886 17456
rect 8440 2128 8760 17456
rect 10314 2128 10634 17456
rect 12188 2128 12508 17456
rect 14062 2128 14382 17456
<< obsm4 >>
rect 8891 9691 8957 11253
<< labels >>
rlabel metal2 s 1214 19200 1270 20000 6 IO_ISOL_N
port 1 nsew signal input
rlabel metal4 s 4692 2128 5012 17456 6 VGND
port 2 nsew ground bidirectional
rlabel metal4 s 8440 2128 8760 17456 6 VGND
port 2 nsew ground bidirectional
rlabel metal4 s 12188 2128 12508 17456 6 VGND
port 2 nsew ground bidirectional
rlabel metal4 s 2818 2128 3138 17456 6 VPWR
port 3 nsew power bidirectional
rlabel metal4 s 6566 2128 6886 17456 6 VPWR
port 3 nsew power bidirectional
rlabel metal4 s 10314 2128 10634 17456 6 VPWR
port 3 nsew power bidirectional
rlabel metal4 s 14062 2128 14382 17456 6 VPWR
port 3 nsew power bidirectional
rlabel metal3 s 0 18096 800 18216 6 ccff_head
port 4 nsew signal input
rlabel metal3 s 16400 12384 17200 12504 6 ccff_tail
port 5 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 chany_bottom_in[0]
port 6 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 chany_bottom_in[10]
port 7 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 chany_bottom_in[11]
port 8 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 chany_bottom_in[12]
port 9 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 chany_bottom_in[13]
port 10 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 chany_bottom_in[14]
port 11 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 chany_bottom_in[15]
port 12 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 chany_bottom_in[16]
port 13 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 chany_bottom_in[17]
port 14 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 chany_bottom_in[18]
port 15 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 chany_bottom_in[19]
port 16 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 chany_bottom_in[1]
port 17 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 chany_bottom_in[2]
port 18 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 chany_bottom_in[3]
port 19 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 chany_bottom_in[4]
port 20 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 chany_bottom_in[5]
port 21 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 chany_bottom_in[6]
port 22 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 chany_bottom_in[7]
port 23 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 chany_bottom_in[8]
port 24 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 chany_bottom_in[9]
port 25 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 chany_bottom_out[0]
port 26 nsew signal output
rlabel metal2 s 5078 0 5134 800 6 chany_bottom_out[10]
port 27 nsew signal output
rlabel metal2 s 5446 0 5502 800 6 chany_bottom_out[11]
port 28 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 chany_bottom_out[12]
port 29 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 chany_bottom_out[13]
port 30 nsew signal output
rlabel metal2 s 6550 0 6606 800 6 chany_bottom_out[14]
port 31 nsew signal output
rlabel metal2 s 6918 0 6974 800 6 chany_bottom_out[15]
port 32 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 chany_bottom_out[16]
port 33 nsew signal output
rlabel metal2 s 7654 0 7710 800 6 chany_bottom_out[17]
port 34 nsew signal output
rlabel metal2 s 8022 0 8078 800 6 chany_bottom_out[18]
port 35 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 chany_bottom_out[19]
port 36 nsew signal output
rlabel metal2 s 1766 0 1822 800 6 chany_bottom_out[1]
port 37 nsew signal output
rlabel metal2 s 2134 0 2190 800 6 chany_bottom_out[2]
port 38 nsew signal output
rlabel metal2 s 2502 0 2558 800 6 chany_bottom_out[3]
port 39 nsew signal output
rlabel metal2 s 2870 0 2926 800 6 chany_bottom_out[4]
port 40 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 chany_bottom_out[5]
port 41 nsew signal output
rlabel metal2 s 3606 0 3662 800 6 chany_bottom_out[6]
port 42 nsew signal output
rlabel metal2 s 3974 0 4030 800 6 chany_bottom_out[7]
port 43 nsew signal output
rlabel metal2 s 4342 0 4398 800 6 chany_bottom_out[8]
port 44 nsew signal output
rlabel metal2 s 4710 0 4766 800 6 chany_bottom_out[9]
port 45 nsew signal output
rlabel metal2 s 8942 19200 8998 20000 6 chany_top_in[0]
port 46 nsew signal input
rlabel metal2 s 12622 19200 12678 20000 6 chany_top_in[10]
port 47 nsew signal input
rlabel metal2 s 12990 19200 13046 20000 6 chany_top_in[11]
port 48 nsew signal input
rlabel metal2 s 13358 19200 13414 20000 6 chany_top_in[12]
port 49 nsew signal input
rlabel metal2 s 13726 19200 13782 20000 6 chany_top_in[13]
port 50 nsew signal input
rlabel metal2 s 14094 19200 14150 20000 6 chany_top_in[14]
port 51 nsew signal input
rlabel metal2 s 14462 19200 14518 20000 6 chany_top_in[15]
port 52 nsew signal input
rlabel metal2 s 14830 19200 14886 20000 6 chany_top_in[16]
port 53 nsew signal input
rlabel metal2 s 15198 19200 15254 20000 6 chany_top_in[17]
port 54 nsew signal input
rlabel metal2 s 15566 19200 15622 20000 6 chany_top_in[18]
port 55 nsew signal input
rlabel metal2 s 15934 19200 15990 20000 6 chany_top_in[19]
port 56 nsew signal input
rlabel metal2 s 9310 19200 9366 20000 6 chany_top_in[1]
port 57 nsew signal input
rlabel metal2 s 9678 19200 9734 20000 6 chany_top_in[2]
port 58 nsew signal input
rlabel metal2 s 10046 19200 10102 20000 6 chany_top_in[3]
port 59 nsew signal input
rlabel metal2 s 10414 19200 10470 20000 6 chany_top_in[4]
port 60 nsew signal input
rlabel metal2 s 10782 19200 10838 20000 6 chany_top_in[5]
port 61 nsew signal input
rlabel metal2 s 11150 19200 11206 20000 6 chany_top_in[6]
port 62 nsew signal input
rlabel metal2 s 11518 19200 11574 20000 6 chany_top_in[7]
port 63 nsew signal input
rlabel metal2 s 11886 19200 11942 20000 6 chany_top_in[8]
port 64 nsew signal input
rlabel metal2 s 12254 19200 12310 20000 6 chany_top_in[9]
port 65 nsew signal input
rlabel metal2 s 1582 19200 1638 20000 6 chany_top_out[0]
port 66 nsew signal output
rlabel metal2 s 5262 19200 5318 20000 6 chany_top_out[10]
port 67 nsew signal output
rlabel metal2 s 5630 19200 5686 20000 6 chany_top_out[11]
port 68 nsew signal output
rlabel metal2 s 5998 19200 6054 20000 6 chany_top_out[12]
port 69 nsew signal output
rlabel metal2 s 6366 19200 6422 20000 6 chany_top_out[13]
port 70 nsew signal output
rlabel metal2 s 6734 19200 6790 20000 6 chany_top_out[14]
port 71 nsew signal output
rlabel metal2 s 7102 19200 7158 20000 6 chany_top_out[15]
port 72 nsew signal output
rlabel metal2 s 7470 19200 7526 20000 6 chany_top_out[16]
port 73 nsew signal output
rlabel metal2 s 7838 19200 7894 20000 6 chany_top_out[17]
port 74 nsew signal output
rlabel metal2 s 8206 19200 8262 20000 6 chany_top_out[18]
port 75 nsew signal output
rlabel metal2 s 8574 19200 8630 20000 6 chany_top_out[19]
port 76 nsew signal output
rlabel metal2 s 1950 19200 2006 20000 6 chany_top_out[1]
port 77 nsew signal output
rlabel metal2 s 2318 19200 2374 20000 6 chany_top_out[2]
port 78 nsew signal output
rlabel metal2 s 2686 19200 2742 20000 6 chany_top_out[3]
port 79 nsew signal output
rlabel metal2 s 3054 19200 3110 20000 6 chany_top_out[4]
port 80 nsew signal output
rlabel metal2 s 3422 19200 3478 20000 6 chany_top_out[5]
port 81 nsew signal output
rlabel metal2 s 3790 19200 3846 20000 6 chany_top_out[6]
port 82 nsew signal output
rlabel metal2 s 4158 19200 4214 20000 6 chany_top_out[7]
port 83 nsew signal output
rlabel metal2 s 4526 19200 4582 20000 6 chany_top_out[8]
port 84 nsew signal output
rlabel metal2 s 4894 19200 4950 20000 6 chany_top_out[9]
port 85 nsew signal output
rlabel metal3 s 0 8304 800 8424 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 86 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 87 nsew signal input
rlabel metal3 s 0 14832 800 14952 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 88 nsew signal output
rlabel metal3 s 0 5040 800 5160 6 left_grid_pin_0_
port 89 nsew signal output
rlabel metal3 s 16400 7488 17200 7608 6 prog_clk_0_E_in
port 90 nsew signal input
rlabel metal3 s 0 1776 800 1896 6 right_width_0_height_0__pin_0_
port 91 nsew signal input
rlabel metal3 s 16400 2592 17200 2712 6 right_width_0_height_0__pin_1_lower
port 92 nsew signal output
rlabel metal3 s 16400 17280 17200 17400 6 right_width_0_height_0__pin_1_upper
port 93 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 17200 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 452934
string GDS_FILE /home/marwan/clear_signoff_final/openlane/cby_0__1_/runs/cby_0__1_/results/signoff/cby_0__1_.magic.gds
string GDS_START 84912
<< end >>

